module dtc_split05_bm78 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node84;

	assign outp = (inp[3]) ? node62 : node1;
		assign node1 = (inp[4]) ? node27 : node2;
			assign node2 = (inp[0]) ? 3'b111 : node3;
				assign node3 = (inp[6]) ? node17 : node4;
					assign node4 = (inp[1]) ? node10 : node5;
						assign node5 = (inp[5]) ? node7 : 3'b010;
							assign node7 = (inp[10]) ? 3'b010 : 3'b000;
						assign node10 = (inp[5]) ? node14 : node11;
							assign node11 = (inp[2]) ? 3'b101 : 3'b001;
							assign node14 = (inp[11]) ? 3'b010 : 3'b100;
					assign node17 = (inp[9]) ? node21 : node18;
						assign node18 = (inp[1]) ? 3'b011 : 3'b010;
						assign node21 = (inp[11]) ? node23 : 3'b111;
							assign node23 = (inp[2]) ? 3'b011 : 3'b111;
			assign node27 = (inp[0]) ? node45 : node28;
				assign node28 = (inp[9]) ? node30 : 3'b000;
					assign node30 = (inp[2]) ? node38 : node31;
						assign node31 = (inp[5]) ? node35 : node32;
							assign node32 = (inp[1]) ? 3'b010 : 3'b000;
							assign node35 = (inp[1]) ? 3'b000 : 3'b100;
						assign node38 = (inp[8]) ? node42 : node39;
							assign node39 = (inp[1]) ? 3'b010 : 3'b000;
							assign node42 = (inp[7]) ? 3'b000 : 3'b000;
				assign node45 = (inp[9]) ? node53 : node46;
					assign node46 = (inp[6]) ? 3'b000 : node47;
						assign node47 = (inp[7]) ? 3'b110 : node48;
							assign node48 = (inp[5]) ? 3'b000 : 3'b001;
					assign node53 = (inp[1]) ? node59 : node54;
						assign node54 = (inp[6]) ? 3'b111 : node55;
							assign node55 = (inp[7]) ? 3'b101 : 3'b010;
						assign node59 = (inp[5]) ? 3'b101 : 3'b111;
		assign node62 = (inp[4]) ? 3'b000 : node63;
			assign node63 = (inp[0]) ? node71 : node64;
				assign node64 = (inp[11]) ? node66 : 3'b000;
					assign node66 = (inp[5]) ? node68 : 3'b000;
						assign node68 = (inp[9]) ? 3'b100 : 3'b000;
				assign node71 = (inp[9]) ? node77 : node72;
					assign node72 = (inp[6]) ? 3'b000 : node73;
						assign node73 = (inp[7]) ? 3'b100 : 3'b000;
					assign node77 = (inp[5]) ? node83 : node78;
						assign node78 = (inp[8]) ? node80 : 3'b101;
							assign node80 = (inp[1]) ? 3'b011 : 3'b010;
						assign node83 = (inp[10]) ? 3'b110 : node84;
							assign node84 = (inp[6]) ? 3'b101 : 3'b100;

endmodule