module dtc_split5_bm90 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node227;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node247;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node271;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node290;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node305;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node318;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node332;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node341;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node350;
	wire [3-1:0] node353;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node368;
	wire [3-1:0] node371;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node403;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node414;
	wire [3-1:0] node417;
	wire [3-1:0] node419;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node431;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node441;
	wire [3-1:0] node443;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node459;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node465;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node476;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node489;
	wire [3-1:0] node491;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node510;
	wire [3-1:0] node512;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node528;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node535;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node557;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node571;
	wire [3-1:0] node574;
	wire [3-1:0] node576;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node583;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node595;
	wire [3-1:0] node598;
	wire [3-1:0] node601;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node612;
	wire [3-1:0] node613;
	wire [3-1:0] node617;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node624;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node641;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node649;
	wire [3-1:0] node653;
	wire [3-1:0] node654;
	wire [3-1:0] node656;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node666;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node694;
	wire [3-1:0] node695;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node703;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node733;
	wire [3-1:0] node735;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node742;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node760;
	wire [3-1:0] node762;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node772;
	wire [3-1:0] node775;
	wire [3-1:0] node778;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node785;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node793;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node803;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node815;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node822;
	wire [3-1:0] node824;
	wire [3-1:0] node826;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node843;
	wire [3-1:0] node846;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node857;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node870;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node879;
	wire [3-1:0] node883;
	wire [3-1:0] node885;
	wire [3-1:0] node887;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node901;
	wire [3-1:0] node904;
	wire [3-1:0] node906;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node914;
	wire [3-1:0] node915;
	wire [3-1:0] node917;
	wire [3-1:0] node919;
	wire [3-1:0] node922;
	wire [3-1:0] node924;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node930;
	wire [3-1:0] node934;
	wire [3-1:0] node935;
	wire [3-1:0] node938;
	wire [3-1:0] node940;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node945;
	wire [3-1:0] node948;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node955;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node967;
	wire [3-1:0] node968;
	wire [3-1:0] node969;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node979;
	wire [3-1:0] node983;
	wire [3-1:0] node985;
	wire [3-1:0] node987;
	wire [3-1:0] node990;
	wire [3-1:0] node991;
	wire [3-1:0] node992;
	wire [3-1:0] node995;
	wire [3-1:0] node998;
	wire [3-1:0] node1001;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1008;
	wire [3-1:0] node1010;
	wire [3-1:0] node1014;
	wire [3-1:0] node1015;
	wire [3-1:0] node1016;
	wire [3-1:0] node1017;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1026;
	wire [3-1:0] node1028;
	wire [3-1:0] node1031;
	wire [3-1:0] node1032;
	wire [3-1:0] node1033;
	wire [3-1:0] node1034;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1041;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1047;
	wire [3-1:0] node1049;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1057;
	wire [3-1:0] node1058;
	wire [3-1:0] node1059;
	wire [3-1:0] node1061;
	wire [3-1:0] node1063;
	wire [3-1:0] node1066;
	wire [3-1:0] node1067;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1078;
	wire [3-1:0] node1081;
	wire [3-1:0] node1082;
	wire [3-1:0] node1083;
	wire [3-1:0] node1087;
	wire [3-1:0] node1089;
	wire [3-1:0] node1092;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1095;
	wire [3-1:0] node1096;
	wire [3-1:0] node1099;
	wire [3-1:0] node1100;
	wire [3-1:0] node1103;
	wire [3-1:0] node1106;
	wire [3-1:0] node1107;
	wire [3-1:0] node1110;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1115;
	wire [3-1:0] node1116;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1123;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1130;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1138;
	wire [3-1:0] node1139;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1147;
	wire [3-1:0] node1150;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1156;
	wire [3-1:0] node1157;
	wire [3-1:0] node1161;
	wire [3-1:0] node1162;
	wire [3-1:0] node1165;
	wire [3-1:0] node1168;
	wire [3-1:0] node1169;
	wire [3-1:0] node1170;
	wire [3-1:0] node1172;
	wire [3-1:0] node1175;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1181;
	wire [3-1:0] node1184;
	wire [3-1:0] node1185;
	wire [3-1:0] node1187;
	wire [3-1:0] node1190;
	wire [3-1:0] node1192;
	wire [3-1:0] node1195;
	wire [3-1:0] node1196;
	wire [3-1:0] node1197;
	wire [3-1:0] node1198;
	wire [3-1:0] node1199;
	wire [3-1:0] node1204;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1207;
	wire [3-1:0] node1209;
	wire [3-1:0] node1212;
	wire [3-1:0] node1215;
	wire [3-1:0] node1216;
	wire [3-1:0] node1218;
	wire [3-1:0] node1219;
	wire [3-1:0] node1222;
	wire [3-1:0] node1226;
	wire [3-1:0] node1228;
	wire [3-1:0] node1230;
	wire [3-1:0] node1231;
	wire [3-1:0] node1235;
	wire [3-1:0] node1236;
	wire [3-1:0] node1237;
	wire [3-1:0] node1238;
	wire [3-1:0] node1240;
	wire [3-1:0] node1243;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1251;
	wire [3-1:0] node1252;
	wire [3-1:0] node1256;
	wire [3-1:0] node1257;
	wire [3-1:0] node1259;
	wire [3-1:0] node1261;
	wire [3-1:0] node1263;
	wire [3-1:0] node1266;
	wire [3-1:0] node1268;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1274;
	wire [3-1:0] node1275;
	wire [3-1:0] node1276;
	wire [3-1:0] node1279;
	wire [3-1:0] node1283;
	wire [3-1:0] node1285;
	wire [3-1:0] node1286;
	wire [3-1:0] node1290;
	wire [3-1:0] node1291;
	wire [3-1:0] node1294;
	wire [3-1:0] node1295;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1302;
	wire [3-1:0] node1303;
	wire [3-1:0] node1306;
	wire [3-1:0] node1309;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1312;
	wire [3-1:0] node1315;
	wire [3-1:0] node1319;
	wire [3-1:0] node1320;
	wire [3-1:0] node1324;
	wire [3-1:0] node1325;
	wire [3-1:0] node1326;
	wire [3-1:0] node1327;
	wire [3-1:0] node1328;
	wire [3-1:0] node1329;
	wire [3-1:0] node1330;
	wire [3-1:0] node1332;
	wire [3-1:0] node1333;
	wire [3-1:0] node1337;
	wire [3-1:0] node1339;
	wire [3-1:0] node1340;
	wire [3-1:0] node1341;
	wire [3-1:0] node1344;
	wire [3-1:0] node1348;
	wire [3-1:0] node1349;
	wire [3-1:0] node1350;
	wire [3-1:0] node1353;
	wire [3-1:0] node1356;
	wire [3-1:0] node1358;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1363;
	wire [3-1:0] node1364;
	wire [3-1:0] node1367;
	wire [3-1:0] node1369;
	wire [3-1:0] node1372;
	wire [3-1:0] node1374;
	wire [3-1:0] node1376;
	wire [3-1:0] node1378;
	wire [3-1:0] node1381;
	wire [3-1:0] node1382;
	wire [3-1:0] node1384;
	wire [3-1:0] node1388;
	wire [3-1:0] node1389;
	wire [3-1:0] node1390;
	wire [3-1:0] node1391;
	wire [3-1:0] node1392;
	wire [3-1:0] node1396;
	wire [3-1:0] node1397;
	wire [3-1:0] node1398;
	wire [3-1:0] node1402;
	wire [3-1:0] node1403;
	wire [3-1:0] node1407;
	wire [3-1:0] node1409;
	wire [3-1:0] node1410;
	wire [3-1:0] node1411;
	wire [3-1:0] node1414;
	wire [3-1:0] node1418;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1421;
	wire [3-1:0] node1422;
	wire [3-1:0] node1424;
	wire [3-1:0] node1428;
	wire [3-1:0] node1430;
	wire [3-1:0] node1432;
	wire [3-1:0] node1435;
	wire [3-1:0] node1436;
	wire [3-1:0] node1437;
	wire [3-1:0] node1441;
	wire [3-1:0] node1445;
	wire [3-1:0] node1446;
	wire [3-1:0] node1447;
	wire [3-1:0] node1448;
	wire [3-1:0] node1449;
	wire [3-1:0] node1450;
	wire [3-1:0] node1455;
	wire [3-1:0] node1457;
	wire [3-1:0] node1458;
	wire [3-1:0] node1460;
	wire [3-1:0] node1463;
	wire [3-1:0] node1464;
	wire [3-1:0] node1468;
	wire [3-1:0] node1470;
	wire [3-1:0] node1472;
	wire [3-1:0] node1473;
	wire [3-1:0] node1477;
	wire [3-1:0] node1478;
	wire [3-1:0] node1479;
	wire [3-1:0] node1481;
	wire [3-1:0] node1483;
	wire [3-1:0] node1484;
	wire [3-1:0] node1488;
	wire [3-1:0] node1489;
	wire [3-1:0] node1490;
	wire [3-1:0] node1493;
	wire [3-1:0] node1494;
	wire [3-1:0] node1495;
	wire [3-1:0] node1500;
	wire [3-1:0] node1501;
	wire [3-1:0] node1502;
	wire [3-1:0] node1506;
	wire [3-1:0] node1507;
	wire [3-1:0] node1511;
	wire [3-1:0] node1512;
	wire [3-1:0] node1513;
	wire [3-1:0] node1514;
	wire [3-1:0] node1516;
	wire [3-1:0] node1519;
	wire [3-1:0] node1522;
	wire [3-1:0] node1524;
	wire [3-1:0] node1527;
	wire [3-1:0] node1528;
	wire [3-1:0] node1529;
	wire [3-1:0] node1530;
	wire [3-1:0] node1531;
	wire [3-1:0] node1536;
	wire [3-1:0] node1539;
	wire [3-1:0] node1540;
	wire [3-1:0] node1543;
	wire [3-1:0] node1544;
	wire [3-1:0] node1547;
	wire [3-1:0] node1550;
	wire [3-1:0] node1551;
	wire [3-1:0] node1552;
	wire [3-1:0] node1553;
	wire [3-1:0] node1555;
	wire [3-1:0] node1556;
	wire [3-1:0] node1560;
	wire [3-1:0] node1561;
	wire [3-1:0] node1562;
	wire [3-1:0] node1563;
	wire [3-1:0] node1566;
	wire [3-1:0] node1569;
	wire [3-1:0] node1570;
	wire [3-1:0] node1573;
	wire [3-1:0] node1575;
	wire [3-1:0] node1578;
	wire [3-1:0] node1580;
	wire [3-1:0] node1581;
	wire [3-1:0] node1586;
	wire [3-1:0] node1587;
	wire [3-1:0] node1588;
	wire [3-1:0] node1589;
	wire [3-1:0] node1590;
	wire [3-1:0] node1595;
	wire [3-1:0] node1596;
	wire [3-1:0] node1597;
	wire [3-1:0] node1599;
	wire [3-1:0] node1600;
	wire [3-1:0] node1604;
	wire [3-1:0] node1605;
	wire [3-1:0] node1609;
	wire [3-1:0] node1610;
	wire [3-1:0] node1612;
	wire [3-1:0] node1616;
	wire [3-1:0] node1617;
	wire [3-1:0] node1618;
	wire [3-1:0] node1619;
	wire [3-1:0] node1621;
	wire [3-1:0] node1624;
	wire [3-1:0] node1626;
	wire [3-1:0] node1627;
	wire [3-1:0] node1631;
	wire [3-1:0] node1632;
	wire [3-1:0] node1633;
	wire [3-1:0] node1634;
	wire [3-1:0] node1638;
	wire [3-1:0] node1640;
	wire [3-1:0] node1643;
	wire [3-1:0] node1644;
	wire [3-1:0] node1645;
	wire [3-1:0] node1649;
	wire [3-1:0] node1651;
	wire [3-1:0] node1652;
	wire [3-1:0] node1655;
	wire [3-1:0] node1658;
	wire [3-1:0] node1659;
	wire [3-1:0] node1661;
	wire [3-1:0] node1662;
	wire [3-1:0] node1663;
	wire [3-1:0] node1664;
	wire [3-1:0] node1667;
	wire [3-1:0] node1672;
	wire [3-1:0] node1673;
	wire [3-1:0] node1674;
	wire [3-1:0] node1675;
	wire [3-1:0] node1676;
	wire [3-1:0] node1681;
	wire [3-1:0] node1682;
	wire [3-1:0] node1684;
	wire [3-1:0] node1688;
	wire [3-1:0] node1689;
	wire [3-1:0] node1692;
	wire [3-1:0] node1694;

	assign outp = (inp[0]) ? node720 : node1;
		assign node1 = (inp[6]) ? node57 : node2;
			assign node2 = (inp[3]) ? node14 : node3;
				assign node3 = (inp[7]) ? node5 : 3'b011;
					assign node5 = (inp[4]) ? node7 : 3'b011;
						assign node7 = (inp[8]) ? node9 : 3'b111;
							assign node9 = (inp[1]) ? node11 : 3'b111;
								assign node11 = (inp[2]) ? 3'b011 : 3'b111;
				assign node14 = (inp[7]) ? node16 : 3'b111;
					assign node16 = (inp[9]) ? 3'b111 : node17;
						assign node17 = (inp[1]) ? node25 : node18;
							assign node18 = (inp[4]) ? 3'b111 : node19;
								assign node19 = (inp[2]) ? node21 : 3'b111;
									assign node21 = (inp[8]) ? 3'b011 : 3'b111;
							assign node25 = (inp[4]) ? node43 : node26;
								assign node26 = (inp[8]) ? node34 : node27;
									assign node27 = (inp[5]) ? node29 : 3'b101;
										assign node29 = (inp[2]) ? 3'b101 : node30;
											assign node30 = (inp[10]) ? 3'b111 : 3'b011;
									assign node34 = (inp[11]) ? node38 : node35;
										assign node35 = (inp[2]) ? 3'b001 : 3'b101;
										assign node38 = (inp[2]) ? node40 : 3'b001;
											assign node40 = (inp[5]) ? 3'b001 : 3'b101;
								assign node43 = (inp[2]) ? node49 : node44;
									assign node44 = (inp[8]) ? node46 : 3'b111;
										assign node46 = (inp[5]) ? 3'b111 : 3'b011;
									assign node49 = (inp[5]) ? node53 : node50;
										assign node50 = (inp[8]) ? 3'b101 : 3'b011;
										assign node53 = (inp[8]) ? 3'b011 : 3'b111;
			assign node57 = (inp[3]) ? node393 : node58;
				assign node58 = (inp[7]) ? node230 : node59;
					assign node59 = (inp[4]) ? node167 : node60;
						assign node60 = (inp[1]) ? node112 : node61;
							assign node61 = (inp[11]) ? node89 : node62;
								assign node62 = (inp[2]) ? node68 : node63;
									assign node63 = (inp[9]) ? node65 : 3'b101;
										assign node65 = (inp[5]) ? 3'b001 : 3'b101;
									assign node68 = (inp[9]) ? node82 : node69;
										assign node69 = (inp[5]) ? node77 : node70;
											assign node70 = (inp[10]) ? node74 : node71;
												assign node71 = (inp[8]) ? 3'b101 : 3'b001;
												assign node74 = (inp[8]) ? 3'b001 : 3'b101;
											assign node77 = (inp[10]) ? node79 : 3'b101;
												assign node79 = (inp[8]) ? 3'b101 : 3'b001;
										assign node82 = (inp[8]) ? node84 : 3'b101;
											assign node84 = (inp[5]) ? node86 : 3'b101;
												assign node86 = (inp[10]) ? 3'b101 : 3'b001;
								assign node89 = (inp[10]) ? node95 : node90;
									assign node90 = (inp[5]) ? node92 : 3'b101;
										assign node92 = (inp[2]) ? 3'b101 : 3'b001;
									assign node95 = (inp[9]) ? node105 : node96;
										assign node96 = (inp[2]) ? node100 : node97;
											assign node97 = (inp[5]) ? 3'b101 : 3'b001;
											assign node100 = (inp[8]) ? node102 : 3'b001;
												assign node102 = (inp[5]) ? 3'b001 : 3'b101;
										assign node105 = (inp[8]) ? node107 : 3'b001;
											assign node107 = (inp[2]) ? node109 : 3'b001;
												assign node109 = (inp[5]) ? 3'b001 : 3'b101;
							assign node112 = (inp[2]) ? node138 : node113;
								assign node113 = (inp[9]) ? node127 : node114;
									assign node114 = (inp[11]) ? node118 : node115;
										assign node115 = (inp[10]) ? 3'b001 : 3'b101;
										assign node118 = (inp[10]) ? node122 : node119;
											assign node119 = (inp[8]) ? 3'b101 : 3'b001;
											assign node122 = (inp[5]) ? 3'b101 : node123;
												assign node123 = (inp[8]) ? 3'b001 : 3'b101;
									assign node127 = (inp[5]) ? node129 : 3'b001;
										assign node129 = (inp[8]) ? node133 : node130;
											assign node130 = (inp[11]) ? 3'b101 : 3'b001;
											assign node133 = (inp[10]) ? 3'b001 : node134;
												assign node134 = (inp[11]) ? 3'b001 : 3'b101;
								assign node138 = (inp[8]) ? node154 : node139;
									assign node139 = (inp[10]) ? node143 : node140;
										assign node140 = (inp[5]) ? 3'b101 : 3'b001;
										assign node143 = (inp[5]) ? node149 : node144;
											assign node144 = (inp[11]) ? node146 : 3'b101;
												assign node146 = (inp[9]) ? 3'b001 : 3'b101;
											assign node149 = (inp[11]) ? 3'b001 : node150;
												assign node150 = (inp[9]) ? 3'b101 : 3'b001;
									assign node154 = (inp[11]) ? node162 : node155;
										assign node155 = (inp[5]) ? node159 : node156;
											assign node156 = (inp[10]) ? 3'b010 : 3'b110;
											assign node159 = (inp[10]) ? 3'b110 : 3'b010;
										assign node162 = (inp[10]) ? 3'b110 : node163;
											assign node163 = (inp[9]) ? 3'b010 : 3'b110;
						assign node167 = (inp[9]) ? node207 : node168;
							assign node168 = (inp[1]) ? node186 : node169;
								assign node169 = (inp[5]) ? node183 : node170;
									assign node170 = (inp[10]) ? node176 : node171;
										assign node171 = (inp[2]) ? node173 : 3'b001;
											assign node173 = (inp[8]) ? 3'b111 : 3'b101;
										assign node176 = (inp[8]) ? node180 : node177;
											assign node177 = (inp[2]) ? 3'b001 : 3'b101;
											assign node180 = (inp[2]) ? 3'b101 : 3'b001;
									assign node183 = (inp[8]) ? 3'b001 : 3'b011;
								assign node186 = (inp[10]) ? node196 : node187;
									assign node187 = (inp[5]) ? node193 : node188;
										assign node188 = (inp[8]) ? 3'b011 : node189;
											assign node189 = (inp[2]) ? 3'b011 : 3'b111;
										assign node193 = (inp[2]) ? 3'b101 : 3'b111;
									assign node196 = (inp[8]) ? node204 : node197;
										assign node197 = (inp[2]) ? 3'b001 : node198;
											assign node198 = (inp[11]) ? 3'b001 : node199;
												assign node199 = (inp[5]) ? 3'b001 : 3'b011;
										assign node204 = (inp[11]) ? 3'b111 : 3'b011;
							assign node207 = (inp[1]) ? node213 : node208;
								assign node208 = (inp[10]) ? 3'b111 : node209;
									assign node209 = (inp[2]) ? 3'b011 : 3'b111;
								assign node213 = (inp[2]) ? node219 : node214;
									assign node214 = (inp[8]) ? node216 : 3'b111;
										assign node216 = (inp[10]) ? 3'b001 : 3'b111;
									assign node219 = (inp[5]) ? node227 : node220;
										assign node220 = (inp[11]) ? node222 : 3'b101;
											assign node222 = (inp[8]) ? 3'b001 : node223;
												assign node223 = (inp[10]) ? 3'b101 : 3'b001;
										assign node227 = (inp[11]) ? 3'b011 : 3'b001;
					assign node230 = (inp[9]) ? node308 : node231;
						assign node231 = (inp[4]) ? node253 : node232;
							assign node232 = (inp[1]) ? 3'b000 : node233;
								assign node233 = (inp[2]) ? node241 : node234;
									assign node234 = (inp[5]) ? node238 : node235;
										assign node235 = (inp[8]) ? 3'b000 : 3'b100;
										assign node238 = (inp[8]) ? 3'b100 : 3'b000;
									assign node241 = (inp[10]) ? 3'b100 : node242;
										assign node242 = (inp[8]) ? 3'b100 : node243;
											assign node243 = (inp[5]) ? node247 : node244;
												assign node244 = (inp[11]) ? 3'b100 : 3'b000;
												assign node247 = (inp[11]) ? 3'b000 : 3'b100;
							assign node253 = (inp[1]) ? node285 : node254;
								assign node254 = (inp[10]) ? node274 : node255;
									assign node255 = (inp[2]) ? node267 : node256;
										assign node256 = (inp[8]) ? node260 : node257;
											assign node257 = (inp[5]) ? 3'b011 : 3'b111;
											assign node260 = (inp[11]) ? node264 : node261;
												assign node261 = (inp[5]) ? 3'b110 : 3'b010;
												assign node264 = (inp[5]) ? 3'b111 : 3'b110;
										assign node267 = (inp[5]) ? node271 : node268;
											assign node268 = (inp[8]) ? 3'b100 : 3'b010;
											assign node271 = (inp[8]) ? 3'b010 : 3'b110;
									assign node274 = (inp[8]) ? node280 : node275;
										assign node275 = (inp[5]) ? node277 : 3'b001;
											assign node277 = (inp[2]) ? 3'b001 : 3'b101;
										assign node280 = (inp[2]) ? node282 : 3'b001;
											assign node282 = (inp[11]) ? 3'b111 : 3'b010;
								assign node285 = (inp[10]) ? node295 : node286;
									assign node286 = (inp[2]) ? 3'b000 : node287;
										assign node287 = (inp[11]) ? 3'b000 : node288;
											assign node288 = (inp[8]) ? node290 : 3'b100;
												assign node290 = (inp[5]) ? 3'b100 : 3'b000;
									assign node295 = (inp[2]) ? node303 : node296;
										assign node296 = (inp[5]) ? node298 : 3'b100;
											assign node298 = (inp[8]) ? node300 : 3'b010;
												assign node300 = (inp[11]) ? 3'b010 : 3'b100;
										assign node303 = (inp[8]) ? node305 : 3'b100;
											assign node305 = (inp[5]) ? 3'b100 : 3'b000;
						assign node308 = (inp[1]) ? node358 : node309;
							assign node309 = (inp[4]) ? node335 : node310;
								assign node310 = (inp[10]) ? node326 : node311;
									assign node311 = (inp[2]) ? node323 : node312;
										assign node312 = (inp[8]) ? node318 : node313;
											assign node313 = (inp[5]) ? 3'b011 : node314;
												assign node314 = (inp[11]) ? 3'b101 : 3'b100;
											assign node318 = (inp[5]) ? node320 : 3'b000;
												assign node320 = (inp[11]) ? 3'b101 : 3'b100;
										assign node323 = (inp[8]) ? 3'b100 : 3'b000;
									assign node326 = (inp[8]) ? node332 : node327;
										assign node327 = (inp[5]) ? 3'b011 : node328;
											assign node328 = (inp[2]) ? 3'b001 : 3'b101;
										assign node332 = (inp[11]) ? 3'b001 : 3'b000;
								assign node335 = (inp[5]) ? node345 : node336;
									assign node336 = (inp[8]) ? 3'b101 : node337;
										assign node337 = (inp[2]) ? node341 : node338;
											assign node338 = (inp[10]) ? 3'b011 : 3'b101;
											assign node341 = (inp[10]) ? 3'b101 : 3'b001;
									assign node345 = (inp[8]) ? node353 : node346;
										assign node346 = (inp[2]) ? node350 : node347;
											assign node347 = (inp[10]) ? 3'b111 : 3'b001;
											assign node350 = (inp[10]) ? 3'b011 : 3'b111;
										assign node353 = (inp[2]) ? node355 : 3'b011;
											assign node355 = (inp[10]) ? 3'b101 : 3'b001;
							assign node358 = (inp[5]) ? node374 : node359;
								assign node359 = (inp[10]) ? node363 : node360;
									assign node360 = (inp[8]) ? 3'b010 : 3'b110;
									assign node363 = (inp[8]) ? node371 : node364;
										assign node364 = (inp[4]) ? node368 : node365;
											assign node365 = (inp[2]) ? 3'b010 : 3'b110;
											assign node368 = (inp[2]) ? 3'b110 : 3'b001;
										assign node371 = (inp[4]) ? 3'b110 : 3'b100;
								assign node374 = (inp[10]) ? node384 : node375;
									assign node375 = (inp[4]) ? node379 : node376;
										assign node376 = (inp[8]) ? 3'b000 : 3'b001;
										assign node379 = (inp[2]) ? node381 : 3'b110;
											assign node381 = (inp[8]) ? 3'b010 : 3'b011;
									assign node384 = (inp[4]) ? node388 : node385;
										assign node385 = (inp[2]) ? 3'b100 : 3'b110;
										assign node388 = (inp[8]) ? 3'b001 : node389;
											assign node389 = (inp[2]) ? 3'b001 : 3'b101;
				assign node393 = (inp[1]) ? node539 : node394;
					assign node394 = (inp[9]) ? node480 : node395;
						assign node395 = (inp[7]) ? node435 : node396;
							assign node396 = (inp[4]) ? node424 : node397;
								assign node397 = (inp[8]) ? node411 : node398;
									assign node398 = (inp[10]) ? node406 : node399;
										assign node399 = (inp[2]) ? node403 : node400;
											assign node400 = (inp[11]) ? 3'b111 : 3'b011;
											assign node403 = (inp[5]) ? 3'b011 : 3'b101;
										assign node406 = (inp[11]) ? 3'b011 : node407;
											assign node407 = (inp[5]) ? 3'b111 : 3'b011;
									assign node411 = (inp[5]) ? node417 : node412;
										assign node412 = (inp[10]) ? node414 : 3'b111;
											assign node414 = (inp[11]) ? 3'b111 : 3'b011;
										assign node417 = (inp[11]) ? node419 : 3'b111;
											assign node419 = (inp[10]) ? node421 : 3'b011;
												assign node421 = (inp[2]) ? 3'b111 : 3'b011;
								assign node424 = (inp[5]) ? node428 : node425;
									assign node425 = (inp[8]) ? 3'b101 : 3'b111;
									assign node428 = (inp[10]) ? 3'b111 : node429;
										assign node429 = (inp[8]) ? node431 : 3'b111;
											assign node431 = (inp[2]) ? 3'b011 : 3'b111;
							assign node435 = (inp[11]) ? node455 : node436;
								assign node436 = (inp[4]) ? node446 : node437;
									assign node437 = (inp[2]) ? node441 : node438;
										assign node438 = (inp[10]) ? 3'b011 : 3'b001;
										assign node441 = (inp[10]) ? node443 : 3'b110;
											assign node443 = (inp[8]) ? 3'b001 : 3'b010;
									assign node446 = (inp[10]) ? node450 : node447;
										assign node447 = (inp[2]) ? 3'b001 : 3'b011;
										assign node450 = (inp[2]) ? 3'b101 : node451;
											assign node451 = (inp[8]) ? 3'b011 : 3'b101;
								assign node455 = (inp[2]) ? node469 : node456;
									assign node456 = (inp[10]) ? node462 : node457;
										assign node457 = (inp[8]) ? node459 : 3'b101;
											assign node459 = (inp[5]) ? 3'b101 : 3'b001;
										assign node462 = (inp[5]) ? 3'b011 : node463;
											assign node463 = (inp[4]) ? node465 : 3'b101;
												assign node465 = (inp[8]) ? 3'b011 : 3'b111;
									assign node469 = (inp[4]) ? node473 : node470;
										assign node470 = (inp[10]) ? 3'b101 : 3'b010;
										assign node473 = (inp[5]) ? 3'b111 : node474;
											assign node474 = (inp[8]) ? node476 : 3'b011;
												assign node476 = (inp[10]) ? 3'b101 : 3'b001;
						assign node480 = (inp[11]) ? node516 : node481;
							assign node481 = (inp[8]) ? node495 : node482;
								assign node482 = (inp[5]) ? 3'b111 : node483;
									assign node483 = (inp[2]) ? node485 : 3'b111;
										assign node485 = (inp[10]) ? node489 : node486;
											assign node486 = (inp[4]) ? 3'b011 : 3'b101;
											assign node489 = (inp[7]) ? node491 : 3'b111;
												assign node491 = (inp[4]) ? 3'b111 : 3'b011;
								assign node495 = (inp[10]) ? node507 : node496;
									assign node496 = (inp[2]) ? node502 : node497;
										assign node497 = (inp[4]) ? 3'b101 : node498;
											assign node498 = (inp[7]) ? 3'b011 : 3'b111;
										assign node502 = (inp[7]) ? node504 : 3'b101;
											assign node504 = (inp[5]) ? 3'b101 : 3'b001;
									assign node507 = (inp[5]) ? 3'b111 : node508;
										assign node508 = (inp[2]) ? node510 : 3'b101;
											assign node510 = (inp[7]) ? node512 : 3'b111;
												assign node512 = (inp[4]) ? 3'b111 : 3'b101;
							assign node516 = (inp[2]) ? node532 : node517;
								assign node517 = (inp[5]) ? node525 : node518;
									assign node518 = (inp[8]) ? node520 : 3'b111;
										assign node520 = (inp[7]) ? 3'b111 : node521;
											assign node521 = (inp[4]) ? 3'b101 : 3'b111;
									assign node525 = (inp[8]) ? 3'b111 : node526;
										assign node526 = (inp[7]) ? node528 : 3'b111;
											assign node528 = (inp[10]) ? 3'b111 : 3'b101;
								assign node532 = (inp[10]) ? 3'b111 : node533;
									assign node533 = (inp[7]) ? node535 : 3'b111;
										assign node535 = (inp[4]) ? 3'b111 : 3'b011;
					assign node539 = (inp[9]) ? node627 : node540;
						assign node540 = (inp[7]) ? node590 : node541;
							assign node541 = (inp[8]) ? node565 : node542;
								assign node542 = (inp[2]) ? node554 : node543;
									assign node543 = (inp[10]) ? node549 : node544;
										assign node544 = (inp[5]) ? 3'b011 : node545;
											assign node545 = (inp[4]) ? 3'b101 : 3'b001;
										assign node549 = (inp[4]) ? 3'b111 : node550;
											assign node550 = (inp[5]) ? 3'b010 : 3'b110;
									assign node554 = (inp[5]) ? node560 : node555;
										assign node555 = (inp[11]) ? node557 : 3'b001;
											assign node557 = (inp[4]) ? 3'b001 : 3'b101;
										assign node560 = (inp[10]) ? 3'b101 : node561;
											assign node561 = (inp[4]) ? 3'b101 : 3'b001;
								assign node565 = (inp[5]) ? node579 : node566;
									assign node566 = (inp[4]) ? node574 : node567;
										assign node567 = (inp[11]) ? node571 : node568;
											assign node568 = (inp[2]) ? 3'b110 : 3'b010;
											assign node571 = (inp[10]) ? 3'b001 : 3'b010;
										assign node574 = (inp[10]) ? node576 : 3'b110;
											assign node576 = (inp[11]) ? 3'b110 : 3'b010;
									assign node579 = (inp[11]) ? node583 : node580;
										assign node580 = (inp[10]) ? 3'b101 : 3'b110;
										assign node583 = (inp[4]) ? node585 : 3'b001;
											assign node585 = (inp[10]) ? 3'b001 : node586;
												assign node586 = (inp[2]) ? 3'b001 : 3'b101;
							assign node590 = (inp[4]) ? node608 : node591;
								assign node591 = (inp[8]) ? node601 : node592;
									assign node592 = (inp[10]) ? node598 : node593;
										assign node593 = (inp[2]) ? node595 : 3'b110;
											assign node595 = (inp[11]) ? 3'b110 : 3'b100;
										assign node598 = (inp[2]) ? 3'b010 : 3'b110;
									assign node601 = (inp[10]) ? node603 : 3'b000;
										assign node603 = (inp[5]) ? 3'b110 : node604;
											assign node604 = (inp[11]) ? 3'b110 : 3'b000;
								assign node608 = (inp[2]) ? node622 : node609;
									assign node609 = (inp[8]) ? node617 : node610;
										assign node610 = (inp[10]) ? node612 : 3'b001;
											assign node612 = (inp[11]) ? 3'b101 : node613;
												assign node613 = (inp[5]) ? 3'b101 : 3'b001;
										assign node617 = (inp[10]) ? node619 : 3'b110;
											assign node619 = (inp[11]) ? 3'b101 : 3'b001;
									assign node622 = (inp[11]) ? node624 : 3'b110;
										assign node624 = (inp[10]) ? 3'b001 : 3'b110;
						assign node627 = (inp[7]) ? node671 : node628;
							assign node628 = (inp[4]) ? node644 : node629;
								assign node629 = (inp[2]) ? node635 : node630;
									assign node630 = (inp[10]) ? 3'b111 : node631;
										assign node631 = (inp[8]) ? 3'b101 : 3'b111;
									assign node635 = (inp[10]) ? node641 : node636;
										assign node636 = (inp[8]) ? 3'b101 : node637;
											assign node637 = (inp[5]) ? 3'b101 : 3'b001;
										assign node641 = (inp[8]) ? 3'b001 : 3'b111;
								assign node644 = (inp[2]) ? node660 : node645;
									assign node645 = (inp[11]) ? node653 : node646;
										assign node646 = (inp[5]) ? 3'b011 : node647;
											assign node647 = (inp[10]) ? node649 : 3'b111;
												assign node649 = (inp[8]) ? 3'b111 : 3'b011;
										assign node653 = (inp[10]) ? 3'b001 : node654;
											assign node654 = (inp[8]) ? node656 : 3'b011;
												assign node656 = (inp[5]) ? 3'b111 : 3'b011;
									assign node660 = (inp[10]) ? 3'b111 : node661;
										assign node661 = (inp[11]) ? 3'b111 : node662;
											assign node662 = (inp[5]) ? node666 : node663;
												assign node663 = (inp[8]) ? 3'b111 : 3'b011;
												assign node666 = (inp[8]) ? 3'b011 : 3'b111;
							assign node671 = (inp[2]) ? node699 : node672;
								assign node672 = (inp[8]) ? node684 : node673;
									assign node673 = (inp[5]) ? node679 : node674;
										assign node674 = (inp[10]) ? 3'b011 : node675;
											assign node675 = (inp[11]) ? 3'b101 : 3'b001;
										assign node679 = (inp[10]) ? 3'b111 : node680;
											assign node680 = (inp[11]) ? 3'b111 : 3'b011;
									assign node684 = (inp[11]) ? node690 : node685;
										assign node685 = (inp[5]) ? 3'b101 : node686;
											assign node686 = (inp[4]) ? 3'b101 : 3'b001;
										assign node690 = (inp[4]) ? node694 : node691;
											assign node691 = (inp[10]) ? 3'b101 : 3'b001;
											assign node694 = (inp[10]) ? 3'b011 : node695;
												assign node695 = (inp[5]) ? 3'b011 : 3'b101;
								assign node699 = (inp[4]) ? node715 : node700;
									assign node700 = (inp[10]) ? node706 : node701;
										assign node701 = (inp[8]) ? node703 : 3'b010;
											assign node703 = (inp[5]) ? 3'b110 : 3'b010;
										assign node706 = (inp[11]) ? node712 : node707;
											assign node707 = (inp[5]) ? node709 : 3'b001;
												assign node709 = (inp[8]) ? 3'b001 : 3'b000;
											assign node712 = (inp[5]) ? 3'b100 : 3'b101;
									assign node715 = (inp[5]) ? 3'b101 : node716;
										assign node716 = (inp[8]) ? 3'b001 : 3'b101;
		assign node720 = (inp[6]) ? node1324 : node721;
			assign node721 = (inp[3]) ? node1001 : node722;
				assign node722 = (inp[4]) ? node890 : node723;
					assign node723 = (inp[9]) ? node819 : node724;
						assign node724 = (inp[7]) ? node766 : node725;
							assign node725 = (inp[1]) ? node747 : node726;
								assign node726 = (inp[8]) ? node738 : node727;
									assign node727 = (inp[11]) ? node733 : node728;
										assign node728 = (inp[2]) ? 3'b010 : node729;
											assign node729 = (inp[5]) ? 3'b110 : 3'b010;
										assign node733 = (inp[2]) ? node735 : 3'b110;
											assign node735 = (inp[10]) ? 3'b010 : 3'b110;
									assign node738 = (inp[2]) ? node742 : node739;
										assign node739 = (inp[10]) ? 3'b010 : 3'b110;
										assign node742 = (inp[5]) ? node744 : 3'b100;
											assign node744 = (inp[11]) ? 3'b010 : 3'b100;
								assign node747 = (inp[8]) ? node755 : node748;
									assign node748 = (inp[10]) ? node752 : node749;
										assign node749 = (inp[2]) ? 3'b000 : 3'b100;
										assign node752 = (inp[2]) ? 3'b110 : 3'b010;
									assign node755 = (inp[5]) ? 3'b000 : node756;
										assign node756 = (inp[10]) ? node760 : node757;
											assign node757 = (inp[2]) ? 3'b110 : 3'b000;
											assign node760 = (inp[2]) ? node762 : 3'b100;
												assign node762 = (inp[11]) ? 3'b000 : 3'b100;
							assign node766 = (inp[1]) ? node796 : node767;
								assign node767 = (inp[8]) ? node781 : node768;
									assign node768 = (inp[10]) ? node778 : node769;
										assign node769 = (inp[2]) ? node775 : node770;
											assign node770 = (inp[11]) ? node772 : 3'b100;
												assign node772 = (inp[5]) ? 3'b010 : 3'b000;
											assign node775 = (inp[11]) ? 3'b100 : 3'b000;
										assign node778 = (inp[5]) ? 3'b010 : 3'b000;
									assign node781 = (inp[2]) ? node789 : node782;
										assign node782 = (inp[5]) ? 3'b100 : node783;
											assign node783 = (inp[11]) ? node785 : 3'b000;
												assign node785 = (inp[10]) ? 3'b000 : 3'b100;
										assign node789 = (inp[5]) ? node793 : node790;
											assign node790 = (inp[11]) ? 3'b100 : 3'b110;
											assign node793 = (inp[10]) ? 3'b100 : 3'b000;
								assign node796 = (inp[10]) ? node806 : node797;
									assign node797 = (inp[2]) ? node803 : node798;
										assign node798 = (inp[5]) ? 3'b110 : node799;
											assign node799 = (inp[8]) ? 3'b010 : 3'b110;
										assign node803 = (inp[8]) ? 3'b100 : 3'b010;
									assign node806 = (inp[8]) ? 3'b010 : node807;
										assign node807 = (inp[2]) ? node811 : node808;
											assign node808 = (inp[5]) ? 3'b000 : 3'b010;
											assign node811 = (inp[11]) ? node815 : node812;
												assign node812 = (inp[5]) ? 3'b100 : 3'b000;
												assign node815 = (inp[5]) ? 3'b000 : 3'b100;
						assign node819 = (inp[1]) ? node829 : node820;
							assign node820 = (inp[2]) ? node822 : 3'b110;
								assign node822 = (inp[7]) ? node824 : 3'b110;
									assign node824 = (inp[10]) ? node826 : 3'b010;
										assign node826 = (inp[8]) ? 3'b010 : 3'b110;
							assign node829 = (inp[7]) ? node857 : node830;
								assign node830 = (inp[10]) ? node850 : node831;
									assign node831 = (inp[2]) ? node841 : node832;
										assign node832 = (inp[8]) ? node836 : node833;
											assign node833 = (inp[11]) ? 3'b110 : 3'b010;
											assign node836 = (inp[5]) ? 3'b010 : node837;
												assign node837 = (inp[11]) ? 3'b010 : 3'b110;
										assign node841 = (inp[5]) ? 3'b010 : node842;
											assign node842 = (inp[11]) ? node846 : node843;
												assign node843 = (inp[8]) ? 3'b010 : 3'b100;
												assign node846 = (inp[8]) ? 3'b100 : 3'b010;
									assign node850 = (inp[5]) ? 3'b110 : node851;
										assign node851 = (inp[11]) ? 3'b010 : node852;
											assign node852 = (inp[2]) ? 3'b110 : 3'b010;
								assign node857 = (inp[2]) ? node873 : node858;
									assign node858 = (inp[10]) ? node862 : node859;
										assign node859 = (inp[11]) ? 3'b000 : 3'b010;
										assign node862 = (inp[8]) ? node866 : node863;
											assign node863 = (inp[11]) ? 3'b010 : 3'b110;
											assign node866 = (inp[5]) ? node870 : node867;
												assign node867 = (inp[11]) ? 3'b100 : 3'b110;
												assign node870 = (inp[11]) ? 3'b010 : 3'b000;
									assign node873 = (inp[8]) ? node883 : node874;
										assign node874 = (inp[10]) ? 3'b100 : node875;
											assign node875 = (inp[11]) ? node879 : node876;
												assign node876 = (inp[5]) ? 3'b000 : 3'b110;
												assign node879 = (inp[5]) ? 3'b100 : 3'b000;
										assign node883 = (inp[5]) ? node885 : 3'b000;
											assign node885 = (inp[11]) ? node887 : 3'b000;
												assign node887 = (inp[10]) ? 3'b100 : 3'b000;
					assign node890 = (inp[1]) ? node958 : node891;
						assign node891 = (inp[7]) ? node927 : node892;
							assign node892 = (inp[11]) ? node914 : node893;
								assign node893 = (inp[9]) ? node909 : node894;
									assign node894 = (inp[8]) ? node904 : node895;
										assign node895 = (inp[10]) ? node897 : 3'b001;
											assign node897 = (inp[5]) ? node901 : node898;
												assign node898 = (inp[2]) ? 3'b110 : 3'b001;
												assign node901 = (inp[2]) ? 3'b001 : 3'b110;
										assign node904 = (inp[5]) ? node906 : 3'b001;
											assign node906 = (inp[2]) ? 3'b001 : 3'b110;
									assign node909 = (inp[8]) ? 3'b110 : node910;
										assign node910 = (inp[10]) ? 3'b001 : 3'b110;
								assign node914 = (inp[5]) ? node922 : node915;
									assign node915 = (inp[2]) ? node917 : 3'b001;
										assign node917 = (inp[9]) ? node919 : 3'b110;
											assign node919 = (inp[8]) ? 3'b001 : 3'b110;
									assign node922 = (inp[2]) ? node924 : 3'b110;
										assign node924 = (inp[10]) ? 3'b001 : 3'b110;
							assign node927 = (inp[5]) ? node943 : node928;
								assign node928 = (inp[10]) ? node934 : node929;
									assign node929 = (inp[8]) ? 3'b101 : node930;
										assign node930 = (inp[2]) ? 3'b101 : 3'b001;
									assign node934 = (inp[2]) ? node938 : node935;
										assign node935 = (inp[8]) ? 3'b001 : 3'b101;
										assign node938 = (inp[8]) ? node940 : 3'b001;
											assign node940 = (inp[11]) ? 3'b001 : 3'b101;
								assign node943 = (inp[2]) ? node951 : node944;
									assign node944 = (inp[8]) ? node948 : node945;
										assign node945 = (inp[10]) ? 3'b011 : 3'b111;
										assign node948 = (inp[10]) ? 3'b101 : 3'b001;
									assign node951 = (inp[10]) ? node955 : node952;
										assign node952 = (inp[8]) ? 3'b101 : 3'b001;
										assign node955 = (inp[8]) ? 3'b001 : 3'b101;
						assign node958 = (inp[9]) ? node974 : node959;
							assign node959 = (inp[7]) ? node967 : node960;
								assign node960 = (inp[10]) ? node962 : 3'b001;
									assign node962 = (inp[2]) ? 3'b001 : node963;
										assign node963 = (inp[8]) ? 3'b001 : 3'b110;
								assign node967 = (inp[8]) ? 3'b000 : node968;
									assign node968 = (inp[2]) ? 3'b000 : node969;
										assign node969 = (inp[5]) ? 3'b001 : 3'b000;
							assign node974 = (inp[7]) ? node990 : node975;
								assign node975 = (inp[2]) ? node983 : node976;
									assign node976 = (inp[5]) ? 3'b110 : node977;
										assign node977 = (inp[11]) ? node979 : 3'b001;
											assign node979 = (inp[8]) ? 3'b110 : 3'b001;
									assign node983 = (inp[11]) ? node985 : 3'b001;
										assign node985 = (inp[8]) ? node987 : 3'b001;
											assign node987 = (inp[10]) ? 3'b110 : 3'b001;
								assign node990 = (inp[8]) ? node998 : node991;
									assign node991 = (inp[5]) ? node995 : node992;
										assign node992 = (inp[2]) ? 3'b010 : 3'b110;
										assign node995 = (inp[2]) ? 3'b110 : 3'b001;
									assign node998 = (inp[2]) ? 3'b100 : 3'b110;
				assign node1001 = (inp[9]) ? node1195 : node1002;
					assign node1002 = (inp[7]) ? node1092 : node1003;
						assign node1003 = (inp[1]) ? node1031 : node1004;
							assign node1004 = (inp[4]) ? node1014 : node1005;
								assign node1005 = (inp[10]) ? 3'b111 : node1006;
									assign node1006 = (inp[2]) ? node1008 : 3'b111;
										assign node1008 = (inp[11]) ? node1010 : 3'b011;
											assign node1010 = (inp[5]) ? 3'b111 : 3'b011;
								assign node1014 = (inp[2]) ? node1026 : node1015;
									assign node1015 = (inp[5]) ? node1021 : node1016;
										assign node1016 = (inp[8]) ? 3'b011 : node1017;
											assign node1017 = (inp[11]) ? 3'b111 : 3'b011;
										assign node1021 = (inp[11]) ? 3'b111 : node1022;
											assign node1022 = (inp[8]) ? 3'b011 : 3'b111;
									assign node1026 = (inp[8]) ? node1028 : 3'b011;
										assign node1028 = (inp[11]) ? 3'b011 : 3'b101;
							assign node1031 = (inp[4]) ? node1057 : node1032;
								assign node1032 = (inp[2]) ? node1044 : node1033;
									assign node1033 = (inp[5]) ? node1037 : node1034;
										assign node1034 = (inp[8]) ? 3'b000 : 3'b010;
										assign node1037 = (inp[8]) ? node1041 : node1038;
											assign node1038 = (inp[10]) ? 3'b111 : 3'b011;
											assign node1041 = (inp[10]) ? 3'b010 : 3'b110;
									assign node1044 = (inp[11]) ? node1052 : node1045;
										assign node1045 = (inp[10]) ? node1047 : 3'b010;
											assign node1047 = (inp[5]) ? node1049 : 3'b110;
												assign node1049 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1052 = (inp[10]) ? 3'b110 : node1053;
											assign node1053 = (inp[5]) ? 3'b110 : 3'b100;
								assign node1057 = (inp[2]) ? node1071 : node1058;
									assign node1058 = (inp[10]) ? node1066 : node1059;
										assign node1059 = (inp[11]) ? node1061 : 3'b001;
											assign node1061 = (inp[8]) ? node1063 : 3'b101;
												assign node1063 = (inp[5]) ? 3'b101 : 3'b001;
										assign node1066 = (inp[11]) ? 3'b011 : node1067;
											assign node1067 = (inp[5]) ? 3'b011 : 3'b101;
									assign node1071 = (inp[11]) ? node1081 : node1072;
										assign node1072 = (inp[10]) ? node1078 : node1073;
											assign node1073 = (inp[8]) ? 3'b110 : node1074;
												assign node1074 = (inp[5]) ? 3'b001 : 3'b110;
											assign node1078 = (inp[5]) ? 3'b000 : 3'b010;
										assign node1081 = (inp[10]) ? node1087 : node1082;
											assign node1082 = (inp[8]) ? 3'b011 : node1083;
												assign node1083 = (inp[5]) ? 3'b001 : 3'b011;
											assign node1087 = (inp[8]) ? node1089 : 3'b111;
												assign node1089 = (inp[5]) ? 3'b101 : 3'b000;
						assign node1092 = (inp[4]) ? node1138 : node1093;
							assign node1093 = (inp[5]) ? node1113 : node1094;
								assign node1094 = (inp[8]) ? node1106 : node1095;
									assign node1095 = (inp[2]) ? node1099 : node1096;
										assign node1096 = (inp[1]) ? 3'b010 : 3'b000;
										assign node1099 = (inp[11]) ? node1103 : node1100;
											assign node1100 = (inp[1]) ? 3'b100 : 3'b110;
											assign node1103 = (inp[1]) ? 3'b010 : 3'b110;
									assign node1106 = (inp[1]) ? node1110 : node1107;
										assign node1107 = (inp[2]) ? 3'b010 : 3'b000;
										assign node1110 = (inp[2]) ? 3'b000 : 3'b010;
								assign node1113 = (inp[1]) ? node1133 : node1114;
									assign node1114 = (inp[2]) ? node1126 : node1115;
										assign node1115 = (inp[8]) ? node1119 : node1116;
											assign node1116 = (inp[10]) ? 3'b101 : 3'b001;
											assign node1119 = (inp[11]) ? node1123 : node1120;
												assign node1120 = (inp[10]) ? 3'b000 : 3'b110;
												assign node1123 = (inp[10]) ? 3'b100 : 3'b000;
										assign node1126 = (inp[10]) ? node1130 : node1127;
											assign node1127 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1130 = (inp[8]) ? 3'b110 : 3'b000;
									assign node1133 = (inp[2]) ? 3'b100 : node1134;
										assign node1134 = (inp[10]) ? 3'b110 : 3'b010;
							assign node1138 = (inp[1]) ? node1168 : node1139;
								assign node1139 = (inp[8]) ? node1153 : node1140;
									assign node1140 = (inp[5]) ? node1144 : node1141;
										assign node1141 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1144 = (inp[10]) ? node1150 : node1145;
											assign node1145 = (inp[2]) ? node1147 : 3'b011;
												assign node1147 = (inp[11]) ? 3'b101 : 3'b001;
											assign node1150 = (inp[2]) ? 3'b011 : 3'b111;
									assign node1153 = (inp[5]) ? node1161 : node1154;
										assign node1154 = (inp[2]) ? node1156 : 3'b001;
											assign node1156 = (inp[11]) ? 3'b010 : node1157;
												assign node1157 = (inp[10]) ? 3'b100 : 3'b110;
										assign node1161 = (inp[10]) ? node1165 : node1162;
											assign node1162 = (inp[2]) ? 3'b001 : 3'b101;
											assign node1165 = (inp[11]) ? 3'b101 : 3'b001;
								assign node1168 = (inp[10]) ? node1178 : node1169;
									assign node1169 = (inp[2]) ? node1175 : node1170;
										assign node1170 = (inp[8]) ? node1172 : 3'b110;
											assign node1172 = (inp[5]) ? 3'b110 : 3'b010;
										assign node1175 = (inp[8]) ? 3'b100 : 3'b010;
									assign node1178 = (inp[5]) ? node1184 : node1179;
										assign node1179 = (inp[8]) ? node1181 : 3'b011;
											assign node1181 = (inp[11]) ? 3'b011 : 3'b010;
										assign node1184 = (inp[8]) ? node1190 : node1185;
											assign node1185 = (inp[2]) ? node1187 : 3'b000;
												assign node1187 = (inp[11]) ? 3'b001 : 3'b101;
											assign node1190 = (inp[2]) ? node1192 : 3'b001;
												assign node1192 = (inp[11]) ? 3'b110 : 3'b010;
					assign node1195 = (inp[1]) ? node1235 : node1196;
						assign node1196 = (inp[7]) ? node1204 : node1197;
							assign node1197 = (inp[5]) ? 3'b111 : node1198;
								assign node1198 = (inp[4]) ? 3'b111 : node1199;
									assign node1199 = (inp[10]) ? 3'b111 : 3'b011;
							assign node1204 = (inp[4]) ? node1226 : node1205;
								assign node1205 = (inp[2]) ? node1215 : node1206;
									assign node1206 = (inp[10]) ? node1212 : node1207;
										assign node1207 = (inp[8]) ? node1209 : 3'b011;
											assign node1209 = (inp[5]) ? 3'b011 : 3'b101;
										assign node1212 = (inp[5]) ? 3'b111 : 3'b011;
									assign node1215 = (inp[11]) ? 3'b101 : node1216;
										assign node1216 = (inp[5]) ? node1218 : 3'b101;
											assign node1218 = (inp[8]) ? node1222 : node1219;
												assign node1219 = (inp[10]) ? 3'b011 : 3'b101;
												assign node1222 = (inp[10]) ? 3'b101 : 3'b001;
								assign node1226 = (inp[2]) ? node1228 : 3'b111;
									assign node1228 = (inp[10]) ? node1230 : 3'b011;
										assign node1230 = (inp[5]) ? 3'b111 : node1231;
											assign node1231 = (inp[8]) ? 3'b011 : 3'b111;
						assign node1235 = (inp[7]) ? node1271 : node1236;
							assign node1236 = (inp[2]) ? node1256 : node1237;
								assign node1237 = (inp[10]) ? node1243 : node1238;
									assign node1238 = (inp[5]) ? node1240 : 3'b011;
										assign node1240 = (inp[8]) ? 3'b111 : 3'b011;
									assign node1243 = (inp[8]) ? node1245 : 3'b111;
										assign node1245 = (inp[4]) ? node1251 : node1246;
											assign node1246 = (inp[5]) ? 3'b011 : node1247;
												assign node1247 = (inp[11]) ? 3'b011 : 3'b111;
											assign node1251 = (inp[11]) ? 3'b111 : node1252;
												assign node1252 = (inp[5]) ? 3'b111 : 3'b011;
								assign node1256 = (inp[11]) ? node1266 : node1257;
									assign node1257 = (inp[5]) ? node1259 : 3'b001;
										assign node1259 = (inp[4]) ? node1261 : 3'b101;
											assign node1261 = (inp[10]) ? node1263 : 3'b101;
												assign node1263 = (inp[8]) ? 3'b011 : 3'b111;
									assign node1266 = (inp[10]) ? node1268 : 3'b011;
										assign node1268 = (inp[4]) ? 3'b111 : 3'b011;
							assign node1271 = (inp[11]) ? node1299 : node1272;
								assign node1272 = (inp[10]) ? node1290 : node1273;
									assign node1273 = (inp[8]) ? node1283 : node1274;
										assign node1274 = (inp[5]) ? 3'b110 : node1275;
											assign node1275 = (inp[2]) ? node1279 : node1276;
												assign node1276 = (inp[4]) ? 3'b010 : 3'b110;
												assign node1279 = (inp[4]) ? 3'b110 : 3'b010;
										assign node1283 = (inp[5]) ? node1285 : 3'b111;
											assign node1285 = (inp[2]) ? 3'b110 : node1286;
												assign node1286 = (inp[4]) ? 3'b010 : 3'b110;
									assign node1290 = (inp[4]) ? node1294 : node1291;
										assign node1291 = (inp[2]) ? 3'b110 : 3'b001;
										assign node1294 = (inp[8]) ? 3'b001 : node1295;
											assign node1295 = (inp[2]) ? 3'b101 : 3'b111;
								assign node1299 = (inp[8]) ? node1309 : node1300;
									assign node1300 = (inp[5]) ? node1302 : 3'b001;
										assign node1302 = (inp[4]) ? node1306 : node1303;
											assign node1303 = (inp[10]) ? 3'b101 : 3'b001;
											assign node1306 = (inp[2]) ? 3'b101 : 3'b111;
									assign node1309 = (inp[4]) ? node1319 : node1310;
										assign node1310 = (inp[2]) ? 3'b110 : node1311;
											assign node1311 = (inp[10]) ? node1315 : node1312;
												assign node1312 = (inp[5]) ? 3'b001 : 3'b110;
												assign node1315 = (inp[5]) ? 3'b101 : 3'b001;
										assign node1319 = (inp[5]) ? 3'b001 : node1320;
											assign node1320 = (inp[2]) ? 3'b001 : 3'b101;
			assign node1324 = (inp[1]) ? node1550 : node1325;
				assign node1325 = (inp[7]) ? node1445 : node1326;
					assign node1326 = (inp[3]) ? node1388 : node1327;
						assign node1327 = (inp[4]) ? node1361 : node1328;
							assign node1328 = (inp[2]) ? node1348 : node1329;
								assign node1329 = (inp[11]) ? node1337 : node1330;
									assign node1330 = (inp[10]) ? node1332 : 3'b110;
										assign node1332 = (inp[5]) ? 3'b010 : node1333;
											assign node1333 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1337 = (inp[5]) ? node1339 : 3'b010;
										assign node1339 = (inp[9]) ? 3'b110 : node1340;
											assign node1340 = (inp[8]) ? node1344 : node1341;
												assign node1341 = (inp[10]) ? 3'b110 : 3'b010;
												assign node1344 = (inp[10]) ? 3'b010 : 3'b110;
								assign node1348 = (inp[10]) ? node1356 : node1349;
									assign node1349 = (inp[8]) ? node1353 : node1350;
										assign node1350 = (inp[5]) ? 3'b100 : 3'b000;
										assign node1353 = (inp[5]) ? 3'b000 : 3'b110;
									assign node1356 = (inp[5]) ? node1358 : 3'b100;
										assign node1358 = (inp[8]) ? 3'b100 : 3'b010;
							assign node1361 = (inp[2]) ? node1381 : node1362;
								assign node1362 = (inp[10]) ? node1372 : node1363;
									assign node1363 = (inp[9]) ? node1367 : node1364;
										assign node1364 = (inp[8]) ? 3'b110 : 3'b100;
										assign node1367 = (inp[8]) ? node1369 : 3'b000;
											assign node1369 = (inp[11]) ? 3'b110 : 3'b000;
									assign node1372 = (inp[8]) ? node1374 : 3'b101;
										assign node1374 = (inp[5]) ? node1376 : 3'b110;
											assign node1376 = (inp[9]) ? node1378 : 3'b101;
												assign node1378 = (inp[11]) ? 3'b001 : 3'b000;
								assign node1381 = (inp[5]) ? 3'b110 : node1382;
									assign node1382 = (inp[9]) ? node1384 : 3'b110;
										assign node1384 = (inp[8]) ? 3'b010 : 3'b110;
						assign node1388 = (inp[9]) ? node1418 : node1389;
							assign node1389 = (inp[2]) ? node1407 : node1390;
								assign node1390 = (inp[4]) ? node1396 : node1391;
									assign node1391 = (inp[5]) ? 3'b010 : node1392;
										assign node1392 = (inp[8]) ? 3'b100 : 3'b010;
									assign node1396 = (inp[5]) ? node1402 : node1397;
										assign node1397 = (inp[8]) ? 3'b010 : node1398;
											assign node1398 = (inp[10]) ? 3'b010 : 3'b110;
										assign node1402 = (inp[8]) ? 3'b110 : node1403;
											assign node1403 = (inp[10]) ? 3'b101 : 3'b001;
								assign node1407 = (inp[4]) ? node1409 : 3'b100;
									assign node1409 = (inp[5]) ? 3'b010 : node1410;
										assign node1410 = (inp[8]) ? node1414 : node1411;
											assign node1411 = (inp[10]) ? 3'b110 : 3'b010;
											assign node1414 = (inp[10]) ? 3'b000 : 3'b100;
							assign node1418 = (inp[4]) ? 3'b101 : node1419;
								assign node1419 = (inp[10]) ? node1435 : node1420;
									assign node1420 = (inp[8]) ? node1428 : node1421;
										assign node1421 = (inp[11]) ? 3'b101 : node1422;
											assign node1422 = (inp[5]) ? node1424 : 3'b100;
												assign node1424 = (inp[2]) ? 3'b100 : 3'b011;
										assign node1428 = (inp[5]) ? node1430 : 3'b010;
											assign node1430 = (inp[2]) ? node1432 : 3'b100;
												assign node1432 = (inp[11]) ? 3'b100 : 3'b000;
									assign node1435 = (inp[5]) ? node1441 : node1436;
										assign node1436 = (inp[2]) ? 3'b001 : node1437;
											assign node1437 = (inp[8]) ? 3'b001 : 3'b101;
										assign node1441 = (inp[2]) ? 3'b001 : 3'b011;
					assign node1445 = (inp[3]) ? node1477 : node1446;
						assign node1446 = (inp[8]) ? node1468 : node1447;
							assign node1447 = (inp[9]) ? node1455 : node1448;
								assign node1448 = (inp[4]) ? 3'b000 : node1449;
									assign node1449 = (inp[2]) ? 3'b000 : node1450;
										assign node1450 = (inp[10]) ? 3'b100 : 3'b000;
								assign node1455 = (inp[4]) ? node1457 : 3'b000;
									assign node1457 = (inp[10]) ? node1463 : node1458;
										assign node1458 = (inp[2]) ? node1460 : 3'b100;
											assign node1460 = (inp[5]) ? 3'b010 : 3'b000;
										assign node1463 = (inp[2]) ? 3'b100 : node1464;
											assign node1464 = (inp[5]) ? 3'b110 : 3'b010;
							assign node1468 = (inp[4]) ? node1470 : 3'b000;
								assign node1470 = (inp[9]) ? node1472 : 3'b000;
									assign node1472 = (inp[5]) ? 3'b000 : node1473;
										assign node1473 = (inp[11]) ? 3'b100 : 3'b000;
						assign node1477 = (inp[9]) ? node1511 : node1478;
							assign node1478 = (inp[4]) ? node1488 : node1479;
								assign node1479 = (inp[10]) ? node1481 : 3'b000;
									assign node1481 = (inp[8]) ? node1483 : 3'b100;
										assign node1483 = (inp[2]) ? 3'b000 : node1484;
											assign node1484 = (inp[11]) ? 3'b100 : 3'b000;
								assign node1488 = (inp[10]) ? node1500 : node1489;
									assign node1489 = (inp[11]) ? node1493 : node1490;
										assign node1490 = (inp[2]) ? 3'b000 : 3'b100;
										assign node1493 = (inp[2]) ? 3'b100 : node1494;
											assign node1494 = (inp[8]) ? 3'b100 : node1495;
												assign node1495 = (inp[5]) ? 3'b110 : 3'b010;
									assign node1500 = (inp[11]) ? node1506 : node1501;
										assign node1501 = (inp[2]) ? 3'b100 : node1502;
											assign node1502 = (inp[5]) ? 3'b110 : 3'b010;
										assign node1506 = (inp[8]) ? 3'b010 : node1507;
											assign node1507 = (inp[2]) ? 3'b010 : 3'b110;
							assign node1511 = (inp[2]) ? node1527 : node1512;
								assign node1512 = (inp[10]) ? node1522 : node1513;
									assign node1513 = (inp[8]) ? node1519 : node1514;
										assign node1514 = (inp[5]) ? node1516 : 3'b011;
											assign node1516 = (inp[4]) ? 3'b001 : 3'b101;
										assign node1519 = (inp[4]) ? 3'b110 : 3'b010;
									assign node1522 = (inp[5]) ? node1524 : 3'b001;
										assign node1524 = (inp[4]) ? 3'b101 : 3'b001;
								assign node1527 = (inp[10]) ? node1539 : node1528;
									assign node1528 = (inp[4]) ? node1536 : node1529;
										assign node1529 = (inp[11]) ? 3'b100 : node1530;
											assign node1530 = (inp[5]) ? 3'b000 : node1531;
												assign node1531 = (inp[8]) ? 3'b000 : 3'b100;
										assign node1536 = (inp[5]) ? 3'b110 : 3'b010;
									assign node1539 = (inp[11]) ? node1543 : node1540;
										assign node1540 = (inp[8]) ? 3'b100 : 3'b110;
										assign node1543 = (inp[4]) ? node1547 : node1544;
											assign node1544 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1547 = (inp[5]) ? 3'b001 : 3'b110;
				assign node1550 = (inp[3]) ? node1586 : node1551;
					assign node1551 = (inp[2]) ? 3'b000 : node1552;
						assign node1552 = (inp[5]) ? node1560 : node1553;
							assign node1553 = (inp[9]) ? node1555 : 3'b000;
								assign node1555 = (inp[7]) ? 3'b000 : node1556;
									assign node1556 = (inp[8]) ? 3'b100 : 3'b000;
							assign node1560 = (inp[8]) ? node1578 : node1561;
								assign node1561 = (inp[10]) ? node1569 : node1562;
									assign node1562 = (inp[7]) ? node1566 : node1563;
										assign node1563 = (inp[4]) ? 3'b000 : 3'b100;
										assign node1566 = (inp[4]) ? 3'b100 : 3'b000;
									assign node1569 = (inp[4]) ? node1573 : node1570;
										assign node1570 = (inp[7]) ? 3'b000 : 3'b100;
										assign node1573 = (inp[7]) ? node1575 : 3'b010;
											assign node1575 = (inp[9]) ? 3'b100 : 3'b000;
								assign node1578 = (inp[4]) ? node1580 : 3'b000;
									assign node1580 = (inp[7]) ? 3'b000 : node1581;
										assign node1581 = (inp[11]) ? 3'b010 : 3'b000;
					assign node1586 = (inp[9]) ? node1616 : node1587;
						assign node1587 = (inp[4]) ? node1595 : node1588;
							assign node1588 = (inp[2]) ? 3'b000 : node1589;
								assign node1589 = (inp[8]) ? 3'b000 : node1590;
									assign node1590 = (inp[5]) ? 3'b010 : 3'b000;
							assign node1595 = (inp[7]) ? node1609 : node1596;
								assign node1596 = (inp[8]) ? node1604 : node1597;
									assign node1597 = (inp[2]) ? node1599 : 3'b010;
										assign node1599 = (inp[11]) ? 3'b010 : node1600;
											assign node1600 = (inp[5]) ? 3'b100 : 3'b000;
									assign node1604 = (inp[5]) ? 3'b100 : node1605;
										assign node1605 = (inp[11]) ? 3'b100 : 3'b000;
								assign node1609 = (inp[2]) ? 3'b000 : node1610;
									assign node1610 = (inp[5]) ? node1612 : 3'b000;
										assign node1612 = (inp[10]) ? 3'b100 : 3'b000;
						assign node1616 = (inp[7]) ? node1658 : node1617;
							assign node1617 = (inp[2]) ? node1631 : node1618;
								assign node1618 = (inp[4]) ? node1624 : node1619;
									assign node1619 = (inp[8]) ? node1621 : 3'b001;
										assign node1621 = (inp[5]) ? 3'b110 : 3'b010;
									assign node1624 = (inp[5]) ? node1626 : 3'b001;
										assign node1626 = (inp[10]) ? 3'b101 : node1627;
											assign node1627 = (inp[8]) ? 3'b101 : 3'b001;
								assign node1631 = (inp[8]) ? node1643 : node1632;
									assign node1632 = (inp[10]) ? node1638 : node1633;
										assign node1633 = (inp[4]) ? 3'b110 : node1634;
											assign node1634 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1638 = (inp[5]) ? node1640 : 3'b110;
											assign node1640 = (inp[4]) ? 3'b001 : 3'b110;
									assign node1643 = (inp[10]) ? node1649 : node1644;
										assign node1644 = (inp[5]) ? 3'b100 : node1645;
											assign node1645 = (inp[4]) ? 3'b100 : 3'b010;
										assign node1649 = (inp[5]) ? node1651 : 3'b010;
											assign node1651 = (inp[11]) ? node1655 : node1652;
												assign node1652 = (inp[4]) ? 3'b110 : 3'b100;
												assign node1655 = (inp[4]) ? 3'b110 : 3'b010;
							assign node1658 = (inp[4]) ? node1672 : node1659;
								assign node1659 = (inp[10]) ? node1661 : 3'b000;
									assign node1661 = (inp[8]) ? 3'b000 : node1662;
										assign node1662 = (inp[11]) ? 3'b100 : node1663;
											assign node1663 = (inp[2]) ? node1667 : node1664;
												assign node1664 = (inp[5]) ? 3'b010 : 3'b100;
												assign node1667 = (inp[5]) ? 3'b100 : 3'b000;
								assign node1672 = (inp[5]) ? node1688 : node1673;
									assign node1673 = (inp[10]) ? node1681 : node1674;
										assign node1674 = (inp[8]) ? 3'b000 : node1675;
											assign node1675 = (inp[11]) ? 3'b100 : node1676;
												assign node1676 = (inp[2]) ? 3'b000 : 3'b100;
										assign node1681 = (inp[8]) ? 3'b100 : node1682;
											assign node1682 = (inp[2]) ? node1684 : 3'b010;
												assign node1684 = (inp[11]) ? 3'b010 : 3'b100;
									assign node1688 = (inp[10]) ? node1692 : node1689;
										assign node1689 = (inp[2]) ? 3'b100 : 3'b010;
										assign node1692 = (inp[11]) ? node1694 : 3'b010;
											assign node1694 = (inp[2]) ? 3'b010 : 3'b110;

endmodule