module dtc_split66_bm90 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node208;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node243;
	wire [3-1:0] node246;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node257;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node272;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node281;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node340;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node352;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node363;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node371;
	wire [3-1:0] node373;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node386;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node396;
	wire [3-1:0] node400;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node408;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node427;
	wire [3-1:0] node429;
	wire [3-1:0] node432;
	wire [3-1:0] node434;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node442;
	wire [3-1:0] node445;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node457;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node471;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node493;
	wire [3-1:0] node496;
	wire [3-1:0] node498;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node517;
	wire [3-1:0] node519;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node530;
	wire [3-1:0] node533;
	wire [3-1:0] node535;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node542;
	wire [3-1:0] node545;
	wire [3-1:0] node547;
	wire [3-1:0] node550;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node564;
	wire [3-1:0] node567;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node573;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node581;
	wire [3-1:0] node583;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node590;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node605;
	wire [3-1:0] node608;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node617;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node651;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node659;
	wire [3-1:0] node661;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node673;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node680;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node686;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node693;
	wire [3-1:0] node696;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node710;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node721;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node728;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node735;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node743;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node759;
	wire [3-1:0] node761;
	wire [3-1:0] node764;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node770;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node777;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node784;
	wire [3-1:0] node787;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node801;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node812;
	wire [3-1:0] node814;
	wire [3-1:0] node817;
	wire [3-1:0] node819;
	wire [3-1:0] node821;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node829;
	wire [3-1:0] node832;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node840;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node854;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node868;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node881;
	wire [3-1:0] node883;
	wire [3-1:0] node884;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node895;
	wire [3-1:0] node899;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node906;
	wire [3-1:0] node908;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node918;
	wire [3-1:0] node919;
	wire [3-1:0] node922;
	wire [3-1:0] node924;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node934;
	wire [3-1:0] node938;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node948;
	wire [3-1:0] node951;
	wire [3-1:0] node953;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node965;
	wire [3-1:0] node967;
	wire [3-1:0] node970;
	wire [3-1:0] node971;
	wire [3-1:0] node972;
	wire [3-1:0] node976;
	wire [3-1:0] node978;
	wire [3-1:0] node981;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node985;
	wire [3-1:0] node990;
	wire [3-1:0] node992;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node998;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1008;
	wire [3-1:0] node1011;
	wire [3-1:0] node1014;
	wire [3-1:0] node1015;
	wire [3-1:0] node1016;
	wire [3-1:0] node1017;
	wire [3-1:0] node1019;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1027;
	wire [3-1:0] node1031;
	wire [3-1:0] node1032;
	wire [3-1:0] node1033;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1041;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1046;
	wire [3-1:0] node1047;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1055;
	wire [3-1:0] node1058;
	wire [3-1:0] node1060;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1066;
	wire [3-1:0] node1068;
	wire [3-1:0] node1070;
	wire [3-1:0] node1072;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1080;
	wire [3-1:0] node1081;
	wire [3-1:0] node1084;
	wire [3-1:0] node1087;
	wire [3-1:0] node1089;
	wire [3-1:0] node1092;
	wire [3-1:0] node1094;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1100;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1108;
	wire [3-1:0] node1109;
	wire [3-1:0] node1110;
	wire [3-1:0] node1113;
	wire [3-1:0] node1117;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1122;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1128;
	wire [3-1:0] node1132;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1135;
	wire [3-1:0] node1136;
	wire [3-1:0] node1138;
	wire [3-1:0] node1139;
	wire [3-1:0] node1141;
	wire [3-1:0] node1144;
	wire [3-1:0] node1147;
	wire [3-1:0] node1148;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1155;
	wire [3-1:0] node1156;
	wire [3-1:0] node1160;
	wire [3-1:0] node1161;
	wire [3-1:0] node1162;
	wire [3-1:0] node1163;
	wire [3-1:0] node1166;
	wire [3-1:0] node1169;
	wire [3-1:0] node1170;
	wire [3-1:0] node1174;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1178;
	wire [3-1:0] node1182;
	wire [3-1:0] node1183;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1191;
	wire [3-1:0] node1193;
	wire [3-1:0] node1197;
	wire [3-1:0] node1199;
	wire [3-1:0] node1200;
	wire [3-1:0] node1204;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1207;
	wire [3-1:0] node1208;
	wire [3-1:0] node1209;
	wire [3-1:0] node1210;
	wire [3-1:0] node1213;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1220;
	wire [3-1:0] node1223;
	wire [3-1:0] node1224;
	wire [3-1:0] node1228;
	wire [3-1:0] node1229;
	wire [3-1:0] node1230;
	wire [3-1:0] node1231;
	wire [3-1:0] node1235;
	wire [3-1:0] node1236;
	wire [3-1:0] node1240;
	wire [3-1:0] node1241;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1248;
	wire [3-1:0] node1251;
	wire [3-1:0] node1254;
	wire [3-1:0] node1255;
	wire [3-1:0] node1259;
	wire [3-1:0] node1261;
	wire [3-1:0] node1262;
	wire [3-1:0] node1265;
	wire [3-1:0] node1268;
	wire [3-1:0] node1269;
	wire [3-1:0] node1270;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1274;
	wire [3-1:0] node1278;
	wire [3-1:0] node1281;
	wire [3-1:0] node1282;
	wire [3-1:0] node1283;
	wire [3-1:0] node1285;
	wire [3-1:0] node1288;
	wire [3-1:0] node1291;
	wire [3-1:0] node1293;
	wire [3-1:0] node1296;
	wire [3-1:0] node1297;
	wire [3-1:0] node1298;
	wire [3-1:0] node1300;
	wire [3-1:0] node1303;
	wire [3-1:0] node1305;
	wire [3-1:0] node1308;
	wire [3-1:0] node1309;
	wire [3-1:0] node1313;
	wire [3-1:0] node1314;
	wire [3-1:0] node1315;
	wire [3-1:0] node1316;
	wire [3-1:0] node1317;
	wire [3-1:0] node1319;
	wire [3-1:0] node1320;
	wire [3-1:0] node1321;
	wire [3-1:0] node1323;
	wire [3-1:0] node1328;
	wire [3-1:0] node1329;
	wire [3-1:0] node1330;
	wire [3-1:0] node1331;
	wire [3-1:0] node1335;
	wire [3-1:0] node1337;
	wire [3-1:0] node1340;
	wire [3-1:0] node1341;
	wire [3-1:0] node1343;
	wire [3-1:0] node1346;
	wire [3-1:0] node1347;
	wire [3-1:0] node1350;
	wire [3-1:0] node1353;
	wire [3-1:0] node1354;
	wire [3-1:0] node1355;
	wire [3-1:0] node1357;
	wire [3-1:0] node1358;
	wire [3-1:0] node1359;
	wire [3-1:0] node1362;
	wire [3-1:0] node1365;
	wire [3-1:0] node1366;
	wire [3-1:0] node1372;
	wire [3-1:0] node1373;
	wire [3-1:0] node1374;
	wire [3-1:0] node1375;
	wire [3-1:0] node1376;
	wire [3-1:0] node1378;
	wire [3-1:0] node1381;
	wire [3-1:0] node1382;
	wire [3-1:0] node1385;
	wire [3-1:0] node1387;
	wire [3-1:0] node1390;
	wire [3-1:0] node1391;
	wire [3-1:0] node1392;
	wire [3-1:0] node1396;
	wire [3-1:0] node1398;
	wire [3-1:0] node1399;
	wire [3-1:0] node1402;
	wire [3-1:0] node1405;
	wire [3-1:0] node1406;
	wire [3-1:0] node1407;
	wire [3-1:0] node1408;
	wire [3-1:0] node1410;
	wire [3-1:0] node1414;
	wire [3-1:0] node1416;
	wire [3-1:0] node1417;
	wire [3-1:0] node1421;
	wire [3-1:0] node1422;
	wire [3-1:0] node1425;
	wire [3-1:0] node1427;
	wire [3-1:0] node1430;
	wire [3-1:0] node1431;
	wire [3-1:0] node1432;
	wire [3-1:0] node1433;
	wire [3-1:0] node1434;
	wire [3-1:0] node1437;
	wire [3-1:0] node1440;
	wire [3-1:0] node1441;
	wire [3-1:0] node1444;
	wire [3-1:0] node1447;
	wire [3-1:0] node1448;
	wire [3-1:0] node1449;
	wire [3-1:0] node1451;
	wire [3-1:0] node1456;
	wire [3-1:0] node1457;
	wire [3-1:0] node1458;
	wire [3-1:0] node1459;
	wire [3-1:0] node1463;
	wire [3-1:0] node1466;
	wire [3-1:0] node1467;
	wire [3-1:0] node1469;
	wire [3-1:0] node1471;
	wire [3-1:0] node1474;
	wire [3-1:0] node1476;
	wire [3-1:0] node1477;
	wire [3-1:0] node1480;
	wire [3-1:0] node1483;
	wire [3-1:0] node1484;
	wire [3-1:0] node1485;
	wire [3-1:0] node1486;
	wire [3-1:0] node1487;
	wire [3-1:0] node1488;
	wire [3-1:0] node1490;
	wire [3-1:0] node1491;
	wire [3-1:0] node1495;
	wire [3-1:0] node1496;
	wire [3-1:0] node1498;
	wire [3-1:0] node1502;
	wire [3-1:0] node1503;
	wire [3-1:0] node1504;
	wire [3-1:0] node1507;
	wire [3-1:0] node1509;
	wire [3-1:0] node1512;
	wire [3-1:0] node1513;
	wire [3-1:0] node1514;
	wire [3-1:0] node1518;
	wire [3-1:0] node1521;
	wire [3-1:0] node1522;
	wire [3-1:0] node1523;
	wire [3-1:0] node1524;
	wire [3-1:0] node1528;
	wire [3-1:0] node1529;
	wire [3-1:0] node1530;
	wire [3-1:0] node1533;
	wire [3-1:0] node1537;
	wire [3-1:0] node1538;
	wire [3-1:0] node1540;
	wire [3-1:0] node1542;
	wire [3-1:0] node1545;
	wire [3-1:0] node1548;
	wire [3-1:0] node1549;
	wire [3-1:0] node1550;
	wire [3-1:0] node1551;
	wire [3-1:0] node1553;
	wire [3-1:0] node1556;
	wire [3-1:0] node1558;
	wire [3-1:0] node1561;
	wire [3-1:0] node1562;
	wire [3-1:0] node1563;
	wire [3-1:0] node1566;
	wire [3-1:0] node1569;
	wire [3-1:0] node1570;
	wire [3-1:0] node1571;
	wire [3-1:0] node1575;
	wire [3-1:0] node1578;
	wire [3-1:0] node1579;
	wire [3-1:0] node1580;
	wire [3-1:0] node1583;
	wire [3-1:0] node1584;
	wire [3-1:0] node1588;
	wire [3-1:0] node1589;
	wire [3-1:0] node1590;
	wire [3-1:0] node1591;
	wire [3-1:0] node1595;
	wire [3-1:0] node1596;
	wire [3-1:0] node1600;
	wire [3-1:0] node1601;
	wire [3-1:0] node1605;
	wire [3-1:0] node1606;
	wire [3-1:0] node1607;
	wire [3-1:0] node1608;
	wire [3-1:0] node1609;
	wire [3-1:0] node1611;
	wire [3-1:0] node1612;
	wire [3-1:0] node1616;
	wire [3-1:0] node1618;
	wire [3-1:0] node1621;
	wire [3-1:0] node1622;
	wire [3-1:0] node1623;
	wire [3-1:0] node1624;
	wire [3-1:0] node1629;
	wire [3-1:0] node1630;
	wire [3-1:0] node1631;
	wire [3-1:0] node1635;
	wire [3-1:0] node1636;
	wire [3-1:0] node1640;
	wire [3-1:0] node1642;
	wire [3-1:0] node1644;
	wire [3-1:0] node1645;
	wire [3-1:0] node1649;
	wire [3-1:0] node1650;
	wire [3-1:0] node1651;
	wire [3-1:0] node1652;
	wire [3-1:0] node1653;
	wire [3-1:0] node1654;
	wire [3-1:0] node1658;
	wire [3-1:0] node1659;
	wire [3-1:0] node1663;
	wire [3-1:0] node1665;
	wire [3-1:0] node1666;
	wire [3-1:0] node1670;
	wire [3-1:0] node1671;
	wire [3-1:0] node1674;
	wire [3-1:0] node1676;
	wire [3-1:0] node1677;
	wire [3-1:0] node1681;
	wire [3-1:0] node1682;
	wire [3-1:0] node1683;
	wire [3-1:0] node1684;
	wire [3-1:0] node1687;
	wire [3-1:0] node1690;
	wire [3-1:0] node1691;
	wire [3-1:0] node1694;
	wire [3-1:0] node1696;
	wire [3-1:0] node1699;
	wire [3-1:0] node1700;
	wire [3-1:0] node1702;
	wire [3-1:0] node1703;
	wire [3-1:0] node1707;
	wire [3-1:0] node1709;
	wire [3-1:0] node1711;
	wire [3-1:0] node1714;
	wire [3-1:0] node1715;
	wire [3-1:0] node1716;
	wire [3-1:0] node1717;
	wire [3-1:0] node1718;
	wire [3-1:0] node1719;
	wire [3-1:0] node1720;
	wire [3-1:0] node1721;
	wire [3-1:0] node1724;
	wire [3-1:0] node1727;
	wire [3-1:0] node1729;
	wire [3-1:0] node1732;
	wire [3-1:0] node1733;
	wire [3-1:0] node1734;
	wire [3-1:0] node1737;
	wire [3-1:0] node1740;
	wire [3-1:0] node1741;
	wire [3-1:0] node1744;
	wire [3-1:0] node1745;
	wire [3-1:0] node1749;
	wire [3-1:0] node1750;
	wire [3-1:0] node1751;
	wire [3-1:0] node1752;
	wire [3-1:0] node1754;
	wire [3-1:0] node1758;
	wire [3-1:0] node1759;
	wire [3-1:0] node1761;
	wire [3-1:0] node1763;
	wire [3-1:0] node1766;
	wire [3-1:0] node1768;
	wire [3-1:0] node1770;
	wire [3-1:0] node1773;
	wire [3-1:0] node1774;
	wire [3-1:0] node1776;
	wire [3-1:0] node1780;
	wire [3-1:0] node1781;
	wire [3-1:0] node1782;
	wire [3-1:0] node1783;
	wire [3-1:0] node1785;
	wire [3-1:0] node1788;
	wire [3-1:0] node1790;
	wire [3-1:0] node1792;
	wire [3-1:0] node1795;
	wire [3-1:0] node1797;
	wire [3-1:0] node1798;
	wire [3-1:0] node1799;
	wire [3-1:0] node1802;
	wire [3-1:0] node1805;
	wire [3-1:0] node1806;
	wire [3-1:0] node1809;
	wire [3-1:0] node1812;
	wire [3-1:0] node1813;
	wire [3-1:0] node1814;
	wire [3-1:0] node1815;
	wire [3-1:0] node1816;
	wire [3-1:0] node1819;
	wire [3-1:0] node1821;
	wire [3-1:0] node1824;
	wire [3-1:0] node1825;
	wire [3-1:0] node1827;
	wire [3-1:0] node1830;
	wire [3-1:0] node1833;
	wire [3-1:0] node1834;
	wire [3-1:0] node1835;
	wire [3-1:0] node1836;
	wire [3-1:0] node1840;
	wire [3-1:0] node1842;
	wire [3-1:0] node1845;
	wire [3-1:0] node1847;
	wire [3-1:0] node1850;
	wire [3-1:0] node1851;
	wire [3-1:0] node1853;
	wire [3-1:0] node1854;
	wire [3-1:0] node1855;
	wire [3-1:0] node1859;
	wire [3-1:0] node1861;
	wire [3-1:0] node1865;
	wire [3-1:0] node1866;
	wire [3-1:0] node1867;
	wire [3-1:0] node1868;
	wire [3-1:0] node1870;
	wire [3-1:0] node1872;
	wire [3-1:0] node1873;
	wire [3-1:0] node1878;
	wire [3-1:0] node1879;
	wire [3-1:0] node1881;
	wire [3-1:0] node1882;
	wire [3-1:0] node1884;
	wire [3-1:0] node1885;
	wire [3-1:0] node1890;
	wire [3-1:0] node1891;
	wire [3-1:0] node1892;
	wire [3-1:0] node1894;
	wire [3-1:0] node1898;
	wire [3-1:0] node1899;
	wire [3-1:0] node1900;
	wire [3-1:0] node1903;
	wire [3-1:0] node1904;
	wire [3-1:0] node1908;
	wire [3-1:0] node1910;
	wire [3-1:0] node1913;
	wire [3-1:0] node1914;
	wire [3-1:0] node1915;
	wire [3-1:0] node1917;
	wire [3-1:0] node1918;
	wire [3-1:0] node1919;
	wire [3-1:0] node1921;
	wire [3-1:0] node1924;
	wire [3-1:0] node1927;
	wire [3-1:0] node1928;
	wire [3-1:0] node1932;
	wire [3-1:0] node1933;
	wire [3-1:0] node1934;
	wire [3-1:0] node1936;
	wire [3-1:0] node1937;
	wire [3-1:0] node1941;
	wire [3-1:0] node1942;
	wire [3-1:0] node1946;
	wire [3-1:0] node1947;
	wire [3-1:0] node1948;
	wire [3-1:0] node1951;
	wire [3-1:0] node1952;
	wire [3-1:0] node1956;
	wire [3-1:0] node1957;
	wire [3-1:0] node1961;
	wire [3-1:0] node1962;
	wire [3-1:0] node1963;
	wire [3-1:0] node1964;
	wire [3-1:0] node1965;
	wire [3-1:0] node1969;
	wire [3-1:0] node1970;
	wire [3-1:0] node1974;
	wire [3-1:0] node1975;
	wire [3-1:0] node1976;
	wire [3-1:0] node1980;
	wire [3-1:0] node1981;
	wire [3-1:0] node1984;
	wire [3-1:0] node1986;
	wire [3-1:0] node1989;
	wire [3-1:0] node1990;
	wire [3-1:0] node1991;
	wire [3-1:0] node1993;
	wire [3-1:0] node1994;
	wire [3-1:0] node1998;
	wire [3-1:0] node1999;
	wire [3-1:0] node2002;
	wire [3-1:0] node2005;
	wire [3-1:0] node2006;
	wire [3-1:0] node2009;
	wire [3-1:0] node2011;
	wire [3-1:0] node2014;
	wire [3-1:0] node2015;
	wire [3-1:0] node2016;
	wire [3-1:0] node2017;
	wire [3-1:0] node2018;
	wire [3-1:0] node2019;
	wire [3-1:0] node2020;
	wire [3-1:0] node2022;
	wire [3-1:0] node2027;
	wire [3-1:0] node2028;
	wire [3-1:0] node2029;
	wire [3-1:0] node2031;
	wire [3-1:0] node2036;
	wire [3-1:0] node2037;
	wire [3-1:0] node2038;
	wire [3-1:0] node2040;
	wire [3-1:0] node2043;
	wire [3-1:0] node2045;
	wire [3-1:0] node2048;
	wire [3-1:0] node2050;
	wire [3-1:0] node2052;
	wire [3-1:0] node2056;
	wire [3-1:0] node2057;
	wire [3-1:0] node2058;
	wire [3-1:0] node2060;
	wire [3-1:0] node2061;
	wire [3-1:0] node2063;
	wire [3-1:0] node2067;
	wire [3-1:0] node2068;
	wire [3-1:0] node2069;
	wire [3-1:0] node2070;
	wire [3-1:0] node2071;
	wire [3-1:0] node2075;
	wire [3-1:0] node2077;
	wire [3-1:0] node2080;
	wire [3-1:0] node2081;
	wire [3-1:0] node2083;
	wire [3-1:0] node2085;
	wire [3-1:0] node2088;
	wire [3-1:0] node2090;
	wire [3-1:0] node2093;
	wire [3-1:0] node2095;
	wire [3-1:0] node2097;
	wire [3-1:0] node2100;
	wire [3-1:0] node2101;
	wire [3-1:0] node2102;
	wire [3-1:0] node2103;
	wire [3-1:0] node2104;
	wire [3-1:0] node2107;
	wire [3-1:0] node2110;
	wire [3-1:0] node2112;
	wire [3-1:0] node2113;
	wire [3-1:0] node2115;
	wire [3-1:0] node2118;
	wire [3-1:0] node2121;
	wire [3-1:0] node2122;
	wire [3-1:0] node2123;
	wire [3-1:0] node2124;
	wire [3-1:0] node2126;
	wire [3-1:0] node2129;
	wire [3-1:0] node2130;
	wire [3-1:0] node2133;
	wire [3-1:0] node2136;
	wire [3-1:0] node2137;
	wire [3-1:0] node2139;
	wire [3-1:0] node2142;
	wire [3-1:0] node2144;
	wire [3-1:0] node2147;
	wire [3-1:0] node2148;
	wire [3-1:0] node2150;
	wire [3-1:0] node2153;
	wire [3-1:0] node2155;
	wire [3-1:0] node2158;
	wire [3-1:0] node2159;
	wire [3-1:0] node2160;
	wire [3-1:0] node2161;
	wire [3-1:0] node2163;
	wire [3-1:0] node2164;
	wire [3-1:0] node2169;
	wire [3-1:0] node2170;
	wire [3-1:0] node2173;
	wire [3-1:0] node2176;
	wire [3-1:0] node2177;
	wire [3-1:0] node2178;
	wire [3-1:0] node2179;
	wire [3-1:0] node2183;
	wire [3-1:0] node2185;
	wire [3-1:0] node2187;
	wire [3-1:0] node2190;
	wire [3-1:0] node2191;
	wire [3-1:0] node2192;
	wire [3-1:0] node2196;
	wire [3-1:0] node2198;
	wire [3-1:0] node2199;
	wire [3-1:0] node2202;

	assign outp = (inp[0]) ? node956 : node1;
		assign node1 = (inp[6]) ? node69 : node2;
			assign node2 = (inp[3]) ? node14 : node3;
				assign node3 = (inp[7]) ? node5 : 3'b011;
					assign node5 = (inp[4]) ? node7 : 3'b011;
						assign node7 = (inp[1]) ? node9 : 3'b111;
							assign node9 = (inp[8]) ? node11 : 3'b111;
								assign node11 = (inp[2]) ? 3'b011 : 3'b111;
				assign node14 = (inp[7]) ? node16 : 3'b111;
					assign node16 = (inp[9]) ? 3'b111 : node17;
						assign node17 = (inp[1]) ? node25 : node18;
							assign node18 = (inp[2]) ? node20 : 3'b111;
								assign node20 = (inp[4]) ? 3'b111 : node21;
									assign node21 = (inp[8]) ? 3'b011 : 3'b111;
							assign node25 = (inp[4]) ? node55 : node26;
								assign node26 = (inp[8]) ? node42 : node27;
									assign node27 = (inp[2]) ? node35 : node28;
										assign node28 = (inp[5]) ? node32 : node29;
											assign node29 = (inp[10]) ? 3'b001 : 3'b101;
											assign node32 = (inp[10]) ? 3'b111 : 3'b011;
										assign node35 = (inp[5]) ? node39 : node36;
											assign node36 = (inp[10]) ? 3'b101 : 3'b001;
											assign node39 = (inp[10]) ? 3'b001 : 3'b101;
									assign node42 = (inp[10]) ? 3'b001 : node43;
										assign node43 = (inp[11]) ? node49 : node44;
											assign node44 = (inp[2]) ? node46 : 3'b001;
												assign node46 = (inp[5]) ? 3'b001 : 3'b101;
											assign node49 = (inp[5]) ? node51 : 3'b001;
												assign node51 = (inp[2]) ? 3'b001 : 3'b101;
								assign node55 = (inp[2]) ? node61 : node56;
									assign node56 = (inp[5]) ? 3'b111 : node57;
										assign node57 = (inp[11]) ? 3'b011 : 3'b111;
									assign node61 = (inp[8]) ? node65 : node62;
										assign node62 = (inp[5]) ? 3'b111 : 3'b011;
										assign node65 = (inp[5]) ? 3'b011 : 3'b101;
			assign node69 = (inp[7]) ? node481 : node70;
				assign node70 = (inp[3]) ? node262 : node71;
					assign node71 = (inp[4]) ? node163 : node72;
						assign node72 = (inp[8]) ? node110 : node73;
							assign node73 = (inp[5]) ? node99 : node74;
								assign node74 = (inp[11]) ? node94 : node75;
									assign node75 = (inp[1]) ? node89 : node76;
										assign node76 = (inp[9]) ? node82 : node77;
											assign node77 = (inp[10]) ? 3'b101 : node78;
												assign node78 = (inp[2]) ? 3'b001 : 3'b101;
											assign node82 = (inp[2]) ? node86 : node83;
												assign node83 = (inp[10]) ? 3'b001 : 3'b101;
												assign node86 = (inp[10]) ? 3'b101 : 3'b001;
										assign node89 = (inp[2]) ? 3'b001 : node90;
											assign node90 = (inp[10]) ? 3'b001 : 3'b101;
									assign node94 = (inp[10]) ? node96 : 3'b001;
										assign node96 = (inp[9]) ? 3'b001 : 3'b101;
								assign node99 = (inp[2]) ? node107 : node100;
									assign node100 = (inp[10]) ? node102 : 3'b001;
										assign node102 = (inp[1]) ? 3'b101 : node103;
											assign node103 = (inp[9]) ? 3'b001 : 3'b101;
									assign node107 = (inp[10]) ? 3'b001 : 3'b101;
							assign node110 = (inp[1]) ? node142 : node111;
								assign node111 = (inp[9]) ? node125 : node112;
									assign node112 = (inp[2]) ? node118 : node113;
										assign node113 = (inp[11]) ? node115 : 3'b101;
											assign node115 = (inp[10]) ? 3'b101 : 3'b001;
										assign node118 = (inp[5]) ? node120 : 3'b001;
											assign node120 = (inp[10]) ? 3'b101 : node121;
												assign node121 = (inp[11]) ? 3'b101 : 3'b001;
									assign node125 = (inp[10]) ? node133 : node126;
										assign node126 = (inp[11]) ? node128 : 3'b001;
											assign node128 = (inp[2]) ? node130 : 3'b101;
												assign node130 = (inp[5]) ? 3'b101 : 3'b001;
										assign node133 = (inp[11]) ? 3'b001 : node134;
											assign node134 = (inp[5]) ? node138 : node135;
												assign node135 = (inp[2]) ? 3'b001 : 3'b101;
												assign node138 = (inp[2]) ? 3'b101 : 3'b001;
								assign node142 = (inp[2]) ? node154 : node143;
									assign node143 = (inp[10]) ? node145 : 3'b101;
										assign node145 = (inp[9]) ? node151 : node146;
											assign node146 = (inp[5]) ? node148 : 3'b101;
												assign node148 = (inp[11]) ? 3'b101 : 3'b001;
											assign node151 = (inp[11]) ? 3'b001 : 3'b101;
									assign node154 = (inp[11]) ? 3'b110 : node155;
										assign node155 = (inp[9]) ? node157 : 3'b010;
											assign node157 = (inp[5]) ? 3'b110 : node158;
												assign node158 = (inp[10]) ? 3'b010 : 3'b110;
						assign node163 = (inp[9]) ? node211 : node164;
							assign node164 = (inp[1]) ? node192 : node165;
								assign node165 = (inp[2]) ? node179 : node166;
									assign node166 = (inp[8]) ? node172 : node167;
										assign node167 = (inp[11]) ? node169 : 3'b101;
											assign node169 = (inp[10]) ? 3'b101 : 3'b001;
										assign node172 = (inp[10]) ? 3'b001 : node173;
											assign node173 = (inp[11]) ? 3'b101 : node174;
												assign node174 = (inp[5]) ? 3'b101 : 3'b001;
									assign node179 = (inp[8]) ? node185 : node180;
										assign node180 = (inp[10]) ? node182 : 3'b001;
											assign node182 = (inp[5]) ? 3'b011 : 3'b001;
										assign node185 = (inp[10]) ? 3'b101 : node186;
											assign node186 = (inp[5]) ? 3'b001 : node187;
												assign node187 = (inp[11]) ? 3'b011 : 3'b111;
								assign node192 = (inp[10]) ? node202 : node193;
									assign node193 = (inp[8]) ? node197 : node194;
										assign node194 = (inp[2]) ? 3'b011 : 3'b111;
										assign node197 = (inp[2]) ? 3'b101 : node198;
											assign node198 = (inp[5]) ? 3'b111 : 3'b011;
									assign node202 = (inp[8]) ? node204 : 3'b001;
										assign node204 = (inp[2]) ? node208 : node205;
											assign node205 = (inp[5]) ? 3'b001 : 3'b011;
											assign node208 = (inp[11]) ? 3'b111 : 3'b011;
							assign node211 = (inp[1]) ? node219 : node212;
								assign node212 = (inp[2]) ? node214 : 3'b111;
									assign node214 = (inp[10]) ? node216 : 3'b011;
										assign node216 = (inp[11]) ? 3'b011 : 3'b111;
								assign node219 = (inp[2]) ? node237 : node220;
									assign node220 = (inp[5]) ? node228 : node221;
										assign node221 = (inp[8]) ? 3'b111 : node222;
											assign node222 = (inp[10]) ? 3'b011 : node223;
												assign node223 = (inp[11]) ? 3'b001 : 3'b011;
										assign node228 = (inp[8]) ? node232 : node229;
											assign node229 = (inp[10]) ? 3'b111 : 3'b101;
											assign node232 = (inp[10]) ? 3'b001 : node233;
												assign node233 = (inp[11]) ? 3'b001 : 3'b011;
									assign node237 = (inp[8]) ? node251 : node238;
										assign node238 = (inp[10]) ? node246 : node239;
											assign node239 = (inp[5]) ? node243 : node240;
												assign node240 = (inp[11]) ? 3'b001 : 3'b111;
												assign node243 = (inp[11]) ? 3'b101 : 3'b001;
											assign node246 = (inp[5]) ? node248 : 3'b101;
												assign node248 = (inp[11]) ? 3'b011 : 3'b101;
										assign node251 = (inp[10]) ? node257 : node252;
											assign node252 = (inp[11]) ? 3'b001 : node253;
												assign node253 = (inp[5]) ? 3'b111 : 3'b101;
											assign node257 = (inp[11]) ? node259 : 3'b001;
												assign node259 = (inp[5]) ? 3'b101 : 3'b001;
					assign node262 = (inp[1]) ? node344 : node263;
						assign node263 = (inp[9]) ? node317 : node264;
							assign node264 = (inp[4]) ? node302 : node265;
								assign node265 = (inp[11]) ? node291 : node266;
									assign node266 = (inp[2]) ? node276 : node267;
										assign node267 = (inp[5]) ? 3'b011 : node268;
											assign node268 = (inp[10]) ? node272 : node269;
												assign node269 = (inp[8]) ? 3'b111 : 3'b011;
												assign node272 = (inp[8]) ? 3'b011 : 3'b111;
										assign node276 = (inp[10]) ? node284 : node277;
											assign node277 = (inp[5]) ? node281 : node278;
												assign node278 = (inp[8]) ? 3'b111 : 3'b101;
												assign node281 = (inp[8]) ? 3'b101 : 3'b011;
											assign node284 = (inp[5]) ? node288 : node285;
												assign node285 = (inp[8]) ? 3'b111 : 3'b011;
												assign node288 = (inp[8]) ? 3'b011 : 3'b111;
									assign node291 = (inp[5]) ? node293 : 3'b011;
										assign node293 = (inp[8]) ? 3'b011 : node294;
											assign node294 = (inp[2]) ? node298 : node295;
												assign node295 = (inp[10]) ? 3'b011 : 3'b111;
												assign node298 = (inp[10]) ? 3'b111 : 3'b011;
								assign node302 = (inp[8]) ? node310 : node303;
									assign node303 = (inp[10]) ? 3'b111 : node304;
										assign node304 = (inp[11]) ? 3'b111 : node305;
											assign node305 = (inp[2]) ? 3'b011 : 3'b111;
									assign node310 = (inp[2]) ? node314 : node311;
										assign node311 = (inp[5]) ? 3'b111 : 3'b101;
										assign node314 = (inp[5]) ? 3'b011 : 3'b001;
							assign node317 = (inp[8]) ? node329 : node318;
								assign node318 = (inp[11]) ? 3'b111 : node319;
									assign node319 = (inp[4]) ? node323 : node320;
										assign node320 = (inp[2]) ? 3'b101 : 3'b111;
										assign node323 = (inp[5]) ? 3'b111 : node324;
											assign node324 = (inp[2]) ? 3'b011 : 3'b111;
								assign node329 = (inp[5]) ? node337 : node330;
									assign node330 = (inp[4]) ? 3'b101 : node331;
										assign node331 = (inp[10]) ? 3'b111 : node332;
											assign node332 = (inp[11]) ? 3'b101 : 3'b111;
									assign node337 = (inp[11]) ? 3'b111 : node338;
										assign node338 = (inp[2]) ? node340 : 3'b111;
											assign node340 = (inp[4]) ? 3'b011 : 3'b101;
						assign node344 = (inp[9]) ? node418 : node345;
							assign node345 = (inp[4]) ? node389 : node346;
								assign node346 = (inp[5]) ? node366 : node347;
									assign node347 = (inp[8]) ? node355 : node348;
										assign node348 = (inp[10]) ? node352 : node349;
											assign node349 = (inp[2]) ? 3'b110 : 3'b001;
											assign node352 = (inp[2]) ? 3'b001 : 3'b110;
										assign node355 = (inp[10]) ? node359 : node356;
											assign node356 = (inp[2]) ? 3'b010 : 3'b110;
											assign node359 = (inp[11]) ? node363 : node360;
												assign node360 = (inp[2]) ? 3'b110 : 3'b010;
												assign node363 = (inp[2]) ? 3'b001 : 3'b101;
									assign node366 = (inp[2]) ? node376 : node367;
										assign node367 = (inp[10]) ? node371 : node368;
											assign node368 = (inp[11]) ? 3'b101 : 3'b001;
											assign node371 = (inp[8]) ? node373 : 3'b010;
												assign node373 = (inp[11]) ? 3'b110 : 3'b101;
										assign node376 = (inp[11]) ? node382 : node377;
											assign node377 = (inp[10]) ? 3'b001 : node378;
												assign node378 = (inp[8]) ? 3'b110 : 3'b001;
											assign node382 = (inp[8]) ? node386 : node383;
												assign node383 = (inp[10]) ? 3'b101 : 3'b001;
												assign node386 = (inp[10]) ? 3'b001 : 3'b101;
								assign node389 = (inp[5]) ? node403 : node390;
									assign node390 = (inp[8]) ? node400 : node391;
										assign node391 = (inp[11]) ? 3'b101 : node392;
											assign node392 = (inp[10]) ? node396 : node393;
												assign node393 = (inp[2]) ? 3'b001 : 3'b101;
												assign node396 = (inp[2]) ? 3'b101 : 3'b001;
										assign node400 = (inp[2]) ? 3'b110 : 3'b001;
									assign node403 = (inp[8]) ? node411 : node404;
										assign node404 = (inp[2]) ? node408 : node405;
											assign node405 = (inp[10]) ? 3'b111 : 3'b011;
											assign node408 = (inp[11]) ? 3'b001 : 3'b101;
										assign node411 = (inp[10]) ? node415 : node412;
											assign node412 = (inp[2]) ? 3'b001 : 3'b101;
											assign node415 = (inp[2]) ? 3'b101 : 3'b001;
							assign node418 = (inp[8]) ? node450 : node419;
								assign node419 = (inp[5]) ? node437 : node420;
									assign node420 = (inp[2]) ? node432 : node421;
										assign node421 = (inp[10]) ? node427 : node422;
											assign node422 = (inp[11]) ? 3'b111 : node423;
												assign node423 = (inp[4]) ? 3'b111 : 3'b101;
											assign node427 = (inp[4]) ? node429 : 3'b111;
												assign node429 = (inp[11]) ? 3'b001 : 3'b011;
										assign node432 = (inp[10]) ? node434 : 3'b011;
											assign node434 = (inp[4]) ? 3'b111 : 3'b011;
									assign node437 = (inp[11]) ? node445 : node438;
										assign node438 = (inp[10]) ? node442 : node439;
											assign node439 = (inp[4]) ? 3'b111 : 3'b101;
											assign node442 = (inp[4]) ? 3'b101 : 3'b111;
										assign node445 = (inp[4]) ? node447 : 3'b111;
											assign node447 = (inp[2]) ? 3'b111 : 3'b011;
								assign node450 = (inp[4]) ? node466 : node451;
									assign node451 = (inp[2]) ? node461 : node452;
										assign node452 = (inp[5]) ? 3'b111 : node453;
											assign node453 = (inp[10]) ? node457 : node454;
												assign node454 = (inp[11]) ? 3'b001 : 3'b011;
												assign node457 = (inp[11]) ? 3'b011 : 3'b001;
										assign node461 = (inp[10]) ? 3'b001 : node462;
											assign node462 = (inp[11]) ? 3'b001 : 3'b011;
									assign node466 = (inp[2]) ? node474 : node467;
										assign node467 = (inp[11]) ? node471 : node468;
											assign node468 = (inp[5]) ? 3'b011 : 3'b111;
											assign node471 = (inp[5]) ? 3'b001 : 3'b011;
										assign node474 = (inp[11]) ? 3'b111 : node475;
											assign node475 = (inp[5]) ? 3'b011 : node476;
												assign node476 = (inp[10]) ? 3'b011 : 3'b111;
				assign node481 = (inp[3]) ? node713 : node482;
					assign node482 = (inp[1]) ? node634 : node483;
						assign node483 = (inp[4]) ? node553 : node484;
							assign node484 = (inp[9]) ? node522 : node485;
								assign node485 = (inp[10]) ? node501 : node486;
									assign node486 = (inp[11]) ? node496 : node487;
										assign node487 = (inp[5]) ? node489 : 3'b000;
											assign node489 = (inp[2]) ? node493 : node490;
												assign node490 = (inp[8]) ? 3'b100 : 3'b000;
												assign node493 = (inp[8]) ? 3'b000 : 3'b100;
										assign node496 = (inp[5]) ? node498 : 3'b100;
											assign node498 = (inp[8]) ? 3'b100 : 3'b000;
									assign node501 = (inp[11]) ? node511 : node502;
										assign node502 = (inp[2]) ? 3'b100 : node503;
											assign node503 = (inp[5]) ? node507 : node504;
												assign node504 = (inp[8]) ? 3'b000 : 3'b100;
												assign node507 = (inp[8]) ? 3'b100 : 3'b000;
										assign node511 = (inp[8]) ? node517 : node512;
											assign node512 = (inp[5]) ? 3'b100 : node513;
												assign node513 = (inp[2]) ? 3'b000 : 3'b100;
											assign node517 = (inp[5]) ? node519 : 3'b000;
												assign node519 = (inp[2]) ? 3'b000 : 3'b100;
								assign node522 = (inp[2]) ? node538 : node523;
									assign node523 = (inp[5]) ? node533 : node524;
										assign node524 = (inp[8]) ? node530 : node525;
											assign node525 = (inp[10]) ? 3'b101 : node526;
												assign node526 = (inp[11]) ? 3'b101 : 3'b100;
											assign node530 = (inp[10]) ? 3'b001 : 3'b000;
										assign node533 = (inp[8]) ? node535 : 3'b011;
											assign node535 = (inp[11]) ? 3'b101 : 3'b100;
									assign node538 = (inp[10]) ? node550 : node539;
										assign node539 = (inp[11]) ? node545 : node540;
											assign node540 = (inp[8]) ? node542 : 3'b000;
												assign node542 = (inp[5]) ? 3'b000 : 3'b010;
											assign node545 = (inp[8]) ? node547 : 3'b100;
												assign node547 = (inp[5]) ? 3'b100 : 3'b010;
										assign node550 = (inp[5]) ? 3'b100 : 3'b110;
							assign node553 = (inp[9]) ? node595 : node554;
								assign node554 = (inp[10]) ? node576 : node555;
									assign node555 = (inp[2]) ? node567 : node556;
										assign node556 = (inp[8]) ? node560 : node557;
											assign node557 = (inp[5]) ? 3'b011 : 3'b111;
											assign node560 = (inp[11]) ? node564 : node561;
												assign node561 = (inp[5]) ? 3'b110 : 3'b010;
												assign node564 = (inp[5]) ? 3'b111 : 3'b110;
										assign node567 = (inp[11]) ? node569 : 3'b100;
											assign node569 = (inp[5]) ? node573 : node570;
												assign node570 = (inp[8]) ? 3'b100 : 3'b010;
												assign node573 = (inp[8]) ? 3'b010 : 3'b110;
									assign node576 = (inp[5]) ? node586 : node577;
										assign node577 = (inp[2]) ? node581 : node578;
											assign node578 = (inp[11]) ? 3'b011 : 3'b111;
											assign node581 = (inp[11]) ? node583 : 3'b010;
												assign node583 = (inp[8]) ? 3'b110 : 3'b111;
										assign node586 = (inp[2]) ? node590 : node587;
											assign node587 = (inp[8]) ? 3'b001 : 3'b101;
											assign node590 = (inp[8]) ? node592 : 3'b001;
												assign node592 = (inp[11]) ? 3'b111 : 3'b110;
								assign node595 = (inp[11]) ? node613 : node596;
									assign node596 = (inp[2]) ? node602 : node597;
										assign node597 = (inp[8]) ? 3'b101 : node598;
											assign node598 = (inp[5]) ? 3'b001 : 3'b101;
										assign node602 = (inp[10]) ? node608 : node603;
											assign node603 = (inp[8]) ? node605 : 3'b001;
												assign node605 = (inp[5]) ? 3'b001 : 3'b101;
											assign node608 = (inp[8]) ? node610 : 3'b101;
												assign node610 = (inp[5]) ? 3'b101 : 3'b001;
									assign node613 = (inp[10]) ? node625 : node614;
										assign node614 = (inp[2]) ? node620 : node615;
											assign node615 = (inp[5]) ? node617 : 3'b101;
												assign node617 = (inp[8]) ? 3'b101 : 3'b001;
											assign node620 = (inp[8]) ? 3'b001 : node621;
												assign node621 = (inp[5]) ? 3'b111 : 3'b001;
										assign node625 = (inp[2]) ? node629 : node626;
											assign node626 = (inp[5]) ? 3'b111 : 3'b011;
											assign node629 = (inp[8]) ? 3'b101 : node630;
												assign node630 = (inp[5]) ? 3'b011 : 3'b101;
						assign node634 = (inp[9]) ? node664 : node635;
							assign node635 = (inp[4]) ? node637 : 3'b000;
								assign node637 = (inp[8]) ? node647 : node638;
									assign node638 = (inp[2]) ? node642 : node639;
										assign node639 = (inp[10]) ? 3'b010 : 3'b000;
										assign node642 = (inp[5]) ? 3'b000 : node643;
											assign node643 = (inp[10]) ? 3'b100 : 3'b000;
									assign node647 = (inp[10]) ? node655 : node648;
										assign node648 = (inp[2]) ? 3'b000 : node649;
											assign node649 = (inp[11]) ? node651 : 3'b100;
												assign node651 = (inp[5]) ? 3'b000 : 3'b100;
										assign node655 = (inp[5]) ? node659 : node656;
											assign node656 = (inp[11]) ? 3'b100 : 3'b000;
											assign node659 = (inp[11]) ? node661 : 3'b100;
												assign node661 = (inp[2]) ? 3'b100 : 3'b010;
							assign node664 = (inp[8]) ? node696 : node665;
								assign node665 = (inp[5]) ? node683 : node666;
									assign node666 = (inp[4]) ? node676 : node667;
										assign node667 = (inp[2]) ? node669 : 3'b110;
											assign node669 = (inp[11]) ? node673 : node670;
												assign node670 = (inp[10]) ? 3'b100 : 3'b000;
												assign node673 = (inp[10]) ? 3'b010 : 3'b100;
										assign node676 = (inp[2]) ? node680 : node677;
											assign node677 = (inp[10]) ? 3'b001 : 3'b110;
											assign node680 = (inp[10]) ? 3'b110 : 3'b010;
									assign node683 = (inp[2]) ? node689 : node684;
										assign node684 = (inp[10]) ? node686 : 3'b110;
											assign node686 = (inp[4]) ? 3'b101 : 3'b001;
										assign node689 = (inp[4]) ? node693 : node690;
											assign node690 = (inp[11]) ? 3'b110 : 3'b010;
											assign node693 = (inp[10]) ? 3'b001 : 3'b011;
								assign node696 = (inp[5]) ? node698 : 3'b010;
									assign node698 = (inp[2]) ? node704 : node699;
										assign node699 = (inp[10]) ? node701 : 3'b110;
											assign node701 = (inp[4]) ? 3'b001 : 3'b110;
										assign node704 = (inp[10]) ? node710 : node705;
											assign node705 = (inp[4]) ? 3'b010 : node706;
												assign node706 = (inp[11]) ? 3'b100 : 3'b000;
											assign node710 = (inp[4]) ? 3'b110 : 3'b010;
					assign node713 = (inp[9]) ? node859 : node714;
						assign node714 = (inp[1]) ? node790 : node715;
							assign node715 = (inp[2]) ? node753 : node716;
								assign node716 = (inp[10]) ? node732 : node717;
									assign node717 = (inp[8]) ? node725 : node718;
										assign node718 = (inp[5]) ? 3'b101 : node719;
											assign node719 = (inp[11]) ? node721 : 3'b001;
												assign node721 = (inp[4]) ? 3'b111 : 3'b101;
										assign node725 = (inp[4]) ? 3'b011 : node726;
											assign node726 = (inp[5]) ? node728 : 3'b001;
												assign node728 = (inp[11]) ? 3'b101 : 3'b001;
									assign node732 = (inp[11]) ? node746 : node733;
										assign node733 = (inp[8]) ? node739 : node734;
											assign node734 = (inp[5]) ? 3'b011 : node735;
												assign node735 = (inp[4]) ? 3'b011 : 3'b101;
											assign node739 = (inp[5]) ? node743 : node740;
												assign node740 = (inp[4]) ? 3'b101 : 3'b001;
												assign node743 = (inp[4]) ? 3'b011 : 3'b101;
										assign node746 = (inp[8]) ? 3'b011 : node747;
											assign node747 = (inp[5]) ? 3'b101 : node748;
												assign node748 = (inp[4]) ? 3'b111 : 3'b011;
								assign node753 = (inp[4]) ? node773 : node754;
									assign node754 = (inp[10]) ? node764 : node755;
										assign node755 = (inp[8]) ? node759 : node756;
											assign node756 = (inp[5]) ? 3'b001 : 3'b010;
											assign node759 = (inp[5]) ? node761 : 3'b110;
												assign node761 = (inp[11]) ? 3'b010 : 3'b110;
										assign node764 = (inp[8]) ? node766 : 3'b110;
											assign node766 = (inp[11]) ? node770 : node767;
												assign node767 = (inp[5]) ? 3'b001 : 3'b101;
												assign node770 = (inp[5]) ? 3'b101 : 3'b001;
									assign node773 = (inp[11]) ? node781 : node774;
										assign node774 = (inp[10]) ? 3'b101 : node775;
											assign node775 = (inp[5]) ? node777 : 3'b001;
												assign node777 = (inp[8]) ? 3'b001 : 3'b111;
										assign node781 = (inp[5]) ? node787 : node782;
											assign node782 = (inp[8]) ? node784 : 3'b011;
												assign node784 = (inp[10]) ? 3'b101 : 3'b001;
											assign node787 = (inp[10]) ? 3'b011 : 3'b111;
							assign node790 = (inp[2]) ? node824 : node791;
								assign node791 = (inp[4]) ? node809 : node792;
									assign node792 = (inp[10]) ? node796 : node793;
										assign node793 = (inp[8]) ? 3'b100 : 3'b110;
										assign node796 = (inp[11]) ? node804 : node797;
											assign node797 = (inp[5]) ? node801 : node798;
												assign node798 = (inp[8]) ? 3'b000 : 3'b110;
												assign node801 = (inp[8]) ? 3'b110 : 3'b001;
											assign node804 = (inp[5]) ? 3'b001 : node805;
												assign node805 = (inp[8]) ? 3'b110 : 3'b001;
									assign node809 = (inp[10]) ? node817 : node810;
										assign node810 = (inp[8]) ? node812 : 3'b001;
											assign node812 = (inp[5]) ? node814 : 3'b110;
												assign node814 = (inp[11]) ? 3'b001 : 3'b110;
										assign node817 = (inp[11]) ? node819 : 3'b001;
											assign node819 = (inp[8]) ? node821 : 3'b101;
												assign node821 = (inp[5]) ? 3'b101 : 3'b001;
								assign node824 = (inp[5]) ? node840 : node825;
									assign node825 = (inp[4]) ? node835 : node826;
										assign node826 = (inp[11]) ? node832 : node827;
											assign node827 = (inp[8]) ? node829 : 3'b100;
												assign node829 = (inp[10]) ? 3'b100 : 3'b000;
											assign node832 = (inp[10]) ? 3'b010 : 3'b110;
										assign node835 = (inp[10]) ? 3'b110 : node836;
											assign node836 = (inp[8]) ? 3'b010 : 3'b110;
									assign node840 = (inp[4]) ? node850 : node841;
										assign node841 = (inp[11]) ? node845 : node842;
											assign node842 = (inp[8]) ? 3'b100 : 3'b010;
											assign node845 = (inp[8]) ? 3'b010 : node846;
												assign node846 = (inp[10]) ? 3'b110 : 3'b010;
										assign node850 = (inp[10]) ? node854 : node851;
											assign node851 = (inp[11]) ? 3'b110 : 3'b010;
											assign node854 = (inp[8]) ? node856 : 3'b001;
												assign node856 = (inp[11]) ? 3'b001 : 3'b110;
						assign node859 = (inp[1]) ? node899 : node860;
							assign node860 = (inp[4]) ? node892 : node861;
								assign node861 = (inp[11]) ? node881 : node862;
									assign node862 = (inp[10]) ? node872 : node863;
										assign node863 = (inp[8]) ? 3'b001 : node864;
											assign node864 = (inp[2]) ? node868 : node865;
												assign node865 = (inp[5]) ? 3'b101 : 3'b011;
												assign node868 = (inp[5]) ? 3'b011 : 3'b101;
										assign node872 = (inp[2]) ? node876 : node873;
											assign node873 = (inp[8]) ? 3'b011 : 3'b111;
											assign node876 = (inp[5]) ? 3'b011 : node877;
												assign node877 = (inp[8]) ? 3'b101 : 3'b011;
									assign node881 = (inp[2]) ? node883 : 3'b111;
										assign node883 = (inp[10]) ? node887 : node884;
											assign node884 = (inp[5]) ? 3'b011 : 3'b101;
											assign node887 = (inp[5]) ? 3'b111 : node888;
												assign node888 = (inp[8]) ? 3'b011 : 3'b111;
								assign node892 = (inp[10]) ? 3'b111 : node893;
									assign node893 = (inp[2]) ? node895 : 3'b111;
										assign node895 = (inp[11]) ? 3'b111 : 3'b011;
							assign node899 = (inp[4]) ? node927 : node900;
								assign node900 = (inp[10]) ? node918 : node901;
									assign node901 = (inp[2]) ? node911 : node902;
										assign node902 = (inp[8]) ? node906 : node903;
											assign node903 = (inp[5]) ? 3'b110 : 3'b001;
											assign node906 = (inp[5]) ? node908 : 3'b110;
												assign node908 = (inp[11]) ? 3'b101 : 3'b001;
										assign node911 = (inp[11]) ? 3'b110 : node912;
											assign node912 = (inp[8]) ? 3'b110 : node913;
												assign node913 = (inp[5]) ? 3'b010 : 3'b110;
									assign node918 = (inp[8]) ? node922 : node919;
										assign node919 = (inp[11]) ? 3'b100 : 3'b111;
										assign node922 = (inp[11]) ? node924 : 3'b001;
											assign node924 = (inp[2]) ? 3'b001 : 3'b101;
								assign node927 = (inp[2]) ? node945 : node928;
									assign node928 = (inp[10]) ? node938 : node929;
										assign node929 = (inp[8]) ? 3'b101 : node930;
											assign node930 = (inp[11]) ? node934 : node931;
												assign node931 = (inp[5]) ? 3'b011 : 3'b101;
												assign node934 = (inp[5]) ? 3'b111 : 3'b011;
										assign node938 = (inp[11]) ? 3'b111 : node939;
											assign node939 = (inp[8]) ? 3'b011 : node940;
												assign node940 = (inp[5]) ? 3'b111 : 3'b011;
									assign node945 = (inp[8]) ? node951 : node946;
										assign node946 = (inp[10]) ? node948 : 3'b101;
											assign node948 = (inp[11]) ? 3'b011 : 3'b101;
										assign node951 = (inp[10]) ? node953 : 3'b001;
											assign node953 = (inp[5]) ? 3'b011 : 3'b101;
		assign node956 = (inp[6]) ? node1714 : node957;
			assign node957 = (inp[3]) ? node1313 : node958;
				assign node958 = (inp[4]) ? node1132 : node959;
					assign node959 = (inp[9]) ? node1063 : node960;
						assign node960 = (inp[7]) ? node1014 : node961;
							assign node961 = (inp[1]) ? node981 : node962;
								assign node962 = (inp[2]) ? node970 : node963;
									assign node963 = (inp[11]) ? node965 : 3'b010;
										assign node965 = (inp[8]) ? node967 : 3'b110;
											assign node967 = (inp[5]) ? 3'b110 : 3'b010;
									assign node970 = (inp[5]) ? node976 : node971;
										assign node971 = (inp[8]) ? 3'b100 : node972;
											assign node972 = (inp[11]) ? 3'b010 : 3'b100;
										assign node976 = (inp[11]) ? node978 : 3'b010;
											assign node978 = (inp[8]) ? 3'b010 : 3'b110;
								assign node981 = (inp[10]) ? node995 : node982;
									assign node982 = (inp[2]) ? node990 : node983;
										assign node983 = (inp[5]) ? 3'b100 : node984;
											assign node984 = (inp[8]) ? 3'b000 : node985;
												assign node985 = (inp[11]) ? 3'b100 : 3'b000;
										assign node990 = (inp[8]) ? node992 : 3'b000;
											assign node992 = (inp[5]) ? 3'b110 : 3'b010;
									assign node995 = (inp[8]) ? node1003 : node996;
										assign node996 = (inp[2]) ? 3'b110 : node997;
											assign node997 = (inp[11]) ? 3'b010 : node998;
												assign node998 = (inp[5]) ? 3'b010 : 3'b100;
										assign node1003 = (inp[11]) ? node1011 : node1004;
											assign node1004 = (inp[5]) ? node1008 : node1005;
												assign node1005 = (inp[2]) ? 3'b100 : 3'b000;
												assign node1008 = (inp[2]) ? 3'b000 : 3'b100;
											assign node1011 = (inp[5]) ? 3'b010 : 3'b000;
							assign node1014 = (inp[1]) ? node1038 : node1015;
								assign node1015 = (inp[2]) ? node1023 : node1016;
									assign node1016 = (inp[8]) ? 3'b000 : node1017;
										assign node1017 = (inp[11]) ? node1019 : 3'b100;
											assign node1019 = (inp[10]) ? 3'b100 : 3'b000;
									assign node1023 = (inp[8]) ? node1031 : node1024;
										assign node1024 = (inp[5]) ? 3'b010 : node1025;
											assign node1025 = (inp[11]) ? node1027 : 3'b000;
												assign node1027 = (inp[10]) ? 3'b000 : 3'b100;
										assign node1031 = (inp[10]) ? 3'b100 : node1032;
											assign node1032 = (inp[5]) ? 3'b000 : node1033;
												assign node1033 = (inp[11]) ? 3'b010 : 3'b110;
								assign node1038 = (inp[10]) ? node1044 : node1039;
									assign node1039 = (inp[2]) ? node1041 : 3'b110;
										assign node1041 = (inp[8]) ? 3'b100 : 3'b010;
									assign node1044 = (inp[8]) ? node1052 : node1045;
										assign node1045 = (inp[2]) ? 3'b100 : node1046;
											assign node1046 = (inp[5]) ? 3'b000 : node1047;
												assign node1047 = (inp[11]) ? 3'b000 : 3'b010;
										assign node1052 = (inp[2]) ? node1058 : node1053;
											assign node1053 = (inp[11]) ? node1055 : 3'b010;
												assign node1055 = (inp[5]) ? 3'b000 : 3'b010;
											assign node1058 = (inp[11]) ? node1060 : 3'b010;
												assign node1060 = (inp[5]) ? 3'b110 : 3'b010;
						assign node1063 = (inp[1]) ? node1075 : node1064;
							assign node1064 = (inp[7]) ? node1066 : 3'b110;
								assign node1066 = (inp[2]) ? node1068 : 3'b110;
									assign node1068 = (inp[10]) ? node1070 : 3'b010;
										assign node1070 = (inp[8]) ? node1072 : 3'b110;
											assign node1072 = (inp[5]) ? 3'b110 : 3'b010;
							assign node1075 = (inp[7]) ? node1097 : node1076;
								assign node1076 = (inp[2]) ? node1078 : 3'b110;
									assign node1078 = (inp[10]) ? node1092 : node1079;
										assign node1079 = (inp[5]) ? node1087 : node1080;
											assign node1080 = (inp[8]) ? node1084 : node1081;
												assign node1081 = (inp[11]) ? 3'b010 : 3'b100;
												assign node1084 = (inp[11]) ? 3'b100 : 3'b010;
											assign node1087 = (inp[8]) ? node1089 : 3'b010;
												assign node1089 = (inp[11]) ? 3'b010 : 3'b100;
										assign node1092 = (inp[11]) ? node1094 : 3'b010;
											assign node1094 = (inp[8]) ? 3'b010 : 3'b110;
								assign node1097 = (inp[11]) ? node1117 : node1098;
									assign node1098 = (inp[10]) ? node1108 : node1099;
										assign node1099 = (inp[5]) ? node1103 : node1100;
											assign node1100 = (inp[2]) ? 3'b110 : 3'b010;
											assign node1103 = (inp[8]) ? 3'b110 : node1104;
												assign node1104 = (inp[2]) ? 3'b000 : 3'b100;
										assign node1108 = (inp[5]) ? 3'b000 : node1109;
											assign node1109 = (inp[2]) ? node1113 : node1110;
												assign node1110 = (inp[8]) ? 3'b110 : 3'b000;
												assign node1113 = (inp[8]) ? 3'b000 : 3'b100;
									assign node1117 = (inp[10]) ? node1125 : node1118;
										assign node1118 = (inp[5]) ? node1122 : node1119;
											assign node1119 = (inp[8]) ? 3'b110 : 3'b000;
											assign node1122 = (inp[8]) ? 3'b000 : 3'b100;
										assign node1125 = (inp[8]) ? 3'b100 : node1126;
											assign node1126 = (inp[5]) ? node1128 : 3'b100;
												assign node1128 = (inp[2]) ? 3'b010 : 3'b110;
					assign node1132 = (inp[9]) ? node1204 : node1133;
						assign node1133 = (inp[1]) ? node1187 : node1134;
							assign node1134 = (inp[7]) ? node1160 : node1135;
								assign node1135 = (inp[5]) ? node1147 : node1136;
									assign node1136 = (inp[2]) ? node1138 : 3'b110;
										assign node1138 = (inp[10]) ? node1144 : node1139;
											assign node1139 = (inp[11]) ? node1141 : 3'b001;
												assign node1141 = (inp[8]) ? 3'b001 : 3'b110;
											assign node1144 = (inp[11]) ? 3'b001 : 3'b110;
									assign node1147 = (inp[10]) ? node1155 : node1148;
										assign node1148 = (inp[2]) ? node1150 : 3'b001;
											assign node1150 = (inp[11]) ? 3'b110 : node1151;
												assign node1151 = (inp[8]) ? 3'b001 : 3'b110;
										assign node1155 = (inp[2]) ? 3'b001 : node1156;
											assign node1156 = (inp[8]) ? 3'b001 : 3'b110;
								assign node1160 = (inp[2]) ? node1174 : node1161;
									assign node1161 = (inp[8]) ? node1169 : node1162;
										assign node1162 = (inp[5]) ? node1166 : node1163;
											assign node1163 = (inp[10]) ? 3'b101 : 3'b001;
											assign node1166 = (inp[10]) ? 3'b011 : 3'b111;
										assign node1169 = (inp[10]) ? 3'b101 : node1170;
											assign node1170 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1174 = (inp[11]) ? node1182 : node1175;
										assign node1175 = (inp[5]) ? 3'b001 : node1176;
											assign node1176 = (inp[10]) ? node1178 : 3'b101;
												assign node1178 = (inp[8]) ? 3'b101 : 3'b001;
										assign node1182 = (inp[8]) ? 3'b001 : node1183;
											assign node1183 = (inp[5]) ? 3'b101 : 3'b001;
							assign node1187 = (inp[7]) ? node1197 : node1188;
								assign node1188 = (inp[2]) ? 3'b001 : node1189;
									assign node1189 = (inp[10]) ? node1191 : 3'b001;
										assign node1191 = (inp[11]) ? node1193 : 3'b001;
											assign node1193 = (inp[5]) ? 3'b110 : 3'b001;
								assign node1197 = (inp[5]) ? node1199 : 3'b000;
									assign node1199 = (inp[2]) ? 3'b000 : node1200;
										assign node1200 = (inp[8]) ? 3'b000 : 3'b001;
						assign node1204 = (inp[1]) ? node1268 : node1205;
							assign node1205 = (inp[7]) ? node1245 : node1206;
								assign node1206 = (inp[5]) ? node1228 : node1207;
									assign node1207 = (inp[10]) ? node1217 : node1208;
										assign node1208 = (inp[8]) ? 3'b110 : node1209;
											assign node1209 = (inp[2]) ? node1213 : node1210;
												assign node1210 = (inp[11]) ? 3'b001 : 3'b110;
												assign node1213 = (inp[11]) ? 3'b110 : 3'b001;
										assign node1217 = (inp[2]) ? node1223 : node1218;
											assign node1218 = (inp[11]) ? node1220 : 3'b001;
												assign node1220 = (inp[8]) ? 3'b001 : 3'b110;
											assign node1223 = (inp[8]) ? 3'b110 : node1224;
												assign node1224 = (inp[11]) ? 3'b001 : 3'b110;
									assign node1228 = (inp[2]) ? node1240 : node1229;
										assign node1229 = (inp[10]) ? node1235 : node1230;
											assign node1230 = (inp[11]) ? 3'b001 : node1231;
												assign node1231 = (inp[8]) ? 3'b110 : 3'b001;
											assign node1235 = (inp[11]) ? 3'b110 : node1236;
												assign node1236 = (inp[8]) ? 3'b001 : 3'b110;
										assign node1240 = (inp[10]) ? 3'b001 : node1241;
											assign node1241 = (inp[8]) ? 3'b001 : 3'b110;
								assign node1245 = (inp[8]) ? node1259 : node1246;
									assign node1246 = (inp[2]) ? node1254 : node1247;
										assign node1247 = (inp[5]) ? node1251 : node1248;
											assign node1248 = (inp[10]) ? 3'b101 : 3'b001;
											assign node1251 = (inp[10]) ? 3'b011 : 3'b111;
										assign node1254 = (inp[5]) ? 3'b101 : node1255;
											assign node1255 = (inp[10]) ? 3'b001 : 3'b101;
									assign node1259 = (inp[5]) ? node1261 : 3'b001;
										assign node1261 = (inp[10]) ? node1265 : node1262;
											assign node1262 = (inp[2]) ? 3'b101 : 3'b001;
											assign node1265 = (inp[2]) ? 3'b001 : 3'b101;
							assign node1268 = (inp[7]) ? node1296 : node1269;
								assign node1269 = (inp[8]) ? node1281 : node1270;
									assign node1270 = (inp[2]) ? node1272 : 3'b110;
										assign node1272 = (inp[10]) ? node1278 : node1273;
											assign node1273 = (inp[11]) ? 3'b110 : node1274;
												assign node1274 = (inp[5]) ? 3'b110 : 3'b001;
											assign node1278 = (inp[5]) ? 3'b001 : 3'b110;
									assign node1281 = (inp[11]) ? node1291 : node1282;
										assign node1282 = (inp[2]) ? node1288 : node1283;
											assign node1283 = (inp[10]) ? node1285 : 3'b110;
												assign node1285 = (inp[5]) ? 3'b001 : 3'b110;
											assign node1288 = (inp[5]) ? 3'b110 : 3'b001;
										assign node1291 = (inp[10]) ? node1293 : 3'b001;
											assign node1293 = (inp[5]) ? 3'b001 : 3'b110;
								assign node1296 = (inp[8]) ? node1308 : node1297;
									assign node1297 = (inp[10]) ? node1303 : node1298;
										assign node1298 = (inp[2]) ? node1300 : 3'b110;
											assign node1300 = (inp[5]) ? 3'b110 : 3'b010;
										assign node1303 = (inp[2]) ? node1305 : 3'b001;
											assign node1305 = (inp[5]) ? 3'b110 : 3'b010;
									assign node1308 = (inp[5]) ? 3'b010 : node1309;
										assign node1309 = (inp[2]) ? 3'b100 : 3'b110;
				assign node1313 = (inp[7]) ? node1483 : node1314;
					assign node1314 = (inp[1]) ? node1372 : node1315;
						assign node1315 = (inp[9]) ? node1353 : node1316;
							assign node1316 = (inp[4]) ? node1328 : node1317;
								assign node1317 = (inp[2]) ? node1319 : 3'b111;
									assign node1319 = (inp[10]) ? 3'b111 : node1320;
										assign node1320 = (inp[5]) ? 3'b111 : node1321;
											assign node1321 = (inp[11]) ? node1323 : 3'b011;
												assign node1323 = (inp[8]) ? 3'b011 : 3'b111;
								assign node1328 = (inp[2]) ? node1340 : node1329;
									assign node1329 = (inp[8]) ? node1335 : node1330;
										assign node1330 = (inp[5]) ? 3'b111 : node1331;
											assign node1331 = (inp[11]) ? 3'b111 : 3'b011;
										assign node1335 = (inp[5]) ? node1337 : 3'b011;
											assign node1337 = (inp[11]) ? 3'b111 : 3'b011;
									assign node1340 = (inp[5]) ? node1346 : node1341;
										assign node1341 = (inp[11]) ? node1343 : 3'b101;
											assign node1343 = (inp[8]) ? 3'b101 : 3'b011;
										assign node1346 = (inp[8]) ? node1350 : node1347;
											assign node1347 = (inp[11]) ? 3'b111 : 3'b011;
											assign node1350 = (inp[11]) ? 3'b011 : 3'b101;
							assign node1353 = (inp[4]) ? 3'b111 : node1354;
								assign node1354 = (inp[10]) ? 3'b111 : node1355;
									assign node1355 = (inp[2]) ? node1357 : 3'b111;
										assign node1357 = (inp[11]) ? node1365 : node1358;
											assign node1358 = (inp[8]) ? node1362 : node1359;
												assign node1359 = (inp[5]) ? 3'b111 : 3'b011;
												assign node1362 = (inp[5]) ? 3'b011 : 3'b111;
											assign node1365 = (inp[5]) ? 3'b111 : node1366;
												assign node1366 = (inp[8]) ? 3'b011 : 3'b111;
						assign node1372 = (inp[9]) ? node1430 : node1373;
							assign node1373 = (inp[4]) ? node1405 : node1374;
								assign node1374 = (inp[5]) ? node1390 : node1375;
									assign node1375 = (inp[8]) ? node1381 : node1376;
										assign node1376 = (inp[10]) ? node1378 : 3'b010;
											assign node1378 = (inp[2]) ? 3'b110 : 3'b010;
										assign node1381 = (inp[10]) ? node1385 : node1382;
											assign node1382 = (inp[2]) ? 3'b100 : 3'b000;
											assign node1385 = (inp[2]) ? node1387 : 3'b100;
												assign node1387 = (inp[11]) ? 3'b100 : 3'b000;
									assign node1390 = (inp[8]) ? node1396 : node1391;
										assign node1391 = (inp[2]) ? 3'b010 : node1392;
											assign node1392 = (inp[10]) ? 3'b111 : 3'b011;
										assign node1396 = (inp[11]) ? node1398 : 3'b010;
											assign node1398 = (inp[2]) ? node1402 : node1399;
												assign node1399 = (inp[10]) ? 3'b010 : 3'b110;
												assign node1402 = (inp[10]) ? 3'b110 : 3'b010;
								assign node1405 = (inp[2]) ? node1421 : node1406;
									assign node1406 = (inp[10]) ? node1414 : node1407;
										assign node1407 = (inp[11]) ? 3'b101 : node1408;
											assign node1408 = (inp[5]) ? node1410 : 3'b001;
												assign node1410 = (inp[8]) ? 3'b001 : 3'b101;
										assign node1414 = (inp[8]) ? node1416 : 3'b011;
											assign node1416 = (inp[11]) ? 3'b101 : node1417;
												assign node1417 = (inp[5]) ? 3'b101 : 3'b001;
									assign node1421 = (inp[11]) ? node1425 : node1422;
										assign node1422 = (inp[5]) ? 3'b000 : 3'b010;
										assign node1425 = (inp[10]) ? node1427 : 3'b011;
											assign node1427 = (inp[8]) ? 3'b101 : 3'b111;
							assign node1430 = (inp[2]) ? node1456 : node1431;
								assign node1431 = (inp[4]) ? node1447 : node1432;
									assign node1432 = (inp[5]) ? node1440 : node1433;
										assign node1433 = (inp[10]) ? node1437 : node1434;
											assign node1434 = (inp[8]) ? 3'b011 : 3'b111;
											assign node1437 = (inp[8]) ? 3'b111 : 3'b011;
										assign node1440 = (inp[8]) ? node1444 : node1441;
											assign node1441 = (inp[10]) ? 3'b111 : 3'b011;
											assign node1444 = (inp[10]) ? 3'b011 : 3'b111;
									assign node1447 = (inp[10]) ? 3'b111 : node1448;
										assign node1448 = (inp[11]) ? 3'b111 : node1449;
											assign node1449 = (inp[8]) ? node1451 : 3'b011;
												assign node1451 = (inp[5]) ? 3'b011 : 3'b111;
								assign node1456 = (inp[4]) ? node1466 : node1457;
									assign node1457 = (inp[8]) ? node1463 : node1458;
										assign node1458 = (inp[10]) ? 3'b011 : node1459;
											assign node1459 = (inp[5]) ? 3'b101 : 3'b001;
										assign node1463 = (inp[10]) ? 3'b101 : 3'b001;
									assign node1466 = (inp[10]) ? node1474 : node1467;
										assign node1467 = (inp[8]) ? node1469 : 3'b011;
											assign node1469 = (inp[5]) ? node1471 : 3'b101;
												assign node1471 = (inp[11]) ? 3'b011 : 3'b101;
										assign node1474 = (inp[8]) ? node1476 : 3'b111;
											assign node1476 = (inp[11]) ? node1480 : node1477;
												assign node1477 = (inp[5]) ? 3'b011 : 3'b111;
												assign node1480 = (inp[5]) ? 3'b111 : 3'b011;
					assign node1483 = (inp[9]) ? node1605 : node1484;
						assign node1484 = (inp[4]) ? node1548 : node1485;
							assign node1485 = (inp[5]) ? node1521 : node1486;
								assign node1486 = (inp[1]) ? node1502 : node1487;
									assign node1487 = (inp[10]) ? node1495 : node1488;
										assign node1488 = (inp[2]) ? node1490 : 3'b110;
											assign node1490 = (inp[8]) ? 3'b010 : node1491;
												assign node1491 = (inp[11]) ? 3'b110 : 3'b010;
										assign node1495 = (inp[8]) ? 3'b110 : node1496;
											assign node1496 = (inp[2]) ? node1498 : 3'b000;
												assign node1498 = (inp[11]) ? 3'b000 : 3'b110;
									assign node1502 = (inp[10]) ? node1512 : node1503;
										assign node1503 = (inp[2]) ? node1507 : node1504;
											assign node1504 = (inp[8]) ? 3'b100 : 3'b010;
											assign node1507 = (inp[11]) ? node1509 : 3'b000;
												assign node1509 = (inp[8]) ? 3'b000 : 3'b100;
										assign node1512 = (inp[2]) ? node1518 : node1513;
											assign node1513 = (inp[8]) ? 3'b010 : node1514;
												assign node1514 = (inp[11]) ? 3'b110 : 3'b010;
											assign node1518 = (inp[11]) ? 3'b010 : 3'b100;
								assign node1521 = (inp[1]) ? node1537 : node1522;
									assign node1522 = (inp[8]) ? node1528 : node1523;
										assign node1523 = (inp[2]) ? 3'b000 : node1524;
											assign node1524 = (inp[10]) ? 3'b101 : 3'b001;
										assign node1528 = (inp[10]) ? 3'b000 : node1529;
											assign node1529 = (inp[2]) ? node1533 : node1530;
												assign node1530 = (inp[11]) ? 3'b000 : 3'b110;
												assign node1533 = (inp[11]) ? 3'b110 : 3'b010;
									assign node1537 = (inp[10]) ? node1545 : node1538;
										assign node1538 = (inp[2]) ? node1540 : 3'b010;
											assign node1540 = (inp[8]) ? node1542 : 3'b100;
												assign node1542 = (inp[11]) ? 3'b100 : 3'b000;
										assign node1545 = (inp[2]) ? 3'b010 : 3'b110;
							assign node1548 = (inp[1]) ? node1578 : node1549;
								assign node1549 = (inp[2]) ? node1561 : node1550;
									assign node1550 = (inp[8]) ? node1556 : node1551;
										assign node1551 = (inp[11]) ? node1553 : 3'b101;
											assign node1553 = (inp[5]) ? 3'b111 : 3'b101;
										assign node1556 = (inp[11]) ? node1558 : 3'b001;
											assign node1558 = (inp[10]) ? 3'b001 : 3'b101;
									assign node1561 = (inp[8]) ? node1569 : node1562;
										assign node1562 = (inp[10]) ? node1566 : node1563;
											assign node1563 = (inp[11]) ? 3'b101 : 3'b001;
											assign node1566 = (inp[5]) ? 3'b011 : 3'b001;
										assign node1569 = (inp[5]) ? node1575 : node1570;
											assign node1570 = (inp[10]) ? 3'b100 : node1571;
												assign node1571 = (inp[11]) ? 3'b010 : 3'b110;
											assign node1575 = (inp[10]) ? 3'b101 : 3'b001;
								assign node1578 = (inp[10]) ? node1588 : node1579;
									assign node1579 = (inp[8]) ? node1583 : node1580;
										assign node1580 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1583 = (inp[2]) ? 3'b100 : node1584;
											assign node1584 = (inp[5]) ? 3'b110 : 3'b010;
									assign node1588 = (inp[8]) ? node1600 : node1589;
										assign node1589 = (inp[2]) ? node1595 : node1590;
											assign node1590 = (inp[5]) ? 3'b000 : node1591;
												assign node1591 = (inp[11]) ? 3'b001 : 3'b011;
											assign node1595 = (inp[5]) ? 3'b101 : node1596;
												assign node1596 = (inp[11]) ? 3'b100 : 3'b000;
										assign node1600 = (inp[2]) ? 3'b010 : node1601;
											assign node1601 = (inp[11]) ? 3'b011 : 3'b010;
						assign node1605 = (inp[1]) ? node1649 : node1606;
							assign node1606 = (inp[4]) ? node1640 : node1607;
								assign node1607 = (inp[2]) ? node1621 : node1608;
									assign node1608 = (inp[8]) ? node1616 : node1609;
										assign node1609 = (inp[10]) ? node1611 : 3'b011;
											assign node1611 = (inp[5]) ? 3'b111 : node1612;
												assign node1612 = (inp[11]) ? 3'b111 : 3'b011;
										assign node1616 = (inp[10]) ? node1618 : 3'b101;
											assign node1618 = (inp[11]) ? 3'b111 : 3'b011;
									assign node1621 = (inp[10]) ? node1629 : node1622;
										assign node1622 = (inp[11]) ? 3'b101 : node1623;
											assign node1623 = (inp[8]) ? 3'b001 : node1624;
												assign node1624 = (inp[5]) ? 3'b101 : 3'b001;
										assign node1629 = (inp[8]) ? node1635 : node1630;
											assign node1630 = (inp[5]) ? 3'b011 : node1631;
												assign node1631 = (inp[11]) ? 3'b011 : 3'b101;
											assign node1635 = (inp[11]) ? 3'b101 : node1636;
												assign node1636 = (inp[5]) ? 3'b101 : 3'b001;
								assign node1640 = (inp[2]) ? node1642 : 3'b111;
									assign node1642 = (inp[10]) ? node1644 : 3'b011;
										assign node1644 = (inp[5]) ? 3'b111 : node1645;
											assign node1645 = (inp[8]) ? 3'b011 : 3'b111;
							assign node1649 = (inp[10]) ? node1681 : node1650;
								assign node1650 = (inp[4]) ? node1670 : node1651;
									assign node1651 = (inp[2]) ? node1663 : node1652;
										assign node1652 = (inp[8]) ? node1658 : node1653;
											assign node1653 = (inp[11]) ? 3'b001 : node1654;
												assign node1654 = (inp[5]) ? 3'b001 : 3'b110;
											assign node1658 = (inp[11]) ? 3'b110 : node1659;
												assign node1659 = (inp[5]) ? 3'b110 : 3'b010;
										assign node1663 = (inp[5]) ? node1665 : 3'b010;
											assign node1665 = (inp[11]) ? 3'b110 : node1666;
												assign node1666 = (inp[8]) ? 3'b010 : 3'b110;
									assign node1670 = (inp[8]) ? node1674 : node1671;
										assign node1671 = (inp[5]) ? 3'b101 : 3'b001;
										assign node1674 = (inp[2]) ? node1676 : 3'b110;
											assign node1676 = (inp[11]) ? 3'b001 : node1677;
												assign node1677 = (inp[5]) ? 3'b110 : 3'b101;
								assign node1681 = (inp[8]) ? node1699 : node1682;
									assign node1682 = (inp[4]) ? node1690 : node1683;
										assign node1683 = (inp[11]) ? node1687 : node1684;
											assign node1684 = (inp[2]) ? 3'b110 : 3'b001;
											assign node1687 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1690 = (inp[2]) ? node1694 : node1691;
											assign node1691 = (inp[5]) ? 3'b111 : 3'b011;
											assign node1694 = (inp[5]) ? node1696 : 3'b101;
												assign node1696 = (inp[11]) ? 3'b011 : 3'b101;
									assign node1699 = (inp[4]) ? node1707 : node1700;
										assign node1700 = (inp[2]) ? node1702 : 3'b001;
											assign node1702 = (inp[5]) ? 3'b001 : node1703;
												assign node1703 = (inp[11]) ? 3'b110 : 3'b010;
										assign node1707 = (inp[11]) ? node1709 : 3'b001;
											assign node1709 = (inp[2]) ? node1711 : 3'b101;
												assign node1711 = (inp[5]) ? 3'b101 : 3'b001;
			assign node1714 = (inp[1]) ? node2014 : node1715;
				assign node1715 = (inp[7]) ? node1865 : node1716;
					assign node1716 = (inp[3]) ? node1780 : node1717;
						assign node1717 = (inp[4]) ? node1749 : node1718;
							assign node1718 = (inp[2]) ? node1732 : node1719;
								assign node1719 = (inp[8]) ? node1727 : node1720;
									assign node1720 = (inp[10]) ? node1724 : node1721;
										assign node1721 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1724 = (inp[5]) ? 3'b110 : 3'b010;
									assign node1727 = (inp[5]) ? node1729 : 3'b010;
										assign node1729 = (inp[10]) ? 3'b010 : 3'b110;
								assign node1732 = (inp[8]) ? node1740 : node1733;
									assign node1733 = (inp[10]) ? node1737 : node1734;
										assign node1734 = (inp[5]) ? 3'b100 : 3'b000;
										assign node1737 = (inp[5]) ? 3'b010 : 3'b100;
									assign node1740 = (inp[10]) ? node1744 : node1741;
										assign node1741 = (inp[5]) ? 3'b000 : 3'b110;
										assign node1744 = (inp[5]) ? 3'b100 : node1745;
											assign node1745 = (inp[11]) ? 3'b100 : 3'b000;
							assign node1749 = (inp[2]) ? node1773 : node1750;
								assign node1750 = (inp[5]) ? node1758 : node1751;
									assign node1751 = (inp[8]) ? 3'b110 : node1752;
										assign node1752 = (inp[9]) ? node1754 : 3'b100;
											assign node1754 = (inp[10]) ? 3'b001 : 3'b000;
									assign node1758 = (inp[9]) ? node1766 : node1759;
										assign node1759 = (inp[10]) ? node1761 : 3'b100;
											assign node1761 = (inp[8]) ? node1763 : 3'b101;
												assign node1763 = (inp[11]) ? 3'b101 : 3'b100;
										assign node1766 = (inp[8]) ? node1768 : 3'b100;
											assign node1768 = (inp[10]) ? node1770 : 3'b000;
												assign node1770 = (inp[11]) ? 3'b001 : 3'b000;
								assign node1773 = (inp[5]) ? 3'b110 : node1774;
									assign node1774 = (inp[8]) ? node1776 : 3'b110;
										assign node1776 = (inp[9]) ? 3'b010 : 3'b110;
						assign node1780 = (inp[9]) ? node1812 : node1781;
							assign node1781 = (inp[2]) ? node1795 : node1782;
								assign node1782 = (inp[4]) ? node1788 : node1783;
									assign node1783 = (inp[10]) ? node1785 : 3'b010;
										assign node1785 = (inp[5]) ? 3'b010 : 3'b100;
									assign node1788 = (inp[10]) ? node1790 : 3'b110;
										assign node1790 = (inp[5]) ? node1792 : 3'b010;
											assign node1792 = (inp[8]) ? 3'b010 : 3'b101;
								assign node1795 = (inp[4]) ? node1797 : 3'b100;
									assign node1797 = (inp[5]) ? node1805 : node1798;
										assign node1798 = (inp[8]) ? node1802 : node1799;
											assign node1799 = (inp[10]) ? 3'b110 : 3'b010;
											assign node1802 = (inp[11]) ? 3'b100 : 3'b000;
										assign node1805 = (inp[8]) ? node1809 : node1806;
											assign node1806 = (inp[10]) ? 3'b010 : 3'b110;
											assign node1809 = (inp[10]) ? 3'b110 : 3'b010;
							assign node1812 = (inp[4]) ? node1850 : node1813;
								assign node1813 = (inp[10]) ? node1833 : node1814;
									assign node1814 = (inp[2]) ? node1824 : node1815;
										assign node1815 = (inp[8]) ? node1819 : node1816;
											assign node1816 = (inp[5]) ? 3'b011 : 3'b101;
											assign node1819 = (inp[5]) ? node1821 : 3'b000;
												assign node1821 = (inp[11]) ? 3'b101 : 3'b100;
										assign node1824 = (inp[8]) ? node1830 : node1825;
											assign node1825 = (inp[5]) ? node1827 : 3'b100;
												assign node1827 = (inp[11]) ? 3'b000 : 3'b100;
											assign node1830 = (inp[5]) ? 3'b000 : 3'b010;
									assign node1833 = (inp[11]) ? node1845 : node1834;
										assign node1834 = (inp[8]) ? node1840 : node1835;
											assign node1835 = (inp[5]) ? 3'b001 : node1836;
												assign node1836 = (inp[2]) ? 3'b100 : 3'b101;
											assign node1840 = (inp[5]) ? node1842 : 3'b000;
												assign node1842 = (inp[2]) ? 3'b100 : 3'b101;
										assign node1845 = (inp[5]) ? node1847 : 3'b001;
											assign node1847 = (inp[2]) ? 3'b001 : 3'b101;
								assign node1850 = (inp[2]) ? 3'b101 : node1851;
									assign node1851 = (inp[10]) ? node1853 : 3'b101;
										assign node1853 = (inp[11]) ? node1859 : node1854;
											assign node1854 = (inp[8]) ? 3'b101 : node1855;
												assign node1855 = (inp[5]) ? 3'b111 : 3'b101;
											assign node1859 = (inp[8]) ? node1861 : 3'b111;
												assign node1861 = (inp[5]) ? 3'b111 : 3'b101;
					assign node1865 = (inp[3]) ? node1913 : node1866;
						assign node1866 = (inp[9]) ? node1878 : node1867;
							assign node1867 = (inp[4]) ? 3'b000 : node1868;
								assign node1868 = (inp[10]) ? node1870 : 3'b000;
									assign node1870 = (inp[5]) ? node1872 : 3'b000;
										assign node1872 = (inp[2]) ? 3'b000 : node1873;
											assign node1873 = (inp[8]) ? 3'b000 : 3'b100;
							assign node1878 = (inp[4]) ? node1890 : node1879;
								assign node1879 = (inp[10]) ? node1881 : 3'b000;
									assign node1881 = (inp[2]) ? 3'b000 : node1882;
										assign node1882 = (inp[11]) ? node1884 : 3'b000;
											assign node1884 = (inp[5]) ? 3'b100 : node1885;
												assign node1885 = (inp[8]) ? 3'b000 : 3'b100;
								assign node1890 = (inp[5]) ? node1898 : node1891;
									assign node1891 = (inp[2]) ? 3'b000 : node1892;
										assign node1892 = (inp[8]) ? node1894 : 3'b100;
											assign node1894 = (inp[10]) ? 3'b100 : 3'b000;
									assign node1898 = (inp[8]) ? node1908 : node1899;
										assign node1899 = (inp[2]) ? node1903 : node1900;
											assign node1900 = (inp[10]) ? 3'b110 : 3'b100;
											assign node1903 = (inp[11]) ? 3'b010 : node1904;
												assign node1904 = (inp[10]) ? 3'b110 : 3'b010;
										assign node1908 = (inp[10]) ? node1910 : 3'b100;
											assign node1910 = (inp[2]) ? 3'b100 : 3'b010;
						assign node1913 = (inp[9]) ? node1961 : node1914;
							assign node1914 = (inp[4]) ? node1932 : node1915;
								assign node1915 = (inp[10]) ? node1917 : 3'b000;
									assign node1917 = (inp[2]) ? node1927 : node1918;
										assign node1918 = (inp[5]) ? node1924 : node1919;
											assign node1919 = (inp[8]) ? node1921 : 3'b100;
												assign node1921 = (inp[11]) ? 3'b100 : 3'b000;
											assign node1924 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1927 = (inp[8]) ? 3'b000 : node1928;
											assign node1928 = (inp[5]) ? 3'b100 : 3'b000;
								assign node1932 = (inp[10]) ? node1946 : node1933;
									assign node1933 = (inp[5]) ? node1941 : node1934;
										assign node1934 = (inp[2]) ? node1936 : 3'b100;
											assign node1936 = (inp[8]) ? 3'b000 : node1937;
												assign node1937 = (inp[11]) ? 3'b100 : 3'b000;
										assign node1941 = (inp[8]) ? 3'b100 : node1942;
											assign node1942 = (inp[11]) ? 3'b110 : 3'b010;
									assign node1946 = (inp[11]) ? node1956 : node1947;
										assign node1947 = (inp[2]) ? node1951 : node1948;
											assign node1948 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1951 = (inp[8]) ? 3'b100 : node1952;
												assign node1952 = (inp[5]) ? 3'b010 : 3'b100;
										assign node1956 = (inp[2]) ? 3'b010 : node1957;
											assign node1957 = (inp[8]) ? 3'b010 : 3'b110;
							assign node1961 = (inp[2]) ? node1989 : node1962;
								assign node1962 = (inp[8]) ? node1974 : node1963;
									assign node1963 = (inp[5]) ? node1969 : node1964;
										assign node1964 = (inp[10]) ? 3'b101 : node1965;
											assign node1965 = (inp[4]) ? 3'b001 : 3'b011;
										assign node1969 = (inp[10]) ? 3'b101 : node1970;
											assign node1970 = (inp[4]) ? 3'b001 : 3'b101;
									assign node1974 = (inp[4]) ? node1980 : node1975;
										assign node1975 = (inp[10]) ? 3'b110 : node1976;
											assign node1976 = (inp[11]) ? 3'b010 : 3'b100;
										assign node1980 = (inp[11]) ? node1984 : node1981;
											assign node1981 = (inp[10]) ? 3'b001 : 3'b110;
											assign node1984 = (inp[5]) ? node1986 : 3'b001;
												assign node1986 = (inp[10]) ? 3'b101 : 3'b001;
								assign node1989 = (inp[4]) ? node2005 : node1990;
									assign node1990 = (inp[10]) ? node1998 : node1991;
										assign node1991 = (inp[11]) ? node1993 : 3'b000;
											assign node1993 = (inp[8]) ? 3'b100 : node1994;
												assign node1994 = (inp[5]) ? 3'b000 : 3'b100;
										assign node1998 = (inp[5]) ? node2002 : node1999;
											assign node1999 = (inp[8]) ? 3'b100 : 3'b010;
											assign node2002 = (inp[8]) ? 3'b010 : 3'b110;
									assign node2005 = (inp[8]) ? node2009 : node2006;
										assign node2006 = (inp[10]) ? 3'b001 : 3'b110;
										assign node2009 = (inp[10]) ? node2011 : 3'b010;
											assign node2011 = (inp[11]) ? 3'b110 : 3'b010;
				assign node2014 = (inp[3]) ? node2056 : node2015;
					assign node2015 = (inp[2]) ? 3'b000 : node2016;
						assign node2016 = (inp[5]) ? node2036 : node2017;
							assign node2017 = (inp[8]) ? node2027 : node2018;
								assign node2018 = (inp[9]) ? 3'b000 : node2019;
									assign node2019 = (inp[7]) ? 3'b000 : node2020;
										assign node2020 = (inp[10]) ? node2022 : 3'b000;
											assign node2022 = (inp[11]) ? 3'b010 : 3'b000;
								assign node2027 = (inp[11]) ? 3'b000 : node2028;
									assign node2028 = (inp[7]) ? 3'b000 : node2029;
										assign node2029 = (inp[9]) ? node2031 : 3'b000;
											assign node2031 = (inp[4]) ? 3'b100 : 3'b000;
							assign node2036 = (inp[8]) ? node2048 : node2037;
								assign node2037 = (inp[7]) ? node2043 : node2038;
									assign node2038 = (inp[4]) ? node2040 : 3'b100;
										assign node2040 = (inp[10]) ? 3'b010 : 3'b000;
									assign node2043 = (inp[4]) ? node2045 : 3'b000;
										assign node2045 = (inp[9]) ? 3'b100 : 3'b000;
								assign node2048 = (inp[10]) ? node2050 : 3'b000;
									assign node2050 = (inp[4]) ? node2052 : 3'b000;
										assign node2052 = (inp[7]) ? 3'b000 : 3'b010;
					assign node2056 = (inp[9]) ? node2100 : node2057;
						assign node2057 = (inp[4]) ? node2067 : node2058;
							assign node2058 = (inp[7]) ? node2060 : 3'b000;
								assign node2060 = (inp[2]) ? 3'b000 : node2061;
									assign node2061 = (inp[5]) ? node2063 : 3'b000;
										assign node2063 = (inp[8]) ? 3'b000 : 3'b010;
							assign node2067 = (inp[7]) ? node2093 : node2068;
								assign node2068 = (inp[8]) ? node2080 : node2069;
									assign node2069 = (inp[5]) ? node2075 : node2070;
										assign node2070 = (inp[2]) ? 3'b000 : node2071;
											assign node2071 = (inp[10]) ? 3'b100 : 3'b010;
										assign node2075 = (inp[2]) ? node2077 : 3'b010;
											assign node2077 = (inp[10]) ? 3'b010 : 3'b100;
									assign node2080 = (inp[5]) ? node2088 : node2081;
										assign node2081 = (inp[11]) ? node2083 : 3'b000;
											assign node2083 = (inp[2]) ? node2085 : 3'b100;
												assign node2085 = (inp[10]) ? 3'b100 : 3'b000;
										assign node2088 = (inp[11]) ? node2090 : 3'b100;
											assign node2090 = (inp[10]) ? 3'b100 : 3'b000;
								assign node2093 = (inp[10]) ? node2095 : 3'b000;
									assign node2095 = (inp[11]) ? node2097 : 3'b000;
										assign node2097 = (inp[5]) ? 3'b100 : 3'b000;
						assign node2100 = (inp[7]) ? node2158 : node2101;
							assign node2101 = (inp[2]) ? node2121 : node2102;
								assign node2102 = (inp[4]) ? node2110 : node2103;
									assign node2103 = (inp[5]) ? node2107 : node2104;
										assign node2104 = (inp[8]) ? 3'b010 : 3'b110;
										assign node2107 = (inp[8]) ? 3'b110 : 3'b001;
									assign node2110 = (inp[11]) ? node2112 : 3'b001;
										assign node2112 = (inp[10]) ? node2118 : node2113;
											assign node2113 = (inp[5]) ? node2115 : 3'b101;
												assign node2115 = (inp[8]) ? 3'b101 : 3'b001;
											assign node2118 = (inp[8]) ? 3'b001 : 3'b101;
								assign node2121 = (inp[4]) ? node2147 : node2122;
									assign node2122 = (inp[8]) ? node2136 : node2123;
										assign node2123 = (inp[5]) ? node2129 : node2124;
											assign node2124 = (inp[11]) ? node2126 : 3'b100;
												assign node2126 = (inp[10]) ? 3'b010 : 3'b100;
											assign node2129 = (inp[11]) ? node2133 : node2130;
												assign node2130 = (inp[10]) ? 3'b010 : 3'b110;
												assign node2133 = (inp[10]) ? 3'b110 : 3'b010;
										assign node2136 = (inp[10]) ? node2142 : node2137;
											assign node2137 = (inp[5]) ? node2139 : 3'b010;
												assign node2139 = (inp[11]) ? 3'b100 : 3'b000;
											assign node2142 = (inp[5]) ? node2144 : 3'b100;
												assign node2144 = (inp[11]) ? 3'b010 : 3'b100;
									assign node2147 = (inp[5]) ? node2153 : node2148;
										assign node2148 = (inp[10]) ? node2150 : 3'b010;
											assign node2150 = (inp[11]) ? 3'b110 : 3'b010;
										assign node2153 = (inp[10]) ? node2155 : 3'b110;
											assign node2155 = (inp[8]) ? 3'b110 : 3'b001;
							assign node2158 = (inp[4]) ? node2176 : node2159;
								assign node2159 = (inp[5]) ? node2169 : node2160;
									assign node2160 = (inp[2]) ? 3'b000 : node2161;
										assign node2161 = (inp[10]) ? node2163 : 3'b000;
											assign node2163 = (inp[11]) ? 3'b100 : node2164;
												assign node2164 = (inp[8]) ? 3'b000 : 3'b100;
									assign node2169 = (inp[2]) ? node2173 : node2170;
										assign node2170 = (inp[8]) ? 3'b000 : 3'b010;
										assign node2173 = (inp[8]) ? 3'b000 : 3'b100;
								assign node2176 = (inp[10]) ? node2190 : node2177;
									assign node2177 = (inp[2]) ? node2183 : node2178;
										assign node2178 = (inp[5]) ? 3'b010 : node2179;
											assign node2179 = (inp[11]) ? 3'b100 : 3'b000;
										assign node2183 = (inp[8]) ? node2185 : 3'b100;
											assign node2185 = (inp[11]) ? node2187 : 3'b000;
												assign node2187 = (inp[5]) ? 3'b100 : 3'b000;
									assign node2190 = (inp[8]) ? node2196 : node2191;
										assign node2191 = (inp[2]) ? 3'b010 : node2192;
											assign node2192 = (inp[11]) ? 3'b110 : 3'b010;
										assign node2196 = (inp[11]) ? node2198 : 3'b100;
											assign node2198 = (inp[2]) ? node2202 : node2199;
												assign node2199 = (inp[5]) ? 3'b110 : 3'b010;
												assign node2202 = (inp[5]) ? 3'b010 : 3'b100;

endmodule