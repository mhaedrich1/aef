module dtc_split5_bm64 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node14;
	wire [4-1:0] node16;
	wire [4-1:0] node20;
	wire [4-1:0] node21;
	wire [4-1:0] node26;
	wire [4-1:0] node28;
	wire [4-1:0] node29;
	wire [4-1:0] node30;
	wire [4-1:0] node34;
	wire [4-1:0] node36;
	wire [4-1:0] node40;
	wire [4-1:0] node42;
	wire [4-1:0] node43;
	wire [4-1:0] node44;
	wire [4-1:0] node45;
	wire [4-1:0] node47;
	wire [4-1:0] node52;
	wire [4-1:0] node54;
	wire [4-1:0] node55;
	wire [4-1:0] node56;
	wire [4-1:0] node58;
	wire [4-1:0] node64;
	wire [4-1:0] node66;
	wire [4-1:0] node67;
	wire [4-1:0] node68;
	wire [4-1:0] node69;
	wire [4-1:0] node70;
	wire [4-1:0] node71;
	wire [4-1:0] node72;
	wire [4-1:0] node76;
	wire [4-1:0] node78;
	wire [4-1:0] node82;
	wire [4-1:0] node84;
	wire [4-1:0] node85;
	wire [4-1:0] node87;
	wire [4-1:0] node90;
	wire [4-1:0] node92;
	wire [4-1:0] node94;
	wire [4-1:0] node98;
	wire [4-1:0] node100;
	wire [4-1:0] node101;
	wire [4-1:0] node102;
	wire [4-1:0] node103;
	wire [4-1:0] node105;
	wire [4-1:0] node108;
	wire [4-1:0] node110;
	wire [4-1:0] node112;
	wire [4-1:0] node116;
	wire [4-1:0] node118;
	wire [4-1:0] node119;
	wire [4-1:0] node121;
	wire [4-1:0] node124;
	wire [4-1:0] node125;
	wire [4-1:0] node130;
	wire [4-1:0] node131;
	wire [4-1:0] node132;
	wire [4-1:0] node133;
	wire [4-1:0] node134;
	wire [4-1:0] node135;
	wire [4-1:0] node136;
	wire [4-1:0] node137;
	wire [4-1:0] node138;
	wire [4-1:0] node140;
	wire [4-1:0] node144;
	wire [4-1:0] node146;
	wire [4-1:0] node148;
	wire [4-1:0] node152;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node156;
	wire [4-1:0] node158;
	wire [4-1:0] node162;
	wire [4-1:0] node163;
	wire [4-1:0] node168;
	wire [4-1:0] node170;
	wire [4-1:0] node171;
	wire [4-1:0] node172;
	wire [4-1:0] node173;
	wire [4-1:0] node174;
	wire [4-1:0] node175;
	wire [4-1:0] node180;
	wire [4-1:0] node182;
	wire [4-1:0] node184;
	wire [4-1:0] node188;
	wire [4-1:0] node190;
	wire [4-1:0] node191;
	wire [4-1:0] node192;
	wire [4-1:0] node194;
	wire [4-1:0] node198;
	wire [4-1:0] node200;
	wire [4-1:0] node202;
	wire [4-1:0] node205;
	wire [4-1:0] node206;
	wire [4-1:0] node207;
	wire [4-1:0] node208;
	wire [4-1:0] node210;
	wire [4-1:0] node211;
	wire [4-1:0] node212;
	wire [4-1:0] node213;
	wire [4-1:0] node218;
	wire [4-1:0] node220;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node229;
	wire [4-1:0] node230;
	wire [4-1:0] node231;
	wire [4-1:0] node233;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node236;
	wire [4-1:0] node240;
	wire [4-1:0] node241;
	wire [4-1:0] node247;
	wire [4-1:0] node248;
	wire [4-1:0] node249;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node253;
	wire [4-1:0] node255;
	wire [4-1:0] node259;
	wire [4-1:0] node261;
	wire [4-1:0] node265;
	wire [4-1:0] node266;
	wire [4-1:0] node268;
	wire [4-1:0] node269;
	wire [4-1:0] node270;
	wire [4-1:0] node275;
	wire [4-1:0] node276;
	wire [4-1:0] node278;
	wire [4-1:0] node279;
	wire [4-1:0] node283;
	wire [4-1:0] node284;
	wire [4-1:0] node286;
	wire [4-1:0] node290;
	wire [4-1:0] node292;
	wire [4-1:0] node293;
	wire [4-1:0] node294;
	wire [4-1:0] node295;
	wire [4-1:0] node296;
	wire [4-1:0] node297;
	wire [4-1:0] node298;
	wire [4-1:0] node300;
	wire [4-1:0] node306;
	wire [4-1:0] node308;
	wire [4-1:0] node309;
	wire [4-1:0] node310;
	wire [4-1:0] node312;
	wire [4-1:0] node316;
	wire [4-1:0] node318;
	wire [4-1:0] node320;
	wire [4-1:0] node324;
	wire [4-1:0] node326;
	wire [4-1:0] node327;
	wire [4-1:0] node328;
	wire [4-1:0] node329;
	wire [4-1:0] node330;
	wire [4-1:0] node332;
	wire [4-1:0] node336;
	wire [4-1:0] node337;
	wire [4-1:0] node339;
	wire [4-1:0] node344;
	wire [4-1:0] node346;
	wire [4-1:0] node347;
	wire [4-1:0] node348;
	wire [4-1:0] node350;
	wire [4-1:0] node354;
	wire [4-1:0] node355;
	wire [4-1:0] node357;
	wire [4-1:0] node361;
	wire [4-1:0] node362;
	wire [4-1:0] node364;
	wire [4-1:0] node365;
	wire [4-1:0] node366;
	wire [4-1:0] node367;
	wire [4-1:0] node368;
	wire [4-1:0] node369;
	wire [4-1:0] node370;
	wire [4-1:0] node371;
	wire [4-1:0] node372;
	wire [4-1:0] node376;
	wire [4-1:0] node378;
	wire [4-1:0] node382;
	wire [4-1:0] node383;
	wire [4-1:0] node385;
	wire [4-1:0] node386;
	wire [4-1:0] node392;
	wire [4-1:0] node394;
	wire [4-1:0] node395;
	wire [4-1:0] node396;
	wire [4-1:0] node397;
	wire [4-1:0] node402;
	wire [4-1:0] node404;
	wire [4-1:0] node405;
	wire [4-1:0] node406;
	wire [4-1:0] node408;
	wire [4-1:0] node412;
	wire [4-1:0] node413;
	wire [4-1:0] node418;
	wire [4-1:0] node420;
	wire [4-1:0] node421;
	wire [4-1:0] node422;
	wire [4-1:0] node423;
	wire [4-1:0] node425;
	wire [4-1:0] node426;
	wire [4-1:0] node430;
	wire [4-1:0] node432;
	wire [4-1:0] node433;
	wire [4-1:0] node434;
	wire [4-1:0] node438;
	wire [4-1:0] node440;
	wire [4-1:0] node442;
	wire [4-1:0] node446;
	wire [4-1:0] node448;
	wire [4-1:0] node449;
	wire [4-1:0] node450;
	wire [4-1:0] node451;
	wire [4-1:0] node452;
	wire [4-1:0] node456;
	wire [4-1:0] node458;
	wire [4-1:0] node460;
	wire [4-1:0] node464;
	wire [4-1:0] node466;
	wire [4-1:0] node467;
	wire [4-1:0] node468;
	wire [4-1:0] node472;
	wire [4-1:0] node474;
	wire [4-1:0] node476;
	wire [4-1:0] node479;
	wire [4-1:0] node480;
	wire [4-1:0] node481;
	wire [4-1:0] node482;
	wire [4-1:0] node483;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node486;
	wire [4-1:0] node487;
	wire [4-1:0] node492;
	wire [4-1:0] node494;
	wire [4-1:0] node496;
	wire [4-1:0] node500;
	wire [4-1:0] node501;
	wire [4-1:0] node503;
	wire [4-1:0] node504;
	wire [4-1:0] node505;
	wire [4-1:0] node506;
	wire [4-1:0] node508;
	wire [4-1:0] node514;
	wire [4-1:0] node515;
	wire [4-1:0] node516;
	wire [4-1:0] node518;
	wire [4-1:0] node522;
	wire [4-1:0] node524;
	wire [4-1:0] node525;
	wire [4-1:0] node529;
	wire [4-1:0] node530;
	wire [4-1:0] node531;
	wire [4-1:0] node532;
	wire [4-1:0] node533;
	wire [4-1:0] node534;
	wire [4-1:0] node537;
	wire [4-1:0] node539;
	wire [4-1:0] node543;
	wire [4-1:0] node544;
	wire [4-1:0] node546;
	wire [4-1:0] node548;
	wire [4-1:0] node552;
	wire [4-1:0] node554;
	wire [4-1:0] node556;
	wire [4-1:0] node557;
	wire [4-1:0] node558;
	wire [4-1:0] node563;
	wire [4-1:0] node565;
	wire [4-1:0] node566;
	wire [4-1:0] node567;
	wire [4-1:0] node568;
	wire [4-1:0] node570;
	wire [4-1:0] node574;
	wire [4-1:0] node575;
	wire [4-1:0] node580;
	wire [4-1:0] node581;
	wire [4-1:0] node582;
	wire [4-1:0] node583;
	wire [4-1:0] node584;
	wire [4-1:0] node585;
	wire [4-1:0] node586;
	wire [4-1:0] node590;
	wire [4-1:0] node593;
	wire [4-1:0] node595;
	wire [4-1:0] node597;
	wire [4-1:0] node599;
	wire [4-1:0] node602;
	wire [4-1:0] node603;
	wire [4-1:0] node604;
	wire [4-1:0] node605;
	wire [4-1:0] node607;
	wire [4-1:0] node609;
	wire [4-1:0] node612;
	wire [4-1:0] node615;
	wire [4-1:0] node616;
	wire [4-1:0] node617;
	wire [4-1:0] node619;
	wire [4-1:0] node622;
	wire [4-1:0] node623;
	wire [4-1:0] node627;
	wire [4-1:0] node628;
	wire [4-1:0] node631;
	wire [4-1:0] node634;
	wire [4-1:0] node635;
	wire [4-1:0] node637;
	wire [4-1:0] node640;
	wire [4-1:0] node643;
	wire [4-1:0] node644;
	wire [4-1:0] node645;
	wire [4-1:0] node646;
	wire [4-1:0] node647;
	wire [4-1:0] node650;
	wire [4-1:0] node651;
	wire [4-1:0] node652;
	wire [4-1:0] node656;
	wire [4-1:0] node657;
	wire [4-1:0] node661;
	wire [4-1:0] node662;
	wire [4-1:0] node664;
	wire [4-1:0] node665;
	wire [4-1:0] node669;
	wire [4-1:0] node670;
	wire [4-1:0] node672;
	wire [4-1:0] node676;
	wire [4-1:0] node677;
	wire [4-1:0] node678;
	wire [4-1:0] node680;
	wire [4-1:0] node683;
	wire [4-1:0] node684;
	wire [4-1:0] node685;
	wire [4-1:0] node686;
	wire [4-1:0] node689;
	wire [4-1:0] node694;
	wire [4-1:0] node695;
	wire [4-1:0] node696;
	wire [4-1:0] node699;
	wire [4-1:0] node700;
	wire [4-1:0] node705;
	wire [4-1:0] node706;
	wire [4-1:0] node707;
	wire [4-1:0] node708;
	wire [4-1:0] node711;
	wire [4-1:0] node714;
	wire [4-1:0] node715;
	wire [4-1:0] node716;
	wire [4-1:0] node717;
	wire [4-1:0] node721;
	wire [4-1:0] node724;
	wire [4-1:0] node725;
	wire [4-1:0] node728;
	wire [4-1:0] node731;
	wire [4-1:0] node732;
	wire [4-1:0] node733;
	wire [4-1:0] node734;
	wire [4-1:0] node739;
	wire [4-1:0] node740;
	wire [4-1:0] node742;
	wire [4-1:0] node744;
	wire [4-1:0] node747;
	wire [4-1:0] node749;
	wire [4-1:0] node752;
	wire [4-1:0] node753;
	wire [4-1:0] node754;
	wire [4-1:0] node755;
	wire [4-1:0] node756;
	wire [4-1:0] node757;
	wire [4-1:0] node758;
	wire [4-1:0] node762;
	wire [4-1:0] node764;
	wire [4-1:0] node767;
	wire [4-1:0] node768;
	wire [4-1:0] node770;
	wire [4-1:0] node773;
	wire [4-1:0] node776;
	wire [4-1:0] node777;
	wire [4-1:0] node779;
	wire [4-1:0] node782;
	wire [4-1:0] node784;
	wire [4-1:0] node785;
	wire [4-1:0] node789;
	wire [4-1:0] node790;
	wire [4-1:0] node791;
	wire [4-1:0] node793;
	wire [4-1:0] node794;
	wire [4-1:0] node799;
	wire [4-1:0] node800;
	wire [4-1:0] node802;
	wire [4-1:0] node803;
	wire [4-1:0] node807;
	wire [4-1:0] node810;
	wire [4-1:0] node811;
	wire [4-1:0] node812;
	wire [4-1:0] node813;
	wire [4-1:0] node814;
	wire [4-1:0] node817;
	wire [4-1:0] node820;
	wire [4-1:0] node821;
	wire [4-1:0] node824;
	wire [4-1:0] node825;
	wire [4-1:0] node829;
	wire [4-1:0] node830;
	wire [4-1:0] node832;
	wire [4-1:0] node834;
	wire [4-1:0] node837;
	wire [4-1:0] node838;
	wire [4-1:0] node840;
	wire [4-1:0] node844;
	wire [4-1:0] node845;
	wire [4-1:0] node846;
	wire [4-1:0] node848;
	wire [4-1:0] node851;
	wire [4-1:0] node853;
	wire [4-1:0] node854;
	wire [4-1:0] node858;
	wire [4-1:0] node861;
	wire [4-1:0] node862;
	wire [4-1:0] node863;
	wire [4-1:0] node864;
	wire [4-1:0] node865;
	wire [4-1:0] node866;
	wire [4-1:0] node867;
	wire [4-1:0] node869;
	wire [4-1:0] node871;
	wire [4-1:0] node875;
	wire [4-1:0] node876;
	wire [4-1:0] node877;
	wire [4-1:0] node879;
	wire [4-1:0] node881;
	wire [4-1:0] node885;
	wire [4-1:0] node886;
	wire [4-1:0] node888;
	wire [4-1:0] node892;
	wire [4-1:0] node893;
	wire [4-1:0] node894;
	wire [4-1:0] node895;
	wire [4-1:0] node898;
	wire [4-1:0] node900;
	wire [4-1:0] node902;
	wire [4-1:0] node905;
	wire [4-1:0] node908;
	wire [4-1:0] node909;
	wire [4-1:0] node910;
	wire [4-1:0] node912;
	wire [4-1:0] node915;
	wire [4-1:0] node916;
	wire [4-1:0] node917;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node926;
	wire [4-1:0] node929;
	wire [4-1:0] node930;
	wire [4-1:0] node931;
	wire [4-1:0] node932;
	wire [4-1:0] node933;
	wire [4-1:0] node934;
	wire [4-1:0] node939;
	wire [4-1:0] node942;
	wire [4-1:0] node943;
	wire [4-1:0] node947;
	wire [4-1:0] node948;
	wire [4-1:0] node949;
	wire [4-1:0] node950;
	wire [4-1:0] node952;
	wire [4-1:0] node956;
	wire [4-1:0] node958;
	wire [4-1:0] node961;
	wire [4-1:0] node963;
	wire [4-1:0] node966;
	wire [4-1:0] node967;
	wire [4-1:0] node968;
	wire [4-1:0] node969;
	wire [4-1:0] node970;
	wire [4-1:0] node971;
	wire [4-1:0] node976;
	wire [4-1:0] node978;
	wire [4-1:0] node979;
	wire [4-1:0] node983;
	wire [4-1:0] node984;
	wire [4-1:0] node985;
	wire [4-1:0] node987;
	wire [4-1:0] node989;
	wire [4-1:0] node993;
	wire [4-1:0] node995;
	wire [4-1:0] node996;
	wire [4-1:0] node997;
	wire [4-1:0] node998;
	wire [4-1:0] node1004;
	wire [4-1:0] node1005;
	wire [4-1:0] node1007;
	wire [4-1:0] node1008;
	wire [4-1:0] node1010;
	wire [4-1:0] node1011;
	wire [4-1:0] node1016;
	wire [4-1:0] node1017;
	wire [4-1:0] node1018;
	wire [4-1:0] node1019;
	wire [4-1:0] node1024;
	wire [4-1:0] node1025;
	wire [4-1:0] node1027;
	wire [4-1:0] node1031;
	wire [4-1:0] node1032;
	wire [4-1:0] node1033;
	wire [4-1:0] node1034;
	wire [4-1:0] node1035;
	wire [4-1:0] node1036;
	wire [4-1:0] node1037;
	wire [4-1:0] node1038;
	wire [4-1:0] node1039;
	wire [4-1:0] node1044;
	wire [4-1:0] node1045;
	wire [4-1:0] node1049;
	wire [4-1:0] node1050;
	wire [4-1:0] node1051;
	wire [4-1:0] node1052;
	wire [4-1:0] node1057;
	wire [4-1:0] node1059;
	wire [4-1:0] node1062;
	wire [4-1:0] node1063;
	wire [4-1:0] node1064;
	wire [4-1:0] node1066;
	wire [4-1:0] node1068;
	wire [4-1:0] node1071;
	wire [4-1:0] node1073;
	wire [4-1:0] node1076;
	wire [4-1:0] node1077;
	wire [4-1:0] node1078;
	wire [4-1:0] node1082;
	wire [4-1:0] node1085;
	wire [4-1:0] node1086;
	wire [4-1:0] node1087;
	wire [4-1:0] node1089;
	wire [4-1:0] node1090;
	wire [4-1:0] node1092;
	wire [4-1:0] node1096;
	wire [4-1:0] node1098;
	wire [4-1:0] node1101;
	wire [4-1:0] node1102;
	wire [4-1:0] node1103;
	wire [4-1:0] node1104;
	wire [4-1:0] node1108;
	wire [4-1:0] node1111;
	wire [4-1:0] node1112;
	wire [4-1:0] node1113;
	wire [4-1:0] node1117;
	wire [4-1:0] node1119;
	wire [4-1:0] node1122;
	wire [4-1:0] node1123;
	wire [4-1:0] node1124;
	wire [4-1:0] node1125;
	wire [4-1:0] node1126;
	wire [4-1:0] node1128;
	wire [4-1:0] node1129;
	wire [4-1:0] node1133;
	wire [4-1:0] node1134;
	wire [4-1:0] node1135;
	wire [4-1:0] node1139;
	wire [4-1:0] node1140;
	wire [4-1:0] node1144;
	wire [4-1:0] node1145;
	wire [4-1:0] node1148;
	wire [4-1:0] node1150;
	wire [4-1:0] node1153;
	wire [4-1:0] node1156;
	wire [4-1:0] node1157;
	wire [4-1:0] node1158;
	wire [4-1:0] node1159;
	wire [4-1:0] node1160;
	wire [4-1:0] node1162;
	wire [4-1:0] node1164;
	wire [4-1:0] node1168;
	wire [4-1:0] node1170;
	wire [4-1:0] node1173;
	wire [4-1:0] node1174;
	wire [4-1:0] node1175;
	wire [4-1:0] node1179;
	wire [4-1:0] node1182;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1187;
	wire [4-1:0] node1188;
	wire [4-1:0] node1189;
	wire [4-1:0] node1190;
	wire [4-1:0] node1191;
	wire [4-1:0] node1193;
	wire [4-1:0] node1196;
	wire [4-1:0] node1199;
	wire [4-1:0] node1200;
	wire [4-1:0] node1203;
	wire [4-1:0] node1204;
	wire [4-1:0] node1205;
	wire [4-1:0] node1208;
	wire [4-1:0] node1211;
	wire [4-1:0] node1212;
	wire [4-1:0] node1216;
	wire [4-1:0] node1217;
	wire [4-1:0] node1219;
	wire [4-1:0] node1222;
	wire [4-1:0] node1223;
	wire [4-1:0] node1224;
	wire [4-1:0] node1228;
	wire [4-1:0] node1231;
	wire [4-1:0] node1232;
	wire [4-1:0] node1233;
	wire [4-1:0] node1236;
	wire [4-1:0] node1237;
	wire [4-1:0] node1240;
	wire [4-1:0] node1242;
	wire [4-1:0] node1245;
	wire [4-1:0] node1246;
	wire [4-1:0] node1247;
	wire [4-1:0] node1250;
	wire [4-1:0] node1252;
	wire [4-1:0] node1255;
	wire [4-1:0] node1256;
	wire [4-1:0] node1257;
	wire [4-1:0] node1261;
	wire [4-1:0] node1264;
	wire [4-1:0] node1265;
	wire [4-1:0] node1266;
	wire [4-1:0] node1269;
	wire [4-1:0] node1272;
	wire [4-1:0] node1273;
	wire [4-1:0] node1276;
	wire [4-1:0] node1279;
	wire [4-1:0] node1280;
	wire [4-1:0] node1281;
	wire [4-1:0] node1282;
	wire [4-1:0] node1285;
	wire [4-1:0] node1288;
	wire [4-1:0] node1289;
	wire [4-1:0] node1292;
	wire [4-1:0] node1296;
	wire [4-1:0] node1298;
	wire [4-1:0] node1299;
	wire [4-1:0] node1300;
	wire [4-1:0] node1301;
	wire [4-1:0] node1302;
	wire [4-1:0] node1303;
	wire [4-1:0] node1304;
	wire [4-1:0] node1305;
	wire [4-1:0] node1306;
	wire [4-1:0] node1308;
	wire [4-1:0] node1310;
	wire [4-1:0] node1312;
	wire [4-1:0] node1316;
	wire [4-1:0] node1318;
	wire [4-1:0] node1320;
	wire [4-1:0] node1322;
	wire [4-1:0] node1326;
	wire [4-1:0] node1328;
	wire [4-1:0] node1329;
	wire [4-1:0] node1330;
	wire [4-1:0] node1331;
	wire [4-1:0] node1332;
	wire [4-1:0] node1333;
	wire [4-1:0] node1340;
	wire [4-1:0] node1342;
	wire [4-1:0] node1344;
	wire [4-1:0] node1346;
	wire [4-1:0] node1348;
	wire [4-1:0] node1352;
	wire [4-1:0] node1353;
	wire [4-1:0] node1354;
	wire [4-1:0] node1355;
	wire [4-1:0] node1356;
	wire [4-1:0] node1357;
	wire [4-1:0] node1358;
	wire [4-1:0] node1362;
	wire [4-1:0] node1363;
	wire [4-1:0] node1365;
	wire [4-1:0] node1370;
	wire [4-1:0] node1372;
	wire [4-1:0] node1373;
	wire [4-1:0] node1374;
	wire [4-1:0] node1375;
	wire [4-1:0] node1381;
	wire [4-1:0] node1382;
	wire [4-1:0] node1384;
	wire [4-1:0] node1385;
	wire [4-1:0] node1386;
	wire [4-1:0] node1388;
	wire [4-1:0] node1392;
	wire [4-1:0] node1393;
	wire [4-1:0] node1397;
	wire [4-1:0] node1398;
	wire [4-1:0] node1400;
	wire [4-1:0] node1401;
	wire [4-1:0] node1402;
	wire [4-1:0] node1407;
	wire [4-1:0] node1408;
	wire [4-1:0] node1410;
	wire [4-1:0] node1411;
	wire [4-1:0] node1415;
	wire [4-1:0] node1416;
	wire [4-1:0] node1417;
	wire [4-1:0] node1422;
	wire [4-1:0] node1424;
	wire [4-1:0] node1425;
	wire [4-1:0] node1426;
	wire [4-1:0] node1427;
	wire [4-1:0] node1428;
	wire [4-1:0] node1432;
	wire [4-1:0] node1434;
	wire [4-1:0] node1435;
	wire [4-1:0] node1440;
	wire [4-1:0] node1442;
	wire [4-1:0] node1443;
	wire [4-1:0] node1444;
	wire [4-1:0] node1445;
	wire [4-1:0] node1446;
	wire [4-1:0] node1452;
	wire [4-1:0] node1454;
	wire [4-1:0] node1457;
	wire [4-1:0] node1458;
	wire [4-1:0] node1460;
	wire [4-1:0] node1461;
	wire [4-1:0] node1462;
	wire [4-1:0] node1463;
	wire [4-1:0] node1464;
	wire [4-1:0] node1465;
	wire [4-1:0] node1466;
	wire [4-1:0] node1468;
	wire [4-1:0] node1472;
	wire [4-1:0] node1474;
	wire [4-1:0] node1475;
	wire [4-1:0] node1480;
	wire [4-1:0] node1482;
	wire [4-1:0] node1484;
	wire [4-1:0] node1486;
	wire [4-1:0] node1487;
	wire [4-1:0] node1492;
	wire [4-1:0] node1494;
	wire [4-1:0] node1495;
	wire [4-1:0] node1496;
	wire [4-1:0] node1497;
	wire [4-1:0] node1500;
	wire [4-1:0] node1501;
	wire [4-1:0] node1506;
	wire [4-1:0] node1508;
	wire [4-1:0] node1509;
	wire [4-1:0] node1510;
	wire [4-1:0] node1515;
	wire [4-1:0] node1516;
	wire [4-1:0] node1517;
	wire [4-1:0] node1518;
	wire [4-1:0] node1519;
	wire [4-1:0] node1520;
	wire [4-1:0] node1521;
	wire [4-1:0] node1525;
	wire [4-1:0] node1526;
	wire [4-1:0] node1527;
	wire [4-1:0] node1531;
	wire [4-1:0] node1534;
	wire [4-1:0] node1535;
	wire [4-1:0] node1538;
	wire [4-1:0] node1540;
	wire [4-1:0] node1541;
	wire [4-1:0] node1545;
	wire [4-1:0] node1546;
	wire [4-1:0] node1547;
	wire [4-1:0] node1549;
	wire [4-1:0] node1552;
	wire [4-1:0] node1553;
	wire [4-1:0] node1556;
	wire [4-1:0] node1558;
	wire [4-1:0] node1561;
	wire [4-1:0] node1562;
	wire [4-1:0] node1564;
	wire [4-1:0] node1568;
	wire [4-1:0] node1569;
	wire [4-1:0] node1570;
	wire [4-1:0] node1571;
	wire [4-1:0] node1573;
	wire [4-1:0] node1575;
	wire [4-1:0] node1579;
	wire [4-1:0] node1581;
	wire [4-1:0] node1582;
	wire [4-1:0] node1583;
	wire [4-1:0] node1584;
	wire [4-1:0] node1590;
	wire [4-1:0] node1591;
	wire [4-1:0] node1592;
	wire [4-1:0] node1594;
	wire [4-1:0] node1595;
	wire [4-1:0] node1597;
	wire [4-1:0] node1601;
	wire [4-1:0] node1602;
	wire [4-1:0] node1603;
	wire [4-1:0] node1606;
	wire [4-1:0] node1609;
	wire [4-1:0] node1610;
	wire [4-1:0] node1613;
	wire [4-1:0] node1614;
	wire [4-1:0] node1618;
	wire [4-1:0] node1619;
	wire [4-1:0] node1620;
	wire [4-1:0] node1621;
	wire [4-1:0] node1623;
	wire [4-1:0] node1628;
	wire [4-1:0] node1629;
	wire [4-1:0] node1633;
	wire [4-1:0] node1634;
	wire [4-1:0] node1635;
	wire [4-1:0] node1636;
	wire [4-1:0] node1637;
	wire [4-1:0] node1638;
	wire [4-1:0] node1640;
	wire [4-1:0] node1641;
	wire [4-1:0] node1644;
	wire [4-1:0] node1647;
	wire [4-1:0] node1648;
	wire [4-1:0] node1651;
	wire [4-1:0] node1653;
	wire [4-1:0] node1656;
	wire [4-1:0] node1658;
	wire [4-1:0] node1661;
	wire [4-1:0] node1662;
	wire [4-1:0] node1663;
	wire [4-1:0] node1664;
	wire [4-1:0] node1665;
	wire [4-1:0] node1670;
	wire [4-1:0] node1672;
	wire [4-1:0] node1675;
	wire [4-1:0] node1676;
	wire [4-1:0] node1677;
	wire [4-1:0] node1681;
	wire [4-1:0] node1684;
	wire [4-1:0] node1685;
	wire [4-1:0] node1686;
	wire [4-1:0] node1688;
	wire [4-1:0] node1692;
	wire [4-1:0] node1693;
	wire [4-1:0] node1694;
	wire [4-1:0] node1698;
	wire [4-1:0] node1700;
	wire [4-1:0] node1703;
	wire [4-1:0] node1704;
	wire [4-1:0] node1705;
	wire [4-1:0] node1706;
	wire [4-1:0] node1707;
	wire [4-1:0] node1708;
	wire [4-1:0] node1709;
	wire [4-1:0] node1714;
	wire [4-1:0] node1716;
	wire [4-1:0] node1717;
	wire [4-1:0] node1721;
	wire [4-1:0] node1722;
	wire [4-1:0] node1724;
	wire [4-1:0] node1726;
	wire [4-1:0] node1727;
	wire [4-1:0] node1730;
	wire [4-1:0] node1733;
	wire [4-1:0] node1736;
	wire [4-1:0] node1737;
	wire [4-1:0] node1738;
	wire [4-1:0] node1740;
	wire [4-1:0] node1741;
	wire [4-1:0] node1745;
	wire [4-1:0] node1746;
	wire [4-1:0] node1747;
	wire [4-1:0] node1752;
	wire [4-1:0] node1755;
	wire [4-1:0] node1756;
	wire [4-1:0] node1757;
	wire [4-1:0] node1758;
	wire [4-1:0] node1761;
	wire [4-1:0] node1764;
	wire [4-1:0] node1765;
	wire [4-1:0] node1768;
	wire [4-1:0] node1772;
	wire [4-1:0] node1774;
	wire [4-1:0] node1775;
	wire [4-1:0] node1776;
	wire [4-1:0] node1777;
	wire [4-1:0] node1778;
	wire [4-1:0] node1779;
	wire [4-1:0] node1780;
	wire [4-1:0] node1781;
	wire [4-1:0] node1783;
	wire [4-1:0] node1786;
	wire [4-1:0] node1788;
	wire [4-1:0] node1790;
	wire [4-1:0] node1794;
	wire [4-1:0] node1796;
	wire [4-1:0] node1797;
	wire [4-1:0] node1798;
	wire [4-1:0] node1802;
	wire [4-1:0] node1803;
	wire [4-1:0] node1805;
	wire [4-1:0] node1810;
	wire [4-1:0] node1811;
	wire [4-1:0] node1812;
	wire [4-1:0] node1814;
	wire [4-1:0] node1815;
	wire [4-1:0] node1816;
	wire [4-1:0] node1821;
	wire [4-1:0] node1822;
	wire [4-1:0] node1824;
	wire [4-1:0] node1825;
	wire [4-1:0] node1829;
	wire [4-1:0] node1831;
	wire [4-1:0] node1832;
	wire [4-1:0] node1833;
	wire [4-1:0] node1838;
	wire [4-1:0] node1840;
	wire [4-1:0] node1841;
	wire [4-1:0] node1842;
	wire [4-1:0] node1844;
	wire [4-1:0] node1848;
	wire [4-1:0] node1849;
	wire [4-1:0] node1851;
	wire [4-1:0] node1855;
	wire [4-1:0] node1856;
	wire [4-1:0] node1858;
	wire [4-1:0] node1859;
	wire [4-1:0] node1860;
	wire [4-1:0] node1861;
	wire [4-1:0] node1863;
	wire [4-1:0] node1866;
	wire [4-1:0] node1868;
	wire [4-1:0] node1872;
	wire [4-1:0] node1873;
	wire [4-1:0] node1875;
	wire [4-1:0] node1879;
	wire [4-1:0] node1880;
	wire [4-1:0] node1881;
	wire [4-1:0] node1882;
	wire [4-1:0] node1883;
	wire [4-1:0] node1886;
	wire [4-1:0] node1887;
	wire [4-1:0] node1891;
	wire [4-1:0] node1892;
	wire [4-1:0] node1893;
	wire [4-1:0] node1897;
	wire [4-1:0] node1899;
	wire [4-1:0] node1902;
	wire [4-1:0] node1903;
	wire [4-1:0] node1906;
	wire [4-1:0] node1907;
	wire [4-1:0] node1911;
	wire [4-1:0] node1912;
	wire [4-1:0] node1913;
	wire [4-1:0] node1914;
	wire [4-1:0] node1916;
	wire [4-1:0] node1919;
	wire [4-1:0] node1921;
	wire [4-1:0] node1923;
	wire [4-1:0] node1926;
	wire [4-1:0] node1927;
	wire [4-1:0] node1930;
	wire [4-1:0] node1933;
	wire [4-1:0] node1934;
	wire [4-1:0] node1935;
	wire [4-1:0] node1938;
	wire [4-1:0] node1942;
	wire [4-1:0] node1944;
	wire [4-1:0] node1945;
	wire [4-1:0] node1946;
	wire [4-1:0] node1947;
	wire [4-1:0] node1948;
	wire [4-1:0] node1949;
	wire [4-1:0] node1951;
	wire [4-1:0] node1952;
	wire [4-1:0] node1956;
	wire [4-1:0] node1957;
	wire [4-1:0] node1959;
	wire [4-1:0] node1963;
	wire [4-1:0] node1964;
	wire [4-1:0] node1966;
	wire [4-1:0] node1967;
	wire [4-1:0] node1971;
	wire [4-1:0] node1974;
	wire [4-1:0] node1975;
	wire [4-1:0] node1976;
	wire [4-1:0] node1977;
	wire [4-1:0] node1978;
	wire [4-1:0] node1984;
	wire [4-1:0] node1985;
	wire [4-1:0] node1986;
	wire [4-1:0] node1989;
	wire [4-1:0] node1992;
	wire [4-1:0] node1993;
	wire [4-1:0] node1997;
	wire [4-1:0] node1998;
	wire [4-1:0] node1999;
	wire [4-1:0] node2000;
	wire [4-1:0] node2001;
	wire [4-1:0] node2003;
	wire [4-1:0] node2008;
	wire [4-1:0] node2009;
	wire [4-1:0] node2012;
	wire [4-1:0] node2013;
	wire [4-1:0] node2014;
	wire [4-1:0] node2018;
	wire [4-1:0] node2021;
	wire [4-1:0] node2022;
	wire [4-1:0] node2023;
	wire [4-1:0] node2024;
	wire [4-1:0] node2029;
	wire [4-1:0] node2030;
	wire [4-1:0] node2031;
	wire [4-1:0] node2034;
	wire [4-1:0] node2037;
	wire [4-1:0] node2038;
	wire [4-1:0] node2039;
	wire [4-1:0] node2043;
	wire [4-1:0] node2044;
	wire [4-1:0] node2048;
	wire [4-1:0] node2050;
	wire [4-1:0] node2051;
	wire [4-1:0] node2052;
	wire [4-1:0] node2053;
	wire [4-1:0] node2055;
	wire [4-1:0] node2057;
	wire [4-1:0] node2060;
	wire [4-1:0] node2061;
	wire [4-1:0] node2063;
	wire [4-1:0] node2066;
	wire [4-1:0] node2068;
	wire [4-1:0] node2071;
	wire [4-1:0] node2072;
	wire [4-1:0] node2074;
	wire [4-1:0] node2075;
	wire [4-1:0] node2078;
	wire [4-1:0] node2081;
	wire [4-1:0] node2082;
	wire [4-1:0] node2084;
	wire [4-1:0] node2087;
	wire [4-1:0] node2088;
	wire [4-1:0] node2092;
	wire [4-1:0] node2094;
	wire [4-1:0] node2095;
	wire [4-1:0] node2096;
	wire [4-1:0] node2098;
	wire [4-1:0] node2101;
	wire [4-1:0] node2102;
	wire [4-1:0] node2106;
	wire [4-1:0] node2107;

	assign outp = (inp[14]) ? node2 : 4'b0000;
		assign node2 = (inp[12]) ? node1296 : node3;
			assign node3 = (inp[3]) ? node361 : node4;
				assign node4 = (inp[0]) ? node130 : node5;
					assign node5 = (inp[4]) ? 4'b0000 : node6;
						assign node6 = (inp[11]) ? node64 : node7;
							assign node7 = (inp[7]) ? 4'b0010 : node8;
								assign node8 = (inp[9]) ? node40 : node9;
									assign node9 = (inp[5]) ? 4'b0000 : node10;
										assign node10 = (inp[15]) ? node26 : node11;
											assign node11 = (inp[13]) ? 4'b0010 : node12;
												assign node12 = (inp[1]) ? node20 : node13;
													assign node13 = (inp[8]) ? 4'b0000 : node14;
														assign node14 = (inp[10]) ? node16 : 4'b0010;
															assign node16 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node20 = (inp[6]) ? 4'b0010 : node21;
														assign node21 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node26 = (inp[13]) ? node28 : 4'b0000;
												assign node28 = (inp[1]) ? node34 : node29;
													assign node29 = (inp[8]) ? 4'b0000 : node30;
														assign node30 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node34 = (inp[8]) ? node36 : 4'b0010;
														assign node36 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node40 = (inp[5]) ? node42 : 4'b0010;
										assign node42 = (inp[13]) ? node52 : node43;
											assign node43 = (inp[15]) ? 4'b0000 : node44;
												assign node44 = (inp[1]) ? 4'b0010 : node45;
													assign node45 = (inp[6]) ? node47 : 4'b0000;
														assign node47 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node52 = (inp[15]) ? node54 : 4'b0010;
												assign node54 = (inp[1]) ? 4'b0010 : node55;
													assign node55 = (inp[8]) ? 4'b0000 : node56;
														assign node56 = (inp[10]) ? node58 : 4'b0010;
															assign node58 = (inp[6]) ? 4'b0010 : 4'b0000;
							assign node64 = (inp[7]) ? node66 : 4'b0000;
								assign node66 = (inp[5]) ? node98 : node67;
									assign node67 = (inp[9]) ? 4'b0010 : node68;
										assign node68 = (inp[13]) ? node82 : node69;
											assign node69 = (inp[15]) ? 4'b0000 : node70;
												assign node70 = (inp[8]) ? node76 : node71;
													assign node71 = (inp[1]) ? 4'b0010 : node72;
														assign node72 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node76 = (inp[1]) ? node78 : 4'b0000;
														assign node78 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node82 = (inp[15]) ? node84 : 4'b0010;
												assign node84 = (inp[8]) ? node90 : node85;
													assign node85 = (inp[10]) ? node87 : 4'b0010;
														assign node87 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node90 = (inp[1]) ? node92 : 4'b0000;
														assign node92 = (inp[10]) ? node94 : 4'b0010;
															assign node94 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node98 = (inp[9]) ? node100 : 4'b0000;
										assign node100 = (inp[13]) ? node116 : node101;
											assign node101 = (inp[15]) ? 4'b0000 : node102;
												assign node102 = (inp[10]) ? node108 : node103;
													assign node103 = (inp[8]) ? node105 : 4'b0010;
														assign node105 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node108 = (inp[1]) ? node110 : 4'b0000;
														assign node110 = (inp[8]) ? node112 : 4'b0010;
															assign node112 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node116 = (inp[15]) ? node118 : 4'b0010;
												assign node118 = (inp[1]) ? node124 : node119;
													assign node119 = (inp[2]) ? node121 : 4'b0000;
														assign node121 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node124 = (inp[6]) ? 4'b0010 : node125;
														assign node125 = (inp[2]) ? 4'b0000 : 4'b0010;
					assign node130 = (inp[4]) ? node290 : node131;
						assign node131 = (inp[7]) ? node205 : node132;
							assign node132 = (inp[9]) ? node168 : node133;
								assign node133 = (inp[11]) ? 4'b0010 : node134;
									assign node134 = (inp[13]) ? node152 : node135;
										assign node135 = (inp[5]) ? 4'b0010 : node136;
											assign node136 = (inp[15]) ? node144 : node137;
												assign node137 = (inp[1]) ? 4'b0000 : node138;
													assign node138 = (inp[8]) ? node140 : 4'b0000;
														assign node140 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node144 = (inp[1]) ? node146 : 4'b0010;
													assign node146 = (inp[8]) ? node148 : 4'b0000;
														assign node148 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node152 = (inp[5]) ? node154 : 4'b0000;
											assign node154 = (inp[1]) ? node162 : node155;
												assign node155 = (inp[15]) ? 4'b0010 : node156;
													assign node156 = (inp[8]) ? node158 : 4'b0000;
														assign node158 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node162 = (inp[6]) ? 4'b0000 : node163;
													assign node163 = (inp[15]) ? 4'b0010 : 4'b0000;
								assign node168 = (inp[11]) ? node170 : 4'b0000;
									assign node170 = (inp[13]) ? node188 : node171;
										assign node171 = (inp[5]) ? 4'b0010 : node172;
											assign node172 = (inp[15]) ? node180 : node173;
												assign node173 = (inp[6]) ? 4'b0000 : node174;
													assign node174 = (inp[1]) ? 4'b0000 : node175;
														assign node175 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node180 = (inp[1]) ? node182 : 4'b0010;
													assign node182 = (inp[8]) ? node184 : 4'b0000;
														assign node184 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node188 = (inp[5]) ? node190 : 4'b0000;
											assign node190 = (inp[15]) ? node198 : node191;
												assign node191 = (inp[6]) ? 4'b0000 : node192;
													assign node192 = (inp[8]) ? node194 : 4'b0000;
														assign node194 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node198 = (inp[1]) ? node200 : 4'b0010;
													assign node200 = (inp[8]) ? node202 : 4'b0000;
														assign node202 = (inp[10]) ? 4'b0010 : 4'b0000;
							assign node205 = (inp[9]) ? node229 : node206;
								assign node206 = (inp[5]) ? 4'b0000 : node207;
									assign node207 = (inp[11]) ? 4'b0000 : node208;
										assign node208 = (inp[13]) ? node210 : 4'b0000;
											assign node210 = (inp[1]) ? node218 : node211;
												assign node211 = (inp[8]) ? 4'b0000 : node212;
													assign node212 = (inp[15]) ? 4'b0000 : node213;
														assign node213 = (inp[2]) ? 4'b0000 : 4'b0010;
												assign node218 = (inp[15]) ? node220 : 4'b0010;
													assign node220 = (inp[6]) ? 4'b0010 : node221;
														assign node221 = (inp[8]) ? 4'b0000 : node222;
															assign node222 = (inp[2]) ? 4'b0010 : 4'b0000;
								assign node229 = (inp[11]) ? node247 : node230;
									assign node230 = (inp[1]) ? 4'b0010 : node231;
										assign node231 = (inp[5]) ? node233 : 4'b0010;
											assign node233 = (inp[13]) ? 4'b0010 : node234;
												assign node234 = (inp[15]) ? node240 : node235;
													assign node235 = (inp[2]) ? 4'b0010 : node236;
														assign node236 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node240 = (inp[8]) ? 4'b0000 : node241;
														assign node241 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node247 = (inp[13]) ? node265 : node248;
										assign node248 = (inp[5]) ? 4'b0000 : node249;
											assign node249 = (inp[1]) ? node251 : 4'b0000;
												assign node251 = (inp[10]) ? node259 : node252;
													assign node252 = (inp[15]) ? 4'b0000 : node253;
														assign node253 = (inp[2]) ? node255 : 4'b0010;
															assign node255 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node259 = (inp[6]) ? node261 : 4'b0000;
														assign node261 = (inp[15]) ? 4'b0000 : 4'b0010;
										assign node265 = (inp[5]) ? node275 : node266;
											assign node266 = (inp[8]) ? node268 : 4'b0010;
												assign node268 = (inp[1]) ? 4'b0010 : node269;
													assign node269 = (inp[6]) ? 4'b0010 : node270;
														assign node270 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node275 = (inp[1]) ? node283 : node276;
												assign node276 = (inp[10]) ? node278 : 4'b0000;
													assign node278 = (inp[8]) ? 4'b0000 : node279;
														assign node279 = (inp[6]) ? 4'b0010 : 4'b0000;
												assign node283 = (inp[6]) ? 4'b0010 : node284;
													assign node284 = (inp[15]) ? node286 : 4'b0010;
														assign node286 = (inp[8]) ? 4'b0000 : 4'b0010;
						assign node290 = (inp[7]) ? node292 : 4'b0010;
							assign node292 = (inp[11]) ? node324 : node293;
								assign node293 = (inp[9]) ? 4'b0000 : node294;
									assign node294 = (inp[13]) ? node306 : node295;
										assign node295 = (inp[5]) ? 4'b0010 : node296;
											assign node296 = (inp[1]) ? 4'b0000 : node297;
												assign node297 = (inp[15]) ? 4'b0010 : node298;
													assign node298 = (inp[8]) ? node300 : 4'b0000;
														assign node300 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node306 = (inp[5]) ? node308 : 4'b0000;
											assign node308 = (inp[15]) ? node316 : node309;
												assign node309 = (inp[1]) ? 4'b0000 : node310;
													assign node310 = (inp[8]) ? node312 : 4'b0000;
														assign node312 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node316 = (inp[1]) ? node318 : 4'b0010;
													assign node318 = (inp[8]) ? node320 : 4'b0000;
														assign node320 = (inp[6]) ? 4'b0000 : 4'b0010;
								assign node324 = (inp[9]) ? node326 : 4'b0010;
									assign node326 = (inp[13]) ? node344 : node327;
										assign node327 = (inp[5]) ? 4'b0010 : node328;
											assign node328 = (inp[1]) ? node336 : node329;
												assign node329 = (inp[15]) ? 4'b0010 : node330;
													assign node330 = (inp[8]) ? node332 : 4'b0000;
														assign node332 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node336 = (inp[6]) ? 4'b0000 : node337;
													assign node337 = (inp[15]) ? node339 : 4'b0000;
														assign node339 = (inp[10]) ? 4'b0000 : 4'b0010;
										assign node344 = (inp[5]) ? node346 : 4'b0000;
											assign node346 = (inp[1]) ? node354 : node347;
												assign node347 = (inp[15]) ? 4'b0010 : node348;
													assign node348 = (inp[8]) ? node350 : 4'b0000;
														assign node350 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node354 = (inp[6]) ? 4'b0000 : node355;
													assign node355 = (inp[15]) ? node357 : 4'b0000;
														assign node357 = (inp[8]) ? 4'b0010 : 4'b0000;
				assign node361 = (inp[0]) ? node479 : node362;
					assign node362 = (inp[4]) ? node364 : 4'b0010;
						assign node364 = (inp[7]) ? node418 : node365;
							assign node365 = (inp[11]) ? 4'b0000 : node366;
								assign node366 = (inp[9]) ? node392 : node367;
									assign node367 = (inp[5]) ? 4'b0000 : node368;
										assign node368 = (inp[13]) ? node382 : node369;
											assign node369 = (inp[15]) ? 4'b0000 : node370;
												assign node370 = (inp[8]) ? node376 : node371;
													assign node371 = (inp[6]) ? 4'b0010 : node372;
														assign node372 = (inp[2]) ? 4'b0010 : 4'b0000;
													assign node376 = (inp[1]) ? node378 : 4'b0000;
														assign node378 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node382 = (inp[1]) ? 4'b0010 : node383;
												assign node383 = (inp[15]) ? node385 : 4'b0010;
													assign node385 = (inp[8]) ? 4'b0000 : node386;
														assign node386 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node392 = (inp[5]) ? node394 : 4'b0010;
										assign node394 = (inp[15]) ? node402 : node395;
											assign node395 = (inp[1]) ? 4'b0010 : node396;
												assign node396 = (inp[13]) ? 4'b0010 : node397;
													assign node397 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node402 = (inp[13]) ? node404 : 4'b0000;
												assign node404 = (inp[6]) ? node412 : node405;
													assign node405 = (inp[10]) ? 4'b0000 : node406;
														assign node406 = (inp[8]) ? node408 : 4'b0010;
															assign node408 = (inp[2]) ? 4'b0010 : 4'b0000;
													assign node412 = (inp[10]) ? 4'b0010 : node413;
														assign node413 = (inp[1]) ? 4'b0010 : 4'b0000;
							assign node418 = (inp[11]) ? node420 : 4'b0010;
								assign node420 = (inp[5]) ? node446 : node421;
									assign node421 = (inp[9]) ? 4'b0010 : node422;
										assign node422 = (inp[15]) ? node430 : node423;
											assign node423 = (inp[8]) ? node425 : 4'b0010;
												assign node425 = (inp[13]) ? 4'b0010 : node426;
													assign node426 = (inp[1]) ? 4'b0010 : 4'b0000;
											assign node430 = (inp[13]) ? node432 : 4'b0000;
												assign node432 = (inp[1]) ? node438 : node433;
													assign node433 = (inp[8]) ? 4'b0000 : node434;
														assign node434 = (inp[2]) ? 4'b0000 : 4'b0010;
													assign node438 = (inp[8]) ? node440 : 4'b0010;
														assign node440 = (inp[10]) ? node442 : 4'b0010;
															assign node442 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node446 = (inp[9]) ? node448 : 4'b0000;
										assign node448 = (inp[15]) ? node464 : node449;
											assign node449 = (inp[13]) ? 4'b0010 : node450;
												assign node450 = (inp[1]) ? node456 : node451;
													assign node451 = (inp[8]) ? 4'b0000 : node452;
														assign node452 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node456 = (inp[8]) ? node458 : 4'b0010;
														assign node458 = (inp[10]) ? node460 : 4'b0010;
															assign node460 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node464 = (inp[13]) ? node466 : 4'b0000;
												assign node466 = (inp[8]) ? node472 : node467;
													assign node467 = (inp[2]) ? 4'b0010 : node468;
														assign node468 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node472 = (inp[1]) ? node474 : 4'b0000;
														assign node474 = (inp[10]) ? node476 : 4'b0010;
															assign node476 = (inp[6]) ? 4'b0010 : 4'b0000;
					assign node479 = (inp[9]) ? node861 : node480;
						assign node480 = (inp[7]) ? node580 : node481;
							assign node481 = (inp[4]) ? node529 : node482;
								assign node482 = (inp[13]) ? node500 : node483;
									assign node483 = (inp[11]) ? 4'b0010 : node484;
										assign node484 = (inp[1]) ? node492 : node485;
											assign node485 = (inp[5]) ? 4'b0010 : node486;
												assign node486 = (inp[6]) ? 4'b1000 : node487;
													assign node487 = (inp[15]) ? 4'b0010 : 4'b1000;
											assign node492 = (inp[5]) ? node494 : 4'b1000;
												assign node494 = (inp[15]) ? node496 : 4'b1000;
													assign node496 = (inp[6]) ? 4'b1000 : 4'b0010;
									assign node500 = (inp[11]) ? node514 : node501;
										assign node501 = (inp[1]) ? node503 : 4'b1000;
											assign node503 = (inp[5]) ? 4'b1000 : node504;
												assign node504 = (inp[6]) ? 4'b1010 : node505;
													assign node505 = (inp[15]) ? 4'b1000 : node506;
														assign node506 = (inp[8]) ? node508 : 4'b1010;
															assign node508 = (inp[2]) ? 4'b1000 : 4'b1010;
										assign node514 = (inp[1]) ? node522 : node515;
											assign node515 = (inp[5]) ? 4'b0010 : node516;
												assign node516 = (inp[15]) ? node518 : 4'b1000;
													assign node518 = (inp[6]) ? 4'b1000 : 4'b0010;
											assign node522 = (inp[5]) ? node524 : 4'b1000;
												assign node524 = (inp[6]) ? 4'b1000 : node525;
													assign node525 = (inp[15]) ? 4'b0010 : 4'b1000;
								assign node529 = (inp[11]) ? node563 : node530;
									assign node530 = (inp[13]) ? node552 : node531;
										assign node531 = (inp[5]) ? node543 : node532;
											assign node532 = (inp[1]) ? 4'b0010 : node533;
												assign node533 = (inp[15]) ? node537 : node534;
													assign node534 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node537 = (inp[6]) ? node539 : 4'b0000;
														assign node539 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node543 = (inp[15]) ? 4'b0000 : node544;
												assign node544 = (inp[1]) ? node546 : 4'b0000;
													assign node546 = (inp[8]) ? node548 : 4'b0010;
														assign node548 = (inp[6]) ? 4'b0010 : 4'b0000;
										assign node552 = (inp[5]) ? node554 : 4'b0010;
											assign node554 = (inp[15]) ? node556 : 4'b0010;
												assign node556 = (inp[6]) ? 4'b0010 : node557;
													assign node557 = (inp[2]) ? 4'b0010 : node558;
														assign node558 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node563 = (inp[13]) ? node565 : 4'b0000;
										assign node565 = (inp[5]) ? 4'b0000 : node566;
											assign node566 = (inp[1]) ? node574 : node567;
												assign node567 = (inp[15]) ? 4'b0000 : node568;
													assign node568 = (inp[6]) ? node570 : 4'b0000;
														assign node570 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node574 = (inp[6]) ? 4'b0010 : node575;
													assign node575 = (inp[10]) ? 4'b0000 : 4'b0010;
							assign node580 = (inp[13]) ? node752 : node581;
								assign node581 = (inp[4]) ? node643 : node582;
									assign node582 = (inp[1]) ? node602 : node583;
										assign node583 = (inp[11]) ? node593 : node584;
											assign node584 = (inp[5]) ? node590 : node585;
												assign node585 = (inp[15]) ? 4'b0000 : node586;
													assign node586 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node590 = (inp[6]) ? 4'b0000 : 4'b1010;
											assign node593 = (inp[5]) ? node595 : 4'b1010;
												assign node595 = (inp[6]) ? node597 : 4'b1000;
													assign node597 = (inp[8]) ? node599 : 4'b1010;
														assign node599 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node602 = (inp[11]) ? node634 : node603;
											assign node603 = (inp[15]) ? node615 : node604;
												assign node604 = (inp[6]) ? node612 : node605;
													assign node605 = (inp[5]) ? node607 : 4'b0010;
														assign node607 = (inp[8]) ? node609 : 4'b0010;
															assign node609 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node612 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node615 = (inp[10]) ? node627 : node616;
													assign node616 = (inp[8]) ? node622 : node617;
														assign node617 = (inp[6]) ? node619 : 4'b0000;
															assign node619 = (inp[2]) ? 4'b0000 : 4'b0010;
														assign node622 = (inp[6]) ? 4'b0000 : node623;
															assign node623 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node627 = (inp[5]) ? node631 : node628;
														assign node628 = (inp[6]) ? 4'b0000 : 4'b0010;
														assign node631 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node634 = (inp[5]) ? node640 : node635;
												assign node635 = (inp[6]) ? node637 : 4'b0000;
													assign node637 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node640 = (inp[6]) ? 4'b0000 : 4'b1010;
									assign node643 = (inp[10]) ? node705 : node644;
										assign node644 = (inp[8]) ? node676 : node645;
											assign node645 = (inp[1]) ? node661 : node646;
												assign node646 = (inp[5]) ? node650 : node647;
													assign node647 = (inp[11]) ? 4'b1010 : 4'b1000;
													assign node650 = (inp[11]) ? node656 : node651;
														assign node651 = (inp[15]) ? 4'b1010 : node652;
															assign node652 = (inp[6]) ? 4'b1000 : 4'b1010;
														assign node656 = (inp[2]) ? 4'b1000 : node657;
															assign node657 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node661 = (inp[11]) ? node669 : node662;
													assign node662 = (inp[5]) ? node664 : 4'b1010;
														assign node664 = (inp[15]) ? 4'b1000 : node665;
															assign node665 = (inp[6]) ? 4'b1010 : 4'b1000;
													assign node669 = (inp[5]) ? 4'b1010 : node670;
														assign node670 = (inp[15]) ? node672 : 4'b1000;
															assign node672 = (inp[6]) ? 4'b1000 : 4'b1010;
											assign node676 = (inp[6]) ? node694 : node677;
												assign node677 = (inp[5]) ? node683 : node678;
													assign node678 = (inp[2]) ? node680 : 4'b1010;
														assign node680 = (inp[1]) ? 4'b1000 : 4'b1010;
													assign node683 = (inp[2]) ? 4'b1010 : node684;
														assign node684 = (inp[15]) ? 4'b1000 : node685;
															assign node685 = (inp[11]) ? node689 : node686;
																assign node686 = (inp[1]) ? 4'b1000 : 4'b1010;
																assign node689 = (inp[1]) ? 4'b1010 : 4'b1000;
												assign node694 = (inp[15]) ? 4'b1010 : node695;
													assign node695 = (inp[1]) ? node699 : node696;
														assign node696 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node699 = (inp[5]) ? 4'b1010 : node700;
															assign node700 = (inp[11]) ? 4'b1000 : 4'b1010;
										assign node705 = (inp[5]) ? node731 : node706;
											assign node706 = (inp[15]) ? node714 : node707;
												assign node707 = (inp[1]) ? node711 : node708;
													assign node708 = (inp[11]) ? 4'b1010 : 4'b1000;
													assign node711 = (inp[11]) ? 4'b1000 : 4'b1010;
												assign node714 = (inp[1]) ? node724 : node715;
													assign node715 = (inp[6]) ? node721 : node716;
														assign node716 = (inp[11]) ? 4'b1000 : node717;
															assign node717 = (inp[8]) ? 4'b1010 : 4'b1000;
														assign node721 = (inp[11]) ? 4'b1010 : 4'b1000;
													assign node724 = (inp[11]) ? node728 : node725;
														assign node725 = (inp[6]) ? 4'b1010 : 4'b1000;
														assign node728 = (inp[6]) ? 4'b1000 : 4'b1010;
											assign node731 = (inp[1]) ? node739 : node732;
												assign node732 = (inp[11]) ? 4'b1000 : node733;
													assign node733 = (inp[15]) ? 4'b1010 : node734;
														assign node734 = (inp[6]) ? 4'b1000 : 4'b1010;
												assign node739 = (inp[6]) ? node747 : node740;
													assign node740 = (inp[11]) ? node742 : 4'b1000;
														assign node742 = (inp[15]) ? node744 : 4'b1010;
															assign node744 = (inp[8]) ? 4'b1000 : 4'b1010;
													assign node747 = (inp[15]) ? node749 : 4'b1010;
														assign node749 = (inp[11]) ? 4'b1010 : 4'b1000;
								assign node752 = (inp[5]) ? node810 : node753;
									assign node753 = (inp[6]) ? node789 : node754;
										assign node754 = (inp[4]) ? node776 : node755;
											assign node755 = (inp[1]) ? node767 : node756;
												assign node756 = (inp[15]) ? node762 : node757;
													assign node757 = (inp[8]) ? 4'b0010 : node758;
														assign node758 = (inp[11]) ? 4'b0000 : 4'b0010;
													assign node762 = (inp[8]) ? node764 : 4'b0010;
														assign node764 = (inp[11]) ? 4'b0010 : 4'b0000;
												assign node767 = (inp[15]) ? node773 : node768;
													assign node768 = (inp[8]) ? node770 : 4'b1000;
														assign node770 = (inp[11]) ? 4'b1000 : 4'b1010;
													assign node773 = (inp[11]) ? 4'b0010 : 4'b1010;
											assign node776 = (inp[1]) ? node782 : node777;
												assign node777 = (inp[11]) ? node779 : 4'b0000;
													assign node779 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node782 = (inp[8]) ? node784 : 4'b0000;
													assign node784 = (inp[11]) ? 4'b0000 : node785;
														assign node785 = (inp[15]) ? 4'b0010 : 4'b0000;
										assign node789 = (inp[4]) ? node799 : node790;
											assign node790 = (inp[1]) ? 4'b1010 : node791;
												assign node791 = (inp[11]) ? node793 : 4'b1000;
													assign node793 = (inp[8]) ? 4'b0000 : node794;
														assign node794 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node799 = (inp[11]) ? node807 : node800;
												assign node800 = (inp[8]) ? node802 : 4'b0010;
													assign node802 = (inp[1]) ? 4'b0010 : node803;
														assign node803 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node807 = (inp[1]) ? 4'b0010 : 4'b1010;
									assign node810 = (inp[6]) ? node844 : node811;
										assign node811 = (inp[4]) ? node829 : node812;
											assign node812 = (inp[15]) ? node820 : node813;
												assign node813 = (inp[1]) ? node817 : node814;
													assign node814 = (inp[11]) ? 4'b0010 : 4'b0000;
													assign node817 = (inp[11]) ? 4'b0010 : 4'b1010;
												assign node820 = (inp[11]) ? node824 : node821;
													assign node821 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node824 = (inp[10]) ? 4'b0000 : node825;
														assign node825 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node829 = (inp[11]) ? node837 : node830;
												assign node830 = (inp[1]) ? node832 : 4'b1010;
													assign node832 = (inp[10]) ? node834 : 4'b0010;
														assign node834 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node837 = (inp[1]) ? 4'b1010 : node838;
													assign node838 = (inp[8]) ? node840 : 4'b1000;
														assign node840 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node844 = (inp[1]) ? node858 : node845;
											assign node845 = (inp[4]) ? node851 : node846;
												assign node846 = (inp[11]) ? node848 : 4'b0010;
													assign node848 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node851 = (inp[11]) ? node853 : 4'b0000;
													assign node853 = (inp[8]) ? 4'b1000 : node854;
														assign node854 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node858 = (inp[4]) ? 4'b0000 : 4'b1000;
						assign node861 = (inp[7]) ? node1031 : node862;
							assign node862 = (inp[4]) ? node966 : node863;
								assign node863 = (inp[1]) ? node929 : node864;
									assign node864 = (inp[2]) ? node892 : node865;
										assign node865 = (inp[13]) ? node875 : node866;
											assign node866 = (inp[11]) ? 4'b1000 : node867;
												assign node867 = (inp[5]) ? node869 : 4'b1010;
													assign node869 = (inp[15]) ? node871 : 4'b1010;
														assign node871 = (inp[6]) ? 4'b1010 : 4'b1000;
											assign node875 = (inp[11]) ? node885 : node876;
												assign node876 = (inp[6]) ? 4'b1000 : node877;
													assign node877 = (inp[8]) ? node879 : 4'b1000;
														assign node879 = (inp[15]) ? node881 : 4'b1000;
															assign node881 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node885 = (inp[5]) ? 4'b1010 : node886;
													assign node886 = (inp[6]) ? node888 : 4'b1010;
														assign node888 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node892 = (inp[6]) ? node908 : node893;
											assign node893 = (inp[11]) ? node905 : node894;
												assign node894 = (inp[13]) ? node898 : node895;
													assign node895 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node898 = (inp[15]) ? node900 : 4'b1000;
														assign node900 = (inp[8]) ? node902 : 4'b1000;
															assign node902 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node905 = (inp[13]) ? 4'b1010 : 4'b1000;
											assign node908 = (inp[15]) ? node922 : node909;
												assign node909 = (inp[11]) ? node915 : node910;
													assign node910 = (inp[13]) ? node912 : 4'b1010;
														assign node912 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node915 = (inp[8]) ? 4'b1000 : node916;
														assign node916 = (inp[5]) ? 4'b1000 : node917;
															assign node917 = (inp[10]) ? 4'b1010 : 4'b1000;
												assign node922 = (inp[11]) ? node926 : node923;
													assign node923 = (inp[13]) ? 4'b1000 : 4'b1010;
													assign node926 = (inp[13]) ? 4'b1010 : 4'b1000;
									assign node929 = (inp[11]) ? node947 : node930;
										assign node930 = (inp[6]) ? node942 : node931;
											assign node931 = (inp[5]) ? node939 : node932;
												assign node932 = (inp[13]) ? 4'b1010 : node933;
													assign node933 = (inp[15]) ? 4'b1010 : node934;
														assign node934 = (inp[2]) ? 4'b1000 : 4'b1010;
												assign node939 = (inp[13]) ? 4'b1000 : 4'b1010;
											assign node942 = (inp[5]) ? 4'b1010 : node943;
												assign node943 = (inp[13]) ? 4'b1010 : 4'b1000;
										assign node947 = (inp[13]) ? node961 : node948;
											assign node948 = (inp[5]) ? node956 : node949;
												assign node949 = (inp[6]) ? 4'b1010 : node950;
													assign node950 = (inp[15]) ? node952 : 4'b1010;
														assign node952 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node956 = (inp[6]) ? node958 : 4'b1000;
													assign node958 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node961 = (inp[5]) ? node963 : 4'b1000;
												assign node963 = (inp[6]) ? 4'b1000 : 4'b1010;
								assign node966 = (inp[11]) ? node1004 : node967;
									assign node967 = (inp[13]) ? node983 : node968;
										assign node968 = (inp[1]) ? node976 : node969;
											assign node969 = (inp[5]) ? 4'b0010 : node970;
												assign node970 = (inp[6]) ? 4'b1000 : node971;
													assign node971 = (inp[15]) ? 4'b0010 : 4'b1000;
											assign node976 = (inp[15]) ? node978 : 4'b1000;
												assign node978 = (inp[6]) ? 4'b1000 : node979;
													assign node979 = (inp[5]) ? 4'b0010 : 4'b1000;
										assign node983 = (inp[1]) ? node993 : node984;
											assign node984 = (inp[5]) ? 4'b1000 : node985;
												assign node985 = (inp[6]) ? node987 : 4'b1000;
													assign node987 = (inp[8]) ? node989 : 4'b1010;
														assign node989 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node993 = (inp[5]) ? node995 : 4'b1010;
												assign node995 = (inp[6]) ? 4'b1010 : node996;
													assign node996 = (inp[15]) ? 4'b1000 : node997;
														assign node997 = (inp[2]) ? 4'b1010 : node998;
															assign node998 = (inp[8]) ? 4'b1000 : 4'b1010;
									assign node1004 = (inp[13]) ? node1016 : node1005;
										assign node1005 = (inp[15]) ? node1007 : 4'b0010;
											assign node1007 = (inp[1]) ? 4'b0010 : node1008;
												assign node1008 = (inp[5]) ? node1010 : 4'b0010;
													assign node1010 = (inp[8]) ? 4'b0000 : node1011;
														assign node1011 = (inp[6]) ? 4'b0010 : 4'b0000;
										assign node1016 = (inp[1]) ? node1024 : node1017;
											assign node1017 = (inp[5]) ? 4'b0010 : node1018;
												assign node1018 = (inp[6]) ? 4'b1000 : node1019;
													assign node1019 = (inp[15]) ? 4'b0010 : 4'b1000;
											assign node1024 = (inp[6]) ? 4'b1000 : node1025;
												assign node1025 = (inp[5]) ? node1027 : 4'b1000;
													assign node1027 = (inp[15]) ? 4'b0010 : 4'b1000;
							assign node1031 = (inp[13]) ? node1185 : node1032;
								assign node1032 = (inp[1]) ? node1122 : node1033;
									assign node1033 = (inp[4]) ? node1085 : node1034;
										assign node1034 = (inp[11]) ? node1062 : node1035;
											assign node1035 = (inp[5]) ? node1049 : node1036;
												assign node1036 = (inp[6]) ? node1044 : node1037;
													assign node1037 = (inp[2]) ? 4'b0001 : node1038;
														assign node1038 = (inp[15]) ? 4'b0011 : node1039;
															assign node1039 = (inp[8]) ? 4'b0011 : 4'b0001;
													assign node1044 = (inp[15]) ? 4'b1001 : node1045;
														assign node1045 = (inp[8]) ? 4'b1001 : 4'b1011;
												assign node1049 = (inp[6]) ? node1057 : node1050;
													assign node1050 = (inp[10]) ? 4'b0001 : node1051;
														assign node1051 = (inp[8]) ? 4'b0001 : node1052;
															assign node1052 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node1057 = (inp[8]) ? node1059 : 4'b0011;
														assign node1059 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node1062 = (inp[6]) ? node1076 : node1063;
												assign node1063 = (inp[5]) ? node1071 : node1064;
													assign node1064 = (inp[8]) ? node1066 : 4'b1010;
														assign node1066 = (inp[10]) ? node1068 : 4'b1010;
															assign node1068 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node1071 = (inp[8]) ? node1073 : 4'b1000;
														assign node1073 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node1076 = (inp[15]) ? node1082 : node1077;
													assign node1077 = (inp[8]) ? 4'b0001 : node1078;
														assign node1078 = (inp[10]) ? 4'b0011 : 4'b0001;
													assign node1082 = (inp[5]) ? 4'b0001 : 4'b0011;
										assign node1085 = (inp[11]) ? node1101 : node1086;
											assign node1086 = (inp[5]) ? node1096 : node1087;
												assign node1087 = (inp[15]) ? node1089 : 4'b1010;
													assign node1089 = (inp[8]) ? 4'b1000 : node1090;
														assign node1090 = (inp[10]) ? node1092 : 4'b1010;
															assign node1092 = (inp[6]) ? 4'b1010 : 4'b1000;
												assign node1096 = (inp[15]) ? node1098 : 4'b1000;
													assign node1098 = (inp[6]) ? 4'b1010 : 4'b0010;
											assign node1101 = (inp[5]) ? node1111 : node1102;
												assign node1102 = (inp[6]) ? node1108 : node1103;
													assign node1103 = (inp[10]) ? 4'b0000 : node1104;
														assign node1104 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node1108 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node1111 = (inp[15]) ? node1117 : node1112;
													assign node1112 = (inp[6]) ? 4'b0010 : node1113;
														assign node1113 = (inp[8]) ? 4'b0010 : 4'b0000;
													assign node1117 = (inp[8]) ? node1119 : 4'b0010;
														assign node1119 = (inp[6]) ? 4'b0000 : 4'b0010;
									assign node1122 = (inp[15]) ? node1156 : node1123;
										assign node1123 = (inp[6]) ? node1153 : node1124;
											assign node1124 = (inp[11]) ? node1144 : node1125;
												assign node1125 = (inp[10]) ? node1133 : node1126;
													assign node1126 = (inp[8]) ? node1128 : 4'b0011;
														assign node1128 = (inp[2]) ? 4'b0011 : node1129;
															assign node1129 = (inp[4]) ? 4'b0011 : 4'b1011;
													assign node1133 = (inp[4]) ? node1139 : node1134;
														assign node1134 = (inp[5]) ? 4'b1011 : node1135;
															assign node1135 = (inp[8]) ? 4'b0001 : 4'b0011;
														assign node1139 = (inp[8]) ? 4'b0001 : node1140;
															assign node1140 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node1144 = (inp[4]) ? node1148 : node1145;
													assign node1145 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node1148 = (inp[5]) ? node1150 : 4'b1010;
														assign node1150 = (inp[8]) ? 4'b1010 : 4'b1000;
											assign node1153 = (inp[11]) ? 4'b0011 : 4'b1011;
										assign node1156 = (inp[6]) ? node1182 : node1157;
											assign node1157 = (inp[11]) ? node1173 : node1158;
												assign node1158 = (inp[10]) ? node1168 : node1159;
													assign node1159 = (inp[5]) ? 4'b1011 : node1160;
														assign node1160 = (inp[2]) ? node1162 : 4'b0011;
															assign node1162 = (inp[8]) ? node1164 : 4'b0001;
																assign node1164 = (inp[4]) ? 4'b0011 : 4'b0001;
													assign node1168 = (inp[5]) ? node1170 : 4'b0001;
														assign node1170 = (inp[4]) ? 4'b0001 : 4'b1001;
												assign node1173 = (inp[4]) ? node1179 : node1174;
													assign node1174 = (inp[5]) ? 4'b0011 : node1175;
														assign node1175 = (inp[8]) ? 4'b1001 : 4'b1011;
													assign node1179 = (inp[10]) ? 4'b1000 : 4'b1010;
											assign node1182 = (inp[11]) ? 4'b0001 : 4'b1001;
								assign node1185 = (inp[6]) ? node1279 : node1186;
									assign node1186 = (inp[1]) ? node1264 : node1187;
										assign node1187 = (inp[4]) ? node1231 : node1188;
											assign node1188 = (inp[11]) ? node1216 : node1189;
												assign node1189 = (inp[5]) ? node1199 : node1190;
													assign node1190 = (inp[8]) ? node1196 : node1191;
														assign node1191 = (inp[15]) ? node1193 : 4'b0000;
															assign node1193 = (inp[2]) ? 4'b0000 : 4'b0010;
														assign node1196 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node1199 = (inp[10]) ? node1203 : node1200;
														assign node1200 = (inp[8]) ? 4'b1010 : 4'b1000;
														assign node1203 = (inp[2]) ? node1211 : node1204;
															assign node1204 = (inp[8]) ? node1208 : node1205;
																assign node1205 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node1208 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node1211 = (inp[8]) ? 4'b1000 : node1212;
																assign node1212 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node1216 = (inp[5]) ? node1222 : node1217;
													assign node1217 = (inp[15]) ? node1219 : 4'b1000;
														assign node1219 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1222 = (inp[8]) ? node1228 : node1223;
														assign node1223 = (inp[10]) ? 4'b0000 : node1224;
															assign node1224 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node1228 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node1231 = (inp[15]) ? node1245 : node1232;
												assign node1232 = (inp[11]) ? node1236 : node1233;
													assign node1233 = (inp[8]) ? 4'b1001 : 4'b1011;
													assign node1236 = (inp[5]) ? node1240 : node1237;
														assign node1237 = (inp[8]) ? 4'b0011 : 4'b0001;
														assign node1240 = (inp[8]) ? node1242 : 4'b1011;
															assign node1242 = (inp[2]) ? 4'b1001 : 4'b1011;
												assign node1245 = (inp[11]) ? node1255 : node1246;
													assign node1246 = (inp[5]) ? node1250 : node1247;
														assign node1247 = (inp[8]) ? 4'b1011 : 4'b1001;
														assign node1250 = (inp[8]) ? node1252 : 4'b0011;
															assign node1252 = (inp[10]) ? 4'b0001 : 4'b0011;
													assign node1255 = (inp[5]) ? node1261 : node1256;
														assign node1256 = (inp[8]) ? 4'b0001 : node1257;
															assign node1257 = (inp[10]) ? 4'b0001 : 4'b0011;
														assign node1261 = (inp[8]) ? 4'b1011 : 4'b1001;
										assign node1264 = (inp[10]) ? node1272 : node1265;
											assign node1265 = (inp[11]) ? node1269 : node1266;
												assign node1266 = (inp[15]) ? 4'b0111 : 4'b1111;
												assign node1269 = (inp[15]) ? 4'b0110 : 4'b1110;
											assign node1272 = (inp[15]) ? node1276 : node1273;
												assign node1273 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node1276 = (inp[11]) ? 4'b0100 : 4'b0101;
									assign node1279 = (inp[1]) ? 4'b0000 : node1280;
										assign node1280 = (inp[8]) ? node1288 : node1281;
											assign node1281 = (inp[4]) ? node1285 : node1282;
												assign node1282 = (inp[5]) ? 4'b0011 : 4'b1011;
												assign node1285 = (inp[5]) ? 4'b0010 : 4'b1010;
											assign node1288 = (inp[5]) ? node1292 : node1289;
												assign node1289 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node1292 = (inp[4]) ? 4'b0000 : 4'b0001;
			assign node1296 = (inp[0]) ? node1298 : 4'b0000;
				assign node1298 = (inp[4]) ? node1772 : node1299;
					assign node1299 = (inp[7]) ? node1457 : node1300;
						assign node1300 = (inp[3]) ? node1352 : node1301;
							assign node1301 = (inp[11]) ? 4'b0000 : node1302;
								assign node1302 = (inp[9]) ? node1326 : node1303;
									assign node1303 = (inp[5]) ? 4'b0000 : node1304;
										assign node1304 = (inp[15]) ? node1316 : node1305;
											assign node1305 = (inp[13]) ? 4'b0010 : node1306;
												assign node1306 = (inp[8]) ? node1308 : 4'b0010;
													assign node1308 = (inp[1]) ? node1310 : 4'b0000;
														assign node1310 = (inp[2]) ? node1312 : 4'b0010;
															assign node1312 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node1316 = (inp[13]) ? node1318 : 4'b0000;
												assign node1318 = (inp[8]) ? node1320 : 4'b0010;
													assign node1320 = (inp[1]) ? node1322 : 4'b0000;
														assign node1322 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node1326 = (inp[5]) ? node1328 : 4'b0010;
										assign node1328 = (inp[15]) ? node1340 : node1329;
											assign node1329 = (inp[1]) ? 4'b0010 : node1330;
												assign node1330 = (inp[13]) ? 4'b0010 : node1331;
													assign node1331 = (inp[8]) ? 4'b0000 : node1332;
														assign node1332 = (inp[6]) ? 4'b0010 : node1333;
															assign node1333 = (inp[2]) ? 4'b0010 : 4'b0000;
											assign node1340 = (inp[13]) ? node1342 : 4'b0000;
												assign node1342 = (inp[8]) ? node1344 : 4'b0010;
													assign node1344 = (inp[1]) ? node1346 : 4'b0000;
														assign node1346 = (inp[10]) ? node1348 : 4'b0010;
															assign node1348 = (inp[6]) ? 4'b0010 : 4'b0000;
							assign node1352 = (inp[11]) ? node1422 : node1353;
								assign node1353 = (inp[13]) ? node1381 : node1354;
									assign node1354 = (inp[9]) ? node1370 : node1355;
										assign node1355 = (inp[5]) ? 4'b0010 : node1356;
											assign node1356 = (inp[1]) ? node1362 : node1357;
												assign node1357 = (inp[15]) ? 4'b0010 : node1358;
													assign node1358 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node1362 = (inp[6]) ? 4'b0000 : node1363;
													assign node1363 = (inp[8]) ? node1365 : 4'b0000;
														assign node1365 = (inp[10]) ? 4'b0010 : 4'b0000;
										assign node1370 = (inp[1]) ? node1372 : 4'b0000;
											assign node1372 = (inp[5]) ? 4'b0000 : node1373;
												assign node1373 = (inp[15]) ? 4'b0000 : node1374;
													assign node1374 = (inp[6]) ? 4'b0010 : node1375;
														assign node1375 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node1381 = (inp[9]) ? node1397 : node1382;
										assign node1382 = (inp[5]) ? node1384 : 4'b0000;
											assign node1384 = (inp[1]) ? node1392 : node1385;
												assign node1385 = (inp[15]) ? 4'b0010 : node1386;
													assign node1386 = (inp[8]) ? node1388 : 4'b0000;
														assign node1388 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node1392 = (inp[6]) ? 4'b0000 : node1393;
													assign node1393 = (inp[15]) ? 4'b0010 : 4'b0000;
										assign node1397 = (inp[5]) ? node1407 : node1398;
											assign node1398 = (inp[10]) ? node1400 : 4'b0010;
												assign node1400 = (inp[2]) ? 4'b0010 : node1401;
													assign node1401 = (inp[6]) ? 4'b0010 : node1402;
														assign node1402 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node1407 = (inp[1]) ? node1415 : node1408;
												assign node1408 = (inp[6]) ? node1410 : 4'b0000;
													assign node1410 = (inp[15]) ? 4'b0000 : node1411;
														assign node1411 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node1415 = (inp[6]) ? 4'b0010 : node1416;
													assign node1416 = (inp[2]) ? 4'b0010 : node1417;
														assign node1417 = (inp[15]) ? 4'b0000 : 4'b0010;
								assign node1422 = (inp[9]) ? node1424 : 4'b0010;
									assign node1424 = (inp[13]) ? node1440 : node1425;
										assign node1425 = (inp[5]) ? 4'b0010 : node1426;
											assign node1426 = (inp[1]) ? node1432 : node1427;
												assign node1427 = (inp[15]) ? 4'b0010 : node1428;
													assign node1428 = (inp[2]) ? 4'b0000 : 4'b0010;
												assign node1432 = (inp[8]) ? node1434 : 4'b0000;
													assign node1434 = (inp[6]) ? 4'b0000 : node1435;
														assign node1435 = (inp[15]) ? 4'b0010 : 4'b0000;
										assign node1440 = (inp[5]) ? node1442 : 4'b0000;
											assign node1442 = (inp[15]) ? node1452 : node1443;
												assign node1443 = (inp[2]) ? 4'b0000 : node1444;
													assign node1444 = (inp[1]) ? 4'b0000 : node1445;
														assign node1445 = (inp[6]) ? 4'b0000 : node1446;
															assign node1446 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node1452 = (inp[1]) ? node1454 : 4'b0010;
													assign node1454 = (inp[10]) ? 4'b0010 : 4'b0000;
						assign node1457 = (inp[3]) ? node1515 : node1458;
							assign node1458 = (inp[11]) ? node1460 : 4'b0010;
								assign node1460 = (inp[5]) ? node1492 : node1461;
									assign node1461 = (inp[9]) ? 4'b0010 : node1462;
										assign node1462 = (inp[13]) ? node1480 : node1463;
											assign node1463 = (inp[15]) ? 4'b0000 : node1464;
												assign node1464 = (inp[8]) ? node1472 : node1465;
													assign node1465 = (inp[6]) ? 4'b0010 : node1466;
														assign node1466 = (inp[10]) ? node1468 : 4'b0010;
															assign node1468 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node1472 = (inp[1]) ? node1474 : 4'b0000;
														assign node1474 = (inp[6]) ? 4'b0010 : node1475;
															assign node1475 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node1480 = (inp[8]) ? node1482 : 4'b0010;
												assign node1482 = (inp[15]) ? node1484 : 4'b0010;
													assign node1484 = (inp[1]) ? node1486 : 4'b0000;
														assign node1486 = (inp[6]) ? 4'b0010 : node1487;
															assign node1487 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node1492 = (inp[9]) ? node1494 : 4'b0000;
										assign node1494 = (inp[15]) ? node1506 : node1495;
											assign node1495 = (inp[13]) ? 4'b0010 : node1496;
												assign node1496 = (inp[1]) ? node1500 : node1497;
													assign node1497 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1500 = (inp[6]) ? 4'b0010 : node1501;
														assign node1501 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node1506 = (inp[13]) ? node1508 : 4'b0000;
												assign node1508 = (inp[1]) ? 4'b0010 : node1509;
													assign node1509 = (inp[8]) ? 4'b0000 : node1510;
														assign node1510 = (inp[2]) ? 4'b0000 : 4'b0010;
							assign node1515 = (inp[13]) ? node1633 : node1516;
								assign node1516 = (inp[11]) ? node1568 : node1517;
									assign node1517 = (inp[1]) ? node1545 : node1518;
										assign node1518 = (inp[5]) ? node1534 : node1519;
											assign node1519 = (inp[9]) ? node1525 : node1520;
												assign node1520 = (inp[6]) ? 4'b1000 : node1521;
													assign node1521 = (inp[15]) ? 4'b0010 : 4'b1000;
												assign node1525 = (inp[6]) ? node1531 : node1526;
													assign node1526 = (inp[10]) ? 4'b0000 : node1527;
														assign node1527 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1531 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node1534 = (inp[6]) ? node1538 : node1535;
												assign node1535 = (inp[9]) ? 4'b1010 : 4'b0010;
												assign node1538 = (inp[9]) ? node1540 : 4'b0010;
													assign node1540 = (inp[15]) ? 4'b0000 : node1541;
														assign node1541 = (inp[8]) ? 4'b0000 : 4'b0010;
										assign node1545 = (inp[6]) ? node1561 : node1546;
											assign node1546 = (inp[15]) ? node1552 : node1547;
												assign node1547 = (inp[5]) ? node1549 : 4'b1000;
													assign node1549 = (inp[9]) ? 4'b0010 : 4'b1000;
												assign node1552 = (inp[9]) ? node1556 : node1553;
													assign node1553 = (inp[5]) ? 4'b0010 : 4'b1000;
													assign node1556 = (inp[5]) ? node1558 : 4'b0010;
														assign node1558 = (inp[8]) ? 4'b0010 : 4'b0000;
											assign node1561 = (inp[15]) ? 4'b1000 : node1562;
												assign node1562 = (inp[5]) ? node1564 : 4'b1010;
													assign node1564 = (inp[9]) ? 4'b1010 : 4'b1000;
									assign node1568 = (inp[9]) ? node1590 : node1569;
										assign node1569 = (inp[5]) ? node1579 : node1570;
											assign node1570 = (inp[1]) ? 4'b0010 : node1571;
												assign node1571 = (inp[15]) ? node1573 : 4'b0010;
													assign node1573 = (inp[6]) ? node1575 : 4'b0000;
														assign node1575 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node1579 = (inp[1]) ? node1581 : 4'b0000;
												assign node1581 = (inp[15]) ? 4'b0000 : node1582;
													assign node1582 = (inp[2]) ? 4'b0010 : node1583;
														assign node1583 = (inp[10]) ? 4'b0000 : node1584;
															assign node1584 = (inp[8]) ? 4'b0000 : 4'b0010;
										assign node1590 = (inp[1]) ? node1618 : node1591;
											assign node1591 = (inp[2]) ? node1601 : node1592;
												assign node1592 = (inp[8]) ? node1594 : 4'b1010;
													assign node1594 = (inp[10]) ? 4'b1010 : node1595;
														assign node1595 = (inp[6]) ? node1597 : 4'b1000;
															assign node1597 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node1601 = (inp[15]) ? node1609 : node1602;
													assign node1602 = (inp[5]) ? node1606 : node1603;
														assign node1603 = (inp[6]) ? 4'b1010 : 4'b1000;
														assign node1606 = (inp[6]) ? 4'b1000 : 4'b1010;
													assign node1609 = (inp[10]) ? node1613 : node1610;
														assign node1610 = (inp[8]) ? 4'b1000 : 4'b1010;
														assign node1613 = (inp[6]) ? 4'b1010 : node1614;
															assign node1614 = (inp[8]) ? 4'b1010 : 4'b1000;
											assign node1618 = (inp[15]) ? node1628 : node1619;
												assign node1619 = (inp[6]) ? 4'b0010 : node1620;
													assign node1620 = (inp[5]) ? 4'b1010 : node1621;
														assign node1621 = (inp[10]) ? node1623 : 4'b0010;
															assign node1623 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node1628 = (inp[6]) ? 4'b0000 : node1629;
													assign node1629 = (inp[5]) ? 4'b1000 : 4'b0000;
								assign node1633 = (inp[9]) ? node1703 : node1634;
									assign node1634 = (inp[11]) ? node1684 : node1635;
										assign node1635 = (inp[5]) ? node1661 : node1636;
											assign node1636 = (inp[15]) ? node1656 : node1637;
												assign node1637 = (inp[10]) ? node1647 : node1638;
													assign node1638 = (inp[8]) ? node1640 : 4'b1010;
														assign node1640 = (inp[6]) ? node1644 : node1641;
															assign node1641 = (inp[1]) ? 4'b1000 : 4'b1010;
															assign node1644 = (inp[1]) ? 4'b1010 : 4'b1000;
													assign node1647 = (inp[2]) ? node1651 : node1648;
														assign node1648 = (inp[6]) ? 4'b1000 : 4'b1010;
														assign node1651 = (inp[6]) ? node1653 : 4'b1000;
															assign node1653 = (inp[1]) ? 4'b1010 : 4'b1000;
												assign node1656 = (inp[1]) ? node1658 : 4'b1010;
													assign node1658 = (inp[6]) ? 4'b1010 : 4'b1000;
											assign node1661 = (inp[8]) ? node1675 : node1662;
												assign node1662 = (inp[1]) ? node1670 : node1663;
													assign node1663 = (inp[6]) ? 4'b1010 : node1664;
														assign node1664 = (inp[10]) ? 4'b1000 : node1665;
															assign node1665 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node1670 = (inp[15]) ? node1672 : 4'b1000;
														assign node1672 = (inp[6]) ? 4'b1000 : 4'b1010;
												assign node1675 = (inp[1]) ? node1681 : node1676;
													assign node1676 = (inp[15]) ? 4'b1000 : node1677;
														assign node1677 = (inp[6]) ? 4'b1010 : 4'b1000;
													assign node1681 = (inp[6]) ? 4'b1000 : 4'b1010;
										assign node1684 = (inp[1]) ? node1692 : node1685;
											assign node1685 = (inp[5]) ? 4'b0010 : node1686;
												assign node1686 = (inp[15]) ? node1688 : 4'b1000;
													assign node1688 = (inp[6]) ? 4'b1000 : 4'b0010;
											assign node1692 = (inp[5]) ? node1698 : node1693;
												assign node1693 = (inp[6]) ? 4'b1010 : node1694;
													assign node1694 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node1698 = (inp[15]) ? node1700 : 4'b1000;
													assign node1700 = (inp[6]) ? 4'b1000 : 4'b0010;
									assign node1703 = (inp[1]) ? node1755 : node1704;
										assign node1704 = (inp[5]) ? node1736 : node1705;
											assign node1705 = (inp[11]) ? node1721 : node1706;
												assign node1706 = (inp[8]) ? node1714 : node1707;
													assign node1707 = (inp[6]) ? 4'b1011 : node1708;
														assign node1708 = (inp[15]) ? 4'b0011 : node1709;
															assign node1709 = (inp[10]) ? 4'b1001 : 4'b1011;
													assign node1714 = (inp[15]) ? node1716 : 4'b1001;
														assign node1716 = (inp[6]) ? 4'b1001 : node1717;
															assign node1717 = (inp[10]) ? 4'b0001 : 4'b0011;
												assign node1721 = (inp[6]) ? node1733 : node1722;
													assign node1722 = (inp[10]) ? node1724 : 4'b1010;
														assign node1724 = (inp[2]) ? node1726 : 4'b1000;
															assign node1726 = (inp[8]) ? node1730 : node1727;
																assign node1727 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node1730 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node1733 = (inp[8]) ? 4'b1001 : 4'b1011;
											assign node1736 = (inp[6]) ? node1752 : node1737;
												assign node1737 = (inp[11]) ? node1745 : node1738;
													assign node1738 = (inp[15]) ? node1740 : 4'b0011;
														assign node1740 = (inp[10]) ? 4'b0001 : node1741;
															assign node1741 = (inp[8]) ? 4'b0001 : 4'b0011;
													assign node1745 = (inp[15]) ? 4'b0010 : node1746;
														assign node1746 = (inp[10]) ? 4'b1000 : node1747;
															assign node1747 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node1752 = (inp[8]) ? 4'b0001 : 4'b0011;
										assign node1755 = (inp[6]) ? 4'b0000 : node1756;
											assign node1756 = (inp[15]) ? node1764 : node1757;
												assign node1757 = (inp[10]) ? node1761 : node1758;
													assign node1758 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node1761 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node1764 = (inp[10]) ? node1768 : node1765;
													assign node1765 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node1768 = (inp[11]) ? 4'b0000 : 4'b0001;
					assign node1772 = (inp[3]) ? node1774 : 4'b0000;
						assign node1774 = (inp[11]) ? node1942 : node1775;
							assign node1775 = (inp[9]) ? node1855 : node1776;
								assign node1776 = (inp[7]) ? node1810 : node1777;
									assign node1777 = (inp[5]) ? 4'b0000 : node1778;
										assign node1778 = (inp[13]) ? node1794 : node1779;
											assign node1779 = (inp[15]) ? 4'b0000 : node1780;
												assign node1780 = (inp[1]) ? node1786 : node1781;
													assign node1781 = (inp[6]) ? node1783 : 4'b0000;
														assign node1783 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1786 = (inp[8]) ? node1788 : 4'b0010;
														assign node1788 = (inp[10]) ? node1790 : 4'b0010;
															assign node1790 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node1794 = (inp[15]) ? node1796 : 4'b0010;
												assign node1796 = (inp[1]) ? node1802 : node1797;
													assign node1797 = (inp[8]) ? 4'b0000 : node1798;
														assign node1798 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1802 = (inp[6]) ? 4'b0010 : node1803;
														assign node1803 = (inp[8]) ? node1805 : 4'b0010;
															assign node1805 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node1810 = (inp[5]) ? node1838 : node1811;
										assign node1811 = (inp[15]) ? node1821 : node1812;
											assign node1812 = (inp[13]) ? node1814 : 4'b0000;
												assign node1814 = (inp[1]) ? 4'b0010 : node1815;
													assign node1815 = (inp[8]) ? 4'b0000 : node1816;
														assign node1816 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node1821 = (inp[13]) ? node1829 : node1822;
												assign node1822 = (inp[1]) ? node1824 : 4'b0010;
													assign node1824 = (inp[6]) ? 4'b0000 : node1825;
														assign node1825 = (inp[10]) ? 4'b0010 : 4'b0000;
												assign node1829 = (inp[1]) ? node1831 : 4'b0000;
													assign node1831 = (inp[6]) ? 4'b0010 : node1832;
														assign node1832 = (inp[10]) ? 4'b0000 : node1833;
															assign node1833 = (inp[8]) ? 4'b0000 : 4'b0010;
										assign node1838 = (inp[13]) ? node1840 : 4'b0010;
											assign node1840 = (inp[1]) ? node1848 : node1841;
												assign node1841 = (inp[15]) ? 4'b0010 : node1842;
													assign node1842 = (inp[8]) ? node1844 : 4'b0000;
														assign node1844 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node1848 = (inp[6]) ? 4'b0000 : node1849;
													assign node1849 = (inp[15]) ? node1851 : 4'b0000;
														assign node1851 = (inp[8]) ? 4'b0010 : 4'b0000;
								assign node1855 = (inp[7]) ? node1879 : node1856;
									assign node1856 = (inp[5]) ? node1858 : 4'b0010;
										assign node1858 = (inp[13]) ? node1872 : node1859;
											assign node1859 = (inp[15]) ? 4'b0000 : node1860;
												assign node1860 = (inp[8]) ? node1866 : node1861;
													assign node1861 = (inp[10]) ? node1863 : 4'b0010;
														assign node1863 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1866 = (inp[1]) ? node1868 : 4'b0000;
														assign node1868 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node1872 = (inp[1]) ? 4'b0010 : node1873;
												assign node1873 = (inp[8]) ? node1875 : 4'b0010;
													assign node1875 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node1879 = (inp[13]) ? node1911 : node1880;
										assign node1880 = (inp[1]) ? node1902 : node1881;
											assign node1881 = (inp[5]) ? node1891 : node1882;
												assign node1882 = (inp[6]) ? node1886 : node1883;
													assign node1883 = (inp[15]) ? 4'b0010 : 4'b1000;
													assign node1886 = (inp[15]) ? 4'b1000 : node1887;
														assign node1887 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node1891 = (inp[6]) ? node1897 : node1892;
													assign node1892 = (inp[10]) ? 4'b0000 : node1893;
														assign node1893 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node1897 = (inp[8]) ? node1899 : 4'b0010;
														assign node1899 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node1902 = (inp[15]) ? node1906 : node1903;
												assign node1903 = (inp[6]) ? 4'b1010 : 4'b1000;
												assign node1906 = (inp[6]) ? 4'b1000 : node1907;
													assign node1907 = (inp[5]) ? 4'b0010 : 4'b1010;
										assign node1911 = (inp[6]) ? node1933 : node1912;
											assign node1912 = (inp[1]) ? node1926 : node1913;
												assign node1913 = (inp[5]) ? node1919 : node1914;
													assign node1914 = (inp[8]) ? node1916 : 4'b0000;
														assign node1916 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node1919 = (inp[10]) ? node1921 : 4'b1010;
														assign node1921 = (inp[15]) ? node1923 : 4'b1000;
															assign node1923 = (inp[8]) ? 4'b1010 : 4'b1000;
												assign node1926 = (inp[15]) ? node1930 : node1927;
													assign node1927 = (inp[10]) ? 4'b1001 : 4'b1011;
													assign node1930 = (inp[10]) ? 4'b0001 : 4'b0011;
											assign node1933 = (inp[1]) ? 4'b0000 : node1934;
												assign node1934 = (inp[8]) ? node1938 : node1935;
													assign node1935 = (inp[5]) ? 4'b0010 : 4'b1010;
													assign node1938 = (inp[5]) ? 4'b0000 : 4'b1000;
							assign node1942 = (inp[7]) ? node1944 : 4'b0000;
								assign node1944 = (inp[5]) ? node2048 : node1945;
									assign node1945 = (inp[10]) ? node1997 : node1946;
										assign node1946 = (inp[6]) ? node1974 : node1947;
											assign node1947 = (inp[13]) ? node1963 : node1948;
												assign node1948 = (inp[1]) ? node1956 : node1949;
													assign node1949 = (inp[2]) ? node1951 : 4'b0010;
														assign node1951 = (inp[8]) ? 4'b0010 : node1952;
															assign node1952 = (inp[9]) ? 4'b0000 : 4'b0010;
													assign node1956 = (inp[15]) ? 4'b0000 : node1957;
														assign node1957 = (inp[8]) ? node1959 : 4'b0010;
															assign node1959 = (inp[9]) ? 4'b0000 : 4'b0010;
												assign node1963 = (inp[9]) ? node1971 : node1964;
													assign node1964 = (inp[15]) ? node1966 : 4'b0010;
														assign node1966 = (inp[1]) ? 4'b0010 : node1967;
															assign node1967 = (inp[2]) ? 4'b0000 : 4'b0010;
													assign node1971 = (inp[15]) ? 4'b0010 : 4'b1010;
											assign node1974 = (inp[9]) ? node1984 : node1975;
												assign node1975 = (inp[13]) ? 4'b0010 : node1976;
													assign node1976 = (inp[15]) ? 4'b0000 : node1977;
														assign node1977 = (inp[1]) ? 4'b0010 : node1978;
															assign node1978 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node1984 = (inp[13]) ? node1992 : node1985;
													assign node1985 = (inp[15]) ? node1989 : node1986;
														assign node1986 = (inp[1]) ? 4'b0010 : 4'b0000;
														assign node1989 = (inp[1]) ? 4'b0000 : 4'b0010;
													assign node1992 = (inp[1]) ? 4'b0000 : node1993;
														assign node1993 = (inp[8]) ? 4'b1000 : 4'b1010;
										assign node1997 = (inp[13]) ? node2021 : node1998;
											assign node1998 = (inp[9]) ? node2008 : node1999;
												assign node1999 = (inp[15]) ? 4'b0000 : node2000;
													assign node2000 = (inp[6]) ? 4'b0010 : node2001;
														assign node2001 = (inp[1]) ? node2003 : 4'b0000;
															assign node2003 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node2008 = (inp[1]) ? node2012 : node2009;
													assign node2009 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node2012 = (inp[8]) ? node2018 : node2013;
														assign node2013 = (inp[15]) ? 4'b0000 : node2014;
															assign node2014 = (inp[6]) ? 4'b0010 : 4'b0000;
														assign node2018 = (inp[6]) ? 4'b0000 : 4'b0010;
											assign node2021 = (inp[9]) ? node2029 : node2022;
												assign node2022 = (inp[1]) ? 4'b0010 : node2023;
													assign node2023 = (inp[8]) ? 4'b0000 : node2024;
														assign node2024 = (inp[6]) ? 4'b0010 : 4'b0000;
												assign node2029 = (inp[8]) ? node2037 : node2030;
													assign node2030 = (inp[1]) ? node2034 : node2031;
														assign node2031 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node2034 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node2037 = (inp[1]) ? node2043 : node2038;
														assign node2038 = (inp[6]) ? 4'b1000 : node2039;
															assign node2039 = (inp[15]) ? 4'b0000 : 4'b1000;
														assign node2043 = (inp[6]) ? 4'b0000 : node2044;
															assign node2044 = (inp[15]) ? 4'b0000 : 4'b1000;
									assign node2048 = (inp[9]) ? node2050 : 4'b0000;
										assign node2050 = (inp[15]) ? node2092 : node2051;
											assign node2051 = (inp[2]) ? node2071 : node2052;
												assign node2052 = (inp[8]) ? node2060 : node2053;
													assign node2053 = (inp[13]) ? node2055 : 4'b0010;
														assign node2055 = (inp[10]) ? node2057 : 4'b1010;
															assign node2057 = (inp[1]) ? 4'b0000 : 4'b0010;
													assign node2060 = (inp[6]) ? node2066 : node2061;
														assign node2061 = (inp[10]) ? node2063 : 4'b0010;
															assign node2063 = (inp[13]) ? 4'b0010 : 4'b0000;
														assign node2066 = (inp[1]) ? node2068 : 4'b0000;
															assign node2068 = (inp[13]) ? 4'b0000 : 4'b0010;
												assign node2071 = (inp[1]) ? node2081 : node2072;
													assign node2072 = (inp[13]) ? node2074 : 4'b0000;
														assign node2074 = (inp[6]) ? node2078 : node2075;
															assign node2075 = (inp[8]) ? 4'b0010 : 4'b0000;
															assign node2078 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node2081 = (inp[13]) ? node2087 : node2082;
														assign node2082 = (inp[10]) ? node2084 : 4'b0010;
															assign node2084 = (inp[6]) ? 4'b0010 : 4'b0000;
														assign node2087 = (inp[6]) ? 4'b0000 : node2088;
															assign node2088 = (inp[10]) ? 4'b1000 : 4'b1010;
											assign node2092 = (inp[13]) ? node2094 : 4'b0000;
												assign node2094 = (inp[10]) ? node2106 : node2095;
													assign node2095 = (inp[6]) ? node2101 : node2096;
														assign node2096 = (inp[8]) ? node2098 : 4'b0010;
															assign node2098 = (inp[1]) ? 4'b0010 : 4'b0000;
														assign node2101 = (inp[8]) ? 4'b0000 : node2102;
															assign node2102 = (inp[2]) ? 4'b0000 : 4'b0010;
													assign node2106 = (inp[1]) ? 4'b0000 : node2107;
														assign node2107 = (inp[6]) ? 4'b0010 : 4'b0000;

endmodule