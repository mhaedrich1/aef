module dtc_split25_bm86 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node101;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node197;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node205;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node219;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node234;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node239;
	wire [3-1:0] node242;
	wire [3-1:0] node243;

	assign outp = (inp[3]) ? node178 : node1;
		assign node1 = (inp[0]) ? node81 : node2;
			assign node2 = (inp[4]) ? node62 : node3;
				assign node3 = (inp[6]) ? 3'b000 : node4;
					assign node4 = (inp[9]) ? node38 : node5;
						assign node5 = (inp[7]) ? node23 : node6;
							assign node6 = (inp[1]) ? node12 : node7;
								assign node7 = (inp[2]) ? node9 : 3'b000;
									assign node9 = (inp[5]) ? 3'b000 : 3'b100;
								assign node12 = (inp[2]) ? node16 : node13;
									assign node13 = (inp[5]) ? 3'b000 : 3'b100;
									assign node16 = (inp[5]) ? node20 : node17;
										assign node17 = (inp[10]) ? 3'b110 : 3'b010;
										assign node20 = (inp[8]) ? 3'b000 : 3'b100;
							assign node23 = (inp[1]) ? node31 : node24;
								assign node24 = (inp[8]) ? node26 : 3'b010;
									assign node26 = (inp[2]) ? node28 : 3'b010;
										assign node28 = (inp[11]) ? 3'b000 : 3'b010;
								assign node31 = (inp[5]) ? node35 : node32;
									assign node32 = (inp[11]) ? 3'b100 : 3'b110;
									assign node35 = (inp[10]) ? 3'b010 : 3'b110;
						assign node38 = (inp[7]) ? node56 : node39;
							assign node39 = (inp[1]) ? node45 : node40;
								assign node40 = (inp[11]) ? node42 : 3'b110;
									assign node42 = (inp[5]) ? 3'b001 : 3'b110;
								assign node45 = (inp[5]) ? node49 : node46;
									assign node46 = (inp[8]) ? 3'b001 : 3'b101;
									assign node49 = (inp[10]) ? node53 : node50;
										assign node50 = (inp[8]) ? 3'b110 : 3'b010;
										assign node53 = (inp[2]) ? 3'b001 : 3'b000;
							assign node56 = (inp[11]) ? node58 : 3'b011;
								assign node58 = (inp[2]) ? 3'b111 : 3'b011;
				assign node62 = (inp[10]) ? node64 : 3'b000;
					assign node64 = (inp[8]) ? node66 : 3'b000;
						assign node66 = (inp[6]) ? 3'b000 : node67;
							assign node67 = (inp[5]) ? node73 : node68;
								assign node68 = (inp[2]) ? node70 : 3'b000;
									assign node70 = (inp[7]) ? 3'b000 : 3'b010;
								assign node73 = (inp[1]) ? node75 : 3'b000;
									assign node75 = (inp[11]) ? 3'b000 : node76;
										assign node76 = (inp[9]) ? 3'b100 : 3'b000;
			assign node81 = (inp[6]) ? node173 : node82;
				assign node82 = (inp[4]) ? node106 : node83;
					assign node83 = (inp[7]) ? 3'b111 : node84;
						assign node84 = (inp[1]) ? node94 : node85;
							assign node85 = (inp[2]) ? node91 : node86;
								assign node86 = (inp[5]) ? 3'b010 : node87;
									assign node87 = (inp[8]) ? 3'b011 : 3'b001;
								assign node91 = (inp[10]) ? 3'b011 : 3'b101;
							assign node94 = (inp[9]) ? node98 : node95;
								assign node95 = (inp[5]) ? 3'b101 : 3'b111;
								assign node98 = (inp[10]) ? 3'b111 : node99;
									assign node99 = (inp[11]) ? node101 : 3'b111;
										assign node101 = (inp[5]) ? 3'b011 : 3'b111;
					assign node106 = (inp[9]) ? node144 : node107;
						assign node107 = (inp[5]) ? node121 : node108;
							assign node108 = (inp[1]) ? node116 : node109;
								assign node109 = (inp[2]) ? node111 : 3'b100;
									assign node111 = (inp[10]) ? node113 : 3'b100;
										assign node113 = (inp[7]) ? 3'b100 : 3'b110;
								assign node116 = (inp[8]) ? 3'b110 : node117;
									assign node117 = (inp[7]) ? 3'b110 : 3'b000;
							assign node121 = (inp[11]) ? node131 : node122;
								assign node122 = (inp[8]) ? node128 : node123;
									assign node123 = (inp[1]) ? node125 : 3'b100;
										assign node125 = (inp[2]) ? 3'b110 : 3'b100;
									assign node128 = (inp[7]) ? 3'b100 : 3'b000;
								assign node131 = (inp[2]) ? node137 : node132;
									assign node132 = (inp[7]) ? 3'b100 : node133;
										assign node133 = (inp[8]) ? 3'b100 : 3'b010;
									assign node137 = (inp[10]) ? node141 : node138;
										assign node138 = (inp[8]) ? 3'b000 : 3'b000;
										assign node141 = (inp[7]) ? 3'b000 : 3'b100;
						assign node144 = (inp[7]) ? node166 : node145;
							assign node145 = (inp[5]) ? node155 : node146;
								assign node146 = (inp[8]) ? 3'b111 : node147;
									assign node147 = (inp[2]) ? node151 : node148;
										assign node148 = (inp[11]) ? 3'b110 : 3'b101;
										assign node151 = (inp[11]) ? 3'b101 : 3'b001;
								assign node155 = (inp[10]) ? node159 : node156;
									assign node156 = (inp[2]) ? 3'b010 : 3'b110;
									assign node159 = (inp[11]) ? node163 : node160;
										assign node160 = (inp[1]) ? 3'b001 : 3'b000;
										assign node163 = (inp[8]) ? 3'b010 : 3'b110;
							assign node166 = (inp[5]) ? node168 : 3'b111;
								assign node168 = (inp[11]) ? node170 : 3'b101;
									assign node170 = (inp[2]) ? 3'b011 : 3'b101;
				assign node173 = (inp[4]) ? 3'b000 : node174;
					assign node174 = (inp[9]) ? 3'b111 : 3'b000;
		assign node178 = (inp[0]) ? node180 : 3'b000;
			assign node180 = (inp[9]) ? node182 : 3'b000;
				assign node182 = (inp[4]) ? node230 : node183;
					assign node183 = (inp[6]) ? node217 : node184;
						assign node184 = (inp[7]) ? node202 : node185;
							assign node185 = (inp[5]) ? node195 : node186;
								assign node186 = (inp[1]) ? node190 : node187;
									assign node187 = (inp[10]) ? 3'b100 : 3'b000;
									assign node190 = (inp[10]) ? node192 : 3'b010;
										assign node192 = (inp[8]) ? 3'b010 : 3'b110;
								assign node195 = (inp[11]) ? node197 : 3'b000;
									assign node197 = (inp[8]) ? node199 : 3'b100;
										assign node199 = (inp[10]) ? 3'b010 : 3'b000;
							assign node202 = (inp[5]) ? node210 : node203;
								assign node203 = (inp[10]) ? node205 : 3'b101;
									assign node205 = (inp[11]) ? node207 : 3'b110;
										assign node207 = (inp[2]) ? 3'b000 : 3'b010;
								assign node210 = (inp[2]) ? node212 : 3'b010;
									assign node212 = (inp[11]) ? node214 : 3'b010;
										assign node214 = (inp[1]) ? 3'b110 : 3'b010;
						assign node217 = (inp[1]) ? node219 : 3'b000;
							assign node219 = (inp[5]) ? node221 : 3'b000;
								assign node221 = (inp[8]) ? node225 : node222;
									assign node222 = (inp[2]) ? 3'b001 : 3'b000;
									assign node225 = (inp[10]) ? 3'b000 : node226;
										assign node226 = (inp[7]) ? 3'b001 : 3'b000;
					assign node230 = (inp[6]) ? node232 : 3'b000;
						assign node232 = (inp[1]) ? node234 : 3'b000;
							assign node234 = (inp[2]) ? node236 : 3'b000;
								assign node236 = (inp[10]) ? node242 : node237;
									assign node237 = (inp[7]) ? node239 : 3'b000;
										assign node239 = (inp[11]) ? 3'b010 : 3'b100;
									assign node242 = (inp[11]) ? 3'b100 : node243;
										assign node243 = (inp[7]) ? 3'b000 : 3'b000;

endmodule