module dtc_split5_bm45 (
	input  wire [16-1:0] inp,
	output wire [46-1:0] outp
);

	wire [46-1:0] node1;
	wire [46-1:0] node2;
	wire [46-1:0] node5;
	wire [46-1:0] node6;
	wire [46-1:0] node7;
	wire [46-1:0] node9;
	wire [46-1:0] node11;
	wire [46-1:0] node13;
	wire [46-1:0] node15;
	wire [46-1:0] node17;
	wire [46-1:0] node18;
	wire [46-1:0] node20;
	wire [46-1:0] node22;
	wire [46-1:0] node24;
	wire [46-1:0] node27;
	wire [46-1:0] node28;
	wire [46-1:0] node30;
	wire [46-1:0] node32;
	wire [46-1:0] node36;
	wire [46-1:0] node38;
	wire [46-1:0] node39;
	wire [46-1:0] node41;
	wire [46-1:0] node43;
	wire [46-1:0] node45;
	wire [46-1:0] node47;
	wire [46-1:0] node48;
	wire [46-1:0] node52;
	wire [46-1:0] node54;
	wire [46-1:0] node56;
	wire [46-1:0] node58;
	wire [46-1:0] node60;
	wire [46-1:0] node62;
	wire [46-1:0] node64;
	wire [46-1:0] node65;
	wire [46-1:0] node69;
	wire [46-1:0] node70;
	wire [46-1:0] node71;
	wire [46-1:0] node72;
	wire [46-1:0] node73;
	wire [46-1:0] node77;
	wire [46-1:0] node79;
	wire [46-1:0] node81;
	wire [46-1:0] node82;
	wire [46-1:0] node84;
	wire [46-1:0] node85;
	wire [46-1:0] node86;
	wire [46-1:0] node88;
	wire [46-1:0] node91;
	wire [46-1:0] node92;
	wire [46-1:0] node96;
	wire [46-1:0] node97;
	wire [46-1:0] node99;
	wire [46-1:0] node102;
	wire [46-1:0] node103;
	wire [46-1:0] node106;
	wire [46-1:0] node110;
	wire [46-1:0] node111;
	wire [46-1:0] node112;
	wire [46-1:0] node116;
	wire [46-1:0] node117;
	wire [46-1:0] node120;
	wire [46-1:0] node123;
	wire [46-1:0] node124;
	wire [46-1:0] node125;
	wire [46-1:0] node126;
	wire [46-1:0] node129;
	wire [46-1:0] node131;
	wire [46-1:0] node133;
	wire [46-1:0] node134;
	wire [46-1:0] node136;
	wire [46-1:0] node138;
	wire [46-1:0] node140;
	wire [46-1:0] node143;
	wire [46-1:0] node144;
	wire [46-1:0] node146;
	wire [46-1:0] node148;
	wire [46-1:0] node151;
	wire [46-1:0] node152;
	wire [46-1:0] node154;
	wire [46-1:0] node157;
	wire [46-1:0] node158;
	wire [46-1:0] node162;
	wire [46-1:0] node163;
	wire [46-1:0] node165;
	wire [46-1:0] node166;
	wire [46-1:0] node168;
	wire [46-1:0] node170;
	wire [46-1:0] node172;
	wire [46-1:0] node174;
	wire [46-1:0] node178;
	wire [46-1:0] node180;
	wire [46-1:0] node182;
	wire [46-1:0] node184;
	wire [46-1:0] node185;
	wire [46-1:0] node187;
	wire [46-1:0] node188;
	wire [46-1:0] node192;
	wire [46-1:0] node193;
	wire [46-1:0] node195;
	wire [46-1:0] node198;
	wire [46-1:0] node199;
	wire [46-1:0] node202;
	wire [46-1:0] node205;
	wire [46-1:0] node207;
	wire [46-1:0] node209;
	wire [46-1:0] node211;
	wire [46-1:0] node212;
	wire [46-1:0] node214;
	wire [46-1:0] node216;
	wire [46-1:0] node218;
	wire [46-1:0] node220;
	wire [46-1:0] node223;
	wire [46-1:0] node224;
	wire [46-1:0] node225;
	wire [46-1:0] node226;
	wire [46-1:0] node228;
	wire [46-1:0] node231;
	wire [46-1:0] node232;
	wire [46-1:0] node237;
	wire [46-1:0] node238;
	wire [46-1:0] node240;
	wire [46-1:0] node241;
	wire [46-1:0] node245;
	wire [46-1:0] node246;
	wire [46-1:0] node247;
	wire [46-1:0] node250;
	wire [46-1:0] node253;
	wire [46-1:0] node254;
	wire [46-1:0] node257;
	wire [46-1:0] node260;
	wire [46-1:0] node261;
	wire [46-1:0] node262;
	wire [46-1:0] node265;
	wire [46-1:0] node266;
	wire [46-1:0] node267;
	wire [46-1:0] node268;
	wire [46-1:0] node269;
	wire [46-1:0] node272;
	wire [46-1:0] node275;
	wire [46-1:0] node276;
	wire [46-1:0] node279;
	wire [46-1:0] node282;
	wire [46-1:0] node283;
	wire [46-1:0] node284;
	wire [46-1:0] node287;
	wire [46-1:0] node290;
	wire [46-1:0] node291;
	wire [46-1:0] node294;
	wire [46-1:0] node297;
	wire [46-1:0] node298;
	wire [46-1:0] node299;
	wire [46-1:0] node300;
	wire [46-1:0] node303;
	wire [46-1:0] node306;
	wire [46-1:0] node307;
	wire [46-1:0] node310;
	wire [46-1:0] node313;
	wire [46-1:0] node314;
	wire [46-1:0] node315;
	wire [46-1:0] node318;
	wire [46-1:0] node321;
	wire [46-1:0] node322;
	wire [46-1:0] node325;
	wire [46-1:0] node328;
	wire [46-1:0] node329;
	wire [46-1:0] node332;
	wire [46-1:0] node334;
	wire [46-1:0] node335;
	wire [46-1:0] node336;
	wire [46-1:0] node337;
	wire [46-1:0] node338;
	wire [46-1:0] node339;
	wire [46-1:0] node340;
	wire [46-1:0] node341;
	wire [46-1:0] node342;
	wire [46-1:0] node343;
	wire [46-1:0] node346;
	wire [46-1:0] node349;
	wire [46-1:0] node350;
	wire [46-1:0] node353;
	wire [46-1:0] node356;
	wire [46-1:0] node357;
	wire [46-1:0] node358;
	wire [46-1:0] node361;
	wire [46-1:0] node364;
	wire [46-1:0] node365;
	wire [46-1:0] node368;
	wire [46-1:0] node371;
	wire [46-1:0] node372;
	wire [46-1:0] node373;
	wire [46-1:0] node374;
	wire [46-1:0] node377;
	wire [46-1:0] node380;
	wire [46-1:0] node381;
	wire [46-1:0] node384;
	wire [46-1:0] node387;
	wire [46-1:0] node388;
	wire [46-1:0] node389;
	wire [46-1:0] node392;
	wire [46-1:0] node395;
	wire [46-1:0] node396;
	wire [46-1:0] node399;
	wire [46-1:0] node402;
	wire [46-1:0] node403;
	wire [46-1:0] node404;
	wire [46-1:0] node405;
	wire [46-1:0] node406;
	wire [46-1:0] node409;
	wire [46-1:0] node412;
	wire [46-1:0] node413;
	wire [46-1:0] node416;
	wire [46-1:0] node419;
	wire [46-1:0] node420;
	wire [46-1:0] node422;
	wire [46-1:0] node425;
	wire [46-1:0] node426;
	wire [46-1:0] node429;
	wire [46-1:0] node432;
	wire [46-1:0] node433;
	wire [46-1:0] node434;
	wire [46-1:0] node435;
	wire [46-1:0] node438;
	wire [46-1:0] node441;
	wire [46-1:0] node442;
	wire [46-1:0] node445;
	wire [46-1:0] node448;
	wire [46-1:0] node449;
	wire [46-1:0] node450;
	wire [46-1:0] node453;
	wire [46-1:0] node456;
	wire [46-1:0] node457;
	wire [46-1:0] node460;
	wire [46-1:0] node463;
	wire [46-1:0] node464;
	wire [46-1:0] node465;
	wire [46-1:0] node466;
	wire [46-1:0] node467;
	wire [46-1:0] node468;
	wire [46-1:0] node471;
	wire [46-1:0] node474;
	wire [46-1:0] node475;
	wire [46-1:0] node478;
	wire [46-1:0] node481;
	wire [46-1:0] node482;
	wire [46-1:0] node483;
	wire [46-1:0] node486;
	wire [46-1:0] node489;
	wire [46-1:0] node490;
	wire [46-1:0] node493;
	wire [46-1:0] node496;
	wire [46-1:0] node497;
	wire [46-1:0] node498;
	wire [46-1:0] node499;
	wire [46-1:0] node502;
	wire [46-1:0] node505;
	wire [46-1:0] node506;
	wire [46-1:0] node509;
	wire [46-1:0] node512;
	wire [46-1:0] node513;
	wire [46-1:0] node514;
	wire [46-1:0] node517;
	wire [46-1:0] node520;
	wire [46-1:0] node521;
	wire [46-1:0] node524;
	wire [46-1:0] node527;
	wire [46-1:0] node528;
	wire [46-1:0] node529;
	wire [46-1:0] node530;
	wire [46-1:0] node532;
	wire [46-1:0] node535;
	wire [46-1:0] node536;
	wire [46-1:0] node539;
	wire [46-1:0] node542;
	wire [46-1:0] node543;
	wire [46-1:0] node544;
	wire [46-1:0] node547;
	wire [46-1:0] node550;
	wire [46-1:0] node551;
	wire [46-1:0] node554;
	wire [46-1:0] node557;
	wire [46-1:0] node558;
	wire [46-1:0] node559;
	wire [46-1:0] node560;
	wire [46-1:0] node563;
	wire [46-1:0] node566;
	wire [46-1:0] node567;
	wire [46-1:0] node570;
	wire [46-1:0] node573;
	wire [46-1:0] node574;
	wire [46-1:0] node575;
	wire [46-1:0] node578;
	wire [46-1:0] node581;
	wire [46-1:0] node582;
	wire [46-1:0] node585;
	wire [46-1:0] node588;
	wire [46-1:0] node589;
	wire [46-1:0] node590;
	wire [46-1:0] node591;
	wire [46-1:0] node593;
	wire [46-1:0] node594;
	wire [46-1:0] node595;
	wire [46-1:0] node598;
	wire [46-1:0] node601;
	wire [46-1:0] node602;
	wire [46-1:0] node606;
	wire [46-1:0] node607;
	wire [46-1:0] node608;
	wire [46-1:0] node609;
	wire [46-1:0] node613;
	wire [46-1:0] node614;
	wire [46-1:0] node617;
	wire [46-1:0] node621;
	wire [46-1:0] node622;
	wire [46-1:0] node623;
	wire [46-1:0] node625;
	wire [46-1:0] node627;
	wire [46-1:0] node630;
	wire [46-1:0] node631;
	wire [46-1:0] node632;
	wire [46-1:0] node639;
	wire [46-1:0] node640;
	wire [46-1:0] node641;
	wire [46-1:0] node643;
	wire [46-1:0] node645;
	wire [46-1:0] node646;
	wire [46-1:0] node648;
	wire [46-1:0] node649;
	wire [46-1:0] node652;
	wire [46-1:0] node655;
	wire [46-1:0] node656;
	wire [46-1:0] node657;
	wire [46-1:0] node660;
	wire [46-1:0] node664;
	wire [46-1:0] node665;
	wire [46-1:0] node666;
	wire [46-1:0] node667;
	wire [46-1:0] node668;
	wire [46-1:0] node669;
	wire [46-1:0] node672;
	wire [46-1:0] node675;
	wire [46-1:0] node676;
	wire [46-1:0] node679;
	wire [46-1:0] node682;
	wire [46-1:0] node683;
	wire [46-1:0] node684;
	wire [46-1:0] node687;
	wire [46-1:0] node690;
	wire [46-1:0] node691;
	wire [46-1:0] node694;
	wire [46-1:0] node697;
	wire [46-1:0] node698;
	wire [46-1:0] node699;
	wire [46-1:0] node700;
	wire [46-1:0] node703;
	wire [46-1:0] node706;
	wire [46-1:0] node707;
	wire [46-1:0] node710;
	wire [46-1:0] node713;
	wire [46-1:0] node714;
	wire [46-1:0] node715;
	wire [46-1:0] node718;
	wire [46-1:0] node721;
	wire [46-1:0] node722;
	wire [46-1:0] node725;
	wire [46-1:0] node728;
	wire [46-1:0] node729;
	wire [46-1:0] node730;
	wire [46-1:0] node731;
	wire [46-1:0] node732;
	wire [46-1:0] node735;
	wire [46-1:0] node738;
	wire [46-1:0] node739;
	wire [46-1:0] node742;
	wire [46-1:0] node745;
	wire [46-1:0] node746;
	wire [46-1:0] node747;
	wire [46-1:0] node750;
	wire [46-1:0] node753;
	wire [46-1:0] node754;
	wire [46-1:0] node757;
	wire [46-1:0] node760;
	wire [46-1:0] node761;
	wire [46-1:0] node762;
	wire [46-1:0] node764;
	wire [46-1:0] node767;
	wire [46-1:0] node768;
	wire [46-1:0] node771;
	wire [46-1:0] node774;
	wire [46-1:0] node775;
	wire [46-1:0] node776;
	wire [46-1:0] node779;
	wire [46-1:0] node782;
	wire [46-1:0] node783;
	wire [46-1:0] node786;
	wire [46-1:0] node789;
	wire [46-1:0] node790;
	wire [46-1:0] node791;
	wire [46-1:0] node792;
	wire [46-1:0] node793;
	wire [46-1:0] node794;
	wire [46-1:0] node795;
	wire [46-1:0] node798;
	wire [46-1:0] node801;
	wire [46-1:0] node802;
	wire [46-1:0] node805;
	wire [46-1:0] node808;
	wire [46-1:0] node809;
	wire [46-1:0] node810;
	wire [46-1:0] node813;
	wire [46-1:0] node816;
	wire [46-1:0] node817;
	wire [46-1:0] node820;
	wire [46-1:0] node823;
	wire [46-1:0] node824;
	wire [46-1:0] node825;
	wire [46-1:0] node826;
	wire [46-1:0] node829;
	wire [46-1:0] node832;
	wire [46-1:0] node833;
	wire [46-1:0] node836;
	wire [46-1:0] node839;
	wire [46-1:0] node840;
	wire [46-1:0] node841;
	wire [46-1:0] node844;
	wire [46-1:0] node847;
	wire [46-1:0] node848;
	wire [46-1:0] node851;
	wire [46-1:0] node854;
	wire [46-1:0] node855;
	wire [46-1:0] node856;
	wire [46-1:0] node857;
	wire [46-1:0] node858;
	wire [46-1:0] node861;
	wire [46-1:0] node864;
	wire [46-1:0] node865;
	wire [46-1:0] node868;
	wire [46-1:0] node871;
	wire [46-1:0] node872;
	wire [46-1:0] node873;
	wire [46-1:0] node876;
	wire [46-1:0] node879;
	wire [46-1:0] node880;
	wire [46-1:0] node883;
	wire [46-1:0] node886;
	wire [46-1:0] node887;
	wire [46-1:0] node888;
	wire [46-1:0] node890;
	wire [46-1:0] node893;
	wire [46-1:0] node894;
	wire [46-1:0] node897;
	wire [46-1:0] node900;
	wire [46-1:0] node901;
	wire [46-1:0] node902;
	wire [46-1:0] node905;
	wire [46-1:0] node908;
	wire [46-1:0] node909;
	wire [46-1:0] node912;
	wire [46-1:0] node915;
	wire [46-1:0] node916;
	wire [46-1:0] node917;
	wire [46-1:0] node918;
	wire [46-1:0] node919;
	wire [46-1:0] node920;
	wire [46-1:0] node923;
	wire [46-1:0] node926;
	wire [46-1:0] node927;
	wire [46-1:0] node930;
	wire [46-1:0] node933;
	wire [46-1:0] node934;
	wire [46-1:0] node935;
	wire [46-1:0] node938;
	wire [46-1:0] node941;
	wire [46-1:0] node942;
	wire [46-1:0] node945;
	wire [46-1:0] node948;
	wire [46-1:0] node949;
	wire [46-1:0] node950;
	wire [46-1:0] node951;
	wire [46-1:0] node954;
	wire [46-1:0] node957;
	wire [46-1:0] node958;
	wire [46-1:0] node961;
	wire [46-1:0] node964;
	wire [46-1:0] node965;
	wire [46-1:0] node967;
	wire [46-1:0] node970;
	wire [46-1:0] node971;
	wire [46-1:0] node974;
	wire [46-1:0] node977;
	wire [46-1:0] node978;
	wire [46-1:0] node979;
	wire [46-1:0] node980;
	wire [46-1:0] node981;
	wire [46-1:0] node984;
	wire [46-1:0] node987;
	wire [46-1:0] node988;
	wire [46-1:0] node991;
	wire [46-1:0] node994;
	wire [46-1:0] node995;
	wire [46-1:0] node996;
	wire [46-1:0] node999;
	wire [46-1:0] node1002;
	wire [46-1:0] node1003;
	wire [46-1:0] node1006;
	wire [46-1:0] node1009;
	wire [46-1:0] node1010;
	wire [46-1:0] node1011;
	wire [46-1:0] node1012;
	wire [46-1:0] node1015;
	wire [46-1:0] node1018;
	wire [46-1:0] node1019;
	wire [46-1:0] node1022;
	wire [46-1:0] node1025;
	wire [46-1:0] node1026;
	wire [46-1:0] node1027;
	wire [46-1:0] node1030;
	wire [46-1:0] node1033;
	wire [46-1:0] node1034;
	wire [46-1:0] node1037;
	wire [46-1:0] node1040;
	wire [46-1:0] node1041;
	wire [46-1:0] node1042;
	wire [46-1:0] node1043;
	wire [46-1:0] node1045;
	wire [46-1:0] node1047;
	wire [46-1:0] node1049;
	wire [46-1:0] node1051;
	wire [46-1:0] node1052;
	wire [46-1:0] node1055;
	wire [46-1:0] node1058;
	wire [46-1:0] node1059;
	wire [46-1:0] node1061;
	wire [46-1:0] node1063;
	wire [46-1:0] node1065;
	wire [46-1:0] node1066;
	wire [46-1:0] node1069;
	wire [46-1:0] node1072;
	wire [46-1:0] node1073;
	wire [46-1:0] node1074;
	wire [46-1:0] node1075;
	wire [46-1:0] node1076;
	wire [46-1:0] node1079;
	wire [46-1:0] node1082;
	wire [46-1:0] node1083;
	wire [46-1:0] node1086;
	wire [46-1:0] node1089;
	wire [46-1:0] node1090;
	wire [46-1:0] node1091;
	wire [46-1:0] node1094;
	wire [46-1:0] node1097;
	wire [46-1:0] node1098;
	wire [46-1:0] node1101;
	wire [46-1:0] node1104;
	wire [46-1:0] node1105;
	wire [46-1:0] node1106;
	wire [46-1:0] node1108;
	wire [46-1:0] node1111;
	wire [46-1:0] node1112;
	wire [46-1:0] node1116;
	wire [46-1:0] node1117;
	wire [46-1:0] node1119;
	wire [46-1:0] node1122;
	wire [46-1:0] node1123;
	wire [46-1:0] node1127;
	wire [46-1:0] node1128;
	wire [46-1:0] node1129;
	wire [46-1:0] node1130;
	wire [46-1:0] node1131;
	wire [46-1:0] node1132;
	wire [46-1:0] node1133;
	wire [46-1:0] node1136;
	wire [46-1:0] node1139;
	wire [46-1:0] node1140;
	wire [46-1:0] node1143;
	wire [46-1:0] node1146;
	wire [46-1:0] node1147;
	wire [46-1:0] node1148;
	wire [46-1:0] node1151;
	wire [46-1:0] node1154;
	wire [46-1:0] node1155;
	wire [46-1:0] node1158;
	wire [46-1:0] node1161;
	wire [46-1:0] node1162;
	wire [46-1:0] node1163;
	wire [46-1:0] node1164;
	wire [46-1:0] node1167;
	wire [46-1:0] node1170;
	wire [46-1:0] node1171;
	wire [46-1:0] node1174;
	wire [46-1:0] node1177;
	wire [46-1:0] node1178;
	wire [46-1:0] node1180;
	wire [46-1:0] node1183;
	wire [46-1:0] node1184;
	wire [46-1:0] node1187;
	wire [46-1:0] node1190;
	wire [46-1:0] node1191;
	wire [46-1:0] node1192;
	wire [46-1:0] node1193;
	wire [46-1:0] node1194;
	wire [46-1:0] node1197;
	wire [46-1:0] node1200;
	wire [46-1:0] node1201;
	wire [46-1:0] node1204;
	wire [46-1:0] node1207;
	wire [46-1:0] node1208;
	wire [46-1:0] node1209;
	wire [46-1:0] node1212;
	wire [46-1:0] node1215;
	wire [46-1:0] node1216;
	wire [46-1:0] node1219;
	wire [46-1:0] node1222;
	wire [46-1:0] node1223;
	wire [46-1:0] node1224;
	wire [46-1:0] node1225;
	wire [46-1:0] node1228;
	wire [46-1:0] node1231;
	wire [46-1:0] node1232;
	wire [46-1:0] node1235;
	wire [46-1:0] node1238;
	wire [46-1:0] node1239;
	wire [46-1:0] node1240;
	wire [46-1:0] node1243;
	wire [46-1:0] node1246;
	wire [46-1:0] node1247;
	wire [46-1:0] node1250;
	wire [46-1:0] node1253;
	wire [46-1:0] node1254;
	wire [46-1:0] node1255;
	wire [46-1:0] node1256;
	wire [46-1:0] node1257;
	wire [46-1:0] node1258;
	wire [46-1:0] node1261;
	wire [46-1:0] node1264;
	wire [46-1:0] node1265;
	wire [46-1:0] node1268;
	wire [46-1:0] node1271;
	wire [46-1:0] node1272;
	wire [46-1:0] node1273;
	wire [46-1:0] node1277;
	wire [46-1:0] node1278;
	wire [46-1:0] node1281;
	wire [46-1:0] node1284;
	wire [46-1:0] node1285;
	wire [46-1:0] node1286;
	wire [46-1:0] node1287;
	wire [46-1:0] node1290;
	wire [46-1:0] node1293;
	wire [46-1:0] node1294;
	wire [46-1:0] node1297;
	wire [46-1:0] node1300;
	wire [46-1:0] node1301;
	wire [46-1:0] node1302;
	wire [46-1:0] node1305;
	wire [46-1:0] node1308;
	wire [46-1:0] node1309;
	wire [46-1:0] node1312;
	wire [46-1:0] node1315;
	wire [46-1:0] node1316;
	wire [46-1:0] node1317;
	wire [46-1:0] node1318;
	wire [46-1:0] node1319;
	wire [46-1:0] node1322;
	wire [46-1:0] node1325;
	wire [46-1:0] node1326;
	wire [46-1:0] node1329;
	wire [46-1:0] node1332;
	wire [46-1:0] node1333;
	wire [46-1:0] node1334;
	wire [46-1:0] node1337;
	wire [46-1:0] node1340;
	wire [46-1:0] node1341;
	wire [46-1:0] node1344;
	wire [46-1:0] node1347;
	wire [46-1:0] node1348;
	wire [46-1:0] node1349;
	wire [46-1:0] node1350;
	wire [46-1:0] node1353;
	wire [46-1:0] node1356;
	wire [46-1:0] node1357;
	wire [46-1:0] node1360;
	wire [46-1:0] node1363;
	wire [46-1:0] node1364;
	wire [46-1:0] node1365;
	wire [46-1:0] node1368;
	wire [46-1:0] node1371;
	wire [46-1:0] node1372;
	wire [46-1:0] node1375;
	wire [46-1:0] node1378;
	wire [46-1:0] node1379;
	wire [46-1:0] node1380;
	wire [46-1:0] node1381;
	wire [46-1:0] node1382;
	wire [46-1:0] node1383;
	wire [46-1:0] node1386;
	wire [46-1:0] node1391;
	wire [46-1:0] node1392;
	wire [46-1:0] node1393;
	wire [46-1:0] node1394;
	wire [46-1:0] node1397;
	wire [46-1:0] node1400;
	wire [46-1:0] node1401;
	wire [46-1:0] node1404;
	wire [46-1:0] node1407;
	wire [46-1:0] node1408;
	wire [46-1:0] node1409;
	wire [46-1:0] node1412;
	wire [46-1:0] node1416;
	wire [46-1:0] node1417;
	wire [46-1:0] node1418;
	wire [46-1:0] node1419;
	wire [46-1:0] node1420;
	wire [46-1:0] node1423;
	wire [46-1:0] node1426;
	wire [46-1:0] node1427;
	wire [46-1:0] node1430;
	wire [46-1:0] node1433;
	wire [46-1:0] node1434;
	wire [46-1:0] node1435;
	wire [46-1:0] node1438;
	wire [46-1:0] node1442;
	wire [46-1:0] node1443;
	wire [46-1:0] node1444;
	wire [46-1:0] node1445;
	wire [46-1:0] node1448;

	assign outp = (inp[1]) ? node260 : node1;
		assign node1 = (inp[3]) ? node5 : node2;
			assign node2 = (inp[15]) ? 46'b0000000000000000000000000000001000000000000000 : 46'b0000000000000000000000000000000000000000000000;
			assign node5 = (inp[15]) ? node69 : node6;
				assign node6 = (inp[13]) ? node36 : node7;
					assign node7 = (inp[10]) ? node9 : 46'b0000000000000000000000000000000000000000000000;
						assign node9 = (inp[5]) ? node11 : 46'b0000000000000000000000000000000000000000000000;
							assign node11 = (inp[8]) ? node13 : 46'b0000000000000000000000000000000000000000000000;
								assign node13 = (inp[7]) ? node15 : 46'b0000000000000000000000000000000000000000000000;
									assign node15 = (inp[14]) ? node17 : 46'b0000000000000000000000000000000000000000000000;
										assign node17 = (inp[2]) ? node27 : node18;
											assign node18 = (inp[4]) ? node20 : 46'b0000000000000000000000000000000000000000000000;
												assign node20 = (inp[9]) ? node22 : 46'b0000000000000000000000000000000000000000000000;
													assign node22 = (inp[0]) ? node24 : 46'b0000000000000000000000000000000000000000000000;
														assign node24 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
											assign node27 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : node28;
												assign node28 = (inp[9]) ? node30 : 46'b0000000000000000000000000000000000000000000000;
													assign node30 = (inp[0]) ? node32 : 46'b0000000000000000000000000000000000000000000000;
														assign node32 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000001 : 46'b0000000000000000000000000000000000000000000000;
					assign node36 = (inp[12]) ? node38 : 46'b0000000000000000000000000000000000000000000000;
						assign node38 = (inp[0]) ? node52 : node39;
							assign node39 = (inp[5]) ? node41 : 46'b0000000000000000000000000000000000000000000000;
								assign node41 = (inp[6]) ? node43 : 46'b0000000000000000000000000000000000000000000000;
									assign node43 = (inp[7]) ? node45 : 46'b0000000000000000000000000000000000000000000000;
										assign node45 = (inp[2]) ? node47 : 46'b0000000000000000000000000000000000000000000000;
											assign node47 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : node48;
												assign node48 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000100000000;
							assign node52 = (inp[10]) ? node54 : 46'b0000000000000000000000000000000000000000000000;
								assign node54 = (inp[7]) ? node56 : 46'b0000000000000000000000000000000000000000000000;
									assign node56 = (inp[6]) ? node58 : 46'b0000000000000000000000000000000000000000000000;
										assign node58 = (inp[14]) ? node60 : 46'b0000000000000000000000000000000000000000000000;
											assign node60 = (inp[4]) ? node62 : 46'b0000000000000000000000000000000000000000000000;
												assign node62 = (inp[8]) ? node64 : 46'b0000000000000000000000000000000000000000000000;
													assign node64 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : node65;
														assign node65 = (inp[5]) ? 46'b0000000001000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
				assign node69 = (inp[9]) ? node123 : node70;
					assign node70 = (inp[11]) ? node110 : node71;
						assign node71 = (inp[13]) ? node77 : node72;
							assign node72 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node73;
								assign node73 = (inp[0]) ? 46'b0000000000001000000000000010000000000000000000 : 46'b0000001000001000000000000000000000000000000000;
							assign node77 = (inp[5]) ? node79 : 46'b0000000000000000000000000000000000000000000000;
								assign node79 = (inp[14]) ? node81 : 46'b0000000000000000000000000000000000000000000000;
									assign node81 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node82;
										assign node82 = (inp[6]) ? node84 : 46'b0000000000000000000000000000000000000000000000;
											assign node84 = (inp[2]) ? node96 : node85;
												assign node85 = (inp[12]) ? node91 : node86;
													assign node86 = (inp[7]) ? node88 : 46'b0000000000000000000000000000000000000000000000;
														assign node88 = (inp[10]) ? 46'b0000000000001000010100000000000000000000010000 : 46'b0000000000000000000000000000000000000000000000;
													assign node91 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node92;
														assign node92 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
												assign node96 = (inp[10]) ? node102 : node97;
													assign node97 = (inp[8]) ? node99 : 46'b0000000000000000000000000000000000000000000000;
														assign node99 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
													assign node102 = (inp[12]) ? node106 : node103;
														assign node103 = (inp[7]) ? 46'b0000000000001000010000000000000001000010000000 : 46'b0000000000000000000000000000000000000000000000;
														assign node106 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
						assign node110 = (inp[13]) ? node116 : node111;
							assign node111 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node112;
								assign node112 = (inp[0]) ? 46'b0000010000000000000000000010000000000000000000 : 46'b0000011000000000000000000000000000000000000000;
							assign node116 = (inp[2]) ? node120 : node117;
								assign node117 = (inp[0]) ? 46'b0000001000000000011000000100000000000000010000 : 46'b0000001000000000010000000100000000000000010010;
								assign node120 = (inp[0]) ? 46'b0000001000000000010010000000010000000010000000 : 46'b0000001000000000010010100000000000000010000000;
					assign node123 = (inp[2]) ? node205 : node124;
						assign node124 = (inp[0]) ? node162 : node125;
							assign node125 = (inp[13]) ? node129 : node126;
								assign node126 = (inp[11]) ? 46'b0000010100000000000000000000000000000000000000 : 46'b0000000100001000000000000000000000000000000000;
								assign node129 = (inp[5]) ? node131 : 46'b0000000000000000000000000000000000000000000000;
									assign node131 = (inp[14]) ? node133 : 46'b0000000000000000000000000000000000000000000000;
										assign node133 = (inp[6]) ? node143 : node134;
											assign node134 = (inp[7]) ? node136 : 46'b0000000000000000000000000000000000000000000000;
												assign node136 = (inp[8]) ? node138 : 46'b0000000000000000000000000000000000000000000000;
													assign node138 = (inp[11]) ? node140 : 46'b0000000000000000000000000000000000000000000000;
														assign node140 = (inp[4]) ? 46'b0000000000000000000000000100000000000000000010 : 46'b0000000000000000000000000000000000000000000000;
											assign node143 = (inp[10]) ? node151 : node144;
												assign node144 = (inp[8]) ? node146 : 46'b0000000000000000000000000000000000000000000000;
													assign node146 = (inp[4]) ? node148 : 46'b0000000000000000000000000000000000000000000000;
														assign node148 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000010000000000010000000100000100000000010010;
												assign node151 = (inp[8]) ? node157 : node152;
													assign node152 = (inp[4]) ? node154 : 46'b0000000000000000000000000000000000000000000000;
														assign node154 = (inp[11]) ? 46'b0010000000010000000000000100000000000000010010 : 46'b0000000000010000010000000000000000000000010000;
													assign node157 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : node158;
														assign node158 = (inp[11]) ? 46'b0000000000000000010000010100000000000000010010 : 46'b0000000000000000000000010000000000000000010000;
							assign node162 = (inp[11]) ? node178 : node163;
								assign node163 = (inp[13]) ? node165 : 46'b0010001000000000000000000000000000000000010000;
									assign node165 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node166;
										assign node166 = (inp[6]) ? node168 : 46'b0000000000000000000000000000000000000000000000;
											assign node168 = (inp[10]) ? node170 : 46'b0000000000000000000000000000000000000000000000;
												assign node170 = (inp[5]) ? node172 : 46'b0000000000000000000000000000000000000000000000;
													assign node172 = (inp[14]) ? node174 : 46'b0000000000000000000000000000000000000000000000;
														assign node174 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
								assign node178 = (inp[5]) ? node180 : 46'b0000000000000000000000000000000000000000000000;
									assign node180 = (inp[14]) ? node182 : 46'b0000000000000000000000000000000000000000000000;
										assign node182 = (inp[13]) ? node184 : 46'b0000000000000000000000000000000000000000000000;
											assign node184 = (inp[4]) ? node192 : node185;
												assign node185 = (inp[10]) ? node187 : 46'b0000000000000000000000000000000000000000000000;
													assign node187 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node188;
														assign node188 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
												assign node192 = (inp[6]) ? node198 : node193;
													assign node193 = (inp[8]) ? node195 : 46'b0000000000000000000000000000000000000000000000;
														assign node195 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000001000000100000000000000000000;
													assign node198 = (inp[8]) ? node202 : node199;
														assign node199 = (inp[10]) ? 46'b0000000000010000011000000100000000000000010000 : 46'b0000000000000000000000000000000000000000000000;
														assign node202 = (inp[10]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000001000000100000100000000010000;
						assign node205 = (inp[5]) ? node207 : 46'b0000000000000000000000000000000000000000000000;
							assign node207 = (inp[13]) ? node209 : 46'b0000000000000000000000000000000000000000000000;
								assign node209 = (inp[14]) ? node211 : 46'b0000000000000000000000000000000000000000000000;
									assign node211 = (inp[6]) ? node223 : node212;
										assign node212 = (inp[11]) ? node214 : 46'b0000000000000000000000000000000000000000000000;
											assign node214 = (inp[8]) ? node216 : 46'b0000000000000000000000000000000000000000000000;
												assign node216 = (inp[4]) ? node218 : 46'b0000000000000000000000000000000000000000000000;
													assign node218 = (inp[10]) ? node220 : 46'b0000000000000000000000000000000000000000000000;
														assign node220 = (inp[7]) ? 46'b0000000000000000000010000000000000000000000100 : 46'b0000000000000000000110000000000000000000000000;
										assign node223 = (inp[11]) ? node237 : node224;
											assign node224 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node225;
												assign node225 = (inp[12]) ? node231 : node226;
													assign node226 = (inp[8]) ? node228 : 46'b0000000000011000010000000000000000000010000000;
														assign node228 = (inp[4]) ? 46'b0000000000000000000000000000000100000010000000 : 46'b0000000000000000000000000000000000000000000000;
													assign node231 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node232;
														assign node232 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000010000000000010000010000000000000010000000;
											assign node237 = (inp[8]) ? node245 : node238;
												assign node238 = (inp[4]) ? node240 : 46'b0000000000000000000000000000000000000000000000;
													assign node240 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node241;
														assign node241 = (inp[10]) ? 46'b0000000000011000010010100000000000000010000000 : 46'b0000000000000000000000000000000000000000000000;
												assign node245 = (inp[0]) ? node253 : node246;
													assign node246 = (inp[10]) ? node250 : node247;
														assign node247 = (inp[4]) ? 46'b0000000000000000010010100000000100000010000000 : 46'b0000000000000000000000000000000000000000000000;
														assign node250 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000010110000000000000010000000;
													assign node253 = (inp[4]) ? node257 : node254;
														assign node254 = (inp[12]) ? 46'b0000010000000000010010010000010000000010000000 : 46'b0010000000000000000010010000010000000010000000;
														assign node257 = (inp[10]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0010000000000000000010000000010100000010000000;
		assign node260 = (inp[15]) ? node328 : node261;
			assign node261 = (inp[13]) ? node265 : node262;
				assign node262 = (inp[3]) ? 46'b0000100000000000000000000000001000000000000000 : 46'b0000100000000000000000000000000000000000000000;
				assign node265 = (inp[2]) ? node297 : node266;
					assign node266 = (inp[11]) ? node282 : node267;
						assign node267 = (inp[9]) ? node275 : node268;
							assign node268 = (inp[0]) ? node272 : node269;
								assign node269 = (inp[3]) ? 46'b0000100000001000010000010100001000000000010010 : 46'b0000100000001000010000010100000000000000010010;
								assign node272 = (inp[3]) ? 46'b0000100000001000010000000100001100000000010010 : 46'b0000100000001000010000000100000100000000010010;
							assign node275 = (inp[0]) ? node279 : node276;
								assign node276 = (inp[3]) ? 46'b0000110000000000010000010100001000000000010010 : 46'b0000110000000000010000010100000000000000010010;
								assign node279 = (inp[3]) ? 46'b0000110000000000010000000100001100000000010010 : 46'b0000110000000000010000000100000100000000010010;
						assign node282 = (inp[0]) ? node290 : node283;
							assign node283 = (inp[9]) ? node287 : node284;
								assign node284 = (inp[3]) ? 46'b0000100000001000011000010100001000000000010000 : 46'b0000100000001000011000010100000000000000010000;
								assign node287 = (inp[3]) ? 46'b0000110000000000011000010100001000000000010000 : 46'b0000110000000000011000010100000000000000010000;
							assign node290 = (inp[9]) ? node294 : node291;
								assign node291 = (inp[3]) ? 46'b0000100000001000011000000100001100000000010000 : 46'b0000100000001000011000000100000100000000010000;
								assign node294 = (inp[3]) ? 46'b0000110000000000011000000100001100000000010000 : 46'b0000110000000000011000000100000100000000010000;
					assign node297 = (inp[9]) ? node313 : node298;
						assign node298 = (inp[0]) ? node306 : node299;
							assign node299 = (inp[11]) ? node303 : node300;
								assign node300 = (inp[3]) ? 46'b0000100000001000010010110000001000000010000000 : 46'b0000100000001000010010110000000000000010000000;
								assign node303 = (inp[3]) ? 46'b0000100000001000010010010000011000000010000000 : 46'b0000100000001000010010010000010000000010000000;
							assign node306 = (inp[11]) ? node310 : node307;
								assign node307 = (inp[3]) ? 46'b0000100000001000010010100000001100000010000000 : 46'b0000100000001000010010100000000100000010000000;
								assign node310 = (inp[3]) ? 46'b0000100000001000010010000000011100000010000000 : 46'b0000100000001000010010000000010100000010000000;
						assign node313 = (inp[11]) ? node321 : node314;
							assign node314 = (inp[0]) ? node318 : node315;
								assign node315 = (inp[3]) ? 46'b0000110000000000010010110000001000000010000000 : 46'b0000110000000000010010110000000000000010000000;
								assign node318 = (inp[3]) ? 46'b0000110000000000010010100000001100000010000000 : 46'b0000110000000000010010100000000100000010000000;
							assign node321 = (inp[0]) ? node325 : node322;
								assign node322 = (inp[3]) ? 46'b0000110000000000010010010000011000000010000000 : 46'b0000110000000000010010010000010000000010000000;
								assign node325 = (inp[3]) ? 46'b0000110000000000010010000000011100000010000000 : 46'b0000110000000000010010000000010100000010000000;
			assign node328 = (inp[13]) ? node332 : node329;
				assign node329 = (inp[3]) ? 46'b0000000000000000000000000000000000000000001000 : 46'b0000000000000000000000000000001000000000001000;
				assign node332 = (inp[3]) ? node334 : 46'b0000000000000000000000000000001000000000000000;
					assign node334 = (inp[2]) ? node1040 : node335;
						assign node335 = (inp[11]) ? node639 : node336;
							assign node336 = (inp[9]) ? node588 : node337;
								assign node337 = (inp[6]) ? node463 : node338;
									assign node338 = (inp[0]) ? node402 : node339;
										assign node339 = (inp[5]) ? node371 : node340;
											assign node340 = (inp[4]) ? node356 : node341;
												assign node341 = (inp[10]) ? node349 : node342;
													assign node342 = (inp[12]) ? node346 : node343;
														assign node343 = (inp[7]) ? 46'b0011000000000100000000010000000010110001010000 : 46'b0011000000000100000000010000100010110001010000;
														assign node346 = (inp[14]) ? 46'b0011000000000110000000010000100000110001010000 : 46'b0011000000000100000000010001000000110001010010;
													assign node349 = (inp[14]) ? node353 : node350;
														assign node350 = (inp[8]) ? 46'b0011000000000000000000010001000000110001010010 : 46'b0011000000000100000000010001100010110001010010;
														assign node353 = (inp[7]) ? 46'b0011000000000000001000010001000010110001010010 : 46'b0011000000000000001000010001100000110001010010;
												assign node356 = (inp[7]) ? node364 : node357;
													assign node357 = (inp[10]) ? node361 : node358;
														assign node358 = (inp[12]) ? 46'b0011000000000000001000010001100000110001010000 : 46'b0011000000000000001000010001100010110001010000;
														assign node361 = (inp[14]) ? 46'b0011000000000010001000010001100000110001010000 : 46'b0011000000000110000000010000100000110001010000;
													assign node364 = (inp[12]) ? node368 : node365;
														assign node365 = (inp[14]) ? 46'b0011000000000010001000010001000010110001010000 : 46'b0011000000000110000000010000000010110001010000;
														assign node368 = (inp[14]) ? 46'b0011000000000010001000010001000000110001010000 : 46'b0011000000000000001000010001000000110001010000;
											assign node371 = (inp[4]) ? node387 : node372;
												assign node372 = (inp[12]) ? node380 : node373;
													assign node373 = (inp[7]) ? node377 : node374;
														assign node374 = (inp[14]) ? 46'b0010000000000000001000010001100010110001010010 : 46'b0010000000000100000000010001100010110001010010;
														assign node377 = (inp[10]) ? 46'b0010000000000000000000010001000010110001010010 : 46'b0010000000000100000000010001000010110001010010;
													assign node380 = (inp[14]) ? node384 : node381;
														assign node381 = (inp[7]) ? 46'b0010000000000100000000010001000000110001010010 : 46'b0010000000000100000000010001100000110001010010;
														assign node384 = (inp[10]) ? 46'b0010000000000010000000010001000000110001010010 : 46'b0010000000000100000000010000000000110001010000;
												assign node387 = (inp[10]) ? node395 : node388;
													assign node388 = (inp[7]) ? node392 : node389;
														assign node389 = (inp[14]) ? 46'b0010000000000000001000010001100000110001010000 : 46'b0010000000000100001000010001100000110001010000;
														assign node392 = (inp[12]) ? 46'b0010000000000000001000010001000000110001010000 : 46'b0010000000000000001000010001000010110001010000;
													assign node395 = (inp[12]) ? node399 : node396;
														assign node396 = (inp[14]) ? 46'b0010000000000010000000010000100010110001010000 : 46'b0010000000000010000000010001000010110001010010;
														assign node399 = (inp[7]) ? 46'b0010000000000010000000010000000000110001010000 : 46'b0010000000000010000000010000100000110001010000;
										assign node402 = (inp[12]) ? node432 : node403;
											assign node403 = (inp[5]) ? node419 : node404;
												assign node404 = (inp[10]) ? node412 : node405;
													assign node405 = (inp[7]) ? node409 : node406;
														assign node406 = (inp[8]) ? 46'b0011000000000000000000010001100010110000010010 : 46'b0011000000000100001000010001100010110000010000;
														assign node409 = (inp[8]) ? 46'b0011000000000100000000010000000010110000010000 : 46'b0011000000000100001000010001000010110000010000;
													assign node412 = (inp[4]) ? node416 : node413;
														assign node413 = (inp[8]) ? 46'b0011000000000010000000010001000010110000010010 : 46'b0011000000000000001000010001000010110000010010;
														assign node416 = (inp[7]) ? 46'b0011000000000010001000010001000010110000010000 : 46'b0011000000000010001000010001100010110000010000;
												assign node419 = (inp[4]) ? node425 : node420;
													assign node420 = (inp[7]) ? node422 : 46'b0010000000000100000000010001100010110000010010;
														assign node422 = (inp[10]) ? 46'b0010000000000000000000010001000010110000010010 : 46'b0010000000000100000000010000000010110000010000;
													assign node425 = (inp[7]) ? node429 : node426;
														assign node426 = (inp[10]) ? 46'b0010000000000010000000010000100010110000010000 : 46'b0010000000000000001000010001100010110000010000;
														assign node429 = (inp[8]) ? 46'b0010000000000000001000010001000010110000010010 : 46'b0010000000000000001000010001000010110000010000;
											assign node432 = (inp[7]) ? node448 : node433;
												assign node433 = (inp[5]) ? node441 : node434;
													assign node434 = (inp[8]) ? node438 : node435;
														assign node435 = (inp[10]) ? 46'b0011000000000010000000010000100000110000010000 : 46'b0011000000000100001000010001100000110000010000;
														assign node438 = (inp[14]) ? 46'b0011000000000110000000010000100000110000010000 : 46'b0011000000000000000000010001100000110000010010;
													assign node441 = (inp[10]) ? node445 : node442;
														assign node442 = (inp[4]) ? 46'b0010000000000000001000010001100000110000010000 : 46'b0010000000000100000000010000100000110000010000;
														assign node445 = (inp[4]) ? 46'b0010000000000010000000010000100000110000010000 : 46'b0010000000000000001000010001100000110000010010;
												assign node448 = (inp[5]) ? node456 : node449;
													assign node449 = (inp[14]) ? node453 : node450;
														assign node450 = (inp[4]) ? 46'b0011000000000000001000010001000000110000010010 : 46'b0011000000000100000000010001000000110000010010;
														assign node453 = (inp[10]) ? 46'b0011000000000010000000010000000000110000010000 : 46'b0011000000000100001000010001000000110000010000;
													assign node456 = (inp[10]) ? node460 : node457;
														assign node457 = (inp[8]) ? 46'b0010000000000010001000010001000000110000010000 : 46'b0010000000000100001000010001000000110000010000;
														assign node460 = (inp[4]) ? 46'b0010000000000110000000010000000000110000010000 : 46'b0010000000000000000000010001000000110000010010;
									assign node463 = (inp[7]) ? node527 : node464;
										assign node464 = (inp[12]) ? node496 : node465;
											assign node465 = (inp[5]) ? node481 : node466;
												assign node466 = (inp[0]) ? node474 : node467;
													assign node467 = (inp[8]) ? node471 : node468;
														assign node468 = (inp[10]) ? 46'b0011000000000000001000010001100010010001010010 : 46'b0011000000000100001000010001100010010001010000;
														assign node471 = (inp[14]) ? 46'b0011000000000010000000010000100010010001010000 : 46'b0011000000000000000000010001100010010001010010;
													assign node474 = (inp[8]) ? node478 : node475;
														assign node475 = (inp[14]) ? 46'b0011000000000000001000010001100010010000010000 : 46'b0011000000000110000000010000100010010000010000;
														assign node478 = (inp[10]) ? 46'b0011000000000010000000010001100010010000010010 : 46'b0011000000000010001000010001100010010000010000;
												assign node481 = (inp[14]) ? node489 : node482;
													assign node482 = (inp[10]) ? node486 : node483;
														assign node483 = (inp[4]) ? 46'b0010000000000100001000010001100010010000010000 : 46'b0010000000000100000000010000100010010000010000;
														assign node486 = (inp[8]) ? 46'b0010000000000000000000010001100010010000010010 : 46'b0010000000000100000000010001100010010000010010;
													assign node489 = (inp[8]) ? node493 : node490;
														assign node490 = (inp[10]) ? 46'b0010000000000000001000010001100010010001010010 : 46'b0010000000000100001000010001100010010001010000;
														assign node493 = (inp[0]) ? 46'b0010000000000010000000010000100010010000010000 : 46'b0010000000000010000000010000100010010001010000;
											assign node496 = (inp[5]) ? node512 : node497;
												assign node497 = (inp[14]) ? node505 : node498;
													assign node498 = (inp[8]) ? node502 : node499;
														assign node499 = (inp[0]) ? 46'b0011000000000100000000010000100000010000010000 : 46'b0011000000000100000000010000100000010001010000;
														assign node502 = (inp[4]) ? 46'b0011000000000000001000010001100000010000010010 : 46'b0011000000000000000000010001100000010000010010;
													assign node505 = (inp[4]) ? node509 : node506;
														assign node506 = (inp[10]) ? 46'b0011000000000010000000010001100000010001010010 : 46'b0011000000000110000000010000100000010001010000;
														assign node509 = (inp[0]) ? 46'b0011000000000010001000010001100000010000010000 : 46'b0011000000000010001000010001100000010001010000;
												assign node512 = (inp[0]) ? node520 : node513;
													assign node513 = (inp[4]) ? node517 : node514;
														assign node514 = (inp[8]) ? 46'b0010000000000000000000010001100000010001010010 : 46'b0010000000000100000000010000100000010001010000;
														assign node517 = (inp[14]) ? 46'b0010000000000010000000010000100000010001010000 : 46'b0010000000000110000000010000100000010001010000;
													assign node520 = (inp[4]) ? node524 : node521;
														assign node521 = (inp[10]) ? 46'b0010000000000000000000010001100000010000010010 : 46'b0010000000000110000000010000100000010000010000;
														assign node524 = (inp[14]) ? 46'b0010000000000010001000010001100000010000010000 : 46'b0010000000000010000000010000100000010000010000;
										assign node527 = (inp[5]) ? node557 : node528;
											assign node528 = (inp[12]) ? node542 : node529;
												assign node529 = (inp[0]) ? node535 : node530;
													assign node530 = (inp[14]) ? node532 : 46'b0011000000000000001000010001000010010001010010;
														assign node532 = (inp[8]) ? 46'b0011000000000010000000010000000010010001010000 : 46'b0011000000000000001000010001000010010001010000;
													assign node535 = (inp[10]) ? node539 : node536;
														assign node536 = (inp[14]) ? 46'b0011000000000100000000010000000010010000010000 : 46'b0011000000000100000000010001000010010000010010;
														assign node539 = (inp[4]) ? 46'b0011000000000010001000010001000010010000010000 : 46'b0011000000000000000000010001000010010000010010;
												assign node542 = (inp[0]) ? node550 : node543;
													assign node543 = (inp[8]) ? node547 : node544;
														assign node544 = (inp[14]) ? 46'b0011000000000010001000010001000000010001010000 : 46'b0011000000000100001000010001000000010001010000;
														assign node547 = (inp[10]) ? 46'b0011000000000010000000010001000000010001010010 : 46'b0011000000000000001000010001000000010001010010;
													assign node550 = (inp[4]) ? node554 : node551;
														assign node551 = (inp[8]) ? 46'b0011000000000000000000010001000000010000010010 : 46'b0011000000000000001000010001000000010000010000;
														assign node554 = (inp[10]) ? 46'b0011000000000010000000010000000000010000010000 : 46'b0011000000000000001000010001000000010000010000;
											assign node557 = (inp[12]) ? node573 : node558;
												assign node558 = (inp[4]) ? node566 : node559;
													assign node559 = (inp[0]) ? node563 : node560;
														assign node560 = (inp[14]) ? 46'b0010000000000000000000010001000010010001010010 : 46'b0010000000000100000000010001000010010001010010;
														assign node563 = (inp[14]) ? 46'b0010000000000110000000010000000010010000010000 : 46'b0010000000000000000000010001000010010000010010;
													assign node566 = (inp[10]) ? node570 : node567;
														assign node567 = (inp[8]) ? 46'b0010000000000000001000010001000010010001010000 : 46'b0010000000000000001000010001000010010000010000;
														assign node570 = (inp[14]) ? 46'b0010000000000010000000010000000010010001010000 : 46'b0010000000000110000000010000000010010001010000;
												assign node573 = (inp[0]) ? node581 : node574;
													assign node574 = (inp[4]) ? node578 : node575;
														assign node575 = (inp[10]) ? 46'b0010000000000000000000010001000000010001010010 : 46'b0010000000000110000000010000000000010001010000;
														assign node578 = (inp[10]) ? 46'b0010000000000010000000010000000000010001010000 : 46'b0010000000000000001000010001000000010001010000;
													assign node581 = (inp[8]) ? node585 : node582;
														assign node582 = (inp[4]) ? 46'b0010000000000100000000010000000000010000010000 : 46'b0010000000000100000000010000000000010000010000;
														assign node585 = (inp[10]) ? 46'b0010000000000010000000010000000000010000010000 : 46'b0010000000000010001000010001000000010000010000;
								assign node588 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node589;
									assign node589 = (inp[4]) ? node621 : node590;
										assign node590 = (inp[5]) ? node606 : node591;
											assign node591 = (inp[7]) ? node593 : 46'b0000000000000000000000000000000000000000000000;
												assign node593 = (inp[10]) ? node601 : node594;
													assign node594 = (inp[12]) ? node598 : node595;
														assign node595 = (inp[6]) ? 46'b0001000000000100000000001000000010000000000000 : 46'b0001000000000100000000001000000010100000000000;
														assign node598 = (inp[6]) ? 46'b0001000000000100000000001000000000000000000000 : 46'b0001000000000100000000001000000000100000000000;
													assign node601 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : node602;
														assign node602 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000000100000000001001000000000000000010;
											assign node606 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node607;
												assign node607 = (inp[10]) ? node613 : node608;
													assign node608 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : node609;
														assign node609 = (inp[8]) ? 46'b0000000000000100000000001001100000000000000010 : 46'b0000000000000000000000000000000000000000000000;
													assign node613 = (inp[12]) ? node617 : node614;
														assign node614 = (inp[14]) ? 46'b0000000000000010000000001001100010000000000010 : 46'b0000000000000000000000001001100010100000000010;
														assign node617 = (inp[6]) ? 46'b0000000000000000000000001001100000000000000010 : 46'b0000000000000100000000001001100000100000000010;
										assign node621 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : node622;
											assign node622 = (inp[7]) ? node630 : node623;
												assign node623 = (inp[8]) ? node625 : 46'b0000000000000000000000000000000000000000000000;
													assign node625 = (inp[5]) ? node627 : 46'b0000000000000000000000000000000000000000000000;
														assign node627 = (inp[10]) ? 46'b0000000000000010000000001001100000000000000010 : 46'b0000000000000000001000001001100000000000000010;
												assign node630 = (inp[5]) ? 46'b0000000000000000000000000000000000000000000000 : node631;
													assign node631 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : node632;
														assign node632 = (inp[10]) ? 46'b0001000000000110000000001000000010100000000000 : 46'b0001000000000100001000001001000010100000000000;
							assign node639 = (inp[9]) ? node789 : node640;
								assign node640 = (inp[0]) ? node664 : node641;
									assign node641 = (inp[5]) ? node643 : 46'b0000000000000000000000000000000000000000000000;
										assign node643 = (inp[7]) ? node645 : 46'b0000000000000000000000000000000000000000000000;
											assign node645 = (inp[6]) ? node655 : node646;
												assign node646 = (inp[12]) ? node648 : 46'b0000000000000000000000000000000000000000000000;
													assign node648 = (inp[8]) ? node652 : node649;
														assign node649 = (inp[10]) ? 46'b0000000000000000001001000001000000100000000000 : 46'b0000000000000100001001000001000000100000000000;
														assign node652 = (inp[4]) ? 46'b0000000000000000001001000001000000100000000010 : 46'b0000000000000110000001000000000000100000000000;
												assign node655 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node656;
													assign node656 = (inp[4]) ? node660 : node657;
														assign node657 = (inp[10]) ? 46'b0000000000000000000001000001000010000000000010 : 46'b0000000000000100000001000000000010000000000000;
														assign node660 = (inp[14]) ? 46'b0000000000000010001001000001000010000000000000 : 46'b0000000000000100001001000001000010000000000000;
									assign node664 = (inp[6]) ? node728 : node665;
										assign node665 = (inp[5]) ? node697 : node666;
											assign node666 = (inp[12]) ? node682 : node667;
												assign node667 = (inp[7]) ? node675 : node668;
													assign node668 = (inp[4]) ? node672 : node669;
														assign node669 = (inp[14]) ? 46'b0101000000000110000000000000100010100000000000 : 46'b0101000000000100000000000001100010100000000010;
														assign node672 = (inp[10]) ? 46'b0101000000000010000000000000100010100000000000 : 46'b0101000000000000001000000001100010100000000000;
													assign node675 = (inp[14]) ? node679 : node676;
														assign node676 = (inp[10]) ? 46'b0101000000000010000000000001000010100000000010 : 46'b0101000000000000000000000001000010100000000010;
														assign node679 = (inp[4]) ? 46'b0101000000000010001000000001000010100000000000 : 46'b0101000000000010000000000001000010100000000010;
												assign node682 = (inp[7]) ? node690 : node683;
													assign node683 = (inp[4]) ? node687 : node684;
														assign node684 = (inp[8]) ? 46'b0101000000000000000000000001100000100000000010 : 46'b0101000000000000001000000001100000100000000010;
														assign node687 = (inp[14]) ? 46'b0101000000000010001000000001100000100000000000 : 46'b0101000000000000001000000001100000100000000010;
													assign node690 = (inp[8]) ? node694 : node691;
														assign node691 = (inp[14]) ? 46'b0101000000000000001000000001000000100000000000 : 46'b0101000000000100000000000000000000100000000000;
														assign node694 = (inp[10]) ? 46'b0101000000000010000000000001000000100000000010 : 46'b0101000000000100000000000001000000100000000010;
											assign node697 = (inp[7]) ? node713 : node698;
												assign node698 = (inp[8]) ? node706 : node699;
													assign node699 = (inp[10]) ? node703 : node700;
														assign node700 = (inp[12]) ? 46'b0100000000000100001000000001100000100000000000 : 46'b0100000000000100001000000001100010100000000000;
														assign node703 = (inp[4]) ? 46'b0100000000000110000000000000100000100000000000 : 46'b0100000000000100000000000001100000100000000010;
													assign node706 = (inp[14]) ? node710 : node707;
														assign node707 = (inp[10]) ? 46'b0100000000000000000000000001100000100000000010 : 46'b0100000000000100000000000001100000100000000010;
														assign node710 = (inp[10]) ? 46'b0100000000000010000000000000100000100000000000 : 46'b0100000000000010001000000001100000100000000000;
												assign node713 = (inp[12]) ? node721 : node714;
													assign node714 = (inp[10]) ? node718 : node715;
														assign node715 = (inp[4]) ? 46'b0100000000000000001000000001000010100000000000 : 46'b0100000000000100000000000000000010100000000000;
														assign node718 = (inp[4]) ? 46'b0100000000000010000000000000000010100000000000 : 46'b0100000000000000000000000001000010100000000010;
													assign node721 = (inp[10]) ? node725 : node722;
														assign node722 = (inp[8]) ? 46'b0100000000000100000000000000000000100000000000 : 46'b0100000000000100001000000001000000100000000000;
														assign node725 = (inp[14]) ? 46'b0100000000000000001000000001000000100000000000 : 46'b0100000000000000000000000001000000100000000010;
										assign node728 = (inp[7]) ? node760 : node729;
											assign node729 = (inp[12]) ? node745 : node730;
												assign node730 = (inp[5]) ? node738 : node731;
													assign node731 = (inp[8]) ? node735 : node732;
														assign node732 = (inp[14]) ? 46'b0101000000000010001000000001100010000000000000 : 46'b0101000000000100000000000000100010000000000000;
														assign node735 = (inp[10]) ? 46'b0101000000000010000000000001100010000000000010 : 46'b0101000000000000001000000001100010000000000010;
													assign node738 = (inp[14]) ? node742 : node739;
														assign node739 = (inp[8]) ? 46'b0100000000000100000000000001100010000000000010 : 46'b0100000000000100000000000000100010000000000000;
														assign node742 = (inp[8]) ? 46'b0100000000000010000000000000100010000000000000 : 46'b0100000000000100001000000001100010000000000000;
												assign node745 = (inp[5]) ? node753 : node746;
													assign node746 = (inp[8]) ? node750 : node747;
														assign node747 = (inp[10]) ? 46'b0101000000000000000000000001100000000000000010 : 46'b0101000000000100001000000001100000000000000000;
														assign node750 = (inp[14]) ? 46'b0101000000000010000000000000100000000000000000 : 46'b0101000000000000000000000001100000000000000010;
													assign node753 = (inp[8]) ? node757 : node754;
														assign node754 = (inp[10]) ? 46'b0100000000000010000000000000100000000000000000 : 46'b0100000000000000001000000001100000000000000000;
														assign node757 = (inp[14]) ? 46'b0100000000000010001000000001100000000000000000 : 46'b0100000000000000000000000001100000000000000010;
											assign node760 = (inp[12]) ? node774 : node761;
												assign node761 = (inp[10]) ? node767 : node762;
													assign node762 = (inp[4]) ? node764 : 46'b0100000000000100001000000001000010000000000000;
														assign node764 = (inp[5]) ? 46'b0100000000000000001000000001000010000000000000 : 46'b0101000000000000001000000001000010000000000000;
													assign node767 = (inp[4]) ? node771 : node768;
														assign node768 = (inp[8]) ? 46'b0100000000000000000000000001000010000000000010 : 46'b0100000000000000001000000001000010000000000010;
														assign node771 = (inp[5]) ? 46'b0100000000000010000000000000000010000000000000 : 46'b0101000000000110000000000000000010000000000000;
												assign node774 = (inp[5]) ? node782 : node775;
													assign node775 = (inp[8]) ? node779 : node776;
														assign node776 = (inp[14]) ? 46'b0101000000000010001000000001000000000000000000 : 46'b0101000000000100000000000000000000000000000000;
														assign node779 = (inp[10]) ? 46'b0101000000000010000000000001000000000000000010 : 46'b0101000000000010000000000000000000000000000000;
													assign node782 = (inp[14]) ? node786 : node783;
														assign node783 = (inp[8]) ? 46'b0100000000000000000000000001000000000000000010 : 46'b0100000000000100000000000000000000000000000000;
														assign node786 = (inp[8]) ? 46'b0100000000000010000000000000000000000000000000 : 46'b0100000000000000001000000001000000000000000000;
								assign node789 = (inp[0]) ? node915 : node790;
									assign node790 = (inp[12]) ? node854 : node791;
										assign node791 = (inp[6]) ? node823 : node792;
											assign node792 = (inp[7]) ? node808 : node793;
												assign node793 = (inp[5]) ? node801 : node794;
													assign node794 = (inp[4]) ? node798 : node795;
														assign node795 = (inp[10]) ? 46'b1001000000000000000000000001100010100000000010 : 46'b1001000000000100000000000000100010100000000000;
														assign node798 = (inp[14]) ? 46'b1001000000000010000000000000100010100000000000 : 46'b1001000000000000000000000001100010100000000010;
													assign node801 = (inp[10]) ? node805 : node802;
														assign node802 = (inp[4]) ? 46'b1000000000000000001000000001100010100000000000 : 46'b1000000000000100000000000000100010100000000000;
														assign node805 = (inp[14]) ? 46'b1000000000000010000000000000100010100000000000 : 46'b1000000000000010000000000000100010100000000000;
												assign node808 = (inp[5]) ? node816 : node809;
													assign node809 = (inp[8]) ? node813 : node810;
														assign node810 = (inp[14]) ? 46'b1001000000000000001000000001000010100000000000 : 46'b1001000000000100001000000001000010100000000000;
														assign node813 = (inp[14]) ? 46'b1001000000000010000000000000000010100000000000 : 46'b1001000000000000000000000001000010100000000010;
													assign node816 = (inp[10]) ? node820 : node817;
														assign node817 = (inp[4]) ? 46'b1000000000000000001000000001000010100000000000 : 46'b1000000000000100000000000000000010100000000000;
														assign node820 = (inp[4]) ? 46'b1000000000000010000000000001000010100000000010 : 46'b1000000000000000000000000001000010100000000010;
											assign node823 = (inp[5]) ? node839 : node824;
												assign node824 = (inp[4]) ? node832 : node825;
													assign node825 = (inp[10]) ? node829 : node826;
														assign node826 = (inp[7]) ? 46'b1001000000000100000000000000000010000000000000 : 46'b1001000000000100000000000000100010000000000000;
														assign node829 = (inp[14]) ? 46'b1001000000000000001000000001000010000000000010 : 46'b1001000000000100000000000001000010000000000010;
													assign node832 = (inp[7]) ? node836 : node833;
														assign node833 = (inp[14]) ? 46'b1001000000000010001000000001100010000000000000 : 46'b1001000000000000001000000001100010000000000010;
														assign node836 = (inp[14]) ? 46'b1001000000000000001000000001000010000000000000 : 46'b1001000000000100001000000001000010000000000000;
												assign node839 = (inp[7]) ? node847 : node840;
													assign node840 = (inp[14]) ? node844 : node841;
														assign node841 = (inp[4]) ? 46'b1000000000000010000000000000100010000000000000 : 46'b1000000000000100000000000001100010000000000010;
														assign node844 = (inp[4]) ? 46'b1000000000000000001000000001100010000000000000 : 46'b1000000000000100001000000001100010000000000000;
													assign node847 = (inp[14]) ? node851 : node848;
														assign node848 = (inp[4]) ? 46'b1000000000000110000000000000000010000000000000 : 46'b1000000000000100000000000001000010000000000010;
														assign node851 = (inp[4]) ? 46'b1000000000000010001000000001000010000000000000 : 46'b1000000000000010000000000001000010000000000010;
										assign node854 = (inp[5]) ? node886 : node855;
											assign node855 = (inp[7]) ? node871 : node856;
												assign node856 = (inp[10]) ? node864 : node857;
													assign node857 = (inp[6]) ? node861 : node858;
														assign node858 = (inp[8]) ? 46'b1001000000000010001000000001100000100000000000 : 46'b1001000000000100001000000001100000100000000000;
														assign node861 = (inp[8]) ? 46'b1001000000000010001000000001100000000000000000 : 46'b1001000000000000001000000001100000000000000000;
													assign node864 = (inp[4]) ? node868 : node865;
														assign node865 = (inp[6]) ? 46'b1001000000000000000000000001100000000000000010 : 46'b1001000000000000000000000001100000100000000010;
														assign node868 = (inp[8]) ? 46'b1001000000000010000000000000100000000000000000 : 46'b1001000000000110000000000000100000000000000000;
												assign node871 = (inp[6]) ? node879 : node872;
													assign node872 = (inp[10]) ? node876 : node873;
														assign node873 = (inp[4]) ? 46'b1001000000000000001000000001000000100000000010 : 46'b1001000000000100000000000000000000100000000000;
														assign node876 = (inp[14]) ? 46'b1001000000000000001000000001000000100000000010 : 46'b1001000000000000000000000001000000100000000010;
													assign node879 = (inp[10]) ? node883 : node880;
														assign node880 = (inp[8]) ? 46'b1001000000000010000000000000000000000000000000 : 46'b1001000000000100001000000001000000000000000000;
														assign node883 = (inp[4]) ? 46'b1001000000000010000000000000000000000000000000 : 46'b1001000000000000000000000001000000000000000010;
											assign node886 = (inp[7]) ? node900 : node887;
												assign node887 = (inp[6]) ? node893 : node888;
													assign node888 = (inp[10]) ? node890 : 46'b1000000000000110000000000000100000100000000000;
														assign node890 = (inp[8]) ? 46'b1000000000000010000000000001100000100000000010 : 46'b1000000000000000001000000001100000100000000010;
													assign node893 = (inp[14]) ? node897 : node894;
														assign node894 = (inp[8]) ? 46'b1000000000000000000000000001100000000000000010 : 46'b1000000000000110000000000000100000000000000000;
														assign node897 = (inp[8]) ? 46'b1000000000000010000000000000100000000000000000 : 46'b1000000000000000001000000001100000000000000000;
												assign node900 = (inp[10]) ? node908 : node901;
													assign node901 = (inp[8]) ? node905 : node902;
														assign node902 = (inp[6]) ? 46'b1000000000000100001000000001000000000000000000 : 46'b1000000000000100001000000001000000100000000000;
														assign node905 = (inp[4]) ? 46'b1000000000000010001000000001000000100000000000 : 46'b1000000000000110000000000000000000100000000000;
													assign node908 = (inp[8]) ? node912 : node909;
														assign node909 = (inp[14]) ? 46'b1000000000000000001000000001000000000000000010 : 46'b1000000000000100000000000001000000000000000010;
														assign node912 = (inp[6]) ? 46'b1000000000000010000000000001000000000000000010 : 46'b1000000000000010000000000001000000100000000010;
									assign node915 = (inp[5]) ? node977 : node916;
										assign node916 = (inp[12]) ? node948 : node917;
											assign node917 = (inp[6]) ? node933 : node918;
												assign node918 = (inp[7]) ? node926 : node919;
													assign node919 = (inp[8]) ? node923 : node920;
														assign node920 = (inp[14]) ? 46'b0001000000000000001000000001100010101000000000 : 46'b0001000000000110000000000000100010101000000000;
														assign node923 = (inp[4]) ? 46'b0001000000000010000000000000100010101000000000 : 46'b0001000000000110000000000000100010101000000000;
													assign node926 = (inp[10]) ? node930 : node927;
														assign node927 = (inp[8]) ? 46'b0001000000000000001000000001000010101000000010 : 46'b0001000000000100001000000001000010101000000000;
														assign node930 = (inp[8]) ? 46'b0001000000000010000000000001000010101000000010 : 46'b0001000000000010001000000001000010101000000000;
												assign node933 = (inp[10]) ? node941 : node934;
													assign node934 = (inp[4]) ? node938 : node935;
														assign node935 = (inp[14]) ? 46'b0001000000000110000000000000000010001000000000 : 46'b0001000000000100000000000000000010001000000000;
														assign node938 = (inp[8]) ? 46'b0001000000000000001000000001000010001000000000 : 46'b0001000000000100001000000001000010001000000000;
													assign node941 = (inp[7]) ? node945 : node942;
														assign node942 = (inp[8]) ? 46'b0001000000000010000000000001100010001000000010 : 46'b0001000000000000001000000001100010001000000010;
														assign node945 = (inp[14]) ? 46'b0001000000000000000000000001000010001000000010 : 46'b0001000000000000000000000001000010001000000010;
											assign node948 = (inp[6]) ? node964 : node949;
												assign node949 = (inp[14]) ? node957 : node950;
													assign node950 = (inp[7]) ? node954 : node951;
														assign node951 = (inp[4]) ? 46'b0001000000000000001000000001100000101000000010 : 46'b0001000000000100000000000001100000101000000010;
														assign node954 = (inp[10]) ? 46'b0001000000000100000000000001000000101000000010 : 46'b0001000000000100000000000000000000101000000000;
													assign node957 = (inp[7]) ? node961 : node958;
														assign node958 = (inp[8]) ? 46'b0001000000000010000000000000100000101000000000 : 46'b0001000000000010001000000001100000101000000000;
														assign node961 = (inp[8]) ? 46'b0001000000000010000000000000000000101000000000 : 46'b0001000000000000001000000001000000101000000000;
												assign node964 = (inp[7]) ? node970 : node965;
													assign node965 = (inp[14]) ? node967 : 46'b0001000000000000001000000001100000001000000010;
														assign node967 = (inp[4]) ? 46'b0001000000000010001000000001100000001000000000 : 46'b0001000000000100000000000000100000001000000000;
													assign node970 = (inp[8]) ? node974 : node971;
														assign node971 = (inp[10]) ? 46'b0001000000000000001000000001000000001000000010 : 46'b0001000000000100001000000001000000001000000000;
														assign node974 = (inp[14]) ? 46'b0001000000000010000000000000000000001000000000 : 46'b0001000000000100000000000001000000001000000010;
										assign node977 = (inp[7]) ? node1009 : node978;
											assign node978 = (inp[6]) ? node994 : node979;
												assign node979 = (inp[12]) ? node987 : node980;
													assign node980 = (inp[8]) ? node984 : node981;
														assign node981 = (inp[4]) ? 46'b0000000000000110000000000000100010101000000000 : 46'b0000000000000100001000000001100010101000000010;
														assign node984 = (inp[4]) ? 46'b0000000000000000001000000001100010101000000010 : 46'b0000000000000000000000000001100010101000000010;
													assign node987 = (inp[10]) ? node991 : node988;
														assign node988 = (inp[8]) ? 46'b0000000000000000001000000001100000101000000010 : 46'b0000000000000000001000000001100000101000000000;
														assign node991 = (inp[8]) ? 46'b0000000000000010000000000001100000101000000010 : 46'b0000000000000100000000000001100000101000000010;
												assign node994 = (inp[12]) ? node1002 : node995;
													assign node995 = (inp[4]) ? node999 : node996;
														assign node996 = (inp[8]) ? 46'b0000000000000100000000000001100010001000000010 : 46'b0000000000000000001000000001100010001000000010;
														assign node999 = (inp[14]) ? 46'b0000000000000010001000000001100010001000000000 : 46'b0000000000000100001000000001100010001000000000;
													assign node1002 = (inp[10]) ? node1006 : node1003;
														assign node1003 = (inp[8]) ? 46'b0000000000000000000000000001100000001000000010 : 46'b0000000000000100001000000001100000001000000000;
														assign node1006 = (inp[8]) ? 46'b0000000000000010000000000001100000001000000010 : 46'b0000000000000100000000000001100000001000000010;
											assign node1009 = (inp[6]) ? node1025 : node1010;
												assign node1010 = (inp[8]) ? node1018 : node1011;
													assign node1011 = (inp[10]) ? node1015 : node1012;
														assign node1012 = (inp[12]) ? 46'b0000000000000100001000000001000000101000000000 : 46'b0000000000000000001000000001000010101000000000;
														assign node1015 = (inp[14]) ? 46'b0000000000000010001000000001000000101000000000 : 46'b0000000000000110000000000000000010101000000000;
													assign node1018 = (inp[14]) ? node1022 : node1019;
														assign node1019 = (inp[10]) ? 46'b0000000000000010000000000001000010101000000010 : 46'b0000000000000100000000000001000010101000000010;
														assign node1022 = (inp[12]) ? 46'b0000000000000010000000000000000000101000000000 : 46'b0000000000000010000000000000000010101000000000;
												assign node1025 = (inp[12]) ? node1033 : node1026;
													assign node1026 = (inp[10]) ? node1030 : node1027;
														assign node1027 = (inp[4]) ? 46'b0000000000000100001000000001000010001000000000 : 46'b0000000000000100000000000000000010001000000000;
														assign node1030 = (inp[8]) ? 46'b0000000000000010000000000001000010001000000010 : 46'b0000000000000100000000000001000010001000000010;
													assign node1033 = (inp[14]) ? node1037 : node1034;
														assign node1034 = (inp[4]) ? 46'b0000000000000100000000000000000000001000000000 : 46'b0000000000000100000000000001000000001000000010;
														assign node1037 = (inp[8]) ? 46'b0000000000000010000000000001000000001000000010 : 46'b0000000000000000001000000001000000001000000010;
						assign node1040 = (inp[11]) ? node1378 : node1041;
							assign node1041 = (inp[9]) ? node1127 : node1042;
								assign node1042 = (inp[5]) ? node1058 : node1043;
									assign node1043 = (inp[6]) ? node1045 : 46'b0000000000000000000000000000000000000000000000;
										assign node1045 = (inp[0]) ? node1047 : 46'b0000000000000000000000000000000000000000000000;
											assign node1047 = (inp[12]) ? node1049 : 46'b0000000000000000000000000000000000000000000000;
												assign node1049 = (inp[7]) ? node1051 : 46'b0000000000000000000000000000000000000000000000;
													assign node1051 = (inp[14]) ? node1055 : node1052;
														assign node1052 = (inp[8]) ? 46'b0001000000000001000000000001000000000000100010 : 46'b0001000000000101000000000000000000000000100000;
														assign node1055 = (inp[8]) ? 46'b0001000000000011000000000000000000000000100000 : 46'b0001000000000001001000000001000000000000100000;
									assign node1058 = (inp[7]) ? node1072 : node1059;
										assign node1059 = (inp[6]) ? node1061 : 46'b0000000000000000000000000000000000000000000000;
											assign node1061 = (inp[0]) ? node1063 : 46'b0000000000000000000000000000000000000000000000;
												assign node1063 = (inp[12]) ? node1065 : 46'b0000000000000000000000000000000000000000000000;
													assign node1065 = (inp[14]) ? node1069 : node1066;
														assign node1066 = (inp[8]) ? 46'b0000000000000001000000000001100000000000100010 : 46'b0000000000000101000000000000100000000000100000;
														assign node1069 = (inp[8]) ? 46'b0000000000000011000000000001100000000000100000 : 46'b0000000000000001001000000001100000000000100000;
										assign node1072 = (inp[0]) ? node1104 : node1073;
											assign node1073 = (inp[6]) ? node1089 : node1074;
												assign node1074 = (inp[10]) ? node1082 : node1075;
													assign node1075 = (inp[12]) ? node1079 : node1076;
														assign node1076 = (inp[8]) ? 46'b0000000000100000001001000001000010100000000010 : 46'b0000000000100100001001000001000010100000000000;
														assign node1079 = (inp[8]) ? 46'b0000000000100010001001000001000000100000000000 : 46'b0000000000100100001001000001000000100000000000;
													assign node1082 = (inp[4]) ? node1086 : node1083;
														assign node1083 = (inp[8]) ? 46'b0000000000100010000001000001000000100000000010 : 46'b0000000000100000001001000001000000100000000010;
														assign node1086 = (inp[12]) ? 46'b0000000000100010000001000000000000100000000000 : 46'b0000000000100010000001000000000010100000000000;
												assign node1089 = (inp[12]) ? node1097 : node1090;
													assign node1090 = (inp[8]) ? node1094 : node1091;
														assign node1091 = (inp[4]) ? 46'b0000000000100000001001000001000010000000000000 : 46'b0000000000100000001001000001000010000000000000;
														assign node1094 = (inp[10]) ? 46'b0000000000100010000001000001000010000000000010 : 46'b0000000000100000000001000001000010000000000010;
													assign node1097 = (inp[8]) ? node1101 : node1098;
														assign node1098 = (inp[14]) ? 46'b0000000000100000001001000001000000000000000010 : 46'b0000000000100100000001000000000000000000000000;
														assign node1101 = (inp[14]) ? 46'b0000000000100010000001000000000000000000000000 : 46'b0000000000100010000001000001000000000000000010;
											assign node1104 = (inp[8]) ? node1116 : node1105;
												assign node1105 = (inp[6]) ? node1111 : node1106;
													assign node1106 = (inp[12]) ? node1108 : 46'b0000000000000000000000000000000000000000000000;
														assign node1108 = (inp[14]) ? 46'b0000000000000001001000000001000000100000100000 : 46'b0000000000000101000000000000000000100000100000;
													assign node1111 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node1112;
														assign node1112 = (inp[14]) ? 46'b0000000000000001001000000001000010000000100000 : 46'b0000000000000101000000000001000010000000100000;
												assign node1116 = (inp[12]) ? node1122 : node1117;
													assign node1117 = (inp[6]) ? node1119 : 46'b0000000000000000000000000000000000000000000000;
														assign node1119 = (inp[10]) ? 46'b0000000000000011000000000000000010000000100000 : 46'b0000000000000001001000000001000010000000100000;
													assign node1122 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : node1123;
														assign node1123 = (inp[4]) ? 46'b0000000000000011001000000001000000100000100000 : 46'b0000000000000111000000000000000000100000100000;
								assign node1127 = (inp[5]) ? node1253 : node1128;
									assign node1128 = (inp[0]) ? node1190 : node1129;
										assign node1129 = (inp[12]) ? node1161 : node1130;
											assign node1130 = (inp[6]) ? node1146 : node1131;
												assign node1131 = (inp[7]) ? node1139 : node1132;
													assign node1132 = (inp[10]) ? node1136 : node1133;
														assign node1133 = (inp[14]) ? 46'b0001000000100110000000000000100010100000100000 : 46'b0001000000100100000000000000100010100000100000;
														assign node1136 = (inp[8]) ? 46'b0001000000100010000000000000100010100000100000 : 46'b0001000000100010001000000001100010100000100000;
													assign node1139 = (inp[4]) ? node1143 : node1140;
														assign node1140 = (inp[14]) ? 46'b0001000000100000000000000001000010100000100010 : 46'b0001000000100100000000000001000010100000100010;
														assign node1143 = (inp[10]) ? 46'b0001000000100010000000000000000010100000100000 : 46'b0001000000100000001000000001000010100000100000;
												assign node1146 = (inp[7]) ? node1154 : node1147;
													assign node1147 = (inp[10]) ? node1151 : node1148;
														assign node1148 = (inp[4]) ? 46'b0001000000100000001000000001100010000000100000 : 46'b0001000000100100000000000000100010000000100000;
														assign node1151 = (inp[14]) ? 46'b0001000000100000001000000001100010000000100010 : 46'b0001000000100000000000000001100010000000100010;
													assign node1154 = (inp[4]) ? node1158 : node1155;
														assign node1155 = (inp[14]) ? 46'b0001000000100000001000000001000010000000100010 : 46'b0001000000100100000000000001000010000000100010;
														assign node1158 = (inp[10]) ? 46'b0001000000100010000000000000000010000000100000 : 46'b0001000000100100001000000001000010000000100000;
											assign node1161 = (inp[6]) ? node1177 : node1162;
												assign node1162 = (inp[7]) ? node1170 : node1163;
													assign node1163 = (inp[4]) ? node1167 : node1164;
														assign node1164 = (inp[14]) ? 46'b0001000000100110000000000000100000100000100000 : 46'b0001000000100100000000000001100000100000100010;
														assign node1167 = (inp[10]) ? 46'b0001000000100010000000000000100000100000100000 : 46'b0001000000100000001000000001100000100000100000;
													assign node1170 = (inp[8]) ? node1174 : node1171;
														assign node1171 = (inp[14]) ? 46'b0001000000100000001000000001000000100000100000 : 46'b0001000000100100000000000000000000100000100000;
														assign node1174 = (inp[10]) ? 46'b0001000000100010000000000001000000100000100010 : 46'b0001000000100000001000000001000000100000100010;
												assign node1177 = (inp[7]) ? node1183 : node1178;
													assign node1178 = (inp[14]) ? node1180 : 46'b0001000000100110000000000000100000000000100000;
														assign node1180 = (inp[10]) ? 46'b0001000000100010001000000001100000000000100010 : 46'b0001000000100110000000000000100000000000100000;
													assign node1183 = (inp[14]) ? node1187 : node1184;
														assign node1184 = (inp[4]) ? 46'b0001000000100010000000000000000000000000100000 : 46'b0001000000100100000000000001000000000000100010;
														assign node1187 = (inp[8]) ? 46'b0001000000100010000000000000000000000000100000 : 46'b0001000000100000001000000001000000000000100000;
										assign node1190 = (inp[12]) ? node1222 : node1191;
											assign node1191 = (inp[6]) ? node1207 : node1192;
												assign node1192 = (inp[8]) ? node1200 : node1193;
													assign node1193 = (inp[7]) ? node1197 : node1194;
														assign node1194 = (inp[14]) ? 46'b0001000000000000001000000001100010100000100000 : 46'b0001000000000100000000000000100010100000100000;
														assign node1197 = (inp[4]) ? 46'b0001000000000000001000000001000010100000100000 : 46'b0001000000000100000000000000000010100000100000;
													assign node1200 = (inp[7]) ? node1204 : node1201;
														assign node1201 = (inp[14]) ? 46'b0001000000000010000000000001100010100000100000 : 46'b0001000000000000000000000001100010100000100010;
														assign node1204 = (inp[14]) ? 46'b0001000000000010000000000000000010100000100000 : 46'b0001000000000000000000000001000010100000100010;
												assign node1207 = (inp[7]) ? node1215 : node1208;
													assign node1208 = (inp[8]) ? node1212 : node1209;
														assign node1209 = (inp[14]) ? 46'b0001000000000000001000000001100010000000100000 : 46'b0001000000000100000000000001100010000000100010;
														assign node1212 = (inp[14]) ? 46'b0001000000000010000000000000100010000000100000 : 46'b0001000000000000000000000001100010000000100010;
													assign node1215 = (inp[14]) ? node1219 : node1216;
														assign node1216 = (inp[8]) ? 46'b0001000000000000000000000001000010000000100010 : 46'b0001000000000100000000000000000010000000100000;
														assign node1219 = (inp[4]) ? 46'b0001000000000010001000000001000010000000100000 : 46'b0001000000000010000000000001000010000000100010;
											assign node1222 = (inp[7]) ? node1238 : node1223;
												assign node1223 = (inp[6]) ? node1231 : node1224;
													assign node1224 = (inp[10]) ? node1228 : node1225;
														assign node1225 = (inp[8]) ? 46'b0001000000000000001000000001100000100000100010 : 46'b0001000000000100001000000001100000100000100000;
														assign node1228 = (inp[14]) ? 46'b0001000000000010000000000000100000100000100000 : 46'b0001000000000010000000000000100000100000100000;
													assign node1231 = (inp[4]) ? node1235 : node1232;
														assign node1232 = (inp[10]) ? 46'b0001000000000000001000000001100000000000100010 : 46'b0001000000000100000000000000100000000000100000;
														assign node1235 = (inp[14]) ? 46'b0001000000000010001000000001100000000000100000 : 46'b0001000000000110000000000000100000000000100000;
												assign node1238 = (inp[6]) ? node1246 : node1239;
													assign node1239 = (inp[14]) ? node1243 : node1240;
														assign node1240 = (inp[8]) ? 46'b0001000000000000000000000001000000100000100010 : 46'b0001000000000100000000000000000000100000100000;
														assign node1243 = (inp[4]) ? 46'b0001000000000010001000000001000000100000100000 : 46'b0001000000000010000000000000000000100000100000;
													assign node1246 = (inp[10]) ? node1250 : node1247;
														assign node1247 = (inp[4]) ? 46'b0001000000000000001000000001000000000000100000 : 46'b0001000000000110000000000000000000000000100000;
														assign node1250 = (inp[8]) ? 46'b0001000000000010000000000001000000000000100010 : 46'b0001000000000100000000000000000000000000100000;
									assign node1253 = (inp[0]) ? node1315 : node1254;
										assign node1254 = (inp[6]) ? node1284 : node1255;
											assign node1255 = (inp[7]) ? node1271 : node1256;
												assign node1256 = (inp[10]) ? node1264 : node1257;
													assign node1257 = (inp[4]) ? node1261 : node1258;
														assign node1258 = (inp[12]) ? 46'b0000000000100100000000000000100000100000100000 : 46'b0000000000100100000000000000100010100000100000;
														assign node1261 = (inp[12]) ? 46'b0000000000100000001000000001100000100000100000 : 46'b0000000000100010001000000001100010100000100000;
													assign node1264 = (inp[8]) ? node1268 : node1265;
														assign node1265 = (inp[12]) ? 46'b0000000000100000001000000001100000100000100010 : 46'b0000000000100000001000000001100010100000100010;
														assign node1268 = (inp[12]) ? 46'b0000000000100010000000000001100000100000100010 : 46'b0000000000100010000000000001100010100000100010;
												assign node1271 = (inp[12]) ? node1277 : node1272;
													assign node1272 = (inp[14]) ? 46'b0000000000100010001000000001000010100000100000 : node1273;
														assign node1273 = (inp[10]) ? 46'b0000000000100110000000000000000010100000100000 : 46'b0000000000100100000000000000000010100000100000;
													assign node1277 = (inp[4]) ? node1281 : node1278;
														assign node1278 = (inp[10]) ? 46'b0000000000100000000000000001000000100000100010 : 46'b0000000000100100001000000001000000100000100000;
														assign node1281 = (inp[10]) ? 46'b0000000000100010000000000000000000100000100000 : 46'b0000000000100000001000000001000000100000100010;
											assign node1284 = (inp[7]) ? node1300 : node1285;
												assign node1285 = (inp[12]) ? node1293 : node1286;
													assign node1286 = (inp[4]) ? node1290 : node1287;
														assign node1287 = (inp[14]) ? 46'b0000000000100100000000000000100010000000100000 : 46'b0000000000100100000000000001100010000000100010;
														assign node1290 = (inp[10]) ? 46'b0000000000100010000000000000100010000000100000 : 46'b0000000000100000001000000001100010000000100000;
													assign node1293 = (inp[10]) ? node1297 : node1294;
														assign node1294 = (inp[8]) ? 46'b0000000000100000000000000001100000000000100010 : 46'b0000000000100100001000000001100000000000100000;
														assign node1297 = (inp[4]) ? 46'b0000000000100010000000000000100000000000100000 : 46'b0000000000100000000000000001100000000000100010;
												assign node1300 = (inp[4]) ? node1308 : node1301;
													assign node1301 = (inp[10]) ? node1305 : node1302;
														assign node1302 = (inp[12]) ? 46'b0000000000100100000000000000000000000000100000 : 46'b0000000000100100000000000001000010000000100000;
														assign node1305 = (inp[14]) ? 46'b0000000000100010000000000001000000000000100010 : 46'b0000000000100100000000000001000010000000100010;
													assign node1308 = (inp[12]) ? node1312 : node1309;
														assign node1309 = (inp[14]) ? 46'b0000000000100010001000000001000010000000100000 : 46'b0000000000100000001000000001000010000000100010;
														assign node1312 = (inp[10]) ? 46'b0000000000100010000000000000000000000000100000 : 46'b0000000000100000001000000001000000000000100000;
										assign node1315 = (inp[6]) ? node1347 : node1316;
											assign node1316 = (inp[7]) ? node1332 : node1317;
												assign node1317 = (inp[12]) ? node1325 : node1318;
													assign node1318 = (inp[4]) ? node1322 : node1319;
														assign node1319 = (inp[14]) ? 46'b0000000000000100001000000001100010100000100000 : 46'b0000000000000100000000000001100010100000100010;
														assign node1322 = (inp[10]) ? 46'b0000000000000010000000000000100010100000100000 : 46'b0000000000000000001000000001100010100000100000;
													assign node1325 = (inp[4]) ? node1329 : node1326;
														assign node1326 = (inp[14]) ? 46'b0000000000000110000000000000100000100000100000 : 46'b0000000000000100000000000000100000100000100000;
														assign node1329 = (inp[10]) ? 46'b0000000000000010000000000000100000100000100000 : 46'b0000000000000000001000000001100000100000100000;
												assign node1332 = (inp[12]) ? node1340 : node1333;
													assign node1333 = (inp[4]) ? node1337 : node1334;
														assign node1334 = (inp[8]) ? 46'b0000000000000010000000000001000010100000100010 : 46'b0000000000000000001000000001000010100000100010;
														assign node1337 = (inp[14]) ? 46'b0000000000000010000000000000000010100000100000 : 46'b0000000000000110000000000000000010100000100000;
													assign node1340 = (inp[14]) ? node1344 : node1341;
														assign node1341 = (inp[8]) ? 46'b0000000000000000000000000001000000100000100010 : 46'b0000000000000100000000000000000000100000100000;
														assign node1344 = (inp[8]) ? 46'b0000000000000010000000000000000000100000100000 : 46'b0000000000000000001000000001000000100000100010;
											assign node1347 = (inp[12]) ? node1363 : node1348;
												assign node1348 = (inp[7]) ? node1356 : node1349;
													assign node1349 = (inp[8]) ? node1353 : node1350;
														assign node1350 = (inp[14]) ? 46'b0000000000000000001000000001100010000000100010 : 46'b0000000000000100000000000001100010000000100010;
														assign node1353 = (inp[4]) ? 46'b0000000000000010000000000000100010000000100000 : 46'b0000000000000000000000000001100010000000100010;
													assign node1356 = (inp[10]) ? node1360 : node1357;
														assign node1357 = (inp[4]) ? 46'b0000000000000010001000000001000010000000100000 : 46'b0000000000000100000000000001000010000000100000;
														assign node1360 = (inp[8]) ? 46'b0000000000000010000000000001000010000000100010 : 46'b0000000000000000001000000001000010000000100010;
												assign node1363 = (inp[7]) ? node1371 : node1364;
													assign node1364 = (inp[8]) ? node1368 : node1365;
														assign node1365 = (inp[4]) ? 46'b0000000000000110000000000000100000000000100000 : 46'b0000000000000100000000000001100000000000100000;
														assign node1368 = (inp[14]) ? 46'b0000000000000010000000000000100000000000100000 : 46'b0000000000000000000000000001100000000000100010;
													assign node1371 = (inp[8]) ? node1375 : node1372;
														assign node1372 = (inp[14]) ? 46'b0000000000000100001000000001000000000000100000 : 46'b0000000000000100000000000000000000000000100000;
														assign node1375 = (inp[14]) ? 46'b0000000000000010000000000001000000000000100000 : 46'b0000000000000000000000000001000000000000100010;
							assign node1378 = (inp[7]) ? node1416 : node1379;
								assign node1379 = (inp[5]) ? node1391 : node1380;
									assign node1380 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1381;
										assign node1381 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1382;
											assign node1382 = (inp[6]) ? node1386 : node1383;
												assign node1383 = (inp[12]) ? 46'b0001000000100000001000000001100000100000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1386 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000100010000000000000100010000000100000;
									assign node1391 = (inp[0]) ? node1407 : node1392;
										assign node1392 = (inp[9]) ? node1400 : node1393;
											assign node1393 = (inp[6]) ? node1397 : node1394;
												assign node1394 = (inp[12]) ? 46'b0000000000100000001000000001100000100000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1397 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000100010000000000000100010000000100000;
											assign node1400 = (inp[6]) ? node1404 : node1401;
												assign node1401 = (inp[12]) ? 46'b0000000010000000000000000001100000100001000010 : 46'b0000000010000000000000000001100010100001000010;
												assign node1404 = (inp[12]) ? 46'b0000000010000000000000000001100000000001000010 : 46'b0000000010000000000000000001100010000001000010;
										assign node1407 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1408;
											assign node1408 = (inp[12]) ? node1412 : node1409;
												assign node1409 = (inp[6]) ? 46'b0000000010000000000000000001100010000000000010 : 46'b0000000010000000000000000001100010100000000010;
												assign node1412 = (inp[6]) ? 46'b0000000010000000000000000001100000000000000010 : 46'b0000000010000000000000000001100000100000000010;
								assign node1416 = (inp[5]) ? node1442 : node1417;
									assign node1417 = (inp[9]) ? node1433 : node1418;
										assign node1418 = (inp[0]) ? node1426 : node1419;
											assign node1419 = (inp[6]) ? node1423 : node1420;
												assign node1420 = (inp[12]) ? 46'b0001000000100000001000000001000000100000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1423 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000100010000000000000000010000000100000;
											assign node1426 = (inp[12]) ? node1430 : node1427;
												assign node1427 = (inp[6]) ? 46'b0001000010000100000000000000000010000000000000 : 46'b0001000010000100000000000000000010100000000000;
												assign node1430 = (inp[6]) ? 46'b0001000010000100000000000000000000000000000000 : 46'b0001000010000100000000000000000000100000000000;
										assign node1433 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1434;
											assign node1434 = (inp[6]) ? node1438 : node1435;
												assign node1435 = (inp[12]) ? 46'b0001000010000100000000000000000000100001000000 : 46'b0001000010000100000000000000000010100001000000;
												assign node1438 = (inp[12]) ? 46'b0001000010000100000000000000000000000001000000 : 46'b0001000010000100000000000000000010000001000000;
									assign node1442 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1443;
										assign node1443 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1444;
											assign node1444 = (inp[6]) ? node1448 : node1445;
												assign node1445 = (inp[12]) ? 46'b0000000000100000001000000001000000100000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1448 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000100010000000000000000010000000100000;

endmodule