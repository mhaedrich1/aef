module dtc_split125_bm72 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node221;
	wire [3-1:0] node224;
	wire [3-1:0] node226;

	assign outp = (inp[3]) ? node126 : node1;
		assign node1 = (inp[6]) ? node65 : node2;
			assign node2 = (inp[9]) ? node34 : node3;
				assign node3 = (inp[0]) ? node19 : node4;
					assign node4 = (inp[1]) ? node12 : node5;
						assign node5 = (inp[10]) ? node9 : node6;
							assign node6 = (inp[5]) ? 3'b101 : 3'b011;
							assign node9 = (inp[2]) ? 3'b001 : 3'b101;
						assign node12 = (inp[10]) ? node16 : node13;
							assign node13 = (inp[4]) ? 3'b001 : 3'b001;
							assign node16 = (inp[4]) ? 3'b010 : 3'b001;
					assign node19 = (inp[8]) ? node27 : node20;
						assign node20 = (inp[5]) ? node24 : node21;
							assign node21 = (inp[11]) ? 3'b110 : 3'b010;
							assign node24 = (inp[10]) ? 3'b100 : 3'b110;
						assign node27 = (inp[7]) ? node31 : node28;
							assign node28 = (inp[2]) ? 3'b100 : 3'b000;
							assign node31 = (inp[5]) ? 3'b001 : 3'b001;
				assign node34 = (inp[1]) ? node50 : node35;
					assign node35 = (inp[8]) ? node43 : node36;
						assign node36 = (inp[5]) ? node40 : node37;
							assign node37 = (inp[10]) ? 3'b000 : 3'b010;
							assign node40 = (inp[2]) ? 3'b100 : 3'b110;
						assign node43 = (inp[0]) ? node47 : node44;
							assign node44 = (inp[5]) ? 3'b110 : 3'b001;
							assign node47 = (inp[7]) ? 3'b010 : 3'b000;
					assign node50 = (inp[8]) ? node58 : node51;
						assign node51 = (inp[0]) ? node55 : node52;
							assign node52 = (inp[10]) ? 3'b000 : 3'b010;
							assign node55 = (inp[4]) ? 3'b000 : 3'b100;
						assign node58 = (inp[7]) ? node62 : node59;
							assign node59 = (inp[0]) ? 3'b000 : 3'b100;
							assign node62 = (inp[5]) ? 3'b000 : 3'b010;
			assign node65 = (inp[9]) ? node95 : node66;
				assign node66 = (inp[0]) ? node80 : node67;
					assign node67 = (inp[4]) ? node73 : node68;
						assign node68 = (inp[7]) ? 3'b111 : node69;
							assign node69 = (inp[8]) ? 3'b111 : 3'b011;
						assign node73 = (inp[1]) ? node77 : node74;
							assign node74 = (inp[2]) ? 3'b101 : 3'b111;
							assign node77 = (inp[8]) ? 3'b011 : 3'b101;
					assign node80 = (inp[8]) ? node88 : node81;
						assign node81 = (inp[7]) ? node85 : node82;
							assign node82 = (inp[2]) ? 3'b011 : 3'b001;
							assign node85 = (inp[10]) ? 3'b101 : 3'b111;
						assign node88 = (inp[10]) ? node92 : node89;
							assign node89 = (inp[4]) ? 3'b011 : 3'b011;
							assign node92 = (inp[5]) ? 3'b101 : 3'b011;
				assign node95 = (inp[7]) ? node111 : node96;
					assign node96 = (inp[0]) ? node104 : node97;
						assign node97 = (inp[4]) ? node101 : node98;
							assign node98 = (inp[10]) ? 3'b101 : 3'b011;
							assign node101 = (inp[1]) ? 3'b110 : 3'b001;
						assign node104 = (inp[1]) ? node108 : node105;
							assign node105 = (inp[8]) ? 3'b110 : 3'b010;
							assign node108 = (inp[10]) ? 3'b010 : 3'b000;
					assign node111 = (inp[0]) ? node119 : node112;
						assign node112 = (inp[10]) ? node116 : node113;
							assign node113 = (inp[4]) ? 3'b011 : 3'b111;
							assign node116 = (inp[4]) ? 3'b001 : 3'b011;
						assign node119 = (inp[4]) ? node123 : node120;
							assign node120 = (inp[2]) ? 3'b001 : 3'b101;
							assign node123 = (inp[5]) ? 3'b010 : 3'b001;
		assign node126 = (inp[6]) ? node170 : node127;
			assign node127 = (inp[0]) ? node155 : node128;
				assign node128 = (inp[9]) ? node142 : node129;
					assign node129 = (inp[4]) ? node137 : node130;
						assign node130 = (inp[8]) ? node134 : node131;
							assign node131 = (inp[1]) ? 3'b000 : 3'b010;
							assign node134 = (inp[2]) ? 3'b010 : 3'b101;
						assign node137 = (inp[5]) ? node139 : 3'b100;
							assign node139 = (inp[10]) ? 3'b100 : 3'b000;
					assign node142 = (inp[2]) ? node150 : node143;
						assign node143 = (inp[4]) ? node147 : node144;
							assign node144 = (inp[5]) ? 3'b100 : 3'b010;
							assign node147 = (inp[10]) ? 3'b000 : 3'b000;
						assign node150 = (inp[4]) ? 3'b000 : node151;
							assign node151 = (inp[10]) ? 3'b000 : 3'b000;
				assign node155 = (inp[1]) ? 3'b000 : node156;
					assign node156 = (inp[8]) ? node162 : node157;
						assign node157 = (inp[4]) ? 3'b000 : node158;
							assign node158 = (inp[10]) ? 3'b000 : 3'b010;
						assign node162 = (inp[9]) ? node166 : node163;
							assign node163 = (inp[4]) ? 3'b000 : 3'b100;
							assign node166 = (inp[2]) ? 3'b000 : 3'b000;
			assign node170 = (inp[9]) ? node200 : node171;
				assign node171 = (inp[4]) ? node187 : node172;
					assign node172 = (inp[10]) ? node180 : node173;
						assign node173 = (inp[11]) ? node177 : node174;
							assign node174 = (inp[1]) ? 3'b001 : 3'b101;
							assign node177 = (inp[5]) ? 3'b001 : 3'b001;
						assign node180 = (inp[7]) ? node184 : node181;
							assign node181 = (inp[8]) ? 3'b101 : 3'b110;
							assign node184 = (inp[5]) ? 3'b100 : 3'b001;
					assign node187 = (inp[5]) ? node195 : node188;
						assign node188 = (inp[8]) ? node192 : node189;
							assign node189 = (inp[7]) ? 3'b000 : 3'b110;
							assign node192 = (inp[1]) ? 3'b010 : 3'b001;
						assign node195 = (inp[7]) ? 3'b110 : node196;
							assign node196 = (inp[0]) ? 3'b000 : 3'b110;
				assign node200 = (inp[0]) ? node216 : node201;
					assign node201 = (inp[7]) ? node209 : node202;
						assign node202 = (inp[4]) ? node206 : node203;
							assign node203 = (inp[1]) ? 3'b010 : 3'b110;
							assign node206 = (inp[10]) ? 3'b000 : 3'b100;
						assign node209 = (inp[4]) ? node213 : node210;
							assign node210 = (inp[1]) ? 3'b110 : 3'b101;
							assign node213 = (inp[8]) ? 3'b110 : 3'b010;
					assign node216 = (inp[4]) ? node224 : node217;
						assign node217 = (inp[5]) ? node221 : node218;
							assign node218 = (inp[1]) ? 3'b000 : 3'b010;
							assign node221 = (inp[10]) ? 3'b000 : 3'b100;
						assign node224 = (inp[7]) ? node226 : 3'b000;
							assign node226 = (inp[5]) ? 3'b000 : 3'b000;

endmodule