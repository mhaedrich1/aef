module dtc_split5_bm34 (
	input  wire [9-1:0] inp,
	output wire [5-1:0] outp
);

	wire [5-1:0] node1;
	wire [5-1:0] node2;
	wire [5-1:0] node3;
	wire [5-1:0] node4;
	wire [5-1:0] node5;
	wire [5-1:0] node6;
	wire [5-1:0] node8;
	wire [5-1:0] node10;
	wire [5-1:0] node13;
	wire [5-1:0] node14;
	wire [5-1:0] node16;
	wire [5-1:0] node19;
	wire [5-1:0] node22;
	wire [5-1:0] node23;
	wire [5-1:0] node24;
	wire [5-1:0] node27;
	wire [5-1:0] node30;
	wire [5-1:0] node31;
	wire [5-1:0] node33;
	wire [5-1:0] node37;
	wire [5-1:0] node38;
	wire [5-1:0] node39;
	wire [5-1:0] node40;
	wire [5-1:0] node42;
	wire [5-1:0] node45;
	wire [5-1:0] node49;
	wire [5-1:0] node50;
	wire [5-1:0] node51;
	wire [5-1:0] node53;
	wire [5-1:0] node56;
	wire [5-1:0] node57;
	wire [5-1:0] node61;
	wire [5-1:0] node62;
	wire [5-1:0] node65;
	wire [5-1:0] node67;
	wire [5-1:0] node70;
	wire [5-1:0] node71;
	wire [5-1:0] node72;
	wire [5-1:0] node73;
	wire [5-1:0] node75;
	wire [5-1:0] node78;
	wire [5-1:0] node79;
	wire [5-1:0] node80;
	wire [5-1:0] node85;
	wire [5-1:0] node86;
	wire [5-1:0] node87;
	wire [5-1:0] node90;
	wire [5-1:0] node92;
	wire [5-1:0] node95;
	wire [5-1:0] node97;
	wire [5-1:0] node99;
	wire [5-1:0] node102;
	wire [5-1:0] node103;
	wire [5-1:0] node104;
	wire [5-1:0] node105;
	wire [5-1:0] node108;
	wire [5-1:0] node109;
	wire [5-1:0] node113;
	wire [5-1:0] node114;
	wire [5-1:0] node117;
	wire [5-1:0] node118;
	wire [5-1:0] node121;
	wire [5-1:0] node124;
	wire [5-1:0] node125;
	wire [5-1:0] node127;
	wire [5-1:0] node130;
	wire [5-1:0] node131;
	wire [5-1:0] node133;
	wire [5-1:0] node137;
	wire [5-1:0] node138;
	wire [5-1:0] node139;
	wire [5-1:0] node140;
	wire [5-1:0] node141;
	wire [5-1:0] node143;
	wire [5-1:0] node146;
	wire [5-1:0] node149;
	wire [5-1:0] node150;
	wire [5-1:0] node151;
	wire [5-1:0] node154;
	wire [5-1:0] node157;
	wire [5-1:0] node160;
	wire [5-1:0] node162;
	wire [5-1:0] node164;
	wire [5-1:0] node165;
	wire [5-1:0] node166;
	wire [5-1:0] node170;
	wire [5-1:0] node173;
	wire [5-1:0] node174;
	wire [5-1:0] node175;
	wire [5-1:0] node176;
	wire [5-1:0] node177;
	wire [5-1:0] node180;
	wire [5-1:0] node182;
	wire [5-1:0] node185;
	wire [5-1:0] node186;
	wire [5-1:0] node188;
	wire [5-1:0] node192;
	wire [5-1:0] node193;
	wire [5-1:0] node194;
	wire [5-1:0] node196;
	wire [5-1:0] node199;
	wire [5-1:0] node202;
	wire [5-1:0] node203;
	wire [5-1:0] node206;
	wire [5-1:0] node209;
	wire [5-1:0] node210;
	wire [5-1:0] node211;
	wire [5-1:0] node213;
	wire [5-1:0] node215;
	wire [5-1:0] node218;
	wire [5-1:0] node219;
	wire [5-1:0] node222;
	wire [5-1:0] node224;
	wire [5-1:0] node227;
	wire [5-1:0] node228;
	wire [5-1:0] node229;
	wire [5-1:0] node233;
	wire [5-1:0] node234;
	wire [5-1:0] node236;
	wire [5-1:0] node239;
	wire [5-1:0] node240;
	wire [5-1:0] node243;
	wire [5-1:0] node246;
	wire [5-1:0] node247;
	wire [5-1:0] node248;
	wire [5-1:0] node249;
	wire [5-1:0] node250;
	wire [5-1:0] node251;
	wire [5-1:0] node252;
	wire [5-1:0] node255;
	wire [5-1:0] node258;
	wire [5-1:0] node259;
	wire [5-1:0] node263;
	wire [5-1:0] node264;
	wire [5-1:0] node266;
	wire [5-1:0] node268;
	wire [5-1:0] node271;
	wire [5-1:0] node274;
	wire [5-1:0] node275;
	wire [5-1:0] node276;
	wire [5-1:0] node277;
	wire [5-1:0] node278;
	wire [5-1:0] node283;
	wire [5-1:0] node285;
	wire [5-1:0] node288;
	wire [5-1:0] node289;
	wire [5-1:0] node290;
	wire [5-1:0] node294;
	wire [5-1:0] node297;
	wire [5-1:0] node298;
	wire [5-1:0] node300;
	wire [5-1:0] node302;
	wire [5-1:0] node305;
	wire [5-1:0] node306;
	wire [5-1:0] node308;
	wire [5-1:0] node309;
	wire [5-1:0] node311;
	wire [5-1:0] node314;
	wire [5-1:0] node316;
	wire [5-1:0] node319;
	wire [5-1:0] node320;
	wire [5-1:0] node321;
	wire [5-1:0] node324;
	wire [5-1:0] node326;
	wire [5-1:0] node329;
	wire [5-1:0] node332;
	wire [5-1:0] node333;
	wire [5-1:0] node334;
	wire [5-1:0] node335;
	wire [5-1:0] node336;
	wire [5-1:0] node337;
	wire [5-1:0] node340;
	wire [5-1:0] node343;
	wire [5-1:0] node344;
	wire [5-1:0] node347;
	wire [5-1:0] node350;
	wire [5-1:0] node351;
	wire [5-1:0] node354;
	wire [5-1:0] node355;
	wire [5-1:0] node359;
	wire [5-1:0] node360;
	wire [5-1:0] node361;
	wire [5-1:0] node363;
	wire [5-1:0] node366;
	wire [5-1:0] node367;
	wire [5-1:0] node369;
	wire [5-1:0] node373;
	wire [5-1:0] node374;
	wire [5-1:0] node375;
	wire [5-1:0] node378;
	wire [5-1:0] node379;
	wire [5-1:0] node383;
	wire [5-1:0] node384;
	wire [5-1:0] node385;
	wire [5-1:0] node389;
	wire [5-1:0] node391;
	wire [5-1:0] node394;
	wire [5-1:0] node395;
	wire [5-1:0] node396;
	wire [5-1:0] node398;
	wire [5-1:0] node401;
	wire [5-1:0] node402;
	wire [5-1:0] node405;
	wire [5-1:0] node406;
	wire [5-1:0] node407;
	wire [5-1:0] node412;
	wire [5-1:0] node413;
	wire [5-1:0] node414;
	wire [5-1:0] node416;
	wire [5-1:0] node417;
	wire [5-1:0] node420;
	wire [5-1:0] node424;
	wire [5-1:0] node425;
	wire [5-1:0] node426;
	wire [5-1:0] node427;
	wire [5-1:0] node430;
	wire [5-1:0] node434;
	wire [5-1:0] node435;
	wire [5-1:0] node436;
	wire [5-1:0] node440;

	assign outp = (inp[2]) ? node246 : node1;
		assign node1 = (inp[0]) ? node137 : node2;
			assign node2 = (inp[8]) ? node70 : node3;
				assign node3 = (inp[5]) ? node37 : node4;
					assign node4 = (inp[6]) ? node22 : node5;
						assign node5 = (inp[1]) ? node13 : node6;
							assign node6 = (inp[4]) ? node8 : 5'b00111;
								assign node8 = (inp[3]) ? node10 : 5'b00111;
									assign node10 = (inp[7]) ? 5'b01110 : 5'b00110;
							assign node13 = (inp[7]) ? node19 : node14;
								assign node14 = (inp[3]) ? node16 : 5'b11011;
									assign node16 = (inp[4]) ? 5'b11011 : 5'b10110;
								assign node19 = (inp[3]) ? 5'b11110 : 5'b10110;
						assign node22 = (inp[1]) ? node30 : node23;
							assign node23 = (inp[7]) ? node27 : node24;
								assign node24 = (inp[4]) ? 5'b10110 : 5'b10111;
								assign node27 = (inp[4]) ? 5'b10111 : 5'b11110;
							assign node30 = (inp[7]) ? 5'b00111 : node31;
								assign node31 = (inp[3]) ? node33 : 5'b00110;
									assign node33 = (inp[4]) ? 5'b00110 : 5'b00111;
					assign node37 = (inp[7]) ? node49 : node38;
						assign node38 = (inp[3]) ? 5'b11010 : node39;
							assign node39 = (inp[4]) ? node45 : node40;
								assign node40 = (inp[6]) ? node42 : 5'b10011;
									assign node42 = (inp[1]) ? 5'b01010 : 5'b11010;
								assign node45 = (inp[6]) ? 5'b10011 : 5'b00011;
						assign node49 = (inp[3]) ? node61 : node50;
							assign node50 = (inp[4]) ? node56 : node51;
								assign node51 = (inp[1]) ? node53 : 5'b00110;
									assign node53 = (inp[6]) ? 5'b00110 : 5'b11011;
								assign node56 = (inp[1]) ? 5'b11010 : node57;
									assign node57 = (inp[6]) ? 5'b11011 : 5'b01011;
							assign node61 = (inp[1]) ? node65 : node62;
								assign node62 = (inp[6]) ? 5'b10110 : 5'b00110;
								assign node65 = (inp[6]) ? node67 : 5'b11011;
									assign node67 = (inp[4]) ? 5'b00110 : 5'b00111;
				assign node70 = (inp[7]) ? node102 : node71;
					assign node71 = (inp[5]) ? node85 : node72;
						assign node72 = (inp[6]) ? node78 : node73;
							assign node73 = (inp[3]) ? node75 : 5'b01000;
								assign node75 = (inp[4]) ? 5'b00001 : 5'b01000;
							assign node78 = (inp[1]) ? 5'b00001 : node79;
								assign node79 = (inp[3]) ? 5'b10001 : node80;
									assign node80 = (inp[4]) ? 5'b10001 : 5'b11000;
						assign node85 = (inp[4]) ? node95 : node86;
							assign node86 = (inp[3]) ? node90 : node87;
								assign node87 = (inp[6]) ? 5'b00000 : 5'b10000;
								assign node90 = (inp[1]) ? node92 : 5'b00000;
									assign node92 = (inp[6]) ? 5'b01111 : 5'b11111;
							assign node95 = (inp[1]) ? node97 : 5'b01111;
								assign node97 = (inp[3]) ? node99 : 5'b01111;
									assign node99 = (inp[6]) ? 5'b01110 : 5'b11110;
					assign node102 = (inp[1]) ? node124 : node103;
						assign node103 = (inp[6]) ? node113 : node104;
							assign node104 = (inp[5]) ? node108 : node105;
								assign node105 = (inp[3]) ? 5'b00000 : 5'b00001;
								assign node108 = (inp[3]) ? 5'b00111 : node109;
									assign node109 = (inp[4]) ? 5'b01110 : 5'b01111;
							assign node113 = (inp[5]) ? node117 : node114;
								assign node114 = (inp[3]) ? 5'b11110 : 5'b10000;
								assign node117 = (inp[4]) ? node121 : node118;
									assign node118 = (inp[3]) ? 5'b10111 : 5'b11110;
									assign node121 = (inp[3]) ? 5'b10110 : 5'b10111;
						assign node124 = (inp[6]) ? node130 : node125;
							assign node125 = (inp[3]) ? node127 : 5'b11111;
								assign node127 = (inp[4]) ? 5'b11110 : 5'b11111;
							assign node130 = (inp[5]) ? 5'b00111 : node131;
								assign node131 = (inp[4]) ? node133 : 5'b01111;
									assign node133 = (inp[3]) ? 5'b01110 : 5'b01111;
			assign node137 = (inp[8]) ? node173 : node138;
				assign node138 = (inp[5]) ? node160 : node139;
					assign node139 = (inp[3]) ? node149 : node140;
						assign node140 = (inp[7]) ? node146 : node141;
							assign node141 = (inp[6]) ? node143 : 5'b00010;
								assign node143 = (inp[1]) ? 5'b00010 : 5'b10010;
							assign node146 = (inp[1]) ? 5'b10010 : 5'b00011;
						assign node149 = (inp[4]) ? node157 : node150;
							assign node150 = (inp[6]) ? node154 : node151;
								assign node151 = (inp[1]) ? 5'b11010 : 5'b01011;
								assign node154 = (inp[1]) ? 5'b01011 : 5'b11011;
							assign node157 = (inp[1]) ? 5'b01010 : 5'b11010;
					assign node160 = (inp[7]) ? node162 : 5'b00010;
						assign node162 = (inp[3]) ? node164 : 5'b00010;
							assign node164 = (inp[4]) ? node170 : node165;
								assign node165 = (inp[1]) ? 5'b00011 : node166;
									assign node166 = (inp[6]) ? 5'b10011 : 5'b00011;
								assign node170 = (inp[1]) ? 5'b00010 : 5'b10010;
				assign node173 = (inp[7]) ? node209 : node174;
					assign node174 = (inp[5]) ? node192 : node175;
						assign node175 = (inp[3]) ? node185 : node176;
							assign node176 = (inp[4]) ? node180 : node177;
								assign node177 = (inp[1]) ? 5'b01110 : 5'b01111;
								assign node180 = (inp[6]) ? node182 : 5'b01110;
									assign node182 = (inp[1]) ? 5'b00111 : 5'b10111;
							assign node185 = (inp[6]) ? 5'b00110 : node186;
								assign node186 = (inp[1]) ? node188 : 5'b00111;
									assign node188 = (inp[4]) ? 5'b10110 : 5'b10111;
						assign node192 = (inp[3]) ? node202 : node193;
							assign node193 = (inp[4]) ? node199 : node194;
								assign node194 = (inp[6]) ? node196 : 5'b10110;
									assign node196 = (inp[1]) ? 5'b00110 : 5'b10110;
								assign node199 = (inp[1]) ? 5'b11011 : 5'b00110;
							assign node202 = (inp[1]) ? node206 : node203;
								assign node203 = (inp[6]) ? 5'b11011 : 5'b01011;
								assign node206 = (inp[6]) ? 5'b01010 : 5'b11010;
					assign node209 = (inp[5]) ? node227 : node210;
						assign node210 = (inp[4]) ? node218 : node211;
							assign node211 = (inp[3]) ? node213 : 5'b00110;
								assign node213 = (inp[6]) ? node215 : 5'b00110;
									assign node215 = (inp[1]) ? 5'b01011 : 5'b11011;
							assign node218 = (inp[6]) ? node222 : node219;
								assign node219 = (inp[1]) ? 5'b11011 : 5'b01011;
								assign node222 = (inp[3]) ? node224 : 5'b01011;
									assign node224 = (inp[1]) ? 5'b01010 : 5'b11010;
						assign node227 = (inp[3]) ? node233 : node228;
							assign node228 = (inp[4]) ? 5'b10011 : node229;
								assign node229 = (inp[1]) ? 5'b01010 : 5'b11010;
							assign node233 = (inp[4]) ? node239 : node234;
								assign node234 = (inp[6]) ? node236 : 5'b10011;
									assign node236 = (inp[1]) ? 5'b00011 : 5'b10011;
								assign node239 = (inp[6]) ? node243 : node240;
									assign node240 = (inp[1]) ? 5'b10010 : 5'b00011;
									assign node243 = (inp[1]) ? 5'b00010 : 5'b10010;
		assign node246 = (inp[0]) ? node332 : node247;
			assign node247 = (inp[8]) ? node297 : node248;
				assign node248 = (inp[5]) ? node274 : node249;
					assign node249 = (inp[7]) ? node263 : node250;
						assign node250 = (inp[3]) ? node258 : node251;
							assign node251 = (inp[6]) ? node255 : node252;
								assign node252 = (inp[4]) ? 5'b11000 : 5'b11001;
								assign node255 = (inp[4]) ? 5'b01001 : 5'b00100;
							assign node258 = (inp[4]) ? 5'b10100 : node259;
								assign node259 = (inp[6]) ? 5'b00101 : 5'b10100;
						assign node263 = (inp[6]) ? node271 : node264;
							assign node264 = (inp[1]) ? node266 : 5'b00101;
								assign node266 = (inp[4]) ? node268 : 5'b10101;
									assign node268 = (inp[3]) ? 5'b10101 : 5'b10100;
							assign node271 = (inp[4]) ? 5'b11100 : 5'b11101;
					assign node274 = (inp[7]) ? node288 : node275;
						assign node275 = (inp[4]) ? node283 : node276;
							assign node276 = (inp[6]) ? 5'b01001 : node277;
								assign node277 = (inp[1]) ? 5'b11000 : node278;
									assign node278 = (inp[3]) ? 5'b01001 : 5'b01000;
							assign node283 = (inp[1]) ? node285 : 5'b00001;
								assign node285 = (inp[3]) ? 5'b10001 : 5'b10000;
						assign node288 = (inp[6]) ? node294 : node289;
							assign node289 = (inp[1]) ? 5'b11000 : node290;
								assign node290 = (inp[4]) ? 5'b01001 : 5'b00101;
							assign node294 = (inp[1]) ? 5'b00100 : 5'b10100;
				assign node297 = (inp[7]) ? node305 : node298;
					assign node298 = (inp[3]) ? node300 : 5'b11101;
						assign node300 = (inp[4]) ? node302 : 5'b11101;
							assign node302 = (inp[1]) ? 5'b11100 : 5'b01101;
					assign node305 = (inp[5]) ? node319 : node306;
						assign node306 = (inp[3]) ? node308 : 5'b11101;
							assign node308 = (inp[4]) ? node314 : node309;
								assign node309 = (inp[6]) ? node311 : 5'b11101;
									assign node311 = (inp[1]) ? 5'b01101 : 5'b11101;
								assign node314 = (inp[1]) ? node316 : 5'b11100;
									assign node316 = (inp[6]) ? 5'b01100 : 5'b11100;
						assign node319 = (inp[6]) ? node329 : node320;
							assign node320 = (inp[1]) ? node324 : node321;
								assign node321 = (inp[3]) ? 5'b00101 : 5'b01101;
								assign node324 = (inp[3]) ? node326 : 5'b11100;
									assign node326 = (inp[4]) ? 5'b10100 : 5'b10101;
							assign node329 = (inp[1]) ? 5'b00101 : 5'b10101;
			assign node332 = (inp[7]) ? node394 : node333;
				assign node333 = (inp[8]) ? node359 : node334;
					assign node334 = (inp[5]) ? node350 : node335;
						assign node335 = (inp[3]) ? node343 : node336;
							assign node336 = (inp[4]) ? node340 : node337;
								assign node337 = (inp[1]) ? 5'b11111 : 5'b10000;
								assign node340 = (inp[6]) ? 5'b11111 : 5'b01111;
							assign node343 = (inp[1]) ? node347 : node344;
								assign node344 = (inp[6]) ? 5'b10001 : 5'b00001;
								assign node347 = (inp[4]) ? 5'b00000 : 5'b10000;
						assign node350 = (inp[1]) ? node354 : node351;
							assign node351 = (inp[6]) ? 5'b11111 : 5'b01110;
							assign node354 = (inp[3]) ? 5'b10111 : node355;
								assign node355 = (inp[4]) ? 5'b10110 : 5'b10111;
					assign node359 = (inp[5]) ? node373 : node360;
						assign node360 = (inp[4]) ? node366 : node361;
							assign node361 = (inp[6]) ? node363 : 5'b10101;
								assign node363 = (inp[1]) ? 5'b01100 : 5'b11100;
							assign node366 = (inp[3]) ? 5'b10100 : node367;
								assign node367 = (inp[1]) ? node369 : 5'b10101;
									assign node369 = (inp[6]) ? 5'b00101 : 5'b10101;
						assign node373 = (inp[4]) ? node383 : node374;
							assign node374 = (inp[3]) ? node378 : node375;
								assign node375 = (inp[6]) ? 5'b00100 : 5'b00101;
								assign node378 = (inp[1]) ? 5'b11001 : node379;
									assign node379 = (inp[6]) ? 5'b11001 : 5'b00100;
							assign node383 = (inp[3]) ? node389 : node384;
								assign node384 = (inp[6]) ? 5'b11001 : node385;
									assign node385 = (inp[1]) ? 5'b11001 : 5'b00100;
								assign node389 = (inp[6]) ? node391 : 5'b11000;
									assign node391 = (inp[1]) ? 5'b01000 : 5'b11000;
				assign node394 = (inp[1]) ? node412 : node395;
					assign node395 = (inp[5]) ? node401 : node396;
						assign node396 = (inp[4]) ? node398 : 5'b11001;
							assign node398 = (inp[3]) ? 5'b11000 : 5'b11001;
						assign node401 = (inp[6]) ? node405 : node402;
							assign node402 = (inp[8]) ? 5'b00001 : 5'b00000;
							assign node405 = (inp[8]) ? 5'b10001 : node406;
								assign node406 = (inp[4]) ? 5'b10000 : node407;
									assign node407 = (inp[3]) ? 5'b10001 : 5'b10000;
					assign node412 = (inp[6]) ? node424 : node413;
						assign node413 = (inp[5]) ? 5'b11111 : node414;
							assign node414 = (inp[3]) ? node416 : 5'b10000;
								assign node416 = (inp[4]) ? node420 : node417;
									assign node417 = (inp[8]) ? 5'b11001 : 5'b11000;
									assign node420 = (inp[8]) ? 5'b11000 : 5'b10001;
						assign node424 = (inp[4]) ? node434 : node425;
							assign node425 = (inp[3]) ? 5'b01001 : node426;
								assign node426 = (inp[5]) ? node430 : node427;
									assign node427 = (inp[8]) ? 5'b00100 : 5'b01000;
									assign node430 = (inp[8]) ? 5'b01000 : 5'b00000;
							assign node434 = (inp[3]) ? node440 : node435;
								assign node435 = (inp[5]) ? 5'b01111 : node436;
									assign node436 = (inp[8]) ? 5'b01001 : 5'b00001;
								assign node440 = (inp[8]) ? 5'b00000 : 5'b01000;

endmodule