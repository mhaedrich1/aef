module dtc_split75_bm47 (
	input  wire [16-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node6;
	wire [1-1:0] node7;
	wire [1-1:0] node8;
	wire [1-1:0] node9;
	wire [1-1:0] node11;
	wire [1-1:0] node14;
	wire [1-1:0] node15;
	wire [1-1:0] node19;
	wire [1-1:0] node21;
	wire [1-1:0] node25;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node28;
	wire [1-1:0] node29;
	wire [1-1:0] node33;
	wire [1-1:0] node34;
	wire [1-1:0] node36;
	wire [1-1:0] node39;
	wire [1-1:0] node40;
	wire [1-1:0] node44;
	wire [1-1:0] node46;
	wire [1-1:0] node47;
	wire [1-1:0] node48;
	wire [1-1:0] node49;
	wire [1-1:0] node53;
	wire [1-1:0] node54;
	wire [1-1:0] node58;
	wire [1-1:0] node59;
	wire [1-1:0] node63;
	wire [1-1:0] node65;
	wire [1-1:0] node66;
	wire [1-1:0] node67;
	wire [1-1:0] node68;
	wire [1-1:0] node70;
	wire [1-1:0] node73;
	wire [1-1:0] node74;
	wire [1-1:0] node78;
	wire [1-1:0] node80;
	wire [1-1:0] node84;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node87;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node90;
	wire [1-1:0] node92;
	wire [1-1:0] node93;
	wire [1-1:0] node94;
	wire [1-1:0] node96;
	wire [1-1:0] node99;
	wire [1-1:0] node101;
	wire [1-1:0] node104;
	wire [1-1:0] node105;
	wire [1-1:0] node110;
	wire [1-1:0] node111;
	wire [1-1:0] node112;
	wire [1-1:0] node113;
	wire [1-1:0] node114;
	wire [1-1:0] node115;
	wire [1-1:0] node119;
	wire [1-1:0] node120;
	wire [1-1:0] node124;
	wire [1-1:0] node126;
	wire [1-1:0] node130;
	wire [1-1:0] node131;
	wire [1-1:0] node133;
	wire [1-1:0] node136;
	wire [1-1:0] node137;
	wire [1-1:0] node138;
	wire [1-1:0] node142;
	wire [1-1:0] node143;
	wire [1-1:0] node147;
	wire [1-1:0] node149;
	wire [1-1:0] node150;
	wire [1-1:0] node151;
	wire [1-1:0] node152;
	wire [1-1:0] node156;
	wire [1-1:0] node157;
	wire [1-1:0] node159;
	wire [1-1:0] node162;
	wire [1-1:0] node163;
	wire [1-1:0] node168;
	wire [1-1:0] node169;
	wire [1-1:0] node170;
	wire [1-1:0] node171;
	wire [1-1:0] node173;
	wire [1-1:0] node174;
	wire [1-1:0] node175;
	wire [1-1:0] node177;
	wire [1-1:0] node180;
	wire [1-1:0] node181;
	wire [1-1:0] node182;
	wire [1-1:0] node186;
	wire [1-1:0] node188;
	wire [1-1:0] node192;
	wire [1-1:0] node193;
	wire [1-1:0] node194;
	wire [1-1:0] node195;
	wire [1-1:0] node196;
	wire [1-1:0] node200;
	wire [1-1:0] node201;
	wire [1-1:0] node202;
	wire [1-1:0] node206;
	wire [1-1:0] node207;
	wire [1-1:0] node212;
	wire [1-1:0] node213;
	wire [1-1:0] node214;
	wire [1-1:0] node218;
	wire [1-1:0] node219;
	wire [1-1:0] node220;
	wire [1-1:0] node224;
	wire [1-1:0] node226;
	wire [1-1:0] node229;
	wire [1-1:0] node231;
	wire [1-1:0] node232;
	wire [1-1:0] node233;
	wire [1-1:0] node234;
	wire [1-1:0] node235;
	wire [1-1:0] node239;
	wire [1-1:0] node240;
	wire [1-1:0] node244;
	wire [1-1:0] node245;
	wire [1-1:0] node250;
	wire [1-1:0] node251;
	wire [1-1:0] node252;
	wire [1-1:0] node254;
	wire [1-1:0] node255;
	wire [1-1:0] node256;
	wire [1-1:0] node260;
	wire [1-1:0] node261;
	wire [1-1:0] node263;
	wire [1-1:0] node266;
	wire [1-1:0] node267;
	wire [1-1:0] node272;
	wire [1-1:0] node273;
	wire [1-1:0] node274;
	wire [1-1:0] node275;
	wire [1-1:0] node276;
	wire [1-1:0] node278;
	wire [1-1:0] node281;
	wire [1-1:0] node283;
	wire [1-1:0] node286;
	wire [1-1:0] node287;
	wire [1-1:0] node291;
	wire [1-1:0] node293;
	wire [1-1:0] node295;
	wire [1-1:0] node296;
	wire [1-1:0] node297;
	wire [1-1:0] node301;
	wire [1-1:0] node302;
	wire [1-1:0] node306;
	wire [1-1:0] node307;
	wire [1-1:0] node309;
	wire [1-1:0] node310;
	wire [1-1:0] node311;
	wire [1-1:0] node313;
	wire [1-1:0] node316;
	wire [1-1:0] node317;
	wire [1-1:0] node320;
	wire [1-1:0] node322;
	wire [1-1:0] node325;
	wire [1-1:0] node326;
	wire [1-1:0] node331;
	wire [1-1:0] node332;
	wire [1-1:0] node333;
	wire [1-1:0] node334;
	wire [1-1:0] node335;
	wire [1-1:0] node336;
	wire [1-1:0] node338;
	wire [1-1:0] node339;
	wire [1-1:0] node340;
	wire [1-1:0] node341;
	wire [1-1:0] node347;
	wire [1-1:0] node348;
	wire [1-1:0] node349;
	wire [1-1:0] node350;
	wire [1-1:0] node351;
	wire [1-1:0] node355;
	wire [1-1:0] node356;
	wire [1-1:0] node360;
	wire [1-1:0] node362;
	wire [1-1:0] node365;
	wire [1-1:0] node367;
	wire [1-1:0] node368;
	wire [1-1:0] node369;
	wire [1-1:0] node373;
	wire [1-1:0] node374;
	wire [1-1:0] node375;
	wire [1-1:0] node378;
	wire [1-1:0] node382;
	wire [1-1:0] node384;
	wire [1-1:0] node385;
	wire [1-1:0] node386;
	wire [1-1:0] node387;
	wire [1-1:0] node391;
	wire [1-1:0] node392;
	wire [1-1:0] node393;
	wire [1-1:0] node397;
	wire [1-1:0] node398;
	wire [1-1:0] node403;
	wire [1-1:0] node404;
	wire [1-1:0] node406;
	wire [1-1:0] node407;
	wire [1-1:0] node408;
	wire [1-1:0] node410;
	wire [1-1:0] node413;
	wire [1-1:0] node414;
	wire [1-1:0] node415;
	wire [1-1:0] node418;
	wire [1-1:0] node423;
	wire [1-1:0] node424;
	wire [1-1:0] node425;
	wire [1-1:0] node426;
	wire [1-1:0] node427;
	wire [1-1:0] node429;
	wire [1-1:0] node432;
	wire [1-1:0] node433;
	wire [1-1:0] node437;
	wire [1-1:0] node439;
	wire [1-1:0] node442;
	wire [1-1:0] node444;
	wire [1-1:0] node445;
	wire [1-1:0] node447;
	wire [1-1:0] node450;
	wire [1-1:0] node451;
	wire [1-1:0] node455;
	wire [1-1:0] node456;
	wire [1-1:0] node458;
	wire [1-1:0] node459;
	wire [1-1:0] node460;
	wire [1-1:0] node464;
	wire [1-1:0] node465;
	wire [1-1:0] node467;
	wire [1-1:0] node470;
	wire [1-1:0] node474;
	wire [1-1:0] node475;
	wire [1-1:0] node476;
	wire [1-1:0] node477;
	wire [1-1:0] node479;
	wire [1-1:0] node480;
	wire [1-1:0] node481;
	wire [1-1:0] node485;
	wire [1-1:0] node486;
	wire [1-1:0] node488;
	wire [1-1:0] node491;
	wire [1-1:0] node495;
	wire [1-1:0] node496;
	wire [1-1:0] node497;
	wire [1-1:0] node499;
	wire [1-1:0] node502;
	wire [1-1:0] node503;
	wire [1-1:0] node505;
	wire [1-1:0] node508;
	wire [1-1:0] node509;
	wire [1-1:0] node513;
	wire [1-1:0] node515;
	wire [1-1:0] node516;
	wire [1-1:0] node518;
	wire [1-1:0] node521;
	wire [1-1:0] node522;
	wire [1-1:0] node524;
	wire [1-1:0] node525;
	wire [1-1:0] node529;
	wire [1-1:0] node531;
	wire [1-1:0] node534;
	wire [1-1:0] node536;
	wire [1-1:0] node537;
	wire [1-1:0] node538;
	wire [1-1:0] node539;
	wire [1-1:0] node543;
	wire [1-1:0] node544;
	wire [1-1:0] node546;
	wire [1-1:0] node549;
	wire [1-1:0] node551;
	wire [1-1:0] node555;
	wire [1-1:0] node556;
	wire [1-1:0] node557;
	wire [1-1:0] node558;
	wire [1-1:0] node559;
	wire [1-1:0] node561;
	wire [1-1:0] node562;
	wire [1-1:0] node564;
	wire [1-1:0] node565;
	wire [1-1:0] node567;
	wire [1-1:0] node570;
	wire [1-1:0] node571;
	wire [1-1:0] node576;
	wire [1-1:0] node577;
	wire [1-1:0] node578;
	wire [1-1:0] node580;
	wire [1-1:0] node583;
	wire [1-1:0] node584;
	wire [1-1:0] node585;
	wire [1-1:0] node589;
	wire [1-1:0] node590;
	wire [1-1:0] node594;
	wire [1-1:0] node596;
	wire [1-1:0] node597;
	wire [1-1:0] node598;
	wire [1-1:0] node600;
	wire [1-1:0] node603;
	wire [1-1:0] node607;
	wire [1-1:0] node609;
	wire [1-1:0] node610;
	wire [1-1:0] node611;
	wire [1-1:0] node612;
	wire [1-1:0] node613;
	wire [1-1:0] node617;
	wire [1-1:0] node618;
	wire [1-1:0] node622;
	wire [1-1:0] node624;
	wire [1-1:0] node628;
	wire [1-1:0] node629;
	wire [1-1:0] node630;
	wire [1-1:0] node631;
	wire [1-1:0] node633;
	wire [1-1:0] node634;
	wire [1-1:0] node635;
	wire [1-1:0] node637;
	wire [1-1:0] node640;
	wire [1-1:0] node643;
	wire [1-1:0] node644;
	wire [1-1:0] node649;
	wire [1-1:0] node650;
	wire [1-1:0] node651;
	wire [1-1:0] node653;
	wire [1-1:0] node656;
	wire [1-1:0] node657;
	wire [1-1:0] node659;
	wire [1-1:0] node662;
	wire [1-1:0] node663;
	wire [1-1:0] node667;
	wire [1-1:0] node669;
	wire [1-1:0] node670;
	wire [1-1:0] node672;
	wire [1-1:0] node675;
	wire [1-1:0] node676;
	wire [1-1:0] node678;
	wire [1-1:0] node681;
	wire [1-1:0] node682;
	wire [1-1:0] node686;
	wire [1-1:0] node688;
	wire [1-1:0] node689;
	wire [1-1:0] node690;
	wire [1-1:0] node691;
	wire [1-1:0] node694;
	wire [1-1:0] node696;
	wire [1-1:0] node699;
	wire [1-1:0] node700;
	wire [1-1:0] node705;
	wire [1-1:0] node706;
	wire [1-1:0] node708;
	wire [1-1:0] node709;
	wire [1-1:0] node710;
	wire [1-1:0] node711;
	wire [1-1:0] node713;
	wire [1-1:0] node716;
	wire [1-1:0] node718;
	wire [1-1:0] node721;
	wire [1-1:0] node722;
	wire [1-1:0] node727;
	wire [1-1:0] node728;
	wire [1-1:0] node729;
	wire [1-1:0] node730;
	wire [1-1:0] node731;
	wire [1-1:0] node732;
	wire [1-1:0] node733;
	wire [1-1:0] node737;
	wire [1-1:0] node739;
	wire [1-1:0] node742;
	wire [1-1:0] node744;
	wire [1-1:0] node748;
	wire [1-1:0] node749;
	wire [1-1:0] node750;
	wire [1-1:0] node754;
	wire [1-1:0] node755;
	wire [1-1:0] node756;
	wire [1-1:0] node760;
	wire [1-1:0] node761;
	wire [1-1:0] node765;
	wire [1-1:0] node767;
	wire [1-1:0] node768;
	wire [1-1:0] node769;
	wire [1-1:0] node771;
	wire [1-1:0] node774;
	wire [1-1:0] node775;
	wire [1-1:0] node776;
	wire [1-1:0] node777;
	wire [1-1:0] node781;
	wire [1-1:0] node782;
	wire [1-1:0] node785;
	wire [1-1:0] node790;
	wire [1-1:0] node791;
	wire [1-1:0] node792;
	wire [1-1:0] node794;
	wire [1-1:0] node795;
	wire [1-1:0] node796;
	wire [1-1:0] node798;
	wire [1-1:0] node801;
	wire [1-1:0] node802;
	wire [1-1:0] node803;
	wire [1-1:0] node807;
	wire [1-1:0] node809;
	wire [1-1:0] node813;
	wire [1-1:0] node814;
	wire [1-1:0] node815;
	wire [1-1:0] node816;
	wire [1-1:0] node817;
	wire [1-1:0] node819;
	wire [1-1:0] node822;
	wire [1-1:0] node824;
	wire [1-1:0] node827;
	wire [1-1:0] node828;
	wire [1-1:0] node833;
	wire [1-1:0] node834;
	wire [1-1:0] node835;
	wire [1-1:0] node836;
	wire [1-1:0] node840;
	wire [1-1:0] node841;
	wire [1-1:0] node845;
	wire [1-1:0] node847;
	wire [1-1:0] node850;
	wire [1-1:0] node851;
	wire [1-1:0] node853;
	wire [1-1:0] node854;
	wire [1-1:0] node855;
	wire [1-1:0] node859;
	wire [1-1:0] node860;
	wire [1-1:0] node862;
	wire [1-1:0] node865;
	wire [1-1:0] node866;
	wire [1-1:0] node871;
	wire [1-1:0] node872;
	wire [1-1:0] node873;
	wire [1-1:0] node874;
	wire [1-1:0] node875;
	wire [1-1:0] node876;
	wire [1-1:0] node877;
	wire [1-1:0] node878;
	wire [1-1:0] node880;
	wire [1-1:0] node881;
	wire [1-1:0] node882;
	wire [1-1:0] node883;
	wire [1-1:0] node887;
	wire [1-1:0] node888;
	wire [1-1:0] node890;
	wire [1-1:0] node893;
	wire [1-1:0] node895;
	wire [1-1:0] node899;
	wire [1-1:0] node900;
	wire [1-1:0] node901;
	wire [1-1:0] node902;
	wire [1-1:0] node903;
	wire [1-1:0] node904;
	wire [1-1:0] node908;
	wire [1-1:0] node909;
	wire [1-1:0] node913;
	wire [1-1:0] node915;
	wire [1-1:0] node919;
	wire [1-1:0] node920;
	wire [1-1:0] node921;
	wire [1-1:0] node922;
	wire [1-1:0] node926;
	wire [1-1:0] node927;
	wire [1-1:0] node931;
	wire [1-1:0] node932;
	wire [1-1:0] node936;
	wire [1-1:0] node938;
	wire [1-1:0] node939;
	wire [1-1:0] node940;
	wire [1-1:0] node941;
	wire [1-1:0] node942;
	wire [1-1:0] node946;
	wire [1-1:0] node947;
	wire [1-1:0] node951;
	wire [1-1:0] node953;
	wire [1-1:0] node957;
	wire [1-1:0] node958;
	wire [1-1:0] node959;
	wire [1-1:0] node960;
	wire [1-1:0] node962;
	wire [1-1:0] node963;
	wire [1-1:0] node964;
	wire [1-1:0] node966;
	wire [1-1:0] node967;
	wire [1-1:0] node970;
	wire [1-1:0] node975;
	wire [1-1:0] node976;
	wire [1-1:0] node977;
	wire [1-1:0] node978;
	wire [1-1:0] node979;
	wire [1-1:0] node983;
	wire [1-1:0] node985;
	wire [1-1:0] node989;
	wire [1-1:0] node990;
	wire [1-1:0] node991;
	wire [1-1:0] node992;
	wire [1-1:0] node995;
	wire [1-1:0] node998;
	wire [1-1:0] node1001;
	wire [1-1:0] node1002;
	wire [1-1:0] node1006;
	wire [1-1:0] node1007;
	wire [1-1:0] node1009;
	wire [1-1:0] node1010;
	wire [1-1:0] node1011;
	wire [1-1:0] node1012;
	wire [1-1:0] node1013;
	wire [1-1:0] node1016;
	wire [1-1:0] node1019;
	wire [1-1:0] node1020;
	wire [1-1:0] node1024;
	wire [1-1:0] node1027;
	wire [1-1:0] node1029;
	wire [1-1:0] node1033;
	wire [1-1:0] node1034;
	wire [1-1:0] node1036;
	wire [1-1:0] node1037;
	wire [1-1:0] node1038;
	wire [1-1:0] node1039;
	wire [1-1:0] node1043;
	wire [1-1:0] node1044;
	wire [1-1:0] node1045;
	wire [1-1:0] node1049;
	wire [1-1:0] node1053;
	wire [1-1:0] node1054;
	wire [1-1:0] node1055;
	wire [1-1:0] node1056;
	wire [1-1:0] node1058;
	wire [1-1:0] node1061;
	wire [1-1:0] node1062;
	wire [1-1:0] node1065;
	wire [1-1:0] node1067;
	wire [1-1:0] node1070;
	wire [1-1:0] node1072;
	wire [1-1:0] node1073;
	wire [1-1:0] node1075;
	wire [1-1:0] node1078;
	wire [1-1:0] node1080;
	wire [1-1:0] node1083;
	wire [1-1:0] node1084;
	wire [1-1:0] node1086;
	wire [1-1:0] node1087;
	wire [1-1:0] node1088;
	wire [1-1:0] node1089;
	wire [1-1:0] node1093;
	wire [1-1:0] node1098;
	wire [1-1:0] node1099;
	wire [1-1:0] node1100;
	wire [1-1:0] node1101;
	wire [1-1:0] node1102;
	wire [1-1:0] node1103;
	wire [1-1:0] node1105;
	wire [1-1:0] node1106;
	wire [1-1:0] node1107;
	wire [1-1:0] node1108;
	wire [1-1:0] node1112;
	wire [1-1:0] node1115;
	wire [1-1:0] node1117;
	wire [1-1:0] node1121;
	wire [1-1:0] node1122;
	wire [1-1:0] node1123;
	wire [1-1:0] node1124;
	wire [1-1:0] node1126;
	wire [1-1:0] node1129;
	wire [1-1:0] node1131;
	wire [1-1:0] node1132;
	wire [1-1:0] node1135;
	wire [1-1:0] node1139;
	wire [1-1:0] node1140;
	wire [1-1:0] node1141;
	wire [1-1:0] node1142;
	wire [1-1:0] node1146;
	wire [1-1:0] node1147;
	wire [1-1:0] node1151;
	wire [1-1:0] node1153;
	wire [1-1:0] node1156;
	wire [1-1:0] node1158;
	wire [1-1:0] node1159;
	wire [1-1:0] node1160;
	wire [1-1:0] node1161;
	wire [1-1:0] node1164;
	wire [1-1:0] node1165;
	wire [1-1:0] node1169;
	wire [1-1:0] node1170;
	wire [1-1:0] node1175;
	wire [1-1:0] node1176;
	wire [1-1:0] node1178;
	wire [1-1:0] node1179;
	wire [1-1:0] node1180;
	wire [1-1:0] node1181;
	wire [1-1:0] node1182;
	wire [1-1:0] node1186;
	wire [1-1:0] node1187;
	wire [1-1:0] node1191;
	wire [1-1:0] node1192;
	wire [1-1:0] node1197;
	wire [1-1:0] node1198;
	wire [1-1:0] node1199;
	wire [1-1:0] node1200;
	wire [1-1:0] node1201;
	wire [1-1:0] node1202;
	wire [1-1:0] node1206;
	wire [1-1:0] node1208;
	wire [1-1:0] node1211;
	wire [1-1:0] node1213;
	wire [1-1:0] node1216;
	wire [1-1:0] node1218;
	wire [1-1:0] node1219;
	wire [1-1:0] node1221;
	wire [1-1:0] node1222;
	wire [1-1:0] node1225;
	wire [1-1:0] node1228;
	wire [1-1:0] node1230;
	wire [1-1:0] node1233;
	wire [1-1:0] node1234;
	wire [1-1:0] node1236;
	wire [1-1:0] node1237;
	wire [1-1:0] node1238;
	wire [1-1:0] node1242;
	wire [1-1:0] node1243;
	wire [1-1:0] node1246;
	wire [1-1:0] node1247;
	wire [1-1:0] node1252;
	wire [1-1:0] node1253;
	wire [1-1:0] node1254;
	wire [1-1:0] node1256;
	wire [1-1:0] node1257;
	wire [1-1:0] node1258;
	wire [1-1:0] node1259;
	wire [1-1:0] node1263;
	wire [1-1:0] node1264;
	wire [1-1:0] node1268;
	wire [1-1:0] node1269;
	wire [1-1:0] node1274;
	wire [1-1:0] node1275;
	wire [1-1:0] node1276;
	wire [1-1:0] node1277;
	wire [1-1:0] node1278;
	wire [1-1:0] node1279;
	wire [1-1:0] node1280;
	wire [1-1:0] node1284;
	wire [1-1:0] node1286;
	wire [1-1:0] node1289;
	wire [1-1:0] node1290;
	wire [1-1:0] node1295;
	wire [1-1:0] node1296;
	wire [1-1:0] node1297;
	wire [1-1:0] node1298;
	wire [1-1:0] node1302;
	wire [1-1:0] node1303;
	wire [1-1:0] node1307;
	wire [1-1:0] node1309;
	wire [1-1:0] node1312;
	wire [1-1:0] node1313;
	wire [1-1:0] node1315;
	wire [1-1:0] node1316;
	wire [1-1:0] node1317;
	wire [1-1:0] node1321;
	wire [1-1:0] node1322;
	wire [1-1:0] node1324;
	wire [1-1:0] node1327;
	wire [1-1:0] node1329;
	wire [1-1:0] node1333;
	wire [1-1:0] node1334;
	wire [1-1:0] node1335;
	wire [1-1:0] node1337;
	wire [1-1:0] node1338;
	wire [1-1:0] node1339;
	wire [1-1:0] node1340;
	wire [1-1:0] node1341;
	wire [1-1:0] node1345;
	wire [1-1:0] node1347;
	wire [1-1:0] node1350;
	wire [1-1:0] node1351;
	wire [1-1:0] node1356;
	wire [1-1:0] node1357;
	wire [1-1:0] node1358;
	wire [1-1:0] node1359;
	wire [1-1:0] node1360;
	wire [1-1:0] node1361;
	wire [1-1:0] node1365;
	wire [1-1:0] node1366;
	wire [1-1:0] node1367;
	wire [1-1:0] node1371;
	wire [1-1:0] node1372;
	wire [1-1:0] node1377;
	wire [1-1:0] node1378;
	wire [1-1:0] node1380;
	wire [1-1:0] node1383;
	wire [1-1:0] node1384;
	wire [1-1:0] node1385;
	wire [1-1:0] node1389;
	wire [1-1:0] node1391;
	wire [1-1:0] node1394;
	wire [1-1:0] node1395;
	wire [1-1:0] node1397;
	wire [1-1:0] node1398;
	wire [1-1:0] node1399;
	wire [1-1:0] node1403;
	wire [1-1:0] node1404;
	wire [1-1:0] node1406;
	wire [1-1:0] node1409;
	wire [1-1:0] node1411;
	wire [1-1:0] node1415;
	wire [1-1:0] node1416;
	wire [1-1:0] node1417;
	wire [1-1:0] node1418;
	wire [1-1:0] node1420;
	wire [1-1:0] node1421;
	wire [1-1:0] node1422;
	wire [1-1:0] node1423;
	wire [1-1:0] node1427;
	wire [1-1:0] node1428;
	wire [1-1:0] node1432;
	wire [1-1:0] node1433;
	wire [1-1:0] node1438;
	wire [1-1:0] node1439;
	wire [1-1:0] node1440;
	wire [1-1:0] node1441;
	wire [1-1:0] node1442;
	wire [1-1:0] node1443;
	wire [1-1:0] node1444;
	wire [1-1:0] node1448;
	wire [1-1:0] node1450;
	wire [1-1:0] node1453;
	wire [1-1:0] node1454;
	wire [1-1:0] node1459;
	wire [1-1:0] node1460;
	wire [1-1:0] node1462;
	wire [1-1:0] node1465;
	wire [1-1:0] node1466;
	wire [1-1:0] node1468;
	wire [1-1:0] node1471;
	wire [1-1:0] node1473;
	wire [1-1:0] node1476;
	wire [1-1:0] node1478;
	wire [1-1:0] node1479;
	wire [1-1:0] node1480;
	wire [1-1:0] node1481;
	wire [1-1:0] node1484;
	wire [1-1:0] node1486;
	wire [1-1:0] node1489;
	wire [1-1:0] node1490;
	wire [1-1:0] node1495;
	wire [1-1:0] node1496;
	wire [1-1:0] node1497;
	wire [1-1:0] node1499;
	wire [1-1:0] node1500;
	wire [1-1:0] node1501;
	wire [1-1:0] node1502;
	wire [1-1:0] node1504;
	wire [1-1:0] node1507;
	wire [1-1:0] node1508;
	wire [1-1:0] node1512;
	wire [1-1:0] node1513;
	wire [1-1:0] node1518;
	wire [1-1:0] node1519;
	wire [1-1:0] node1520;
	wire [1-1:0] node1521;
	wire [1-1:0] node1525;
	wire [1-1:0] node1526;
	wire [1-1:0] node1528;
	wire [1-1:0] node1531;
	wire [1-1:0] node1533;
	wire [1-1:0] node1536;
	wire [1-1:0] node1538;
	wire [1-1:0] node1539;
	wire [1-1:0] node1540;
	wire [1-1:0] node1542;
	wire [1-1:0] node1545;
	wire [1-1:0] node1548;
	wire [1-1:0] node1549;
	wire [1-1:0] node1553;
	wire [1-1:0] node1555;
	wire [1-1:0] node1556;
	wire [1-1:0] node1557;
	wire [1-1:0] node1559;
	wire [1-1:0] node1562;
	wire [1-1:0] node1563;
	wire [1-1:0] node1565;
	wire [1-1:0] node1568;
	wire [1-1:0] node1570;
	wire [1-1:0] node1574;
	wire [1-1:0] node1575;
	wire [1-1:0] node1576;
	wire [1-1:0] node1577;
	wire [1-1:0] node1579;
	wire [1-1:0] node1580;
	wire [1-1:0] node1581;
	wire [1-1:0] node1582;
	wire [1-1:0] node1586;
	wire [1-1:0] node1587;
	wire [1-1:0] node1591;
	wire [1-1:0] node1592;
	wire [1-1:0] node1597;
	wire [1-1:0] node1598;
	wire [1-1:0] node1599;
	wire [1-1:0] node1600;
	wire [1-1:0] node1601;
	wire [1-1:0] node1602;
	wire [1-1:0] node1606;
	wire [1-1:0] node1607;
	wire [1-1:0] node1611;
	wire [1-1:0] node1613;
	wire [1-1:0] node1617;
	wire [1-1:0] node1618;
	wire [1-1:0] node1619;
	wire [1-1:0] node1621;
	wire [1-1:0] node1624;
	wire [1-1:0] node1625;
	wire [1-1:0] node1629;
	wire [1-1:0] node1631;
	wire [1-1:0] node1634;
	wire [1-1:0] node1635;
	wire [1-1:0] node1637;
	wire [1-1:0] node1638;
	wire [1-1:0] node1639;
	wire [1-1:0] node1641;
	wire [1-1:0] node1644;
	wire [1-1:0] node1645;
	wire [1-1:0] node1649;
	wire [1-1:0] node1650;
	wire [1-1:0] node1655;
	wire [1-1:0] node1656;
	wire [1-1:0] node1657;
	wire [1-1:0] node1658;
	wire [1-1:0] node1659;
	wire [1-1:0] node1660;
	wire [1-1:0] node1661;
	wire [1-1:0] node1663;
	wire [1-1:0] node1664;
	wire [1-1:0] node1665;
	wire [1-1:0] node1666;
	wire [1-1:0] node1670;
	wire [1-1:0] node1671;
	wire [1-1:0] node1673;
	wire [1-1:0] node1676;
	wire [1-1:0] node1680;
	wire [1-1:0] node1681;
	wire [1-1:0] node1682;
	wire [1-1:0] node1683;
	wire [1-1:0] node1685;
	wire [1-1:0] node1688;
	wire [1-1:0] node1690;
	wire [1-1:0] node1691;
	wire [1-1:0] node1696;
	wire [1-1:0] node1697;
	wire [1-1:0] node1698;
	wire [1-1:0] node1702;
	wire [1-1:0] node1703;
	wire [1-1:0] node1705;
	wire [1-1:0] node1708;
	wire [1-1:0] node1710;
	wire [1-1:0] node1713;
	wire [1-1:0] node1714;
	wire [1-1:0] node1716;
	wire [1-1:0] node1717;
	wire [1-1:0] node1718;
	wire [1-1:0] node1719;
	wire [1-1:0] node1723;
	wire [1-1:0] node1724;
	wire [1-1:0] node1728;
	wire [1-1:0] node1730;
	wire [1-1:0] node1734;
	wire [1-1:0] node1735;
	wire [1-1:0] node1736;
	wire [1-1:0] node1738;
	wire [1-1:0] node1739;
	wire [1-1:0] node1740;
	wire [1-1:0] node1742;
	wire [1-1:0] node1745;
	wire [1-1:0] node1746;
	wire [1-1:0] node1748;
	wire [1-1:0] node1751;
	wire [1-1:0] node1753;
	wire [1-1:0] node1757;
	wire [1-1:0] node1758;
	wire [1-1:0] node1759;
	wire [1-1:0] node1760;
	wire [1-1:0] node1761;
	wire [1-1:0] node1762;
	wire [1-1:0] node1766;
	wire [1-1:0] node1768;
	wire [1-1:0] node1771;
	wire [1-1:0] node1773;
	wire [1-1:0] node1777;
	wire [1-1:0] node1778;
	wire [1-1:0] node1780;
	wire [1-1:0] node1783;
	wire [1-1:0] node1784;
	wire [1-1:0] node1785;
	wire [1-1:0] node1789;
	wire [1-1:0] node1791;
	wire [1-1:0] node1794;
	wire [1-1:0] node1796;
	wire [1-1:0] node1797;
	wire [1-1:0] node1798;
	wire [1-1:0] node1799;
	wire [1-1:0] node1800;
	wire [1-1:0] node1804;
	wire [1-1:0] node1805;
	wire [1-1:0] node1809;
	wire [1-1:0] node1811;
	wire [1-1:0] node1815;
	wire [1-1:0] node1816;
	wire [1-1:0] node1817;
	wire [1-1:0] node1819;
	wire [1-1:0] node1820;
	wire [1-1:0] node1821;
	wire [1-1:0] node1822;
	wire [1-1:0] node1823;
	wire [1-1:0] node1827;
	wire [1-1:0] node1829;
	wire [1-1:0] node1832;
	wire [1-1:0] node1833;
	wire [1-1:0] node1838;
	wire [1-1:0] node1839;
	wire [1-1:0] node1840;
	wire [1-1:0] node1842;
	wire [1-1:0] node1845;
	wire [1-1:0] node1846;
	wire [1-1:0] node1848;
	wire [1-1:0] node1851;
	wire [1-1:0] node1852;
	wire [1-1:0] node1856;
	wire [1-1:0] node1858;
	wire [1-1:0] node1859;
	wire [1-1:0] node1860;
	wire [1-1:0] node1862;
	wire [1-1:0] node1865;
	wire [1-1:0] node1866;
	wire [1-1:0] node1870;
	wire [1-1:0] node1871;
	wire [1-1:0] node1875;
	wire [1-1:0] node1876;
	wire [1-1:0] node1878;
	wire [1-1:0] node1879;
	wire [1-1:0] node1881;
	wire [1-1:0] node1884;
	wire [1-1:0] node1885;
	wire [1-1:0] node1886;
	wire [1-1:0] node1890;
	wire [1-1:0] node1892;
	wire [1-1:0] node1896;
	wire [1-1:0] node1897;
	wire [1-1:0] node1898;
	wire [1-1:0] node1899;
	wire [1-1:0] node1901;
	wire [1-1:0] node1902;
	wire [1-1:0] node1903;
	wire [1-1:0] node1904;
	wire [1-1:0] node1906;
	wire [1-1:0] node1909;
	wire [1-1:0] node1911;
	wire [1-1:0] node1914;
	wire [1-1:0] node1916;
	wire [1-1:0] node1920;
	wire [1-1:0] node1921;
	wire [1-1:0] node1922;
	wire [1-1:0] node1923;
	wire [1-1:0] node1925;
	wire [1-1:0] node1928;
	wire [1-1:0] node1929;
	wire [1-1:0] node1931;
	wire [1-1:0] node1934;
	wire [1-1:0] node1935;
	wire [1-1:0] node1939;
	wire [1-1:0] node1941;
	wire [1-1:0] node1942;
	wire [1-1:0] node1943;
	wire [1-1:0] node1945;
	wire [1-1:0] node1948;
	wire [1-1:0] node1949;
	wire [1-1:0] node1953;
	wire [1-1:0] node1954;
	wire [1-1:0] node1955;
	wire [1-1:0] node1960;
	wire [1-1:0] node1962;
	wire [1-1:0] node1963;
	wire [1-1:0] node1964;
	wire [1-1:0] node1966;
	wire [1-1:0] node1969;
	wire [1-1:0] node1970;
	wire [1-1:0] node1972;
	wire [1-1:0] node1975;
	wire [1-1:0] node1977;
	wire [1-1:0] node1981;
	wire [1-1:0] node1982;
	wire [1-1:0] node1983;
	wire [1-1:0] node1985;
	wire [1-1:0] node1986;
	wire [1-1:0] node1987;
	wire [1-1:0] node1989;
	wire [1-1:0] node1992;
	wire [1-1:0] node1993;
	wire [1-1:0] node1997;
	wire [1-1:0] node1998;
	wire [1-1:0] node2003;
	wire [1-1:0] node2004;
	wire [1-1:0] node2005;
	wire [1-1:0] node2006;
	wire [1-1:0] node2008;
	wire [1-1:0] node2011;
	wire [1-1:0] node2012;
	wire [1-1:0] node2013;
	wire [1-1:0] node2017;
	wire [1-1:0] node2018;
	wire [1-1:0] node2022;
	wire [1-1:0] node2024;
	wire [1-1:0] node2025;
	wire [1-1:0] node2026;
	wire [1-1:0] node2030;
	wire [1-1:0] node2031;
	wire [1-1:0] node2033;
	wire [1-1:0] node2036;
	wire [1-1:0] node2038;
	wire [1-1:0] node2041;
	wire [1-1:0] node2042;
	wire [1-1:0] node2044;
	wire [1-1:0] node2045;
	wire [1-1:0] node2046;
	wire [1-1:0] node2047;
	wire [1-1:0] node2051;
	wire [1-1:0] node2052;
	wire [1-1:0] node2056;
	wire [1-1:0] node2058;
	wire [1-1:0] node2062;
	wire [1-1:0] node2063;
	wire [1-1:0] node2064;
	wire [1-1:0] node2066;
	wire [1-1:0] node2067;
	wire [1-1:0] node2069;
	wire [1-1:0] node2072;
	wire [1-1:0] node2073;
	wire [1-1:0] node2075;
	wire [1-1:0] node2078;
	wire [1-1:0] node2079;
	wire [1-1:0] node2084;
	wire [1-1:0] node2085;
	wire [1-1:0] node2086;
	wire [1-1:0] node2087;
	wire [1-1:0] node2088;
	wire [1-1:0] node2089;
	wire [1-1:0] node2093;
	wire [1-1:0] node2094;
	wire [1-1:0] node2096;
	wire [1-1:0] node2099;
	wire [1-1:0] node2100;
	wire [1-1:0] node2105;
	wire [1-1:0] node2106;
	wire [1-1:0] node2107;
	wire [1-1:0] node2108;
	wire [1-1:0] node2112;
	wire [1-1:0] node2114;
	wire [1-1:0] node2117;
	wire [1-1:0] node2118;
	wire [1-1:0] node2122;
	wire [1-1:0] node2123;
	wire [1-1:0] node2125;
	wire [1-1:0] node2126;
	wire [1-1:0] node2127;
	wire [1-1:0] node2128;
	wire [1-1:0] node2132;
	wire [1-1:0] node2133;
	wire [1-1:0] node2137;
	wire [1-1:0] node2139;
	wire [1-1:0] node2143;
	wire [1-1:0] node2144;
	wire [1-1:0] node2145;
	wire [1-1:0] node2146;
	wire [1-1:0] node2148;
	wire [1-1:0] node2149;
	wire [1-1:0] node2150;
	wire [1-1:0] node2154;
	wire [1-1:0] node2155;
	wire [1-1:0] node2157;
	wire [1-1:0] node2160;
	wire [1-1:0] node2162;
	wire [1-1:0] node2166;
	wire [1-1:0] node2167;
	wire [1-1:0] node2168;
	wire [1-1:0] node2169;
	wire [1-1:0] node2170;
	wire [1-1:0] node2172;
	wire [1-1:0] node2175;
	wire [1-1:0] node2176;
	wire [1-1:0] node2180;
	wire [1-1:0] node2182;
	wire [1-1:0] node2185;
	wire [1-1:0] node2187;
	wire [1-1:0] node2188;
	wire [1-1:0] node2189;
	wire [1-1:0] node2193;
	wire [1-1:0] node2194;
	wire [1-1:0] node2196;
	wire [1-1:0] node2199;
	wire [1-1:0] node2201;
	wire [1-1:0] node2204;
	wire [1-1:0] node2205;
	wire [1-1:0] node2207;
	wire [1-1:0] node2208;
	wire [1-1:0] node2209;
	wire [1-1:0] node2210;
	wire [1-1:0] node2214;
	wire [1-1:0] node2216;
	wire [1-1:0] node2219;
	wire [1-1:0] node2221;
	wire [1-1:0] node2225;
	wire [1-1:0] node2226;
	wire [1-1:0] node2227;
	wire [1-1:0] node2228;
	wire [1-1:0] node2230;
	wire [1-1:0] node2231;
	wire [1-1:0] node2232;
	wire [1-1:0] node2233;
	wire [1-1:0] node2237;
	wire [1-1:0] node2238;
	wire [1-1:0] node2240;
	wire [1-1:0] node2243;
	wire [1-1:0] node2245;
	wire [1-1:0] node2249;
	wire [1-1:0] node2250;
	wire [1-1:0] node2251;
	wire [1-1:0] node2252;
	wire [1-1:0] node2254;
	wire [1-1:0] node2257;
	wire [1-1:0] node2258;
	wire [1-1:0] node2262;
	wire [1-1:0] node2263;
	wire [1-1:0] node2267;
	wire [1-1:0] node2269;
	wire [1-1:0] node2270;
	wire [1-1:0] node2271;
	wire [1-1:0] node2272;
	wire [1-1:0] node2276;
	wire [1-1:0] node2278;
	wire [1-1:0] node2281;
	wire [1-1:0] node2283;
	wire [1-1:0] node2286;
	wire [1-1:0] node2287;
	wire [1-1:0] node2289;
	wire [1-1:0] node2290;
	wire [1-1:0] node2292;
	wire [1-1:0] node2295;
	wire [1-1:0] node2296;
	wire [1-1:0] node2297;
	wire [1-1:0] node2301;
	wire [1-1:0] node2302;
	wire [1-1:0] node2307;
	wire [1-1:0] node2308;
	wire [1-1:0] node2309;
	wire [1-1:0] node2310;
	wire [1-1:0] node2312;
	wire [1-1:0] node2313;
	wire [1-1:0] node2315;
	wire [1-1:0] node2318;
	wire [1-1:0] node2319;
	wire [1-1:0] node2321;
	wire [1-1:0] node2324;
	wire [1-1:0] node2325;
	wire [1-1:0] node2330;
	wire [1-1:0] node2331;
	wire [1-1:0] node2332;
	wire [1-1:0] node2333;
	wire [1-1:0] node2337;
	wire [1-1:0] node2338;
	wire [1-1:0] node2339;
	wire [1-1:0] node2343;
	wire [1-1:0] node2345;
	wire [1-1:0] node2348;
	wire [1-1:0] node2350;
	wire [1-1:0] node2351;
	wire [1-1:0] node2352;
	wire [1-1:0] node2353;
	wire [1-1:0] node2357;
	wire [1-1:0] node2359;
	wire [1-1:0] node2362;
	wire [1-1:0] node2364;
	wire [1-1:0] node2367;
	wire [1-1:0] node2368;
	wire [1-1:0] node2370;
	wire [1-1:0] node2371;
	wire [1-1:0] node2372;
	wire [1-1:0] node2374;
	wire [1-1:0] node2377;
	wire [1-1:0] node2379;
	wire [1-1:0] node2382;
	wire [1-1:0] node2384;
	wire [1-1:0] node2388;
	wire [1-1:0] node2389;
	wire [1-1:0] node2390;
	wire [1-1:0] node2391;
	wire [1-1:0] node2393;
	wire [1-1:0] node2394;
	wire [1-1:0] node2395;
	wire [1-1:0] node2396;
	wire [1-1:0] node2397;
	wire [1-1:0] node2401;
	wire [1-1:0] node2402;
	wire [1-1:0] node2406;
	wire [1-1:0] node2408;
	wire [1-1:0] node2412;
	wire [1-1:0] node2413;
	wire [1-1:0] node2414;
	wire [1-1:0] node2415;
	wire [1-1:0] node2417;
	wire [1-1:0] node2420;
	wire [1-1:0] node2422;
	wire [1-1:0] node2425;
	wire [1-1:0] node2427;
	wire [1-1:0] node2430;
	wire [1-1:0] node2432;
	wire [1-1:0] node2433;
	wire [1-1:0] node2434;
	wire [1-1:0] node2435;
	wire [1-1:0] node2439;
	wire [1-1:0] node2440;
	wire [1-1:0] node2444;
	wire [1-1:0] node2445;
	wire [1-1:0] node2449;
	wire [1-1:0] node2451;
	wire [1-1:0] node2452;
	wire [1-1:0] node2453;
	wire [1-1:0] node2454;
	wire [1-1:0] node2458;
	wire [1-1:0] node2459;
	wire [1-1:0] node2460;
	wire [1-1:0] node2464;
	wire [1-1:0] node2465;
	wire [1-1:0] node2470;
	wire [1-1:0] node2471;
	wire [1-1:0] node2472;
	wire [1-1:0] node2473;
	wire [1-1:0] node2474;
	wire [1-1:0] node2475;
	wire [1-1:0] node2476;
	wire [1-1:0] node2478;
	wire [1-1:0] node2479;
	wire [1-1:0] node2480;
	wire [1-1:0] node2481;
	wire [1-1:0] node2485;
	wire [1-1:0] node2487;
	wire [1-1:0] node2490;
	wire [1-1:0] node2492;
	wire [1-1:0] node2496;
	wire [1-1:0] node2497;
	wire [1-1:0] node2498;
	wire [1-1:0] node2499;
	wire [1-1:0] node2500;
	wire [1-1:0] node2502;
	wire [1-1:0] node2505;
	wire [1-1:0] node2507;
	wire [1-1:0] node2510;
	wire [1-1:0] node2511;
	wire [1-1:0] node2516;
	wire [1-1:0] node2517;
	wire [1-1:0] node2518;
	wire [1-1:0] node2520;
	wire [1-1:0] node2523;
	wire [1-1:0] node2525;
	wire [1-1:0] node2528;
	wire [1-1:0] node2530;
	wire [1-1:0] node2533;
	wire [1-1:0] node2534;
	wire [1-1:0] node2536;
	wire [1-1:0] node2537;
	wire [1-1:0] node2538;
	wire [1-1:0] node2542;
	wire [1-1:0] node2543;
	wire [1-1:0] node2545;
	wire [1-1:0] node2548;
	wire [1-1:0] node2550;
	wire [1-1:0] node2554;
	wire [1-1:0] node2555;
	wire [1-1:0] node2556;
	wire [1-1:0] node2558;
	wire [1-1:0] node2559;
	wire [1-1:0] node2560;
	wire [1-1:0] node2561;
	wire [1-1:0] node2563;
	wire [1-1:0] node2566;
	wire [1-1:0] node2567;
	wire [1-1:0] node2571;
	wire [1-1:0] node2572;
	wire [1-1:0] node2577;
	wire [1-1:0] node2578;
	wire [1-1:0] node2579;
	wire [1-1:0] node2580;
	wire [1-1:0] node2581;
	wire [1-1:0] node2585;
	wire [1-1:0] node2586;
	wire [1-1:0] node2588;
	wire [1-1:0] node2591;
	wire [1-1:0] node2592;
	wire [1-1:0] node2596;
	wire [1-1:0] node2598;
	wire [1-1:0] node2599;
	wire [1-1:0] node2600;
	wire [1-1:0] node2601;
	wire [1-1:0] node2605;
	wire [1-1:0] node2607;
	wire [1-1:0] node2610;
	wire [1-1:0] node2611;
	wire [1-1:0] node2615;
	wire [1-1:0] node2616;
	wire [1-1:0] node2618;
	wire [1-1:0] node2619;
	wire [1-1:0] node2620;
	wire [1-1:0] node2624;
	wire [1-1:0] node2625;
	wire [1-1:0] node2626;
	wire [1-1:0] node2630;
	wire [1-1:0] node2631;
	wire [1-1:0] node2636;
	wire [1-1:0] node2637;
	wire [1-1:0] node2638;
	wire [1-1:0] node2640;
	wire [1-1:0] node2641;
	wire [1-1:0] node2642;
	wire [1-1:0] node2643;
	wire [1-1:0] node2647;
	wire [1-1:0] node2648;
	wire [1-1:0] node2649;
	wire [1-1:0] node2653;
	wire [1-1:0] node2654;
	wire [1-1:0] node2659;
	wire [1-1:0] node2660;
	wire [1-1:0] node2661;
	wire [1-1:0] node2662;
	wire [1-1:0] node2664;
	wire [1-1:0] node2667;
	wire [1-1:0] node2668;
	wire [1-1:0] node2672;
	wire [1-1:0] node2673;
	wire [1-1:0] node2677;
	wire [1-1:0] node2679;
	wire [1-1:0] node2680;
	wire [1-1:0] node2681;
	wire [1-1:0] node2683;
	wire [1-1:0] node2686;
	wire [1-1:0] node2687;
	wire [1-1:0] node2691;
	wire [1-1:0] node2693;
	wire [1-1:0] node2696;
	wire [1-1:0] node2698;
	wire [1-1:0] node2699;
	wire [1-1:0] node2700;
	wire [1-1:0] node2701;
	wire [1-1:0] node2702;
	wire [1-1:0] node2706;
	wire [1-1:0] node2707;
	wire [1-1:0] node2711;
	wire [1-1:0] node2712;
	wire [1-1:0] node2717;
	wire [1-1:0] node2718;
	wire [1-1:0] node2719;
	wire [1-1:0] node2720;
	wire [1-1:0] node2721;
	wire [1-1:0] node2723;
	wire [1-1:0] node2724;
	wire [1-1:0] node2726;
	wire [1-1:0] node2729;
	wire [1-1:0] node2730;
	wire [1-1:0] node2732;
	wire [1-1:0] node2735;
	wire [1-1:0] node2736;
	wire [1-1:0] node2741;
	wire [1-1:0] node2742;
	wire [1-1:0] node2743;
	wire [1-1:0] node2744;
	wire [1-1:0] node2745;
	wire [1-1:0] node2746;
	wire [1-1:0] node2748;
	wire [1-1:0] node2751;
	wire [1-1:0] node2753;
	wire [1-1:0] node2756;
	wire [1-1:0] node2758;
	wire [1-1:0] node2762;
	wire [1-1:0] node2763;
	wire [1-1:0] node2764;
	wire [1-1:0] node2765;
	wire [1-1:0] node2769;
	wire [1-1:0] node2770;
	wire [1-1:0] node2774;
	wire [1-1:0] node2775;
	wire [1-1:0] node2779;
	wire [1-1:0] node2780;
	wire [1-1:0] node2782;
	wire [1-1:0] node2783;
	wire [1-1:0] node2784;
	wire [1-1:0] node2785;
	wire [1-1:0] node2789;
	wire [1-1:0] node2791;
	wire [1-1:0] node2794;
	wire [1-1:0] node2796;
	wire [1-1:0] node2800;
	wire [1-1:0] node2801;
	wire [1-1:0] node2802;
	wire [1-1:0] node2803;
	wire [1-1:0] node2805;
	wire [1-1:0] node2806;
	wire [1-1:0] node2807;
	wire [1-1:0] node2811;
	wire [1-1:0] node2812;
	wire [1-1:0] node2813;
	wire [1-1:0] node2817;
	wire [1-1:0] node2819;
	wire [1-1:0] node2823;
	wire [1-1:0] node2824;
	wire [1-1:0] node2825;
	wire [1-1:0] node2826;
	wire [1-1:0] node2827;
	wire [1-1:0] node2828;
	wire [1-1:0] node2830;
	wire [1-1:0] node2833;
	wire [1-1:0] node2835;
	wire [1-1:0] node2838;
	wire [1-1:0] node2840;
	wire [1-1:0] node2844;
	wire [1-1:0] node2845;
	wire [1-1:0] node2846;
	wire [1-1:0] node2847;
	wire [1-1:0] node2851;
	wire [1-1:0] node2852;
	wire [1-1:0] node2856;
	wire [1-1:0] node2858;
	wire [1-1:0] node2861;
	wire [1-1:0] node2862;
	wire [1-1:0] node2864;
	wire [1-1:0] node2865;
	wire [1-1:0] node2866;
	wire [1-1:0] node2867;
	wire [1-1:0] node2871;
	wire [1-1:0] node2873;
	wire [1-1:0] node2876;
	wire [1-1:0] node2878;
	wire [1-1:0] node2882;
	wire [1-1:0] node2883;
	wire [1-1:0] node2884;
	wire [1-1:0] node2885;
	wire [1-1:0] node2887;
	wire [1-1:0] node2888;
	wire [1-1:0] node2889;
	wire [1-1:0] node2890;
	wire [1-1:0] node2894;
	wire [1-1:0] node2896;
	wire [1-1:0] node2899;
	wire [1-1:0] node2900;
	wire [1-1:0] node2905;
	wire [1-1:0] node2906;
	wire [1-1:0] node2907;
	wire [1-1:0] node2909;
	wire [1-1:0] node2912;
	wire [1-1:0] node2913;
	wire [1-1:0] node2914;
	wire [1-1:0] node2918;
	wire [1-1:0] node2920;
	wire [1-1:0] node2923;
	wire [1-1:0] node2925;
	wire [1-1:0] node2926;
	wire [1-1:0] node2927;
	wire [1-1:0] node2929;
	wire [1-1:0] node2932;
	wire [1-1:0] node2934;
	wire [1-1:0] node2937;
	wire [1-1:0] node2939;
	wire [1-1:0] node2942;
	wire [1-1:0] node2943;
	wire [1-1:0] node2945;
	wire [1-1:0] node2946;
	wire [1-1:0] node2948;
	wire [1-1:0] node2951;
	wire [1-1:0] node2952;
	wire [1-1:0] node2954;
	wire [1-1:0] node2957;
	wire [1-1:0] node2958;
	wire [1-1:0] node2963;
	wire [1-1:0] node2964;
	wire [1-1:0] node2965;
	wire [1-1:0] node2966;
	wire [1-1:0] node2967;
	wire [1-1:0] node2968;
	wire [1-1:0] node2970;
	wire [1-1:0] node2972;
	wire [1-1:0] node2973;
	wire [1-1:0] node2976;
	wire [1-1:0] node2978;
	wire [1-1:0] node2982;
	wire [1-1:0] node2983;
	wire [1-1:0] node2984;
	wire [1-1:0] node2985;
	wire [1-1:0] node2986;
	wire [1-1:0] node2990;
	wire [1-1:0] node2991;
	wire [1-1:0] node2995;
	wire [1-1:0] node2996;
	wire [1-1:0] node3000;
	wire [1-1:0] node3002;
	wire [1-1:0] node3003;
	wire [1-1:0] node3004;
	wire [1-1:0] node3008;
	wire [1-1:0] node3009;
	wire [1-1:0] node3010;
	wire [1-1:0] node3014;
	wire [1-1:0] node3015;
	wire [1-1:0] node3019;
	wire [1-1:0] node3021;
	wire [1-1:0] node3022;
	wire [1-1:0] node3023;
	wire [1-1:0] node3024;
	wire [1-1:0] node3026;
	wire [1-1:0] node3029;
	wire [1-1:0] node3031;
	wire [1-1:0] node3034;
	wire [1-1:0] node3035;
	wire [1-1:0] node3040;
	wire [1-1:0] node3041;
	wire [1-1:0] node3043;
	wire [1-1:0] node3044;
	wire [1-1:0] node3045;
	wire [1-1:0] node3046;
	wire [1-1:0] node3048;
	wire [1-1:0] node3051;
	wire [1-1:0] node3052;
	wire [1-1:0] node3056;
	wire [1-1:0] node3058;
	wire [1-1:0] node3062;
	wire [1-1:0] node3063;
	wire [1-1:0] node3064;
	wire [1-1:0] node3065;
	wire [1-1:0] node3066;
	wire [1-1:0] node3070;
	wire [1-1:0] node3071;
	wire [1-1:0] node3073;
	wire [1-1:0] node3076;
	wire [1-1:0] node3077;
	wire [1-1:0] node3081;
	wire [1-1:0] node3083;
	wire [1-1:0] node3084;
	wire [1-1:0] node3086;
	wire [1-1:0] node3089;
	wire [1-1:0] node3090;
	wire [1-1:0] node3093;
	wire [1-1:0] node3096;
	wire [1-1:0] node3098;
	wire [1-1:0] node3099;
	wire [1-1:0] node3100;
	wire [1-1:0] node3102;
	wire [1-1:0] node3105;
	wire [1-1:0] node3106;
	wire [1-1:0] node3107;
	wire [1-1:0] node3111;
	wire [1-1:0] node3112;
	wire [1-1:0] node3117;
	wire [1-1:0] node3118;
	wire [1-1:0] node3119;
	wire [1-1:0] node3121;
	wire [1-1:0] node3122;
	wire [1-1:0] node3123;
	wire [1-1:0] node3124;
	wire [1-1:0] node3126;
	wire [1-1:0] node3129;
	wire [1-1:0] node3131;
	wire [1-1:0] node3134;
	wire [1-1:0] node3135;
	wire [1-1:0] node3140;
	wire [1-1:0] node3141;
	wire [1-1:0] node3142;
	wire [1-1:0] node3144;
	wire [1-1:0] node3147;
	wire [1-1:0] node3148;
	wire [1-1:0] node3150;
	wire [1-1:0] node3153;
	wire [1-1:0] node3155;
	wire [1-1:0] node3158;
	wire [1-1:0] node3160;
	wire [1-1:0] node3161;
	wire [1-1:0] node3162;
	wire [1-1:0] node3163;
	wire [1-1:0] node3167;
	wire [1-1:0] node3168;
	wire [1-1:0] node3172;
	wire [1-1:0] node3174;
	wire [1-1:0] node3177;
	wire [1-1:0] node3179;
	wire [1-1:0] node3180;
	wire [1-1:0] node3181;
	wire [1-1:0] node3182;
	wire [1-1:0] node3184;
	wire [1-1:0] node3187;
	wire [1-1:0] node3188;
	wire [1-1:0] node3192;
	wire [1-1:0] node3194;
	wire [1-1:0] node3198;
	wire [1-1:0] node3199;
	wire [1-1:0] node3200;
	wire [1-1:0] node3202;
	wire [1-1:0] node3203;
	wire [1-1:0] node3204;
	wire [1-1:0] node3205;
	wire [1-1:0] node3209;
	wire [1-1:0] node3210;
	wire [1-1:0] node3214;
	wire [1-1:0] node3216;
	wire [1-1:0] node3220;
	wire [1-1:0] node3221;
	wire [1-1:0] node3222;
	wire [1-1:0] node3223;
	wire [1-1:0] node3224;
	wire [1-1:0] node3225;
	wire [1-1:0] node3229;
	wire [1-1:0] node3230;
	wire [1-1:0] node3232;
	wire [1-1:0] node3235;
	wire [1-1:0] node3236;
	wire [1-1:0] node3241;
	wire [1-1:0] node3242;
	wire [1-1:0] node3243;
	wire [1-1:0] node3245;
	wire [1-1:0] node3248;
	wire [1-1:0] node3250;
	wire [1-1:0] node3253;
	wire [1-1:0] node3255;
	wire [1-1:0] node3258;
	wire [1-1:0] node3259;
	wire [1-1:0] node3261;
	wire [1-1:0] node3262;
	wire [1-1:0] node3264;
	wire [1-1:0] node3267;
	wire [1-1:0] node3268;
	wire [1-1:0] node3270;
	wire [1-1:0] node3273;
	wire [1-1:0] node3275;

	assign outp = (inp[4]) ? node2388 : node1;
		assign node1 = (inp[0]) ? node871 : node2;
			assign node2 = (inp[1]) ? node84 : node3;
				assign node3 = (inp[12]) ? node25 : node4;
					assign node4 = (inp[6]) ? node6 : 1'b1;
						assign node6 = (inp[5]) ? 1'b1 : node7;
							assign node7 = (inp[7]) ? node19 : node8;
								assign node8 = (inp[3]) ? node14 : node9;
									assign node9 = (inp[9]) ? node11 : 1'b0;
										assign node11 = (inp[10]) ? 1'b0 : 1'b1;
									assign node14 = (inp[10]) ? 1'b1 : node15;
										assign node15 = (inp[9]) ? 1'b0 : 1'b1;
								assign node19 = (inp[9]) ? node21 : 1'b0;
									assign node21 = (inp[10]) ? 1'b0 : 1'b1;
					assign node25 = (inp[15]) ? node63 : node26;
						assign node26 = (inp[6]) ? node44 : node27;
							assign node27 = (inp[9]) ? node33 : node28;
								assign node28 = (inp[7]) ? 1'b0 : node29;
									assign node29 = (inp[3]) ? 1'b1 : 1'b0;
								assign node33 = (inp[10]) ? node39 : node34;
									assign node34 = (inp[3]) ? node36 : 1'b1;
										assign node36 = (inp[7]) ? 1'b1 : 1'b0;
									assign node39 = (inp[7]) ? 1'b0 : node40;
										assign node40 = (inp[3]) ? 1'b1 : 1'b0;
							assign node44 = (inp[5]) ? node46 : 1'b1;
								assign node46 = (inp[10]) ? node58 : node47;
									assign node47 = (inp[9]) ? node53 : node48;
										assign node48 = (inp[7]) ? 1'b0 : node49;
											assign node49 = (inp[3]) ? 1'b1 : 1'b0;
										assign node53 = (inp[7]) ? 1'b1 : node54;
											assign node54 = (inp[3]) ? 1'b0 : 1'b1;
									assign node58 = (inp[7]) ? 1'b0 : node59;
										assign node59 = (inp[3]) ? 1'b1 : 1'b0;
						assign node63 = (inp[6]) ? node65 : 1'b1;
							assign node65 = (inp[5]) ? 1'b1 : node66;
								assign node66 = (inp[10]) ? node78 : node67;
									assign node67 = (inp[9]) ? node73 : node68;
										assign node68 = (inp[3]) ? node70 : 1'b0;
											assign node70 = (inp[7]) ? 1'b0 : 1'b1;
										assign node73 = (inp[7]) ? 1'b1 : node74;
											assign node74 = (inp[3]) ? 1'b0 : 1'b1;
									assign node78 = (inp[3]) ? node80 : 1'b0;
										assign node80 = (inp[7]) ? 1'b0 : 1'b1;
				assign node84 = (inp[8]) ? node790 : node85;
					assign node85 = (inp[14]) ? node331 : node86;
						assign node86 = (inp[13]) ? node168 : node87;
							assign node87 = (inp[15]) ? node147 : node88;
								assign node88 = (inp[12]) ? node110 : node89;
									assign node89 = (inp[5]) ? 1'b0 : node90;
										assign node90 = (inp[6]) ? node92 : 1'b0;
											assign node92 = (inp[10]) ? node104 : node93;
												assign node93 = (inp[9]) ? node99 : node94;
													assign node94 = (inp[3]) ? node96 : 1'b1;
														assign node96 = (inp[7]) ? 1'b1 : 1'b0;
													assign node99 = (inp[3]) ? node101 : 1'b0;
														assign node101 = (inp[7]) ? 1'b0 : 1'b1;
												assign node104 = (inp[7]) ? 1'b1 : node105;
													assign node105 = (inp[3]) ? 1'b0 : 1'b1;
									assign node110 = (inp[5]) ? node130 : node111;
										assign node111 = (inp[6]) ? 1'b0 : node112;
											assign node112 = (inp[10]) ? node124 : node113;
												assign node113 = (inp[9]) ? node119 : node114;
													assign node114 = (inp[7]) ? 1'b1 : node115;
														assign node115 = (inp[3]) ? 1'b0 : 1'b1;
													assign node119 = (inp[7]) ? 1'b0 : node120;
														assign node120 = (inp[3]) ? 1'b1 : 1'b0;
												assign node124 = (inp[3]) ? node126 : 1'b1;
													assign node126 = (inp[7]) ? 1'b1 : 1'b0;
										assign node130 = (inp[9]) ? node136 : node131;
											assign node131 = (inp[3]) ? node133 : 1'b1;
												assign node133 = (inp[7]) ? 1'b1 : 1'b0;
											assign node136 = (inp[10]) ? node142 : node137;
												assign node137 = (inp[7]) ? 1'b0 : node138;
													assign node138 = (inp[3]) ? 1'b1 : 1'b0;
												assign node142 = (inp[7]) ? 1'b1 : node143;
													assign node143 = (inp[3]) ? 1'b0 : 1'b1;
								assign node147 = (inp[6]) ? node149 : 1'b0;
									assign node149 = (inp[5]) ? 1'b0 : node150;
										assign node150 = (inp[9]) ? node156 : node151;
											assign node151 = (inp[7]) ? 1'b1 : node152;
												assign node152 = (inp[3]) ? 1'b0 : 1'b1;
											assign node156 = (inp[10]) ? node162 : node157;
												assign node157 = (inp[3]) ? node159 : 1'b0;
													assign node159 = (inp[7]) ? 1'b0 : 1'b1;
												assign node162 = (inp[7]) ? 1'b1 : node163;
													assign node163 = (inp[3]) ? 1'b0 : 1'b1;
							assign node168 = (inp[11]) ? node250 : node169;
								assign node169 = (inp[5]) ? node229 : node170;
									assign node170 = (inp[6]) ? node192 : node171;
										assign node171 = (inp[12]) ? node173 : 1'b1;
											assign node173 = (inp[15]) ? 1'b1 : node174;
												assign node174 = (inp[3]) ? node180 : node175;
													assign node175 = (inp[9]) ? node177 : 1'b0;
														assign node177 = (inp[10]) ? 1'b0 : 1'b1;
													assign node180 = (inp[7]) ? node186 : node181;
														assign node181 = (inp[10]) ? 1'b1 : node182;
															assign node182 = (inp[9]) ? 1'b0 : 1'b1;
														assign node186 = (inp[9]) ? node188 : 1'b0;
															assign node188 = (inp[10]) ? 1'b0 : 1'b1;
										assign node192 = (inp[15]) ? node212 : node193;
											assign node193 = (inp[12]) ? 1'b1 : node194;
												assign node194 = (inp[3]) ? node200 : node195;
													assign node195 = (inp[10]) ? 1'b0 : node196;
														assign node196 = (inp[9]) ? 1'b1 : 1'b0;
													assign node200 = (inp[7]) ? node206 : node201;
														assign node201 = (inp[10]) ? 1'b1 : node202;
															assign node202 = (inp[9]) ? 1'b0 : 1'b1;
														assign node206 = (inp[10]) ? 1'b0 : node207;
															assign node207 = (inp[9]) ? 1'b1 : 1'b0;
											assign node212 = (inp[9]) ? node218 : node213;
												assign node213 = (inp[7]) ? 1'b0 : node214;
													assign node214 = (inp[3]) ? 1'b1 : 1'b0;
												assign node218 = (inp[10]) ? node224 : node219;
													assign node219 = (inp[7]) ? 1'b1 : node220;
														assign node220 = (inp[3]) ? 1'b0 : 1'b1;
													assign node224 = (inp[3]) ? node226 : 1'b0;
														assign node226 = (inp[7]) ? 1'b0 : 1'b1;
									assign node229 = (inp[12]) ? node231 : 1'b1;
										assign node231 = (inp[15]) ? 1'b1 : node232;
											assign node232 = (inp[7]) ? node244 : node233;
												assign node233 = (inp[3]) ? node239 : node234;
													assign node234 = (inp[10]) ? 1'b0 : node235;
														assign node235 = (inp[9]) ? 1'b1 : 1'b0;
													assign node239 = (inp[10]) ? 1'b1 : node240;
														assign node240 = (inp[9]) ? 1'b0 : 1'b1;
												assign node244 = (inp[10]) ? 1'b0 : node245;
													assign node245 = (inp[9]) ? 1'b1 : 1'b0;
								assign node250 = (inp[12]) ? node272 : node251;
									assign node251 = (inp[5]) ? 1'b0 : node252;
										assign node252 = (inp[6]) ? node254 : 1'b0;
											assign node254 = (inp[9]) ? node260 : node255;
												assign node255 = (inp[7]) ? 1'b1 : node256;
													assign node256 = (inp[3]) ? 1'b0 : 1'b1;
												assign node260 = (inp[10]) ? node266 : node261;
													assign node261 = (inp[3]) ? node263 : 1'b0;
														assign node263 = (inp[7]) ? 1'b0 : 1'b1;
													assign node266 = (inp[7]) ? 1'b1 : node267;
														assign node267 = (inp[3]) ? 1'b0 : 1'b1;
									assign node272 = (inp[15]) ? node306 : node273;
										assign node273 = (inp[6]) ? node291 : node274;
											assign node274 = (inp[10]) ? node286 : node275;
												assign node275 = (inp[9]) ? node281 : node276;
													assign node276 = (inp[3]) ? node278 : 1'b1;
														assign node278 = (inp[7]) ? 1'b1 : 1'b0;
													assign node281 = (inp[3]) ? node283 : 1'b0;
														assign node283 = (inp[7]) ? 1'b0 : 1'b1;
												assign node286 = (inp[7]) ? 1'b1 : node287;
													assign node287 = (inp[3]) ? 1'b0 : 1'b1;
											assign node291 = (inp[5]) ? node293 : 1'b0;
												assign node293 = (inp[9]) ? node295 : 1'b1;
													assign node295 = (inp[10]) ? node301 : node296;
														assign node296 = (inp[7]) ? 1'b0 : node297;
															assign node297 = (inp[3]) ? 1'b1 : 1'b0;
														assign node301 = (inp[7]) ? 1'b1 : node302;
															assign node302 = (inp[3]) ? 1'b0 : 1'b1;
										assign node306 = (inp[5]) ? 1'b0 : node307;
											assign node307 = (inp[6]) ? node309 : 1'b0;
												assign node309 = (inp[10]) ? node325 : node310;
													assign node310 = (inp[2]) ? node316 : node311;
														assign node311 = (inp[9]) ? node313 : 1'b1;
															assign node313 = (inp[7]) ? 1'b0 : 1'b1;
														assign node316 = (inp[9]) ? node320 : node317;
															assign node317 = (inp[7]) ? 1'b1 : 1'b0;
															assign node320 = (inp[3]) ? node322 : 1'b0;
																assign node322 = (inp[7]) ? 1'b0 : 1'b1;
													assign node325 = (inp[7]) ? 1'b1 : node326;
														assign node326 = (inp[3]) ? 1'b0 : 1'b1;
						assign node331 = (inp[2]) ? node555 : node332;
							assign node332 = (inp[11]) ? node474 : node333;
								assign node333 = (inp[13]) ? node403 : node334;
									assign node334 = (inp[15]) ? node382 : node335;
										assign node335 = (inp[12]) ? node347 : node336;
											assign node336 = (inp[6]) ? node338 : 1'b1;
												assign node338 = (inp[5]) ? 1'b1 : node339;
													assign node339 = (inp[7]) ? 1'b0 : node340;
														assign node340 = (inp[3]) ? 1'b1 : node341;
															assign node341 = (inp[10]) ? 1'b0 : 1'b1;
											assign node347 = (inp[6]) ? node365 : node348;
												assign node348 = (inp[10]) ? node360 : node349;
													assign node349 = (inp[9]) ? node355 : node350;
														assign node350 = (inp[7]) ? 1'b0 : node351;
															assign node351 = (inp[3]) ? 1'b1 : 1'b0;
														assign node355 = (inp[7]) ? 1'b1 : node356;
															assign node356 = (inp[3]) ? 1'b0 : 1'b1;
													assign node360 = (inp[3]) ? node362 : 1'b0;
														assign node362 = (inp[7]) ? 1'b0 : 1'b1;
												assign node365 = (inp[5]) ? node367 : 1'b1;
													assign node367 = (inp[9]) ? node373 : node368;
														assign node368 = (inp[7]) ? 1'b0 : node369;
															assign node369 = (inp[3]) ? 1'b1 : 1'b0;
														assign node373 = (inp[7]) ? 1'b1 : node374;
															assign node374 = (inp[3]) ? node378 : node375;
																assign node375 = (inp[10]) ? 1'b0 : 1'b1;
																assign node378 = (inp[10]) ? 1'b1 : 1'b0;
										assign node382 = (inp[6]) ? node384 : 1'b1;
											assign node384 = (inp[5]) ? 1'b1 : node385;
												assign node385 = (inp[9]) ? node391 : node386;
													assign node386 = (inp[7]) ? 1'b0 : node387;
														assign node387 = (inp[3]) ? 1'b1 : 1'b0;
													assign node391 = (inp[10]) ? node397 : node392;
														assign node392 = (inp[7]) ? 1'b1 : node393;
															assign node393 = (inp[3]) ? 1'b0 : 1'b1;
														assign node397 = (inp[7]) ? 1'b0 : node398;
															assign node398 = (inp[3]) ? 1'b1 : 1'b0;
									assign node403 = (inp[6]) ? node423 : node404;
										assign node404 = (inp[12]) ? node406 : 1'b0;
											assign node406 = (inp[15]) ? 1'b0 : node407;
												assign node407 = (inp[3]) ? node413 : node408;
													assign node408 = (inp[9]) ? node410 : 1'b1;
														assign node410 = (inp[10]) ? 1'b1 : 1'b0;
													assign node413 = (inp[10]) ? 1'b0 : node414;
														assign node414 = (inp[7]) ? node418 : node415;
															assign node415 = (inp[9]) ? 1'b1 : 1'b0;
															assign node418 = (inp[9]) ? 1'b0 : 1'b1;
										assign node423 = (inp[5]) ? node455 : node424;
											assign node424 = (inp[12]) ? node442 : node425;
												assign node425 = (inp[7]) ? node437 : node426;
													assign node426 = (inp[3]) ? node432 : node427;
														assign node427 = (inp[9]) ? node429 : 1'b1;
															assign node429 = (inp[10]) ? 1'b1 : 1'b0;
														assign node432 = (inp[10]) ? 1'b0 : node433;
															assign node433 = (inp[9]) ? 1'b1 : 1'b0;
													assign node437 = (inp[9]) ? node439 : 1'b1;
														assign node439 = (inp[10]) ? 1'b1 : 1'b0;
												assign node442 = (inp[15]) ? node444 : 1'b0;
													assign node444 = (inp[10]) ? node450 : node445;
														assign node445 = (inp[9]) ? node447 : 1'b1;
															assign node447 = (inp[3]) ? 1'b1 : 1'b0;
														assign node450 = (inp[7]) ? 1'b1 : node451;
															assign node451 = (inp[3]) ? 1'b0 : 1'b1;
											assign node455 = (inp[15]) ? 1'b0 : node456;
												assign node456 = (inp[12]) ? node458 : 1'b0;
													assign node458 = (inp[3]) ? node464 : node459;
														assign node459 = (inp[10]) ? 1'b1 : node460;
															assign node460 = (inp[9]) ? 1'b0 : 1'b1;
														assign node464 = (inp[7]) ? node470 : node465;
															assign node465 = (inp[9]) ? node467 : 1'b0;
																assign node467 = (inp[10]) ? 1'b0 : 1'b1;
															assign node470 = (inp[9]) ? 1'b0 : 1'b1;
								assign node474 = (inp[5]) ? node534 : node475;
									assign node475 = (inp[6]) ? node495 : node476;
										assign node476 = (inp[15]) ? 1'b1 : node477;
											assign node477 = (inp[12]) ? node479 : 1'b1;
												assign node479 = (inp[3]) ? node485 : node480;
													assign node480 = (inp[10]) ? 1'b0 : node481;
														assign node481 = (inp[9]) ? 1'b1 : 1'b0;
													assign node485 = (inp[7]) ? node491 : node486;
														assign node486 = (inp[9]) ? node488 : 1'b1;
															assign node488 = (inp[10]) ? 1'b1 : 1'b0;
														assign node491 = (inp[9]) ? 1'b1 : 1'b0;
										assign node495 = (inp[12]) ? node513 : node496;
											assign node496 = (inp[9]) ? node502 : node497;
												assign node497 = (inp[3]) ? node499 : 1'b0;
													assign node499 = (inp[7]) ? 1'b0 : 1'b1;
												assign node502 = (inp[10]) ? node508 : node503;
													assign node503 = (inp[3]) ? node505 : 1'b1;
														assign node505 = (inp[7]) ? 1'b1 : 1'b0;
													assign node508 = (inp[7]) ? 1'b0 : node509;
														assign node509 = (inp[3]) ? 1'b1 : 1'b0;
											assign node513 = (inp[15]) ? node515 : 1'b1;
												assign node515 = (inp[9]) ? node521 : node516;
													assign node516 = (inp[3]) ? node518 : 1'b0;
														assign node518 = (inp[7]) ? 1'b0 : 1'b1;
													assign node521 = (inp[10]) ? node529 : node522;
														assign node522 = (inp[13]) ? node524 : 1'b1;
															assign node524 = (inp[7]) ? 1'b1 : node525;
																assign node525 = (inp[3]) ? 1'b0 : 1'b1;
														assign node529 = (inp[3]) ? node531 : 1'b0;
															assign node531 = (inp[7]) ? 1'b0 : 1'b1;
									assign node534 = (inp[12]) ? node536 : 1'b1;
										assign node536 = (inp[15]) ? 1'b1 : node537;
											assign node537 = (inp[3]) ? node543 : node538;
												assign node538 = (inp[10]) ? 1'b0 : node539;
													assign node539 = (inp[9]) ? 1'b1 : 1'b0;
												assign node543 = (inp[7]) ? node549 : node544;
													assign node544 = (inp[9]) ? node546 : 1'b1;
														assign node546 = (inp[10]) ? 1'b1 : 1'b0;
													assign node549 = (inp[9]) ? node551 : 1'b0;
														assign node551 = (inp[10]) ? 1'b0 : 1'b1;
							assign node555 = (inp[11]) ? node705 : node556;
								assign node556 = (inp[13]) ? node628 : node557;
									assign node557 = (inp[5]) ? node607 : node558;
										assign node558 = (inp[6]) ? node576 : node559;
											assign node559 = (inp[12]) ? node561 : 1'b0;
												assign node561 = (inp[15]) ? 1'b0 : node562;
													assign node562 = (inp[9]) ? node564 : 1'b1;
														assign node564 = (inp[10]) ? node570 : node565;
															assign node565 = (inp[3]) ? node567 : 1'b0;
																assign node567 = (inp[7]) ? 1'b0 : 1'b1;
															assign node570 = (inp[7]) ? 1'b1 : node571;
																assign node571 = (inp[3]) ? 1'b0 : 1'b1;
											assign node576 = (inp[12]) ? node594 : node577;
												assign node577 = (inp[3]) ? node583 : node578;
													assign node578 = (inp[9]) ? node580 : 1'b1;
														assign node580 = (inp[10]) ? 1'b1 : 1'b0;
													assign node583 = (inp[7]) ? node589 : node584;
														assign node584 = (inp[10]) ? 1'b0 : node585;
															assign node585 = (inp[9]) ? 1'b1 : 1'b0;
														assign node589 = (inp[10]) ? 1'b1 : node590;
															assign node590 = (inp[9]) ? 1'b0 : 1'b1;
												assign node594 = (inp[15]) ? node596 : 1'b0;
													assign node596 = (inp[7]) ? 1'b1 : node597;
														assign node597 = (inp[10]) ? node603 : node598;
															assign node598 = (inp[9]) ? node600 : 1'b1;
																assign node600 = (inp[3]) ? 1'b1 : 1'b0;
															assign node603 = (inp[3]) ? 1'b0 : 1'b1;
										assign node607 = (inp[12]) ? node609 : 1'b0;
											assign node609 = (inp[15]) ? 1'b0 : node610;
												assign node610 = (inp[7]) ? node622 : node611;
													assign node611 = (inp[3]) ? node617 : node612;
														assign node612 = (inp[10]) ? 1'b1 : node613;
															assign node613 = (inp[9]) ? 1'b0 : 1'b1;
														assign node617 = (inp[10]) ? 1'b0 : node618;
															assign node618 = (inp[9]) ? 1'b1 : 1'b0;
													assign node622 = (inp[9]) ? node624 : 1'b1;
														assign node624 = (inp[10]) ? 1'b1 : 1'b0;
									assign node628 = (inp[15]) ? node686 : node629;
										assign node629 = (inp[12]) ? node649 : node630;
											assign node630 = (inp[5]) ? 1'b1 : node631;
												assign node631 = (inp[6]) ? node633 : 1'b1;
													assign node633 = (inp[10]) ? node643 : node634;
														assign node634 = (inp[9]) ? node640 : node635;
															assign node635 = (inp[3]) ? node637 : 1'b0;
																assign node637 = (inp[7]) ? 1'b0 : 1'b1;
															assign node640 = (inp[7]) ? 1'b1 : 1'b0;
														assign node643 = (inp[7]) ? 1'b0 : node644;
															assign node644 = (inp[3]) ? 1'b1 : 1'b0;
											assign node649 = (inp[6]) ? node667 : node650;
												assign node650 = (inp[3]) ? node656 : node651;
													assign node651 = (inp[9]) ? node653 : 1'b0;
														assign node653 = (inp[10]) ? 1'b0 : 1'b1;
													assign node656 = (inp[7]) ? node662 : node657;
														assign node657 = (inp[9]) ? node659 : 1'b1;
															assign node659 = (inp[10]) ? 1'b1 : 1'b0;
														assign node662 = (inp[10]) ? 1'b0 : node663;
															assign node663 = (inp[9]) ? 1'b1 : 1'b0;
												assign node667 = (inp[5]) ? node669 : 1'b1;
													assign node669 = (inp[3]) ? node675 : node670;
														assign node670 = (inp[9]) ? node672 : 1'b0;
															assign node672 = (inp[10]) ? 1'b0 : 1'b1;
														assign node675 = (inp[7]) ? node681 : node676;
															assign node676 = (inp[9]) ? node678 : 1'b1;
																assign node678 = (inp[10]) ? 1'b1 : 1'b0;
															assign node681 = (inp[10]) ? 1'b0 : node682;
																assign node682 = (inp[9]) ? 1'b1 : 1'b0;
										assign node686 = (inp[6]) ? node688 : 1'b1;
											assign node688 = (inp[5]) ? 1'b1 : node689;
												assign node689 = (inp[7]) ? node699 : node690;
													assign node690 = (inp[9]) ? node694 : node691;
														assign node691 = (inp[3]) ? 1'b1 : 1'b0;
														assign node694 = (inp[3]) ? node696 : 1'b1;
															assign node696 = (inp[10]) ? 1'b1 : 1'b0;
													assign node699 = (inp[10]) ? 1'b0 : node700;
														assign node700 = (inp[9]) ? 1'b1 : 1'b0;
								assign node705 = (inp[6]) ? node727 : node706;
									assign node706 = (inp[12]) ? node708 : 1'b0;
										assign node708 = (inp[15]) ? 1'b0 : node709;
											assign node709 = (inp[10]) ? node721 : node710;
												assign node710 = (inp[9]) ? node716 : node711;
													assign node711 = (inp[3]) ? node713 : 1'b1;
														assign node713 = (inp[7]) ? 1'b1 : 1'b0;
													assign node716 = (inp[3]) ? node718 : 1'b0;
														assign node718 = (inp[7]) ? 1'b0 : 1'b1;
												assign node721 = (inp[7]) ? 1'b1 : node722;
													assign node722 = (inp[3]) ? 1'b0 : 1'b1;
									assign node727 = (inp[5]) ? node765 : node728;
										assign node728 = (inp[15]) ? node748 : node729;
											assign node729 = (inp[12]) ? 1'b0 : node730;
												assign node730 = (inp[10]) ? node742 : node731;
													assign node731 = (inp[9]) ? node737 : node732;
														assign node732 = (inp[7]) ? 1'b1 : node733;
															assign node733 = (inp[3]) ? 1'b0 : 1'b1;
														assign node737 = (inp[3]) ? node739 : 1'b0;
															assign node739 = (inp[7]) ? 1'b0 : 1'b1;
													assign node742 = (inp[3]) ? node744 : 1'b1;
														assign node744 = (inp[7]) ? 1'b1 : 1'b0;
											assign node748 = (inp[9]) ? node754 : node749;
												assign node749 = (inp[7]) ? 1'b1 : node750;
													assign node750 = (inp[3]) ? 1'b0 : 1'b1;
												assign node754 = (inp[10]) ? node760 : node755;
													assign node755 = (inp[7]) ? 1'b0 : node756;
														assign node756 = (inp[3]) ? 1'b1 : 1'b0;
													assign node760 = (inp[7]) ? 1'b1 : node761;
														assign node761 = (inp[3]) ? 1'b0 : 1'b1;
										assign node765 = (inp[12]) ? node767 : 1'b0;
											assign node767 = (inp[15]) ? 1'b0 : node768;
												assign node768 = (inp[3]) ? node774 : node769;
													assign node769 = (inp[9]) ? node771 : 1'b1;
														assign node771 = (inp[10]) ? 1'b1 : 1'b0;
													assign node774 = (inp[10]) ? 1'b0 : node775;
														assign node775 = (inp[13]) ? node781 : node776;
															assign node776 = (inp[7]) ? 1'b1 : node777;
																assign node777 = (inp[9]) ? 1'b1 : 1'b0;
															assign node781 = (inp[7]) ? node785 : node782;
																assign node782 = (inp[9]) ? 1'b1 : 1'b0;
																assign node785 = (inp[9]) ? 1'b0 : 1'b1;
					assign node790 = (inp[5]) ? node850 : node791;
						assign node791 = (inp[6]) ? node813 : node792;
							assign node792 = (inp[12]) ? node794 : 1'b1;
								assign node794 = (inp[15]) ? 1'b1 : node795;
									assign node795 = (inp[3]) ? node801 : node796;
										assign node796 = (inp[9]) ? node798 : 1'b0;
											assign node798 = (inp[10]) ? 1'b0 : 1'b1;
										assign node801 = (inp[7]) ? node807 : node802;
											assign node802 = (inp[10]) ? 1'b1 : node803;
												assign node803 = (inp[9]) ? 1'b0 : 1'b1;
											assign node807 = (inp[9]) ? node809 : 1'b0;
												assign node809 = (inp[10]) ? 1'b0 : 1'b1;
							assign node813 = (inp[15]) ? node833 : node814;
								assign node814 = (inp[12]) ? 1'b1 : node815;
									assign node815 = (inp[10]) ? node827 : node816;
										assign node816 = (inp[9]) ? node822 : node817;
											assign node817 = (inp[3]) ? node819 : 1'b0;
												assign node819 = (inp[7]) ? 1'b0 : 1'b1;
											assign node822 = (inp[3]) ? node824 : 1'b1;
												assign node824 = (inp[7]) ? 1'b1 : 1'b0;
										assign node827 = (inp[7]) ? 1'b0 : node828;
											assign node828 = (inp[3]) ? 1'b1 : 1'b0;
								assign node833 = (inp[10]) ? node845 : node834;
									assign node834 = (inp[9]) ? node840 : node835;
										assign node835 = (inp[7]) ? 1'b0 : node836;
											assign node836 = (inp[3]) ? 1'b1 : 1'b0;
										assign node840 = (inp[7]) ? 1'b1 : node841;
											assign node841 = (inp[3]) ? 1'b0 : 1'b1;
									assign node845 = (inp[3]) ? node847 : 1'b0;
										assign node847 = (inp[7]) ? 1'b0 : 1'b1;
						assign node850 = (inp[15]) ? 1'b1 : node851;
							assign node851 = (inp[12]) ? node853 : 1'b1;
								assign node853 = (inp[3]) ? node859 : node854;
									assign node854 = (inp[10]) ? 1'b0 : node855;
										assign node855 = (inp[9]) ? 1'b1 : 1'b0;
									assign node859 = (inp[7]) ? node865 : node860;
										assign node860 = (inp[9]) ? node862 : 1'b1;
											assign node862 = (inp[10]) ? 1'b1 : 1'b0;
										assign node865 = (inp[10]) ? 1'b0 : node866;
											assign node866 = (inp[9]) ? 1'b1 : 1'b0;
			assign node871 = (inp[8]) ? node1655 : node872;
				assign node872 = (inp[1]) ? node1574 : node873;
					assign node873 = (inp[2]) ? node1333 : node874;
						assign node874 = (inp[14]) ? node1098 : node875;
							assign node875 = (inp[13]) ? node957 : node876;
								assign node876 = (inp[15]) ? node936 : node877;
									assign node877 = (inp[12]) ? node899 : node878;
										assign node878 = (inp[6]) ? node880 : 1'b0;
											assign node880 = (inp[5]) ? 1'b0 : node881;
												assign node881 = (inp[9]) ? node887 : node882;
													assign node882 = (inp[7]) ? 1'b1 : node883;
														assign node883 = (inp[3]) ? 1'b0 : 1'b1;
													assign node887 = (inp[10]) ? node893 : node888;
														assign node888 = (inp[3]) ? node890 : 1'b0;
															assign node890 = (inp[7]) ? 1'b0 : 1'b1;
														assign node893 = (inp[3]) ? node895 : 1'b1;
															assign node895 = (inp[7]) ? 1'b1 : 1'b0;
										assign node899 = (inp[5]) ? node919 : node900;
											assign node900 = (inp[6]) ? 1'b0 : node901;
												assign node901 = (inp[7]) ? node913 : node902;
													assign node902 = (inp[3]) ? node908 : node903;
														assign node903 = (inp[10]) ? 1'b1 : node904;
															assign node904 = (inp[9]) ? 1'b0 : 1'b1;
														assign node908 = (inp[10]) ? 1'b0 : node909;
															assign node909 = (inp[9]) ? 1'b1 : 1'b0;
													assign node913 = (inp[9]) ? node915 : 1'b1;
														assign node915 = (inp[10]) ? 1'b1 : 1'b0;
											assign node919 = (inp[7]) ? node931 : node920;
												assign node920 = (inp[3]) ? node926 : node921;
													assign node921 = (inp[10]) ? 1'b1 : node922;
														assign node922 = (inp[9]) ? 1'b0 : 1'b1;
													assign node926 = (inp[10]) ? 1'b0 : node927;
														assign node927 = (inp[9]) ? 1'b1 : 1'b0;
												assign node931 = (inp[10]) ? 1'b1 : node932;
													assign node932 = (inp[9]) ? 1'b0 : 1'b1;
									assign node936 = (inp[6]) ? node938 : 1'b0;
										assign node938 = (inp[5]) ? 1'b0 : node939;
											assign node939 = (inp[10]) ? node951 : node940;
												assign node940 = (inp[9]) ? node946 : node941;
													assign node941 = (inp[7]) ? 1'b1 : node942;
														assign node942 = (inp[3]) ? 1'b0 : 1'b1;
													assign node946 = (inp[7]) ? 1'b0 : node947;
														assign node947 = (inp[3]) ? 1'b1 : 1'b0;
												assign node951 = (inp[3]) ? node953 : 1'b1;
													assign node953 = (inp[7]) ? 1'b1 : 1'b0;
								assign node957 = (inp[11]) ? node1033 : node958;
									assign node958 = (inp[5]) ? node1006 : node959;
										assign node959 = (inp[6]) ? node975 : node960;
											assign node960 = (inp[12]) ? node962 : 1'b1;
												assign node962 = (inp[15]) ? 1'b1 : node963;
													assign node963 = (inp[7]) ? 1'b0 : node964;
														assign node964 = (inp[9]) ? node966 : 1'b1;
															assign node966 = (inp[10]) ? node970 : node967;
																assign node967 = (inp[3]) ? 1'b0 : 1'b1;
																assign node970 = (inp[3]) ? 1'b1 : 1'b0;
											assign node975 = (inp[15]) ? node989 : node976;
												assign node976 = (inp[12]) ? 1'b1 : node977;
													assign node977 = (inp[3]) ? node983 : node978;
														assign node978 = (inp[10]) ? 1'b0 : node979;
															assign node979 = (inp[9]) ? 1'b1 : 1'b0;
														assign node983 = (inp[7]) ? node985 : 1'b1;
															assign node985 = (inp[9]) ? 1'b1 : 1'b0;
												assign node989 = (inp[10]) ? node1001 : node990;
													assign node990 = (inp[7]) ? node998 : node991;
														assign node991 = (inp[9]) ? node995 : node992;
															assign node992 = (inp[3]) ? 1'b1 : 1'b0;
															assign node995 = (inp[3]) ? 1'b0 : 1'b1;
														assign node998 = (inp[9]) ? 1'b1 : 1'b0;
													assign node1001 = (inp[7]) ? 1'b0 : node1002;
														assign node1002 = (inp[3]) ? 1'b1 : 1'b0;
										assign node1006 = (inp[15]) ? 1'b1 : node1007;
											assign node1007 = (inp[12]) ? node1009 : 1'b1;
												assign node1009 = (inp[10]) ? node1027 : node1010;
													assign node1010 = (inp[7]) ? node1024 : node1011;
														assign node1011 = (inp[6]) ? node1019 : node1012;
															assign node1012 = (inp[9]) ? node1016 : node1013;
																assign node1013 = (inp[3]) ? 1'b1 : 1'b0;
																assign node1016 = (inp[3]) ? 1'b0 : 1'b1;
															assign node1019 = (inp[9]) ? 1'b0 : node1020;
																assign node1020 = (inp[3]) ? 1'b1 : 1'b0;
														assign node1024 = (inp[9]) ? 1'b1 : 1'b0;
													assign node1027 = (inp[3]) ? node1029 : 1'b0;
														assign node1029 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1033 = (inp[12]) ? node1053 : node1034;
										assign node1034 = (inp[6]) ? node1036 : 1'b0;
											assign node1036 = (inp[5]) ? 1'b0 : node1037;
												assign node1037 = (inp[9]) ? node1043 : node1038;
													assign node1038 = (inp[7]) ? 1'b1 : node1039;
														assign node1039 = (inp[3]) ? 1'b0 : 1'b1;
													assign node1043 = (inp[7]) ? node1049 : node1044;
														assign node1044 = (inp[10]) ? 1'b0 : node1045;
															assign node1045 = (inp[3]) ? 1'b1 : 1'b0;
														assign node1049 = (inp[10]) ? 1'b1 : 1'b0;
										assign node1053 = (inp[15]) ? node1083 : node1054;
											assign node1054 = (inp[6]) ? node1070 : node1055;
												assign node1055 = (inp[3]) ? node1061 : node1056;
													assign node1056 = (inp[9]) ? node1058 : 1'b1;
														assign node1058 = (inp[10]) ? 1'b1 : 1'b0;
													assign node1061 = (inp[7]) ? node1065 : node1062;
														assign node1062 = (inp[9]) ? 1'b1 : 1'b0;
														assign node1065 = (inp[9]) ? node1067 : 1'b1;
															assign node1067 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1070 = (inp[5]) ? node1072 : 1'b0;
													assign node1072 = (inp[9]) ? node1078 : node1073;
														assign node1073 = (inp[3]) ? node1075 : 1'b1;
															assign node1075 = (inp[7]) ? 1'b1 : 1'b0;
														assign node1078 = (inp[10]) ? node1080 : 1'b0;
															assign node1080 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1083 = (inp[5]) ? 1'b0 : node1084;
												assign node1084 = (inp[6]) ? node1086 : 1'b0;
													assign node1086 = (inp[7]) ? 1'b1 : node1087;
														assign node1087 = (inp[3]) ? node1093 : node1088;
															assign node1088 = (inp[10]) ? 1'b1 : node1089;
																assign node1089 = (inp[9]) ? 1'b0 : 1'b1;
															assign node1093 = (inp[9]) ? 1'b1 : 1'b0;
							assign node1098 = (inp[11]) ? node1252 : node1099;
								assign node1099 = (inp[13]) ? node1175 : node1100;
									assign node1100 = (inp[15]) ? node1156 : node1101;
										assign node1101 = (inp[12]) ? node1121 : node1102;
											assign node1102 = (inp[5]) ? 1'b1 : node1103;
												assign node1103 = (inp[6]) ? node1105 : 1'b1;
													assign node1105 = (inp[7]) ? node1115 : node1106;
														assign node1106 = (inp[10]) ? node1112 : node1107;
															assign node1107 = (inp[3]) ? 1'b0 : node1108;
																assign node1108 = (inp[9]) ? 1'b1 : 1'b0;
															assign node1112 = (inp[3]) ? 1'b1 : 1'b0;
														assign node1115 = (inp[9]) ? node1117 : 1'b0;
															assign node1117 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1121 = (inp[5]) ? node1139 : node1122;
												assign node1122 = (inp[6]) ? 1'b1 : node1123;
													assign node1123 = (inp[9]) ? node1129 : node1124;
														assign node1124 = (inp[3]) ? node1126 : 1'b0;
															assign node1126 = (inp[7]) ? 1'b0 : 1'b1;
														assign node1129 = (inp[3]) ? node1131 : 1'b1;
															assign node1131 = (inp[10]) ? node1135 : node1132;
																assign node1132 = (inp[7]) ? 1'b1 : 1'b0;
																assign node1135 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1139 = (inp[10]) ? node1151 : node1140;
													assign node1140 = (inp[9]) ? node1146 : node1141;
														assign node1141 = (inp[7]) ? 1'b0 : node1142;
															assign node1142 = (inp[3]) ? 1'b1 : 1'b0;
														assign node1146 = (inp[7]) ? 1'b1 : node1147;
															assign node1147 = (inp[3]) ? 1'b0 : 1'b1;
													assign node1151 = (inp[3]) ? node1153 : 1'b0;
														assign node1153 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1156 = (inp[6]) ? node1158 : 1'b1;
											assign node1158 = (inp[5]) ? 1'b1 : node1159;
												assign node1159 = (inp[10]) ? node1169 : node1160;
													assign node1160 = (inp[3]) ? node1164 : node1161;
														assign node1161 = (inp[9]) ? 1'b1 : 1'b0;
														assign node1164 = (inp[12]) ? 1'b1 : node1165;
															assign node1165 = (inp[9]) ? 1'b0 : 1'b1;
													assign node1169 = (inp[7]) ? 1'b0 : node1170;
														assign node1170 = (inp[3]) ? 1'b1 : 1'b0;
									assign node1175 = (inp[6]) ? node1197 : node1176;
										assign node1176 = (inp[12]) ? node1178 : 1'b0;
											assign node1178 = (inp[15]) ? 1'b0 : node1179;
												assign node1179 = (inp[7]) ? node1191 : node1180;
													assign node1180 = (inp[3]) ? node1186 : node1181;
														assign node1181 = (inp[10]) ? 1'b1 : node1182;
															assign node1182 = (inp[9]) ? 1'b0 : 1'b1;
														assign node1186 = (inp[10]) ? 1'b0 : node1187;
															assign node1187 = (inp[5]) ? 1'b0 : 1'b1;
													assign node1191 = (inp[10]) ? 1'b1 : node1192;
														assign node1192 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1197 = (inp[5]) ? node1233 : node1198;
											assign node1198 = (inp[12]) ? node1216 : node1199;
												assign node1199 = (inp[10]) ? node1211 : node1200;
													assign node1200 = (inp[9]) ? node1206 : node1201;
														assign node1201 = (inp[7]) ? 1'b1 : node1202;
															assign node1202 = (inp[3]) ? 1'b0 : 1'b1;
														assign node1206 = (inp[3]) ? node1208 : 1'b0;
															assign node1208 = (inp[7]) ? 1'b0 : 1'b1;
													assign node1211 = (inp[3]) ? node1213 : 1'b1;
														assign node1213 = (inp[7]) ? 1'b1 : 1'b0;
												assign node1216 = (inp[15]) ? node1218 : 1'b0;
													assign node1218 = (inp[10]) ? node1228 : node1219;
														assign node1219 = (inp[3]) ? node1221 : 1'b0;
															assign node1221 = (inp[7]) ? node1225 : node1222;
																assign node1222 = (inp[9]) ? 1'b1 : 1'b0;
																assign node1225 = (inp[9]) ? 1'b0 : 1'b1;
														assign node1228 = (inp[3]) ? node1230 : 1'b1;
															assign node1230 = (inp[7]) ? 1'b1 : 1'b0;
											assign node1233 = (inp[15]) ? 1'b0 : node1234;
												assign node1234 = (inp[12]) ? node1236 : 1'b0;
													assign node1236 = (inp[3]) ? node1242 : node1237;
														assign node1237 = (inp[10]) ? 1'b1 : node1238;
															assign node1238 = (inp[9]) ? 1'b0 : 1'b1;
														assign node1242 = (inp[7]) ? node1246 : node1243;
															assign node1243 = (inp[10]) ? 1'b0 : 1'b1;
															assign node1246 = (inp[10]) ? 1'b1 : node1247;
																assign node1247 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1252 = (inp[12]) ? node1274 : node1253;
									assign node1253 = (inp[5]) ? 1'b1 : node1254;
										assign node1254 = (inp[6]) ? node1256 : 1'b1;
											assign node1256 = (inp[7]) ? node1268 : node1257;
												assign node1257 = (inp[3]) ? node1263 : node1258;
													assign node1258 = (inp[10]) ? 1'b0 : node1259;
														assign node1259 = (inp[9]) ? 1'b1 : 1'b0;
													assign node1263 = (inp[10]) ? 1'b1 : node1264;
														assign node1264 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1268 = (inp[10]) ? 1'b0 : node1269;
													assign node1269 = (inp[9]) ? 1'b1 : 1'b0;
									assign node1274 = (inp[15]) ? node1312 : node1275;
										assign node1275 = (inp[5]) ? node1295 : node1276;
											assign node1276 = (inp[6]) ? 1'b1 : node1277;
												assign node1277 = (inp[7]) ? node1289 : node1278;
													assign node1278 = (inp[3]) ? node1284 : node1279;
														assign node1279 = (inp[10]) ? 1'b0 : node1280;
															assign node1280 = (inp[9]) ? 1'b1 : 1'b0;
														assign node1284 = (inp[9]) ? node1286 : 1'b1;
															assign node1286 = (inp[10]) ? 1'b1 : 1'b0;
													assign node1289 = (inp[10]) ? 1'b0 : node1290;
														assign node1290 = (inp[9]) ? 1'b1 : 1'b0;
											assign node1295 = (inp[10]) ? node1307 : node1296;
												assign node1296 = (inp[9]) ? node1302 : node1297;
													assign node1297 = (inp[7]) ? 1'b0 : node1298;
														assign node1298 = (inp[3]) ? 1'b1 : 1'b0;
													assign node1302 = (inp[7]) ? 1'b1 : node1303;
														assign node1303 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1307 = (inp[3]) ? node1309 : 1'b0;
													assign node1309 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1312 = (inp[5]) ? 1'b1 : node1313;
											assign node1313 = (inp[6]) ? node1315 : 1'b1;
												assign node1315 = (inp[9]) ? node1321 : node1316;
													assign node1316 = (inp[7]) ? 1'b0 : node1317;
														assign node1317 = (inp[3]) ? 1'b1 : 1'b0;
													assign node1321 = (inp[10]) ? node1327 : node1322;
														assign node1322 = (inp[3]) ? node1324 : 1'b1;
															assign node1324 = (inp[7]) ? 1'b1 : 1'b0;
														assign node1327 = (inp[3]) ? node1329 : 1'b0;
															assign node1329 = (inp[7]) ? 1'b0 : 1'b1;
						assign node1333 = (inp[13]) ? node1415 : node1334;
							assign node1334 = (inp[6]) ? node1356 : node1335;
								assign node1335 = (inp[12]) ? node1337 : 1'b0;
									assign node1337 = (inp[15]) ? 1'b0 : node1338;
										assign node1338 = (inp[10]) ? node1350 : node1339;
											assign node1339 = (inp[9]) ? node1345 : node1340;
												assign node1340 = (inp[7]) ? 1'b1 : node1341;
													assign node1341 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1345 = (inp[3]) ? node1347 : 1'b0;
													assign node1347 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1350 = (inp[7]) ? 1'b1 : node1351;
												assign node1351 = (inp[3]) ? 1'b0 : 1'b1;
								assign node1356 = (inp[5]) ? node1394 : node1357;
									assign node1357 = (inp[15]) ? node1377 : node1358;
										assign node1358 = (inp[12]) ? 1'b0 : node1359;
											assign node1359 = (inp[9]) ? node1365 : node1360;
												assign node1360 = (inp[7]) ? 1'b1 : node1361;
													assign node1361 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1365 = (inp[10]) ? node1371 : node1366;
													assign node1366 = (inp[7]) ? 1'b0 : node1367;
														assign node1367 = (inp[3]) ? 1'b1 : 1'b0;
													assign node1371 = (inp[7]) ? 1'b1 : node1372;
														assign node1372 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1377 = (inp[3]) ? node1383 : node1378;
											assign node1378 = (inp[9]) ? node1380 : 1'b1;
												assign node1380 = (inp[10]) ? 1'b1 : 1'b0;
											assign node1383 = (inp[7]) ? node1389 : node1384;
												assign node1384 = (inp[10]) ? 1'b0 : node1385;
													assign node1385 = (inp[9]) ? 1'b1 : 1'b0;
												assign node1389 = (inp[9]) ? node1391 : 1'b1;
													assign node1391 = (inp[10]) ? 1'b1 : 1'b0;
									assign node1394 = (inp[15]) ? 1'b0 : node1395;
										assign node1395 = (inp[12]) ? node1397 : 1'b0;
											assign node1397 = (inp[3]) ? node1403 : node1398;
												assign node1398 = (inp[10]) ? 1'b1 : node1399;
													assign node1399 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1403 = (inp[7]) ? node1409 : node1404;
													assign node1404 = (inp[9]) ? node1406 : 1'b0;
														assign node1406 = (inp[10]) ? 1'b0 : 1'b1;
													assign node1409 = (inp[9]) ? node1411 : 1'b1;
														assign node1411 = (inp[10]) ? 1'b1 : 1'b0;
							assign node1415 = (inp[11]) ? node1495 : node1416;
								assign node1416 = (inp[6]) ? node1438 : node1417;
									assign node1417 = (inp[15]) ? 1'b1 : node1418;
										assign node1418 = (inp[12]) ? node1420 : 1'b1;
											assign node1420 = (inp[10]) ? node1432 : node1421;
												assign node1421 = (inp[9]) ? node1427 : node1422;
													assign node1422 = (inp[7]) ? 1'b0 : node1423;
														assign node1423 = (inp[3]) ? 1'b1 : 1'b0;
													assign node1427 = (inp[7]) ? 1'b1 : node1428;
														assign node1428 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1432 = (inp[7]) ? 1'b0 : node1433;
													assign node1433 = (inp[3]) ? 1'b1 : 1'b0;
									assign node1438 = (inp[5]) ? node1476 : node1439;
										assign node1439 = (inp[15]) ? node1459 : node1440;
											assign node1440 = (inp[12]) ? 1'b1 : node1441;
												assign node1441 = (inp[10]) ? node1453 : node1442;
													assign node1442 = (inp[9]) ? node1448 : node1443;
														assign node1443 = (inp[7]) ? 1'b0 : node1444;
															assign node1444 = (inp[3]) ? 1'b1 : 1'b0;
														assign node1448 = (inp[3]) ? node1450 : 1'b1;
															assign node1450 = (inp[7]) ? 1'b1 : 1'b0;
													assign node1453 = (inp[7]) ? 1'b0 : node1454;
														assign node1454 = (inp[3]) ? 1'b1 : 1'b0;
											assign node1459 = (inp[9]) ? node1465 : node1460;
												assign node1460 = (inp[3]) ? node1462 : 1'b0;
													assign node1462 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1465 = (inp[10]) ? node1471 : node1466;
													assign node1466 = (inp[3]) ? node1468 : 1'b1;
														assign node1468 = (inp[7]) ? 1'b1 : 1'b0;
													assign node1471 = (inp[3]) ? node1473 : 1'b0;
														assign node1473 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1476 = (inp[12]) ? node1478 : 1'b1;
											assign node1478 = (inp[15]) ? 1'b1 : node1479;
												assign node1479 = (inp[10]) ? node1489 : node1480;
													assign node1480 = (inp[9]) ? node1484 : node1481;
														assign node1481 = (inp[3]) ? 1'b1 : 1'b0;
														assign node1484 = (inp[3]) ? node1486 : 1'b1;
															assign node1486 = (inp[7]) ? 1'b1 : 1'b0;
													assign node1489 = (inp[7]) ? 1'b0 : node1490;
														assign node1490 = (inp[3]) ? 1'b1 : 1'b0;
								assign node1495 = (inp[5]) ? node1553 : node1496;
									assign node1496 = (inp[6]) ? node1518 : node1497;
										assign node1497 = (inp[12]) ? node1499 : 1'b0;
											assign node1499 = (inp[15]) ? 1'b0 : node1500;
												assign node1500 = (inp[7]) ? node1512 : node1501;
													assign node1501 = (inp[3]) ? node1507 : node1502;
														assign node1502 = (inp[9]) ? node1504 : 1'b1;
															assign node1504 = (inp[10]) ? 1'b1 : 1'b0;
														assign node1507 = (inp[10]) ? 1'b0 : node1508;
															assign node1508 = (inp[9]) ? 1'b1 : 1'b0;
													assign node1512 = (inp[10]) ? 1'b1 : node1513;
														assign node1513 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1518 = (inp[12]) ? node1536 : node1519;
											assign node1519 = (inp[9]) ? node1525 : node1520;
												assign node1520 = (inp[7]) ? 1'b1 : node1521;
													assign node1521 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1525 = (inp[10]) ? node1531 : node1526;
													assign node1526 = (inp[3]) ? node1528 : 1'b0;
														assign node1528 = (inp[7]) ? 1'b0 : 1'b1;
													assign node1531 = (inp[3]) ? node1533 : 1'b1;
														assign node1533 = (inp[7]) ? 1'b1 : 1'b0;
											assign node1536 = (inp[15]) ? node1538 : 1'b0;
												assign node1538 = (inp[10]) ? node1548 : node1539;
													assign node1539 = (inp[9]) ? node1545 : node1540;
														assign node1540 = (inp[3]) ? node1542 : 1'b1;
															assign node1542 = (inp[7]) ? 1'b1 : 1'b0;
														assign node1545 = (inp[3]) ? 1'b1 : 1'b0;
													assign node1548 = (inp[7]) ? 1'b1 : node1549;
														assign node1549 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1553 = (inp[12]) ? node1555 : 1'b0;
										assign node1555 = (inp[15]) ? 1'b0 : node1556;
											assign node1556 = (inp[3]) ? node1562 : node1557;
												assign node1557 = (inp[9]) ? node1559 : 1'b1;
													assign node1559 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1562 = (inp[7]) ? node1568 : node1563;
													assign node1563 = (inp[9]) ? node1565 : 1'b0;
														assign node1565 = (inp[10]) ? 1'b0 : 1'b1;
													assign node1568 = (inp[9]) ? node1570 : 1'b1;
														assign node1570 = (inp[10]) ? 1'b1 : 1'b0;
					assign node1574 = (inp[5]) ? node1634 : node1575;
						assign node1575 = (inp[6]) ? node1597 : node1576;
							assign node1576 = (inp[15]) ? 1'b1 : node1577;
								assign node1577 = (inp[12]) ? node1579 : 1'b1;
									assign node1579 = (inp[7]) ? node1591 : node1580;
										assign node1580 = (inp[3]) ? node1586 : node1581;
											assign node1581 = (inp[10]) ? 1'b0 : node1582;
												assign node1582 = (inp[9]) ? 1'b1 : 1'b0;
											assign node1586 = (inp[10]) ? 1'b1 : node1587;
												assign node1587 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1591 = (inp[10]) ? 1'b0 : node1592;
											assign node1592 = (inp[9]) ? 1'b1 : 1'b0;
							assign node1597 = (inp[15]) ? node1617 : node1598;
								assign node1598 = (inp[12]) ? 1'b1 : node1599;
									assign node1599 = (inp[7]) ? node1611 : node1600;
										assign node1600 = (inp[3]) ? node1606 : node1601;
											assign node1601 = (inp[10]) ? 1'b0 : node1602;
												assign node1602 = (inp[9]) ? 1'b1 : 1'b0;
											assign node1606 = (inp[10]) ? 1'b1 : node1607;
												assign node1607 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1611 = (inp[9]) ? node1613 : 1'b0;
											assign node1613 = (inp[10]) ? 1'b0 : 1'b1;
								assign node1617 = (inp[10]) ? node1629 : node1618;
									assign node1618 = (inp[9]) ? node1624 : node1619;
										assign node1619 = (inp[3]) ? node1621 : 1'b0;
											assign node1621 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1624 = (inp[7]) ? 1'b1 : node1625;
											assign node1625 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1629 = (inp[3]) ? node1631 : 1'b0;
										assign node1631 = (inp[7]) ? 1'b0 : 1'b1;
						assign node1634 = (inp[15]) ? 1'b1 : node1635;
							assign node1635 = (inp[12]) ? node1637 : 1'b1;
								assign node1637 = (inp[7]) ? node1649 : node1638;
									assign node1638 = (inp[3]) ? node1644 : node1639;
										assign node1639 = (inp[9]) ? node1641 : 1'b0;
											assign node1641 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1644 = (inp[10]) ? 1'b1 : node1645;
											assign node1645 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1649 = (inp[10]) ? 1'b0 : node1650;
										assign node1650 = (inp[9]) ? 1'b1 : 1'b0;
				assign node1655 = (inp[11]) ? node2143 : node1656;
					assign node1656 = (inp[13]) ? node1896 : node1657;
						assign node1657 = (inp[2]) ? node1815 : node1658;
							assign node1658 = (inp[14]) ? node1734 : node1659;
								assign node1659 = (inp[15]) ? node1713 : node1660;
									assign node1660 = (inp[12]) ? node1680 : node1661;
										assign node1661 = (inp[6]) ? node1663 : 1'b0;
											assign node1663 = (inp[5]) ? 1'b0 : node1664;
												assign node1664 = (inp[9]) ? node1670 : node1665;
													assign node1665 = (inp[7]) ? 1'b1 : node1666;
														assign node1666 = (inp[3]) ? 1'b0 : 1'b1;
													assign node1670 = (inp[10]) ? node1676 : node1671;
														assign node1671 = (inp[3]) ? node1673 : 1'b0;
															assign node1673 = (inp[7]) ? 1'b0 : 1'b1;
														assign node1676 = (inp[7]) ? 1'b1 : 1'b0;
										assign node1680 = (inp[5]) ? node1696 : node1681;
											assign node1681 = (inp[6]) ? 1'b0 : node1682;
												assign node1682 = (inp[9]) ? node1688 : node1683;
													assign node1683 = (inp[3]) ? node1685 : 1'b1;
														assign node1685 = (inp[7]) ? 1'b1 : 1'b0;
													assign node1688 = (inp[10]) ? node1690 : 1'b0;
														assign node1690 = (inp[1]) ? 1'b1 : node1691;
															assign node1691 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1696 = (inp[3]) ? node1702 : node1697;
												assign node1697 = (inp[10]) ? 1'b1 : node1698;
													assign node1698 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1702 = (inp[7]) ? node1708 : node1703;
													assign node1703 = (inp[9]) ? node1705 : 1'b0;
														assign node1705 = (inp[10]) ? 1'b0 : 1'b1;
													assign node1708 = (inp[9]) ? node1710 : 1'b1;
														assign node1710 = (inp[10]) ? 1'b1 : 1'b0;
									assign node1713 = (inp[5]) ? 1'b0 : node1714;
										assign node1714 = (inp[6]) ? node1716 : 1'b0;
											assign node1716 = (inp[10]) ? node1728 : node1717;
												assign node1717 = (inp[9]) ? node1723 : node1718;
													assign node1718 = (inp[7]) ? 1'b1 : node1719;
														assign node1719 = (inp[3]) ? 1'b0 : 1'b1;
													assign node1723 = (inp[7]) ? 1'b0 : node1724;
														assign node1724 = (inp[3]) ? 1'b1 : 1'b0;
												assign node1728 = (inp[3]) ? node1730 : 1'b1;
													assign node1730 = (inp[7]) ? 1'b1 : 1'b0;
								assign node1734 = (inp[15]) ? node1794 : node1735;
									assign node1735 = (inp[12]) ? node1757 : node1736;
										assign node1736 = (inp[6]) ? node1738 : 1'b1;
											assign node1738 = (inp[5]) ? 1'b1 : node1739;
												assign node1739 = (inp[3]) ? node1745 : node1740;
													assign node1740 = (inp[9]) ? node1742 : 1'b0;
														assign node1742 = (inp[10]) ? 1'b0 : 1'b1;
													assign node1745 = (inp[7]) ? node1751 : node1746;
														assign node1746 = (inp[9]) ? node1748 : 1'b1;
															assign node1748 = (inp[10]) ? 1'b1 : 1'b0;
														assign node1751 = (inp[9]) ? node1753 : 1'b0;
															assign node1753 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1757 = (inp[5]) ? node1777 : node1758;
											assign node1758 = (inp[6]) ? 1'b1 : node1759;
												assign node1759 = (inp[10]) ? node1771 : node1760;
													assign node1760 = (inp[9]) ? node1766 : node1761;
														assign node1761 = (inp[7]) ? 1'b0 : node1762;
															assign node1762 = (inp[3]) ? 1'b1 : 1'b0;
														assign node1766 = (inp[3]) ? node1768 : 1'b1;
															assign node1768 = (inp[7]) ? 1'b1 : 1'b0;
													assign node1771 = (inp[3]) ? node1773 : 1'b0;
														assign node1773 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1777 = (inp[3]) ? node1783 : node1778;
												assign node1778 = (inp[9]) ? node1780 : 1'b0;
													assign node1780 = (inp[10]) ? 1'b0 : 1'b1;
												assign node1783 = (inp[7]) ? node1789 : node1784;
													assign node1784 = (inp[10]) ? 1'b1 : node1785;
														assign node1785 = (inp[9]) ? 1'b0 : 1'b1;
													assign node1789 = (inp[9]) ? node1791 : 1'b0;
														assign node1791 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1794 = (inp[6]) ? node1796 : 1'b1;
										assign node1796 = (inp[5]) ? 1'b1 : node1797;
											assign node1797 = (inp[7]) ? node1809 : node1798;
												assign node1798 = (inp[3]) ? node1804 : node1799;
													assign node1799 = (inp[10]) ? 1'b0 : node1800;
														assign node1800 = (inp[9]) ? 1'b1 : 1'b0;
													assign node1804 = (inp[10]) ? 1'b1 : node1805;
														assign node1805 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1809 = (inp[9]) ? node1811 : 1'b0;
													assign node1811 = (inp[10]) ? 1'b0 : 1'b1;
							assign node1815 = (inp[15]) ? node1875 : node1816;
								assign node1816 = (inp[12]) ? node1838 : node1817;
									assign node1817 = (inp[6]) ? node1819 : 1'b0;
										assign node1819 = (inp[5]) ? 1'b0 : node1820;
											assign node1820 = (inp[10]) ? node1832 : node1821;
												assign node1821 = (inp[9]) ? node1827 : node1822;
													assign node1822 = (inp[7]) ? 1'b1 : node1823;
														assign node1823 = (inp[3]) ? 1'b0 : 1'b1;
													assign node1827 = (inp[3]) ? node1829 : 1'b0;
														assign node1829 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1832 = (inp[7]) ? 1'b1 : node1833;
													assign node1833 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1838 = (inp[6]) ? node1856 : node1839;
										assign node1839 = (inp[3]) ? node1845 : node1840;
											assign node1840 = (inp[9]) ? node1842 : 1'b1;
												assign node1842 = (inp[10]) ? 1'b1 : 1'b0;
											assign node1845 = (inp[7]) ? node1851 : node1846;
												assign node1846 = (inp[9]) ? node1848 : 1'b0;
													assign node1848 = (inp[10]) ? 1'b0 : 1'b1;
												assign node1851 = (inp[10]) ? 1'b1 : node1852;
													assign node1852 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1856 = (inp[5]) ? node1858 : 1'b0;
											assign node1858 = (inp[7]) ? node1870 : node1859;
												assign node1859 = (inp[3]) ? node1865 : node1860;
													assign node1860 = (inp[9]) ? node1862 : 1'b1;
														assign node1862 = (inp[10]) ? 1'b1 : 1'b0;
													assign node1865 = (inp[10]) ? 1'b0 : node1866;
														assign node1866 = (inp[9]) ? 1'b1 : 1'b0;
												assign node1870 = (inp[10]) ? 1'b1 : node1871;
													assign node1871 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1875 = (inp[5]) ? 1'b0 : node1876;
									assign node1876 = (inp[6]) ? node1878 : 1'b0;
										assign node1878 = (inp[3]) ? node1884 : node1879;
											assign node1879 = (inp[9]) ? node1881 : 1'b1;
												assign node1881 = (inp[10]) ? 1'b1 : 1'b0;
											assign node1884 = (inp[7]) ? node1890 : node1885;
												assign node1885 = (inp[10]) ? 1'b0 : node1886;
													assign node1886 = (inp[9]) ? 1'b1 : 1'b0;
												assign node1890 = (inp[9]) ? node1892 : 1'b1;
													assign node1892 = (inp[10]) ? 1'b1 : 1'b0;
						assign node1896 = (inp[2]) ? node2062 : node1897;
							assign node1897 = (inp[14]) ? node1981 : node1898;
								assign node1898 = (inp[6]) ? node1920 : node1899;
									assign node1899 = (inp[12]) ? node1901 : 1'b1;
										assign node1901 = (inp[15]) ? 1'b1 : node1902;
											assign node1902 = (inp[7]) ? node1914 : node1903;
												assign node1903 = (inp[3]) ? node1909 : node1904;
													assign node1904 = (inp[9]) ? node1906 : 1'b0;
														assign node1906 = (inp[10]) ? 1'b0 : 1'b1;
													assign node1909 = (inp[9]) ? node1911 : 1'b1;
														assign node1911 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1914 = (inp[9]) ? node1916 : 1'b0;
													assign node1916 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1920 = (inp[5]) ? node1960 : node1921;
										assign node1921 = (inp[12]) ? node1939 : node1922;
											assign node1922 = (inp[3]) ? node1928 : node1923;
												assign node1923 = (inp[9]) ? node1925 : 1'b0;
													assign node1925 = (inp[10]) ? 1'b0 : 1'b1;
												assign node1928 = (inp[7]) ? node1934 : node1929;
													assign node1929 = (inp[9]) ? node1931 : 1'b1;
														assign node1931 = (inp[10]) ? 1'b1 : 1'b0;
													assign node1934 = (inp[10]) ? 1'b0 : node1935;
														assign node1935 = (inp[9]) ? 1'b1 : 1'b0;
											assign node1939 = (inp[15]) ? node1941 : 1'b1;
												assign node1941 = (inp[7]) ? node1953 : node1942;
													assign node1942 = (inp[3]) ? node1948 : node1943;
														assign node1943 = (inp[1]) ? node1945 : 1'b0;
															assign node1945 = (inp[10]) ? 1'b0 : 1'b1;
														assign node1948 = (inp[10]) ? 1'b1 : node1949;
															assign node1949 = (inp[9]) ? 1'b0 : 1'b1;
													assign node1953 = (inp[1]) ? 1'b0 : node1954;
														assign node1954 = (inp[10]) ? 1'b0 : node1955;
															assign node1955 = (inp[9]) ? 1'b1 : 1'b0;
										assign node1960 = (inp[12]) ? node1962 : 1'b1;
											assign node1962 = (inp[15]) ? 1'b1 : node1963;
												assign node1963 = (inp[9]) ? node1969 : node1964;
													assign node1964 = (inp[3]) ? node1966 : 1'b0;
														assign node1966 = (inp[7]) ? 1'b0 : 1'b1;
													assign node1969 = (inp[10]) ? node1975 : node1970;
														assign node1970 = (inp[3]) ? node1972 : 1'b1;
															assign node1972 = (inp[7]) ? 1'b1 : 1'b0;
														assign node1975 = (inp[3]) ? node1977 : 1'b0;
															assign node1977 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1981 = (inp[6]) ? node2003 : node1982;
									assign node1982 = (inp[15]) ? 1'b0 : node1983;
										assign node1983 = (inp[12]) ? node1985 : 1'b0;
											assign node1985 = (inp[10]) ? node1997 : node1986;
												assign node1986 = (inp[9]) ? node1992 : node1987;
													assign node1987 = (inp[3]) ? node1989 : 1'b1;
														assign node1989 = (inp[7]) ? 1'b1 : 1'b0;
													assign node1992 = (inp[7]) ? 1'b0 : node1993;
														assign node1993 = (inp[3]) ? 1'b1 : 1'b0;
												assign node1997 = (inp[7]) ? 1'b1 : node1998;
													assign node1998 = (inp[3]) ? 1'b0 : 1'b1;
									assign node2003 = (inp[5]) ? node2041 : node2004;
										assign node2004 = (inp[12]) ? node2022 : node2005;
											assign node2005 = (inp[3]) ? node2011 : node2006;
												assign node2006 = (inp[9]) ? node2008 : 1'b1;
													assign node2008 = (inp[10]) ? 1'b1 : 1'b0;
												assign node2011 = (inp[7]) ? node2017 : node2012;
													assign node2012 = (inp[10]) ? 1'b0 : node2013;
														assign node2013 = (inp[9]) ? 1'b1 : 1'b0;
													assign node2017 = (inp[10]) ? 1'b1 : node2018;
														assign node2018 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2022 = (inp[15]) ? node2024 : 1'b0;
												assign node2024 = (inp[9]) ? node2030 : node2025;
													assign node2025 = (inp[7]) ? 1'b1 : node2026;
														assign node2026 = (inp[3]) ? 1'b0 : 1'b1;
													assign node2030 = (inp[10]) ? node2036 : node2031;
														assign node2031 = (inp[3]) ? node2033 : 1'b0;
															assign node2033 = (inp[7]) ? 1'b0 : 1'b1;
														assign node2036 = (inp[3]) ? node2038 : 1'b1;
															assign node2038 = (inp[7]) ? 1'b1 : 1'b0;
										assign node2041 = (inp[15]) ? 1'b0 : node2042;
											assign node2042 = (inp[12]) ? node2044 : 1'b0;
												assign node2044 = (inp[10]) ? node2056 : node2045;
													assign node2045 = (inp[9]) ? node2051 : node2046;
														assign node2046 = (inp[7]) ? 1'b1 : node2047;
															assign node2047 = (inp[3]) ? 1'b0 : 1'b1;
														assign node2051 = (inp[7]) ? 1'b0 : node2052;
															assign node2052 = (inp[3]) ? 1'b1 : 1'b0;
													assign node2056 = (inp[3]) ? node2058 : 1'b1;
														assign node2058 = (inp[7]) ? 1'b1 : 1'b0;
							assign node2062 = (inp[12]) ? node2084 : node2063;
								assign node2063 = (inp[5]) ? 1'b1 : node2064;
									assign node2064 = (inp[6]) ? node2066 : 1'b1;
										assign node2066 = (inp[9]) ? node2072 : node2067;
											assign node2067 = (inp[3]) ? node2069 : 1'b0;
												assign node2069 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2072 = (inp[10]) ? node2078 : node2073;
												assign node2073 = (inp[3]) ? node2075 : 1'b1;
													assign node2075 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2078 = (inp[7]) ? 1'b0 : node2079;
													assign node2079 = (inp[3]) ? 1'b1 : 1'b0;
								assign node2084 = (inp[15]) ? node2122 : node2085;
									assign node2085 = (inp[5]) ? node2105 : node2086;
										assign node2086 = (inp[6]) ? 1'b1 : node2087;
											assign node2087 = (inp[9]) ? node2093 : node2088;
												assign node2088 = (inp[7]) ? 1'b0 : node2089;
													assign node2089 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2093 = (inp[10]) ? node2099 : node2094;
													assign node2094 = (inp[3]) ? node2096 : 1'b1;
														assign node2096 = (inp[7]) ? 1'b1 : 1'b0;
													assign node2099 = (inp[7]) ? 1'b0 : node2100;
														assign node2100 = (inp[3]) ? 1'b1 : 1'b0;
										assign node2105 = (inp[10]) ? node2117 : node2106;
											assign node2106 = (inp[9]) ? node2112 : node2107;
												assign node2107 = (inp[7]) ? 1'b0 : node2108;
													assign node2108 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2112 = (inp[3]) ? node2114 : 1'b1;
													assign node2114 = (inp[7]) ? 1'b1 : 1'b0;
											assign node2117 = (inp[7]) ? 1'b0 : node2118;
												assign node2118 = (inp[3]) ? 1'b1 : 1'b0;
									assign node2122 = (inp[5]) ? 1'b1 : node2123;
										assign node2123 = (inp[6]) ? node2125 : 1'b1;
											assign node2125 = (inp[10]) ? node2137 : node2126;
												assign node2126 = (inp[9]) ? node2132 : node2127;
													assign node2127 = (inp[7]) ? 1'b0 : node2128;
														assign node2128 = (inp[3]) ? 1'b1 : 1'b0;
													assign node2132 = (inp[7]) ? 1'b1 : node2133;
														assign node2133 = (inp[3]) ? 1'b0 : 1'b1;
												assign node2137 = (inp[3]) ? node2139 : 1'b0;
													assign node2139 = (inp[7]) ? 1'b0 : 1'b1;
					assign node2143 = (inp[14]) ? node2225 : node2144;
						assign node2144 = (inp[12]) ? node2166 : node2145;
							assign node2145 = (inp[5]) ? 1'b0 : node2146;
								assign node2146 = (inp[6]) ? node2148 : 1'b0;
									assign node2148 = (inp[9]) ? node2154 : node2149;
										assign node2149 = (inp[7]) ? 1'b1 : node2150;
											assign node2150 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2154 = (inp[10]) ? node2160 : node2155;
											assign node2155 = (inp[3]) ? node2157 : 1'b0;
												assign node2157 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2160 = (inp[3]) ? node2162 : 1'b1;
												assign node2162 = (inp[7]) ? 1'b1 : 1'b0;
							assign node2166 = (inp[15]) ? node2204 : node2167;
								assign node2167 = (inp[6]) ? node2185 : node2168;
									assign node2168 = (inp[10]) ? node2180 : node2169;
										assign node2169 = (inp[9]) ? node2175 : node2170;
											assign node2170 = (inp[3]) ? node2172 : 1'b1;
												assign node2172 = (inp[7]) ? 1'b1 : 1'b0;
											assign node2175 = (inp[7]) ? 1'b0 : node2176;
												assign node2176 = (inp[3]) ? 1'b1 : 1'b0;
										assign node2180 = (inp[3]) ? node2182 : 1'b1;
											assign node2182 = (inp[7]) ? 1'b1 : 1'b0;
									assign node2185 = (inp[5]) ? node2187 : 1'b0;
										assign node2187 = (inp[9]) ? node2193 : node2188;
											assign node2188 = (inp[7]) ? 1'b1 : node2189;
												assign node2189 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2193 = (inp[10]) ? node2199 : node2194;
												assign node2194 = (inp[3]) ? node2196 : 1'b0;
													assign node2196 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2199 = (inp[3]) ? node2201 : 1'b1;
													assign node2201 = (inp[7]) ? 1'b1 : 1'b0;
								assign node2204 = (inp[5]) ? 1'b0 : node2205;
									assign node2205 = (inp[6]) ? node2207 : 1'b0;
										assign node2207 = (inp[7]) ? node2219 : node2208;
											assign node2208 = (inp[3]) ? node2214 : node2209;
												assign node2209 = (inp[10]) ? 1'b1 : node2210;
													assign node2210 = (inp[9]) ? 1'b0 : 1'b1;
												assign node2214 = (inp[9]) ? node2216 : 1'b0;
													assign node2216 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2219 = (inp[9]) ? node2221 : 1'b1;
												assign node2221 = (inp[10]) ? 1'b1 : 1'b0;
						assign node2225 = (inp[2]) ? node2307 : node2226;
							assign node2226 = (inp[15]) ? node2286 : node2227;
								assign node2227 = (inp[12]) ? node2249 : node2228;
									assign node2228 = (inp[6]) ? node2230 : 1'b1;
										assign node2230 = (inp[5]) ? 1'b1 : node2231;
											assign node2231 = (inp[3]) ? node2237 : node2232;
												assign node2232 = (inp[10]) ? 1'b0 : node2233;
													assign node2233 = (inp[9]) ? 1'b1 : 1'b0;
												assign node2237 = (inp[7]) ? node2243 : node2238;
													assign node2238 = (inp[9]) ? node2240 : 1'b1;
														assign node2240 = (inp[10]) ? 1'b1 : 1'b0;
													assign node2243 = (inp[9]) ? node2245 : 1'b0;
														assign node2245 = (inp[10]) ? 1'b0 : 1'b1;
									assign node2249 = (inp[6]) ? node2267 : node2250;
										assign node2250 = (inp[10]) ? node2262 : node2251;
											assign node2251 = (inp[9]) ? node2257 : node2252;
												assign node2252 = (inp[3]) ? node2254 : 1'b0;
													assign node2254 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2257 = (inp[7]) ? 1'b1 : node2258;
													assign node2258 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2262 = (inp[7]) ? 1'b0 : node2263;
												assign node2263 = (inp[3]) ? 1'b1 : 1'b0;
										assign node2267 = (inp[5]) ? node2269 : 1'b1;
											assign node2269 = (inp[10]) ? node2281 : node2270;
												assign node2270 = (inp[9]) ? node2276 : node2271;
													assign node2271 = (inp[7]) ? 1'b0 : node2272;
														assign node2272 = (inp[3]) ? 1'b1 : 1'b0;
													assign node2276 = (inp[3]) ? node2278 : 1'b1;
														assign node2278 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2281 = (inp[3]) ? node2283 : 1'b0;
													assign node2283 = (inp[7]) ? 1'b0 : 1'b1;
								assign node2286 = (inp[5]) ? 1'b1 : node2287;
									assign node2287 = (inp[6]) ? node2289 : 1'b1;
										assign node2289 = (inp[9]) ? node2295 : node2290;
											assign node2290 = (inp[3]) ? node2292 : 1'b0;
												assign node2292 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2295 = (inp[10]) ? node2301 : node2296;
												assign node2296 = (inp[7]) ? 1'b1 : node2297;
													assign node2297 = (inp[3]) ? 1'b0 : 1'b1;
												assign node2301 = (inp[7]) ? 1'b0 : node2302;
													assign node2302 = (inp[3]) ? 1'b1 : 1'b0;
							assign node2307 = (inp[15]) ? node2367 : node2308;
								assign node2308 = (inp[12]) ? node2330 : node2309;
									assign node2309 = (inp[5]) ? 1'b0 : node2310;
										assign node2310 = (inp[6]) ? node2312 : 1'b0;
											assign node2312 = (inp[9]) ? node2318 : node2313;
												assign node2313 = (inp[3]) ? node2315 : 1'b1;
													assign node2315 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2318 = (inp[10]) ? node2324 : node2319;
													assign node2319 = (inp[3]) ? node2321 : 1'b0;
														assign node2321 = (inp[7]) ? 1'b0 : 1'b1;
													assign node2324 = (inp[7]) ? 1'b1 : node2325;
														assign node2325 = (inp[3]) ? 1'b0 : 1'b1;
									assign node2330 = (inp[6]) ? node2348 : node2331;
										assign node2331 = (inp[9]) ? node2337 : node2332;
											assign node2332 = (inp[7]) ? 1'b1 : node2333;
												assign node2333 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2337 = (inp[10]) ? node2343 : node2338;
												assign node2338 = (inp[7]) ? 1'b0 : node2339;
													assign node2339 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2343 = (inp[3]) ? node2345 : 1'b1;
													assign node2345 = (inp[7]) ? 1'b1 : 1'b0;
										assign node2348 = (inp[5]) ? node2350 : 1'b0;
											assign node2350 = (inp[10]) ? node2362 : node2351;
												assign node2351 = (inp[9]) ? node2357 : node2352;
													assign node2352 = (inp[7]) ? 1'b1 : node2353;
														assign node2353 = (inp[3]) ? 1'b0 : 1'b1;
													assign node2357 = (inp[3]) ? node2359 : 1'b0;
														assign node2359 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2362 = (inp[3]) ? node2364 : 1'b1;
													assign node2364 = (inp[7]) ? 1'b1 : 1'b0;
								assign node2367 = (inp[5]) ? 1'b0 : node2368;
									assign node2368 = (inp[6]) ? node2370 : 1'b0;
										assign node2370 = (inp[10]) ? node2382 : node2371;
											assign node2371 = (inp[9]) ? node2377 : node2372;
												assign node2372 = (inp[3]) ? node2374 : 1'b1;
													assign node2374 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2377 = (inp[3]) ? node2379 : 1'b0;
													assign node2379 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2382 = (inp[3]) ? node2384 : 1'b1;
												assign node2384 = (inp[7]) ? 1'b1 : 1'b0;
		assign node2388 = (inp[1]) ? node2470 : node2389;
			assign node2389 = (inp[5]) ? node2449 : node2390;
				assign node2390 = (inp[6]) ? node2412 : node2391;
					assign node2391 = (inp[12]) ? node2393 : 1'b1;
						assign node2393 = (inp[15]) ? 1'b1 : node2394;
							assign node2394 = (inp[7]) ? node2406 : node2395;
								assign node2395 = (inp[3]) ? node2401 : node2396;
									assign node2396 = (inp[10]) ? 1'b0 : node2397;
										assign node2397 = (inp[9]) ? 1'b1 : 1'b0;
									assign node2401 = (inp[10]) ? 1'b1 : node2402;
										assign node2402 = (inp[9]) ? 1'b0 : 1'b1;
								assign node2406 = (inp[9]) ? node2408 : 1'b0;
									assign node2408 = (inp[10]) ? 1'b0 : 1'b1;
					assign node2412 = (inp[12]) ? node2430 : node2413;
						assign node2413 = (inp[10]) ? node2425 : node2414;
							assign node2414 = (inp[9]) ? node2420 : node2415;
								assign node2415 = (inp[3]) ? node2417 : 1'b0;
									assign node2417 = (inp[7]) ? 1'b0 : 1'b1;
								assign node2420 = (inp[3]) ? node2422 : 1'b1;
									assign node2422 = (inp[7]) ? 1'b1 : 1'b0;
							assign node2425 = (inp[3]) ? node2427 : 1'b0;
								assign node2427 = (inp[7]) ? 1'b0 : 1'b1;
						assign node2430 = (inp[15]) ? node2432 : 1'b1;
							assign node2432 = (inp[7]) ? node2444 : node2433;
								assign node2433 = (inp[3]) ? node2439 : node2434;
									assign node2434 = (inp[10]) ? 1'b0 : node2435;
										assign node2435 = (inp[9]) ? 1'b1 : 1'b0;
									assign node2439 = (inp[10]) ? 1'b1 : node2440;
										assign node2440 = (inp[9]) ? 1'b0 : 1'b1;
								assign node2444 = (inp[10]) ? 1'b0 : node2445;
									assign node2445 = (inp[9]) ? 1'b1 : 1'b0;
				assign node2449 = (inp[12]) ? node2451 : 1'b1;
					assign node2451 = (inp[15]) ? 1'b1 : node2452;
						assign node2452 = (inp[3]) ? node2458 : node2453;
							assign node2453 = (inp[10]) ? 1'b0 : node2454;
								assign node2454 = (inp[9]) ? 1'b1 : 1'b0;
							assign node2458 = (inp[7]) ? node2464 : node2459;
								assign node2459 = (inp[10]) ? 1'b1 : node2460;
									assign node2460 = (inp[9]) ? 1'b0 : 1'b1;
								assign node2464 = (inp[10]) ? 1'b0 : node2465;
									assign node2465 = (inp[9]) ? 1'b1 : 1'b0;
			assign node2470 = (inp[8]) ? node3198 : node2471;
				assign node2471 = (inp[13]) ? node2717 : node2472;
					assign node2472 = (inp[14]) ? node2554 : node2473;
						assign node2473 = (inp[5]) ? node2533 : node2474;
							assign node2474 = (inp[6]) ? node2496 : node2475;
								assign node2475 = (inp[15]) ? 1'b0 : node2476;
									assign node2476 = (inp[12]) ? node2478 : 1'b0;
										assign node2478 = (inp[7]) ? node2490 : node2479;
											assign node2479 = (inp[3]) ? node2485 : node2480;
												assign node2480 = (inp[10]) ? 1'b1 : node2481;
													assign node2481 = (inp[9]) ? 1'b0 : 1'b1;
												assign node2485 = (inp[9]) ? node2487 : 1'b0;
													assign node2487 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2490 = (inp[9]) ? node2492 : 1'b1;
												assign node2492 = (inp[10]) ? 1'b1 : 1'b0;
								assign node2496 = (inp[15]) ? node2516 : node2497;
									assign node2497 = (inp[12]) ? 1'b0 : node2498;
										assign node2498 = (inp[10]) ? node2510 : node2499;
											assign node2499 = (inp[9]) ? node2505 : node2500;
												assign node2500 = (inp[3]) ? node2502 : 1'b1;
													assign node2502 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2505 = (inp[3]) ? node2507 : 1'b0;
													assign node2507 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2510 = (inp[7]) ? 1'b1 : node2511;
												assign node2511 = (inp[3]) ? 1'b0 : 1'b1;
									assign node2516 = (inp[7]) ? node2528 : node2517;
										assign node2517 = (inp[3]) ? node2523 : node2518;
											assign node2518 = (inp[9]) ? node2520 : 1'b1;
												assign node2520 = (inp[10]) ? 1'b1 : 1'b0;
											assign node2523 = (inp[9]) ? node2525 : 1'b0;
												assign node2525 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2528 = (inp[9]) ? node2530 : 1'b1;
											assign node2530 = (inp[10]) ? 1'b1 : 1'b0;
							assign node2533 = (inp[15]) ? 1'b0 : node2534;
								assign node2534 = (inp[12]) ? node2536 : 1'b0;
									assign node2536 = (inp[9]) ? node2542 : node2537;
										assign node2537 = (inp[7]) ? 1'b1 : node2538;
											assign node2538 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2542 = (inp[10]) ? node2548 : node2543;
											assign node2543 = (inp[3]) ? node2545 : 1'b0;
												assign node2545 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2548 = (inp[3]) ? node2550 : 1'b1;
												assign node2550 = (inp[7]) ? 1'b1 : 1'b0;
						assign node2554 = (inp[2]) ? node2636 : node2555;
							assign node2555 = (inp[6]) ? node2577 : node2556;
								assign node2556 = (inp[12]) ? node2558 : 1'b1;
									assign node2558 = (inp[15]) ? 1'b1 : node2559;
										assign node2559 = (inp[7]) ? node2571 : node2560;
											assign node2560 = (inp[3]) ? node2566 : node2561;
												assign node2561 = (inp[9]) ? node2563 : 1'b0;
													assign node2563 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2566 = (inp[10]) ? 1'b1 : node2567;
													assign node2567 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2571 = (inp[10]) ? 1'b0 : node2572;
												assign node2572 = (inp[9]) ? 1'b1 : 1'b0;
								assign node2577 = (inp[5]) ? node2615 : node2578;
									assign node2578 = (inp[12]) ? node2596 : node2579;
										assign node2579 = (inp[3]) ? node2585 : node2580;
											assign node2580 = (inp[10]) ? 1'b0 : node2581;
												assign node2581 = (inp[9]) ? 1'b1 : 1'b0;
											assign node2585 = (inp[7]) ? node2591 : node2586;
												assign node2586 = (inp[9]) ? node2588 : 1'b1;
													assign node2588 = (inp[10]) ? 1'b1 : 1'b0;
												assign node2591 = (inp[10]) ? 1'b0 : node2592;
													assign node2592 = (inp[9]) ? 1'b1 : 1'b0;
										assign node2596 = (inp[15]) ? node2598 : 1'b1;
											assign node2598 = (inp[10]) ? node2610 : node2599;
												assign node2599 = (inp[9]) ? node2605 : node2600;
													assign node2600 = (inp[7]) ? 1'b0 : node2601;
														assign node2601 = (inp[3]) ? 1'b1 : 1'b0;
													assign node2605 = (inp[3]) ? node2607 : 1'b1;
														assign node2607 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2610 = (inp[7]) ? 1'b0 : node2611;
													assign node2611 = (inp[3]) ? 1'b1 : 1'b0;
									assign node2615 = (inp[15]) ? 1'b1 : node2616;
										assign node2616 = (inp[12]) ? node2618 : 1'b1;
											assign node2618 = (inp[3]) ? node2624 : node2619;
												assign node2619 = (inp[10]) ? 1'b0 : node2620;
													assign node2620 = (inp[9]) ? 1'b1 : 1'b0;
												assign node2624 = (inp[7]) ? node2630 : node2625;
													assign node2625 = (inp[10]) ? 1'b1 : node2626;
														assign node2626 = (inp[9]) ? 1'b0 : 1'b1;
													assign node2630 = (inp[10]) ? 1'b0 : node2631;
														assign node2631 = (inp[9]) ? 1'b1 : 1'b0;
							assign node2636 = (inp[15]) ? node2696 : node2637;
								assign node2637 = (inp[12]) ? node2659 : node2638;
									assign node2638 = (inp[6]) ? node2640 : 1'b0;
										assign node2640 = (inp[5]) ? 1'b0 : node2641;
											assign node2641 = (inp[9]) ? node2647 : node2642;
												assign node2642 = (inp[7]) ? 1'b1 : node2643;
													assign node2643 = (inp[3]) ? 1'b0 : 1'b1;
												assign node2647 = (inp[10]) ? node2653 : node2648;
													assign node2648 = (inp[7]) ? 1'b0 : node2649;
														assign node2649 = (inp[3]) ? 1'b1 : 1'b0;
													assign node2653 = (inp[7]) ? 1'b1 : node2654;
														assign node2654 = (inp[3]) ? 1'b0 : 1'b1;
									assign node2659 = (inp[6]) ? node2677 : node2660;
										assign node2660 = (inp[10]) ? node2672 : node2661;
											assign node2661 = (inp[9]) ? node2667 : node2662;
												assign node2662 = (inp[3]) ? node2664 : 1'b1;
													assign node2664 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2667 = (inp[7]) ? 1'b0 : node2668;
													assign node2668 = (inp[3]) ? 1'b1 : 1'b0;
											assign node2672 = (inp[7]) ? 1'b1 : node2673;
												assign node2673 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2677 = (inp[5]) ? node2679 : 1'b0;
											assign node2679 = (inp[7]) ? node2691 : node2680;
												assign node2680 = (inp[3]) ? node2686 : node2681;
													assign node2681 = (inp[9]) ? node2683 : 1'b1;
														assign node2683 = (inp[10]) ? 1'b1 : 1'b0;
													assign node2686 = (inp[10]) ? 1'b0 : node2687;
														assign node2687 = (inp[9]) ? 1'b1 : 1'b0;
												assign node2691 = (inp[9]) ? node2693 : 1'b1;
													assign node2693 = (inp[10]) ? 1'b1 : 1'b0;
								assign node2696 = (inp[6]) ? node2698 : 1'b0;
									assign node2698 = (inp[5]) ? 1'b0 : node2699;
										assign node2699 = (inp[10]) ? node2711 : node2700;
											assign node2700 = (inp[9]) ? node2706 : node2701;
												assign node2701 = (inp[7]) ? 1'b1 : node2702;
													assign node2702 = (inp[3]) ? 1'b0 : 1'b1;
												assign node2706 = (inp[7]) ? 1'b0 : node2707;
													assign node2707 = (inp[3]) ? 1'b1 : 1'b0;
											assign node2711 = (inp[7]) ? 1'b1 : node2712;
												assign node2712 = (inp[3]) ? 1'b0 : 1'b1;
					assign node2717 = (inp[11]) ? node2963 : node2718;
						assign node2718 = (inp[14]) ? node2800 : node2719;
							assign node2719 = (inp[12]) ? node2741 : node2720;
								assign node2720 = (inp[5]) ? 1'b1 : node2721;
									assign node2721 = (inp[6]) ? node2723 : 1'b1;
										assign node2723 = (inp[9]) ? node2729 : node2724;
											assign node2724 = (inp[3]) ? node2726 : 1'b0;
												assign node2726 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2729 = (inp[10]) ? node2735 : node2730;
												assign node2730 = (inp[3]) ? node2732 : 1'b1;
													assign node2732 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2735 = (inp[7]) ? 1'b0 : node2736;
													assign node2736 = (inp[3]) ? 1'b1 : 1'b0;
								assign node2741 = (inp[15]) ? node2779 : node2742;
									assign node2742 = (inp[5]) ? node2762 : node2743;
										assign node2743 = (inp[6]) ? 1'b1 : node2744;
											assign node2744 = (inp[10]) ? node2756 : node2745;
												assign node2745 = (inp[9]) ? node2751 : node2746;
													assign node2746 = (inp[3]) ? node2748 : 1'b0;
														assign node2748 = (inp[7]) ? 1'b0 : 1'b1;
													assign node2751 = (inp[3]) ? node2753 : 1'b1;
														assign node2753 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2756 = (inp[3]) ? node2758 : 1'b0;
													assign node2758 = (inp[7]) ? 1'b0 : 1'b1;
										assign node2762 = (inp[7]) ? node2774 : node2763;
											assign node2763 = (inp[3]) ? node2769 : node2764;
												assign node2764 = (inp[10]) ? 1'b0 : node2765;
													assign node2765 = (inp[9]) ? 1'b1 : 1'b0;
												assign node2769 = (inp[10]) ? 1'b1 : node2770;
													assign node2770 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2774 = (inp[10]) ? 1'b0 : node2775;
												assign node2775 = (inp[9]) ? 1'b1 : 1'b0;
									assign node2779 = (inp[5]) ? 1'b1 : node2780;
										assign node2780 = (inp[6]) ? node2782 : 1'b1;
											assign node2782 = (inp[7]) ? node2794 : node2783;
												assign node2783 = (inp[3]) ? node2789 : node2784;
													assign node2784 = (inp[10]) ? 1'b0 : node2785;
														assign node2785 = (inp[9]) ? 1'b1 : 1'b0;
													assign node2789 = (inp[9]) ? node2791 : 1'b1;
														assign node2791 = (inp[10]) ? 1'b1 : 1'b0;
												assign node2794 = (inp[9]) ? node2796 : 1'b0;
													assign node2796 = (inp[10]) ? 1'b0 : 1'b1;
							assign node2800 = (inp[2]) ? node2882 : node2801;
								assign node2801 = (inp[6]) ? node2823 : node2802;
									assign node2802 = (inp[15]) ? 1'b0 : node2803;
										assign node2803 = (inp[12]) ? node2805 : 1'b0;
											assign node2805 = (inp[3]) ? node2811 : node2806;
												assign node2806 = (inp[10]) ? 1'b1 : node2807;
													assign node2807 = (inp[9]) ? 1'b0 : 1'b1;
												assign node2811 = (inp[7]) ? node2817 : node2812;
													assign node2812 = (inp[10]) ? 1'b0 : node2813;
														assign node2813 = (inp[9]) ? 1'b1 : 1'b0;
													assign node2817 = (inp[9]) ? node2819 : 1'b1;
														assign node2819 = (inp[10]) ? 1'b1 : 1'b0;
									assign node2823 = (inp[5]) ? node2861 : node2824;
										assign node2824 = (inp[15]) ? node2844 : node2825;
											assign node2825 = (inp[12]) ? 1'b0 : node2826;
												assign node2826 = (inp[10]) ? node2838 : node2827;
													assign node2827 = (inp[9]) ? node2833 : node2828;
														assign node2828 = (inp[3]) ? node2830 : 1'b1;
															assign node2830 = (inp[7]) ? 1'b1 : 1'b0;
														assign node2833 = (inp[3]) ? node2835 : 1'b0;
															assign node2835 = (inp[7]) ? 1'b0 : 1'b1;
													assign node2838 = (inp[3]) ? node2840 : 1'b1;
														assign node2840 = (inp[7]) ? 1'b1 : 1'b0;
											assign node2844 = (inp[7]) ? node2856 : node2845;
												assign node2845 = (inp[3]) ? node2851 : node2846;
													assign node2846 = (inp[10]) ? 1'b1 : node2847;
														assign node2847 = (inp[9]) ? 1'b0 : 1'b1;
													assign node2851 = (inp[10]) ? 1'b0 : node2852;
														assign node2852 = (inp[9]) ? 1'b1 : 1'b0;
												assign node2856 = (inp[9]) ? node2858 : 1'b1;
													assign node2858 = (inp[10]) ? 1'b1 : 1'b0;
										assign node2861 = (inp[15]) ? 1'b0 : node2862;
											assign node2862 = (inp[12]) ? node2864 : 1'b0;
												assign node2864 = (inp[7]) ? node2876 : node2865;
													assign node2865 = (inp[3]) ? node2871 : node2866;
														assign node2866 = (inp[10]) ? 1'b1 : node2867;
															assign node2867 = (inp[9]) ? 1'b0 : 1'b1;
														assign node2871 = (inp[9]) ? node2873 : 1'b0;
															assign node2873 = (inp[10]) ? 1'b0 : 1'b1;
													assign node2876 = (inp[9]) ? node2878 : 1'b1;
														assign node2878 = (inp[10]) ? 1'b1 : 1'b0;
								assign node2882 = (inp[15]) ? node2942 : node2883;
									assign node2883 = (inp[12]) ? node2905 : node2884;
										assign node2884 = (inp[5]) ? 1'b1 : node2885;
											assign node2885 = (inp[6]) ? node2887 : 1'b1;
												assign node2887 = (inp[7]) ? node2899 : node2888;
													assign node2888 = (inp[3]) ? node2894 : node2889;
														assign node2889 = (inp[10]) ? 1'b0 : node2890;
															assign node2890 = (inp[9]) ? 1'b1 : 1'b0;
														assign node2894 = (inp[9]) ? node2896 : 1'b1;
															assign node2896 = (inp[10]) ? 1'b1 : 1'b0;
													assign node2899 = (inp[10]) ? 1'b0 : node2900;
														assign node2900 = (inp[9]) ? 1'b1 : 1'b0;
										assign node2905 = (inp[6]) ? node2923 : node2906;
											assign node2906 = (inp[9]) ? node2912 : node2907;
												assign node2907 = (inp[3]) ? node2909 : 1'b0;
													assign node2909 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2912 = (inp[10]) ? node2918 : node2913;
													assign node2913 = (inp[7]) ? 1'b1 : node2914;
														assign node2914 = (inp[3]) ? 1'b0 : 1'b1;
													assign node2918 = (inp[3]) ? node2920 : 1'b0;
														assign node2920 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2923 = (inp[5]) ? node2925 : 1'b1;
												assign node2925 = (inp[10]) ? node2937 : node2926;
													assign node2926 = (inp[9]) ? node2932 : node2927;
														assign node2927 = (inp[3]) ? node2929 : 1'b0;
															assign node2929 = (inp[7]) ? 1'b0 : 1'b1;
														assign node2932 = (inp[3]) ? node2934 : 1'b1;
															assign node2934 = (inp[7]) ? 1'b1 : 1'b0;
													assign node2937 = (inp[3]) ? node2939 : 1'b0;
														assign node2939 = (inp[7]) ? 1'b0 : 1'b1;
									assign node2942 = (inp[5]) ? 1'b1 : node2943;
										assign node2943 = (inp[6]) ? node2945 : 1'b1;
											assign node2945 = (inp[3]) ? node2951 : node2946;
												assign node2946 = (inp[9]) ? node2948 : 1'b0;
													assign node2948 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2951 = (inp[7]) ? node2957 : node2952;
													assign node2952 = (inp[9]) ? node2954 : 1'b1;
														assign node2954 = (inp[10]) ? 1'b1 : 1'b0;
													assign node2957 = (inp[10]) ? 1'b0 : node2958;
														assign node2958 = (inp[9]) ? 1'b1 : 1'b0;
						assign node2963 = (inp[2]) ? node3117 : node2964;
							assign node2964 = (inp[14]) ? node3040 : node2965;
								assign node2965 = (inp[5]) ? node3019 : node2966;
									assign node2966 = (inp[6]) ? node2982 : node2967;
										assign node2967 = (inp[15]) ? 1'b0 : node2968;
											assign node2968 = (inp[12]) ? node2970 : 1'b0;
												assign node2970 = (inp[3]) ? node2972 : 1'b1;
													assign node2972 = (inp[7]) ? node2976 : node2973;
														assign node2973 = (inp[9]) ? 1'b1 : 1'b0;
														assign node2976 = (inp[9]) ? node2978 : 1'b1;
															assign node2978 = (inp[10]) ? 1'b1 : 1'b0;
										assign node2982 = (inp[12]) ? node3000 : node2983;
											assign node2983 = (inp[10]) ? node2995 : node2984;
												assign node2984 = (inp[9]) ? node2990 : node2985;
													assign node2985 = (inp[7]) ? 1'b1 : node2986;
														assign node2986 = (inp[3]) ? 1'b0 : 1'b1;
													assign node2990 = (inp[7]) ? 1'b0 : node2991;
														assign node2991 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2995 = (inp[7]) ? 1'b1 : node2996;
													assign node2996 = (inp[3]) ? 1'b0 : 1'b1;
											assign node3000 = (inp[15]) ? node3002 : 1'b0;
												assign node3002 = (inp[9]) ? node3008 : node3003;
													assign node3003 = (inp[7]) ? 1'b1 : node3004;
														assign node3004 = (inp[3]) ? 1'b0 : 1'b1;
													assign node3008 = (inp[10]) ? node3014 : node3009;
														assign node3009 = (inp[7]) ? 1'b0 : node3010;
															assign node3010 = (inp[3]) ? 1'b1 : 1'b0;
														assign node3014 = (inp[7]) ? 1'b1 : node3015;
															assign node3015 = (inp[3]) ? 1'b0 : 1'b1;
									assign node3019 = (inp[12]) ? node3021 : 1'b0;
										assign node3021 = (inp[15]) ? 1'b0 : node3022;
											assign node3022 = (inp[7]) ? node3034 : node3023;
												assign node3023 = (inp[3]) ? node3029 : node3024;
													assign node3024 = (inp[9]) ? node3026 : 1'b1;
														assign node3026 = (inp[10]) ? 1'b1 : 1'b0;
													assign node3029 = (inp[9]) ? node3031 : 1'b0;
														assign node3031 = (inp[10]) ? 1'b0 : 1'b1;
												assign node3034 = (inp[10]) ? 1'b1 : node3035;
													assign node3035 = (inp[9]) ? 1'b0 : 1'b1;
								assign node3040 = (inp[6]) ? node3062 : node3041;
									assign node3041 = (inp[12]) ? node3043 : 1'b1;
										assign node3043 = (inp[15]) ? 1'b1 : node3044;
											assign node3044 = (inp[7]) ? node3056 : node3045;
												assign node3045 = (inp[3]) ? node3051 : node3046;
													assign node3046 = (inp[9]) ? node3048 : 1'b0;
														assign node3048 = (inp[10]) ? 1'b0 : 1'b1;
													assign node3051 = (inp[10]) ? 1'b1 : node3052;
														assign node3052 = (inp[9]) ? 1'b0 : 1'b1;
												assign node3056 = (inp[9]) ? node3058 : 1'b0;
													assign node3058 = (inp[10]) ? 1'b0 : 1'b1;
									assign node3062 = (inp[5]) ? node3096 : node3063;
										assign node3063 = (inp[12]) ? node3081 : node3064;
											assign node3064 = (inp[9]) ? node3070 : node3065;
												assign node3065 = (inp[7]) ? 1'b0 : node3066;
													assign node3066 = (inp[3]) ? 1'b1 : 1'b0;
												assign node3070 = (inp[10]) ? node3076 : node3071;
													assign node3071 = (inp[3]) ? node3073 : 1'b1;
														assign node3073 = (inp[7]) ? 1'b1 : 1'b0;
													assign node3076 = (inp[7]) ? 1'b0 : node3077;
														assign node3077 = (inp[3]) ? 1'b1 : 1'b0;
											assign node3081 = (inp[15]) ? node3083 : 1'b1;
												assign node3083 = (inp[3]) ? node3089 : node3084;
													assign node3084 = (inp[9]) ? node3086 : 1'b0;
														assign node3086 = (inp[10]) ? 1'b0 : 1'b1;
													assign node3089 = (inp[7]) ? node3093 : node3090;
														assign node3090 = (inp[9]) ? 1'b0 : 1'b1;
														assign node3093 = (inp[10]) ? 1'b0 : 1'b1;
										assign node3096 = (inp[12]) ? node3098 : 1'b1;
											assign node3098 = (inp[15]) ? 1'b1 : node3099;
												assign node3099 = (inp[9]) ? node3105 : node3100;
													assign node3100 = (inp[3]) ? node3102 : 1'b0;
														assign node3102 = (inp[7]) ? 1'b0 : 1'b1;
													assign node3105 = (inp[10]) ? node3111 : node3106;
														assign node3106 = (inp[7]) ? 1'b1 : node3107;
															assign node3107 = (inp[3]) ? 1'b0 : 1'b1;
														assign node3111 = (inp[7]) ? 1'b0 : node3112;
															assign node3112 = (inp[3]) ? 1'b1 : 1'b0;
							assign node3117 = (inp[15]) ? node3177 : node3118;
								assign node3118 = (inp[12]) ? node3140 : node3119;
									assign node3119 = (inp[6]) ? node3121 : 1'b0;
										assign node3121 = (inp[5]) ? 1'b0 : node3122;
											assign node3122 = (inp[7]) ? node3134 : node3123;
												assign node3123 = (inp[3]) ? node3129 : node3124;
													assign node3124 = (inp[9]) ? node3126 : 1'b1;
														assign node3126 = (inp[10]) ? 1'b1 : 1'b0;
													assign node3129 = (inp[9]) ? node3131 : 1'b0;
														assign node3131 = (inp[10]) ? 1'b0 : 1'b1;
												assign node3134 = (inp[10]) ? 1'b1 : node3135;
													assign node3135 = (inp[9]) ? 1'b0 : 1'b1;
									assign node3140 = (inp[6]) ? node3158 : node3141;
										assign node3141 = (inp[9]) ? node3147 : node3142;
											assign node3142 = (inp[3]) ? node3144 : 1'b1;
												assign node3144 = (inp[7]) ? 1'b1 : 1'b0;
											assign node3147 = (inp[10]) ? node3153 : node3148;
												assign node3148 = (inp[3]) ? node3150 : 1'b0;
													assign node3150 = (inp[7]) ? 1'b0 : 1'b1;
												assign node3153 = (inp[3]) ? node3155 : 1'b1;
													assign node3155 = (inp[7]) ? 1'b1 : 1'b0;
										assign node3158 = (inp[5]) ? node3160 : 1'b0;
											assign node3160 = (inp[10]) ? node3172 : node3161;
												assign node3161 = (inp[9]) ? node3167 : node3162;
													assign node3162 = (inp[7]) ? 1'b1 : node3163;
														assign node3163 = (inp[3]) ? 1'b0 : 1'b1;
													assign node3167 = (inp[7]) ? 1'b0 : node3168;
														assign node3168 = (inp[3]) ? 1'b1 : 1'b0;
												assign node3172 = (inp[3]) ? node3174 : 1'b1;
													assign node3174 = (inp[7]) ? 1'b1 : 1'b0;
								assign node3177 = (inp[6]) ? node3179 : 1'b0;
									assign node3179 = (inp[5]) ? 1'b0 : node3180;
										assign node3180 = (inp[7]) ? node3192 : node3181;
											assign node3181 = (inp[3]) ? node3187 : node3182;
												assign node3182 = (inp[9]) ? node3184 : 1'b1;
													assign node3184 = (inp[10]) ? 1'b1 : 1'b0;
												assign node3187 = (inp[10]) ? 1'b0 : node3188;
													assign node3188 = (inp[9]) ? 1'b1 : 1'b0;
											assign node3192 = (inp[9]) ? node3194 : 1'b1;
												assign node3194 = (inp[10]) ? 1'b1 : 1'b0;
				assign node3198 = (inp[12]) ? node3220 : node3199;
					assign node3199 = (inp[5]) ? 1'b1 : node3200;
						assign node3200 = (inp[6]) ? node3202 : 1'b1;
							assign node3202 = (inp[10]) ? node3214 : node3203;
								assign node3203 = (inp[9]) ? node3209 : node3204;
									assign node3204 = (inp[7]) ? 1'b0 : node3205;
										assign node3205 = (inp[3]) ? 1'b1 : 1'b0;
									assign node3209 = (inp[7]) ? 1'b1 : node3210;
										assign node3210 = (inp[3]) ? 1'b0 : 1'b1;
								assign node3214 = (inp[3]) ? node3216 : 1'b0;
									assign node3216 = (inp[7]) ? 1'b0 : 1'b1;
					assign node3220 = (inp[15]) ? node3258 : node3221;
						assign node3221 = (inp[5]) ? node3241 : node3222;
							assign node3222 = (inp[6]) ? 1'b1 : node3223;
								assign node3223 = (inp[3]) ? node3229 : node3224;
									assign node3224 = (inp[10]) ? 1'b0 : node3225;
										assign node3225 = (inp[9]) ? 1'b1 : 1'b0;
									assign node3229 = (inp[7]) ? node3235 : node3230;
										assign node3230 = (inp[9]) ? node3232 : 1'b1;
											assign node3232 = (inp[10]) ? 1'b1 : 1'b0;
										assign node3235 = (inp[10]) ? 1'b0 : node3236;
											assign node3236 = (inp[9]) ? 1'b1 : 1'b0;
							assign node3241 = (inp[7]) ? node3253 : node3242;
								assign node3242 = (inp[3]) ? node3248 : node3243;
									assign node3243 = (inp[9]) ? node3245 : 1'b0;
										assign node3245 = (inp[10]) ? 1'b0 : 1'b1;
									assign node3248 = (inp[9]) ? node3250 : 1'b1;
										assign node3250 = (inp[10]) ? 1'b1 : 1'b0;
								assign node3253 = (inp[9]) ? node3255 : 1'b0;
									assign node3255 = (inp[10]) ? 1'b0 : 1'b1;
						assign node3258 = (inp[5]) ? 1'b1 : node3259;
							assign node3259 = (inp[6]) ? node3261 : 1'b1;
								assign node3261 = (inp[3]) ? node3267 : node3262;
									assign node3262 = (inp[9]) ? node3264 : 1'b0;
										assign node3264 = (inp[10]) ? 1'b0 : 1'b1;
									assign node3267 = (inp[7]) ? node3273 : node3268;
										assign node3268 = (inp[9]) ? node3270 : 1'b1;
											assign node3270 = (inp[10]) ? 1'b1 : 1'b0;
										assign node3273 = (inp[9]) ? node3275 : 1'b0;
											assign node3275 = (inp[10]) ? 1'b0 : 1'b1;

endmodule