module dtc_split66_bm49 (
	input  wire [7-1:0] inp,
	output wire [10-1:0] outp
);

	wire [10-1:0] node1;
	wire [10-1:0] node2;
	wire [10-1:0] node3;
	wire [10-1:0] node4;
	wire [10-1:0] node5;
	wire [10-1:0] node9;
	wire [10-1:0] node10;
	wire [10-1:0] node11;
	wire [10-1:0] node15;
	wire [10-1:0] node18;
	wire [10-1:0] node19;
	wire [10-1:0] node20;
	wire [10-1:0] node21;
	wire [10-1:0] node25;
	wire [10-1:0] node27;
	wire [10-1:0] node30;
	wire [10-1:0] node31;
	wire [10-1:0] node33;
	wire [10-1:0] node36;
	wire [10-1:0] node37;
	wire [10-1:0] node40;
	wire [10-1:0] node43;
	wire [10-1:0] node44;
	wire [10-1:0] node45;
	wire [10-1:0] node46;
	wire [10-1:0] node47;
	wire [10-1:0] node50;
	wire [10-1:0] node53;
	wire [10-1:0] node54;
	wire [10-1:0] node58;
	wire [10-1:0] node59;
	wire [10-1:0] node60;
	wire [10-1:0] node64;
	wire [10-1:0] node65;
	wire [10-1:0] node69;
	wire [10-1:0] node70;
	wire [10-1:0] node71;
	wire [10-1:0] node74;
	wire [10-1:0] node77;
	wire [10-1:0] node78;
	wire [10-1:0] node79;
	wire [10-1:0] node83;
	wire [10-1:0] node85;
	wire [10-1:0] node88;
	wire [10-1:0] node89;
	wire [10-1:0] node90;
	wire [10-1:0] node91;
	wire [10-1:0] node92;
	wire [10-1:0] node95;
	wire [10-1:0] node97;
	wire [10-1:0] node100;
	wire [10-1:0] node101;
	wire [10-1:0] node104;
	wire [10-1:0] node105;
	wire [10-1:0] node109;
	wire [10-1:0] node110;
	wire [10-1:0] node111;
	wire [10-1:0] node114;
	wire [10-1:0] node115;
	wire [10-1:0] node118;
	wire [10-1:0] node121;
	wire [10-1:0] node122;
	wire [10-1:0] node124;
	wire [10-1:0] node127;
	wire [10-1:0] node129;
	wire [10-1:0] node132;
	wire [10-1:0] node133;
	wire [10-1:0] node134;
	wire [10-1:0] node135;
	wire [10-1:0] node137;
	wire [10-1:0] node141;
	wire [10-1:0] node142;
	wire [10-1:0] node143;
	wire [10-1:0] node146;
	wire [10-1:0] node149;
	wire [10-1:0] node150;
	wire [10-1:0] node153;
	wire [10-1:0] node156;
	wire [10-1:0] node157;
	wire [10-1:0] node160;
	wire [10-1:0] node161;
	wire [10-1:0] node163;
	wire [10-1:0] node166;

	assign outp = (inp[3]) ? node88 : node1;
		assign node1 = (inp[1]) ? node43 : node2;
			assign node2 = (inp[0]) ? node18 : node3;
				assign node3 = (inp[2]) ? node9 : node4;
					assign node4 = (inp[5]) ? 10'b1100000001 : node5;
						assign node5 = (inp[4]) ? 10'b1000001101 : 10'b1100001111;
					assign node9 = (inp[4]) ? node15 : node10;
						assign node10 = (inp[6]) ? 10'b1000011110 : node11;
							assign node11 = (inp[5]) ? 10'b1000000110 : 10'b1101000010;
						assign node15 = (inp[6]) ? 10'b1000010000 : 10'b1100001000;
				assign node18 = (inp[2]) ? node30 : node19;
					assign node19 = (inp[5]) ? node25 : node20;
						assign node20 = (inp[6]) ? 10'b0100010111 : node21;
							assign node21 = (inp[4]) ? 10'b0001000011 : 10'b0101010001;
						assign node25 = (inp[4]) ? node27 : 10'b0000001001;
							assign node27 = (inp[6]) ? 10'b0000010011 : 10'b0100001011;
					assign node30 = (inp[4]) ? node36 : node31;
						assign node31 = (inp[5]) ? node33 : 10'b0101000000;
							assign node33 = (inp[6]) ? 10'b0100010000 : 10'b0000000100;
						assign node36 = (inp[5]) ? node40 : node37;
							assign node37 = (inp[6]) ? 10'b0100000110 : 10'b0100011110;
							assign node40 = (inp[6]) ? 10'b0000000010 : 10'b0000011010;
			assign node43 = (inp[0]) ? node69 : node44;
				assign node44 = (inp[2]) ? node58 : node45;
					assign node45 = (inp[6]) ? node53 : node46;
						assign node46 = (inp[4]) ? node50 : node47;
							assign node47 = (inp[5]) ? 10'b0000110110 : 10'b0101110010;
							assign node50 = (inp[5]) ? 10'b0100111000 : 10'b0001110000;
						assign node53 = (inp[5]) ? 10'b0100100000 : node54;
							assign node54 = (inp[4]) ? 10'b0000101100 : 10'b0100101110;
					assign node58 = (inp[4]) ? node64 : node59;
						assign node59 = (inp[6]) ? 10'b0100110001 : node60;
							assign node60 = (inp[5]) ? 10'b0000100101 : 10'b0101100001;
						assign node64 = (inp[5]) ? 10'b0000111011 : node65;
							assign node65 = (inp[6]) ? 10'b0100100111 : 10'b0100111111;
				assign node69 = (inp[2]) ? node77 : node70;
					assign node70 = (inp[6]) ? node74 : node71;
						assign node71 = (inp[4]) ? 10'b1001100001 : 10'b1101100011;
						assign node74 = (inp[4]) ? 10'b1100110101 : 10'b1100110011;
					assign node77 = (inp[6]) ? node83 : node78;
						assign node78 = (inp[4]) ? 10'b1100111100 : node79;
							assign node79 = (inp[5]) ? 10'b1100111010 : 10'b1001110010;
						assign node83 = (inp[4]) ? node85 : 10'b1000101110;
							assign node85 = (inp[5]) ? 10'b1000100000 : 10'b1100100100;
		assign node88 = (inp[1]) ? node132 : node89;
			assign node89 = (inp[0]) ? node109 : node90;
				assign node90 = (inp[2]) ? node100 : node91;
					assign node91 = (inp[6]) ? node95 : node92;
						assign node92 = (inp[5]) ? 10'b1110111000 : 10'b1011110000;
						assign node95 = (inp[4]) ? node97 : 10'b1010101010;
							assign node97 = (inp[5]) ? 10'b1110100000 : 10'b1010101100;
					assign node100 = (inp[4]) ? node104 : node101;
						assign node101 = (inp[6]) ? 10'b1110110001 : 10'b1010100101;
						assign node104 = (inp[6]) ? 10'b1010100011 : node105;
							assign node105 = (inp[5]) ? 10'b1010111011 : 10'b1110111111;
				assign node109 = (inp[2]) ? node121 : node110;
					assign node110 = (inp[5]) ? node114 : node111;
						assign node111 = (inp[6]) ? 10'b0110110110 : 10'b0111110000;
						assign node114 = (inp[4]) ? node118 : node115;
							assign node115 = (inp[6]) ? 10'b0010101000 : 10'b0010110100;
							assign node118 = (inp[6]) ? 10'b0010110010 : 10'b0110101010;
					assign node121 = (inp[4]) ? node127 : node122;
						assign node122 = (inp[5]) ? node124 : 10'b0011110011;
							assign node124 = (inp[6]) ? 10'b0110100011 : 10'b0110111011;
						assign node127 = (inp[6]) ? node129 : 10'b0110111101;
							assign node129 = (inp[5]) ? 10'b0010100001 : 10'b0110100101;
			assign node132 = (inp[2]) ? node156 : node133;
				assign node133 = (inp[0]) ? node141 : node134;
					assign node134 = (inp[5]) ? 10'b1110001011 : node135;
						assign node135 = (inp[6]) ? node137 : 10'b1111010001;
							assign node137 = (inp[4]) ? 10'b1110010111 : 10'b1110001101;
					assign node141 = (inp[6]) ? node149 : node142;
						assign node142 = (inp[4]) ? node146 : node143;
							assign node143 = (inp[5]) ? 10'b0010000111 : 10'b0111000011;
							assign node146 = (inp[5]) ? 10'b0110001001 : 10'b0011000001;
						assign node149 = (inp[5]) ? node153 : node150;
							assign node150 = (inp[4]) ? 10'b0110010101 : 10'b0010011111;
							assign node153 = (inp[4]) ? 10'b0010010001 : 10'b0110010011;
				assign node156 = (inp[0]) ? node160 : node157;
					assign node157 = (inp[5]) ? 10'b1010011010 : 10'b1010011100;
					assign node160 = (inp[5]) ? node166 : node161;
						assign node161 = (inp[4]) ? node163 : 10'b0010001110;
							assign node163 = (inp[6]) ? 10'b0110000100 : 10'b0110011100;
						assign node166 = (inp[4]) ? 10'b0010000000 : 10'b0110000010;

endmodule