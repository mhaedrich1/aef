module dtc_split875_bm58 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node37;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node52;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node63;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node114;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node120;
	wire [3-1:0] node124;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node147;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node181;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node232;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node246;
	wire [3-1:0] node248;
	wire [3-1:0] node250;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node266;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node282;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node310;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node322;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node330;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node346;

	assign outp = (inp[6]) ? node2 : 3'b000;
		assign node2 = (inp[0]) ? node218 : node3;
			assign node3 = (inp[4]) ? node93 : node4;
				assign node4 = (inp[9]) ? node42 : node5;
					assign node5 = (inp[1]) ? 3'b000 : node6;
						assign node6 = (inp[8]) ? node24 : node7;
							assign node7 = (inp[11]) ? 3'b000 : node8;
								assign node8 = (inp[10]) ? node16 : node9;
									assign node9 = (inp[3]) ? 3'b000 : node10;
										assign node10 = (inp[2]) ? 3'b100 : node11;
											assign node11 = (inp[7]) ? 3'b000 : 3'b100;
									assign node16 = (inp[7]) ? node18 : 3'b100;
										assign node18 = (inp[3]) ? node20 : 3'b100;
											assign node20 = (inp[2]) ? 3'b100 : 3'b000;
							assign node24 = (inp[11]) ? node26 : 3'b100;
								assign node26 = (inp[10]) ? node34 : node27;
									assign node27 = (inp[3]) ? 3'b000 : node28;
										assign node28 = (inp[2]) ? 3'b100 : node29;
											assign node29 = (inp[7]) ? 3'b000 : 3'b100;
									assign node34 = (inp[2]) ? 3'b100 : node35;
										assign node35 = (inp[7]) ? node37 : 3'b100;
											assign node37 = (inp[3]) ? 3'b000 : 3'b100;
					assign node42 = (inp[1]) ? node76 : node43;
						assign node43 = (inp[10]) ? node59 : node44;
							assign node44 = (inp[8]) ? node52 : node45;
								assign node45 = (inp[11]) ? 3'b100 : node46;
									assign node46 = (inp[2]) ? 3'b000 : node47;
										assign node47 = (inp[3]) ? 3'b100 : 3'b000;
								assign node52 = (inp[2]) ? node54 : 3'b000;
									assign node54 = (inp[11]) ? 3'b000 : node55;
										assign node55 = (inp[3]) ? 3'b000 : 3'b100;
							assign node59 = (inp[8]) ? node67 : node60;
								assign node60 = (inp[2]) ? 3'b000 : node61;
									assign node61 = (inp[11]) ? node63 : 3'b000;
										assign node63 = (inp[3]) ? 3'b100 : 3'b000;
								assign node67 = (inp[2]) ? 3'b100 : node68;
									assign node68 = (inp[11]) ? node70 : 3'b100;
										assign node70 = (inp[3]) ? 3'b000 : node71;
											assign node71 = (inp[7]) ? 3'b000 : 3'b100;
						assign node76 = (inp[8]) ? node78 : 3'b100;
							assign node78 = (inp[10]) ? node86 : node79;
								assign node79 = (inp[11]) ? 3'b100 : node80;
									assign node80 = (inp[2]) ? 3'b000 : node81;
										assign node81 = (inp[3]) ? 3'b100 : 3'b000;
								assign node86 = (inp[11]) ? node88 : 3'b000;
									assign node88 = (inp[3]) ? node90 : 3'b000;
										assign node90 = (inp[2]) ? 3'b000 : 3'b100;
				assign node93 = (inp[9]) ? node131 : node94;
					assign node94 = (inp[1]) ? node96 : 3'b100;
						assign node96 = (inp[8]) ? node114 : node97;
							assign node97 = (inp[11]) ? 3'b000 : node98;
								assign node98 = (inp[3]) ? node106 : node99;
									assign node99 = (inp[7]) ? node101 : 3'b100;
										assign node101 = (inp[10]) ? 3'b100 : node102;
											assign node102 = (inp[2]) ? 3'b100 : 3'b000;
									assign node106 = (inp[10]) ? node108 : 3'b000;
										assign node108 = (inp[2]) ? 3'b100 : node109;
											assign node109 = (inp[7]) ? 3'b000 : 3'b100;
							assign node114 = (inp[11]) ? node116 : 3'b100;
								assign node116 = (inp[3]) ? node124 : node117;
									assign node117 = (inp[2]) ? 3'b100 : node118;
										assign node118 = (inp[7]) ? node120 : 3'b100;
											assign node120 = (inp[5]) ? 3'b000 : 3'b100;
									assign node124 = (inp[10]) ? node126 : 3'b000;
										assign node126 = (inp[7]) ? node128 : 3'b100;
											assign node128 = (inp[2]) ? 3'b100 : 3'b000;
					assign node131 = (inp[8]) ? node173 : node132;
						assign node132 = (inp[10]) ? node156 : node133;
							assign node133 = (inp[1]) ? node143 : node134;
								assign node134 = (inp[2]) ? node138 : node135;
									assign node135 = (inp[11]) ? 3'b100 : 3'b001;
									assign node138 = (inp[3]) ? 3'b001 : node139;
										assign node139 = (inp[11]) ? 3'b001 : 3'b101;
								assign node143 = (inp[11]) ? node151 : node144;
									assign node144 = (inp[2]) ? 3'b100 : node145;
										assign node145 = (inp[7]) ? node147 : 3'b100;
											assign node147 = (inp[3]) ? 3'b000 : 3'b100;
									assign node151 = (inp[3]) ? 3'b000 : node152;
										assign node152 = (inp[2]) ? 3'b100 : 3'b000;
							assign node156 = (inp[11]) ? node164 : node157;
								assign node157 = (inp[2]) ? 3'b101 : node158;
									assign node158 = (inp[1]) ? 3'b001 : node159;
										assign node159 = (inp[3]) ? 3'b101 : 3'b001;
								assign node164 = (inp[2]) ? 3'b001 : node165;
									assign node165 = (inp[1]) ? 3'b100 : node166;
										assign node166 = (inp[7]) ? node168 : 3'b101;
											assign node168 = (inp[3]) ? 3'b001 : 3'b101;
						assign node173 = (inp[2]) ? node209 : node174;
							assign node174 = (inp[10]) ? node202 : node175;
								assign node175 = (inp[1]) ? node189 : node176;
									assign node176 = (inp[7]) ? node184 : node177;
										assign node177 = (inp[11]) ? node181 : node178;
											assign node178 = (inp[3]) ? 3'b100 : 3'b000;
											assign node181 = (inp[3]) ? 3'b000 : 3'b100;
										assign node184 = (inp[3]) ? node186 : 3'b000;
											assign node186 = (inp[11]) ? 3'b000 : 3'b100;
									assign node189 = (inp[7]) ? node195 : node190;
										assign node190 = (inp[11]) ? node192 : 3'b101;
											assign node192 = (inp[3]) ? 3'b101 : 3'b001;
										assign node195 = (inp[11]) ? node199 : node196;
											assign node196 = (inp[3]) ? 3'b001 : 3'b101;
											assign node199 = (inp[3]) ? 3'b101 : 3'b001;
								assign node202 = (inp[11]) ? node206 : node203;
									assign node203 = (inp[7]) ? 3'b011 : 3'b111;
									assign node206 = (inp[7]) ? 3'b010 : 3'b110;
							assign node209 = (inp[10]) ? 3'b000 : node210;
								assign node210 = (inp[1]) ? node214 : node211;
									assign node211 = (inp[3]) ? 3'b001 : 3'b101;
									assign node214 = (inp[3]) ? 3'b000 : 3'b100;
			assign node218 = (inp[9]) ? node220 : 3'b000;
				assign node220 = (inp[1]) ? node298 : node221;
					assign node221 = (inp[8]) ? node255 : node222;
						assign node222 = (inp[11]) ? node246 : node223;
							assign node223 = (inp[10]) ? node237 : node224;
								assign node224 = (inp[3]) ? node232 : node225;
									assign node225 = (inp[4]) ? 3'b000 : node226;
										assign node226 = (inp[7]) ? node228 : 3'b100;
											assign node228 = (inp[2]) ? 3'b100 : 3'b000;
									assign node232 = (inp[4]) ? node234 : 3'b000;
										assign node234 = (inp[2]) ? 3'b000 : 3'b100;
								assign node237 = (inp[2]) ? 3'b100 : node238;
									assign node238 = (inp[4]) ? node240 : 3'b100;
										assign node240 = (inp[7]) ? 3'b000 : node241;
											assign node241 = (inp[3]) ? 3'b000 : 3'b100;
							assign node246 = (inp[4]) ? node248 : 3'b000;
								assign node248 = (inp[10]) ? node250 : 3'b100;
									assign node250 = (inp[3]) ? node252 : 3'b000;
										assign node252 = (inp[2]) ? 3'b000 : 3'b100;
						assign node255 = (inp[4]) ? node273 : node256;
							assign node256 = (inp[11]) ? node258 : 3'b100;
								assign node258 = (inp[3]) ? node266 : node259;
									assign node259 = (inp[7]) ? node261 : 3'b100;
										assign node261 = (inp[10]) ? 3'b100 : node262;
											assign node262 = (inp[2]) ? 3'b100 : 3'b000;
									assign node266 = (inp[10]) ? node268 : 3'b000;
										assign node268 = (inp[2]) ? 3'b100 : node269;
											assign node269 = (inp[7]) ? 3'b000 : 3'b100;
							assign node273 = (inp[10]) ? node289 : node274;
								assign node274 = (inp[3]) ? node282 : node275;
									assign node275 = (inp[2]) ? 3'b101 : node276;
										assign node276 = (inp[11]) ? 3'b100 : node277;
											assign node277 = (inp[7]) ? 3'b001 : 3'b101;
									assign node282 = (inp[11]) ? node284 : 3'b001;
										assign node284 = (inp[2]) ? 3'b001 : node285;
											assign node285 = (inp[7]) ? 3'b000 : 3'b100;
								assign node289 = (inp[2]) ? 3'b000 : node290;
									assign node290 = (inp[11]) ? node294 : node291;
										assign node291 = (inp[7]) ? 3'b001 : 3'b101;
										assign node294 = (inp[7]) ? 3'b000 : 3'b100;
					assign node298 = (inp[4]) ? node300 : 3'b000;
						assign node300 = (inp[11]) ? node330 : node301;
							assign node301 = (inp[8]) ? node317 : node302;
								assign node302 = (inp[10]) ? node310 : node303;
									assign node303 = (inp[3]) ? 3'b000 : node304;
										assign node304 = (inp[2]) ? 3'b100 : node305;
											assign node305 = (inp[7]) ? 3'b000 : 3'b100;
									assign node310 = (inp[3]) ? node312 : 3'b100;
										assign node312 = (inp[2]) ? 3'b100 : node313;
											assign node313 = (inp[7]) ? 3'b000 : 3'b100;
								assign node317 = (inp[10]) ? node325 : node318;
									assign node318 = (inp[2]) ? node322 : node319;
										assign node319 = (inp[3]) ? 3'b100 : 3'b000;
										assign node322 = (inp[3]) ? 3'b000 : 3'b100;
									assign node325 = (inp[2]) ? 3'b000 : node326;
										assign node326 = (inp[7]) ? 3'b001 : 3'b101;
							assign node330 = (inp[8]) ? node332 : 3'b000;
								assign node332 = (inp[7]) ? node344 : node333;
									assign node333 = (inp[2]) ? node339 : node334;
										assign node334 = (inp[10]) ? 3'b100 : node335;
											assign node335 = (inp[3]) ? 3'b000 : 3'b100;
										assign node339 = (inp[3]) ? 3'b000 : node340;
											assign node340 = (inp[10]) ? 3'b000 : 3'b100;
									assign node344 = (inp[10]) ? 3'b000 : node345;
										assign node345 = (inp[3]) ? 3'b000 : node346;
											assign node346 = (inp[2]) ? 3'b100 : 3'b000;

endmodule