module dtc_split875_bm98 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node35;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node162;
	wire [3-1:0] node164;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node181;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node205;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node264;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node273;
	wire [3-1:0] node275;
	wire [3-1:0] node278;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node284;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node292;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node317;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node323;
	wire [3-1:0] node325;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node340;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node356;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node363;
	wire [3-1:0] node366;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node382;
	wire [3-1:0] node385;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node390;
	wire [3-1:0] node392;
	wire [3-1:0] node395;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node401;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node426;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node433;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node439;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node446;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node457;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node466;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node473;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node480;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node499;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node514;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node523;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node529;
	wire [3-1:0] node531;
	wire [3-1:0] node534;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node540;
	wire [3-1:0] node543;
	wire [3-1:0] node545;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node552;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node569;
	wire [3-1:0] node572;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node578;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node601;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node607;
	wire [3-1:0] node609;
	wire [3-1:0] node612;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node618;
	wire [3-1:0] node621;
	wire [3-1:0] node624;
	wire [3-1:0] node626;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node632;
	wire [3-1:0] node635;
	wire [3-1:0] node637;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node643;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node661;
	wire [3-1:0] node664;
	wire [3-1:0] node666;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node672;
	wire [3-1:0] node675;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node681;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node692;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node707;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node718;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node734;
	wire [3-1:0] node736;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node743;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node753;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node763;
	wire [3-1:0] node764;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node771;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node778;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node785;
	wire [3-1:0] node787;
	wire [3-1:0] node790;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node797;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node804;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node812;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node819;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node828;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node840;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node847;
	wire [3-1:0] node850;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node869;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node876;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node882;
	wire [3-1:0] node884;
	wire [3-1:0] node887;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node893;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node902;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node915;
	wire [3-1:0] node918;
	wire [3-1:0] node919;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node929;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node936;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node944;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node951;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node957;
	wire [3-1:0] node959;
	wire [3-1:0] node962;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node968;

	assign outp = (inp[0]) ? node404 : node1;
		assign node1 = (inp[6]) ? node3 : 3'b111;
			assign node3 = (inp[9]) ? node119 : node4;
				assign node4 = (inp[3]) ? node88 : node5;
					assign node5 = (inp[4]) ? node7 : 3'b100;
						assign node7 = (inp[1]) ? node45 : node8;
							assign node8 = (inp[7]) ? node10 : 3'b100;
								assign node10 = (inp[2]) ? node32 : node11;
									assign node11 = (inp[10]) ? node17 : node12;
										assign node12 = (inp[11]) ? node14 : 3'b000;
											assign node14 = (inp[5]) ? 3'b100 : 3'b000;
										assign node17 = (inp[8]) ? node25 : node18;
											assign node18 = (inp[5]) ? node22 : node19;
												assign node19 = (inp[11]) ? 3'b100 : 3'b000;
												assign node22 = (inp[11]) ? 3'b000 : 3'b100;
											assign node25 = (inp[11]) ? node29 : node26;
												assign node26 = (inp[5]) ? 3'b100 : 3'b000;
												assign node29 = (inp[5]) ? 3'b000 : 3'b100;
									assign node32 = (inp[5]) ? node38 : node33;
										assign node33 = (inp[11]) ? node35 : 3'b100;
											assign node35 = (inp[10]) ? 3'b000 : 3'b100;
										assign node38 = (inp[11]) ? node42 : node39;
											assign node39 = (inp[10]) ? 3'b000 : 3'b100;
											assign node42 = (inp[10]) ? 3'b100 : 3'b000;
							assign node45 = (inp[7]) ? node47 : 3'b000;
								assign node47 = (inp[2]) ? node67 : node48;
									assign node48 = (inp[10]) ? node54 : node49;
										assign node49 = (inp[5]) ? node51 : 3'b101;
											assign node51 = (inp[11]) ? 3'b100 : 3'b101;
										assign node54 = (inp[8]) ? node62 : node55;
											assign node55 = (inp[11]) ? node59 : node56;
												assign node56 = (inp[5]) ? 3'b100 : 3'b101;
												assign node59 = (inp[5]) ? 3'b101 : 3'b100;
											assign node62 = (inp[11]) ? node64 : 3'b100;
												assign node64 = (inp[5]) ? 3'b101 : 3'b100;
									assign node67 = (inp[5]) ? node73 : node68;
										assign node68 = (inp[10]) ? node70 : 3'b100;
											assign node70 = (inp[11]) ? 3'b101 : 3'b100;
										assign node73 = (inp[8]) ? node81 : node74;
											assign node74 = (inp[10]) ? node78 : node75;
												assign node75 = (inp[11]) ? 3'b101 : 3'b100;
												assign node78 = (inp[11]) ? 3'b100 : 3'b101;
											assign node81 = (inp[11]) ? node85 : node82;
												assign node82 = (inp[10]) ? 3'b101 : 3'b100;
												assign node85 = (inp[10]) ? 3'b100 : 3'b101;
					assign node88 = (inp[4]) ? node90 : 3'b010;
						assign node90 = (inp[7]) ? node92 : 3'b010;
							assign node92 = (inp[1]) ? node94 : 3'b010;
								assign node94 = (inp[2]) ? node106 : node95;
									assign node95 = (inp[11]) ? node101 : node96;
										assign node96 = (inp[8]) ? node98 : 3'b110;
											assign node98 = (inp[10]) ? 3'b010 : 3'b110;
										assign node101 = (inp[5]) ? 3'b010 : node102;
											assign node102 = (inp[10]) ? 3'b010 : 3'b110;
									assign node106 = (inp[10]) ? node112 : node107;
										assign node107 = (inp[5]) ? node109 : 3'b010;
											assign node109 = (inp[11]) ? 3'b110 : 3'b010;
										assign node112 = (inp[11]) ? node116 : node113;
											assign node113 = (inp[5]) ? 3'b110 : 3'b010;
											assign node116 = (inp[5]) ? 3'b010 : 3'b110;
				assign node119 = (inp[3]) ? node331 : node120;
					assign node120 = (inp[1]) ? node232 : node121;
						assign node121 = (inp[4]) ? node157 : node122;
							assign node122 = (inp[2]) ? node132 : node123;
								assign node123 = (inp[7]) ? 3'b001 : node124;
									assign node124 = (inp[11]) ? node128 : node125;
										assign node125 = (inp[5]) ? 3'b101 : 3'b001;
										assign node128 = (inp[5]) ? 3'b001 : 3'b101;
								assign node132 = (inp[7]) ? 3'b101 : node133;
									assign node133 = (inp[8]) ? node149 : node134;
										assign node134 = (inp[10]) ? node142 : node135;
											assign node135 = (inp[5]) ? node139 : node136;
												assign node136 = (inp[11]) ? 3'b101 : 3'b001;
												assign node139 = (inp[11]) ? 3'b001 : 3'b101;
											assign node142 = (inp[5]) ? node146 : node143;
												assign node143 = (inp[11]) ? 3'b101 : 3'b001;
												assign node146 = (inp[11]) ? 3'b001 : 3'b101;
										assign node149 = (inp[5]) ? node153 : node150;
											assign node150 = (inp[11]) ? 3'b101 : 3'b001;
											assign node153 = (inp[11]) ? 3'b001 : 3'b101;
							assign node157 = (inp[2]) ? node197 : node158;
								assign node158 = (inp[7]) ? node176 : node159;
									assign node159 = (inp[5]) ? node167 : node160;
										assign node160 = (inp[10]) ? node162 : 3'b101;
											assign node162 = (inp[8]) ? node164 : 3'b101;
												assign node164 = (inp[11]) ? 3'b111 : 3'b101;
										assign node167 = (inp[8]) ? node169 : 3'b111;
											assign node169 = (inp[11]) ? node173 : node170;
												assign node170 = (inp[10]) ? 3'b111 : 3'b101;
												assign node173 = (inp[10]) ? 3'b101 : 3'b111;
									assign node176 = (inp[10]) ? node184 : node177;
										assign node177 = (inp[5]) ? node181 : node178;
											assign node178 = (inp[11]) ? 3'b111 : 3'b011;
											assign node181 = (inp[11]) ? 3'b011 : 3'b111;
										assign node184 = (inp[8]) ? node192 : node185;
											assign node185 = (inp[11]) ? node189 : node186;
												assign node186 = (inp[5]) ? 3'b111 : 3'b011;
												assign node189 = (inp[5]) ? 3'b011 : 3'b111;
											assign node192 = (inp[5]) ? 3'b011 : node193;
												assign node193 = (inp[11]) ? 3'b111 : 3'b011;
								assign node197 = (inp[7]) ? node219 : node198;
									assign node198 = (inp[11]) ? node208 : node199;
										assign node199 = (inp[8]) ? node203 : node200;
											assign node200 = (inp[10]) ? 3'b101 : 3'b001;
											assign node203 = (inp[10]) ? node205 : 3'b111;
												assign node205 = (inp[5]) ? 3'b001 : 3'b011;
										assign node208 = (inp[8]) ? node212 : node209;
											assign node209 = (inp[10]) ? 3'b111 : 3'b011;
											assign node212 = (inp[10]) ? node216 : node213;
												assign node213 = (inp[5]) ? 3'b101 : 3'b111;
												assign node216 = (inp[5]) ? 3'b011 : 3'b001;
									assign node219 = (inp[11]) ? node223 : node220;
										assign node220 = (inp[8]) ? 3'b101 : 3'b001;
										assign node223 = (inp[8]) ? node225 : 3'b101;
											assign node225 = (inp[10]) ? node229 : node226;
												assign node226 = (inp[5]) ? 3'b001 : 3'b101;
												assign node229 = (inp[5]) ? 3'b101 : 3'b001;
						assign node232 = (inp[4]) ? node268 : node233;
							assign node233 = (inp[2]) ? node243 : node234;
								assign node234 = (inp[7]) ? 3'b001 : node235;
									assign node235 = (inp[11]) ? node239 : node236;
										assign node236 = (inp[5]) ? 3'b100 : 3'b001;
										assign node239 = (inp[5]) ? 3'b001 : 3'b100;
								assign node243 = (inp[7]) ? 3'b100 : node244;
									assign node244 = (inp[8]) ? node254 : node245;
										assign node245 = (inp[10]) ? 3'b100 : node246;
											assign node246 = (inp[11]) ? node250 : node247;
												assign node247 = (inp[5]) ? 3'b100 : 3'b001;
												assign node250 = (inp[5]) ? 3'b001 : 3'b100;
										assign node254 = (inp[10]) ? node262 : node255;
											assign node255 = (inp[5]) ? node259 : node256;
												assign node256 = (inp[11]) ? 3'b100 : 3'b001;
												assign node259 = (inp[11]) ? 3'b001 : 3'b100;
											assign node262 = (inp[11]) ? node264 : 3'b001;
												assign node264 = (inp[5]) ? 3'b001 : 3'b100;
							assign node268 = (inp[7]) ? node304 : node269;
								assign node269 = (inp[2]) ? node287 : node270;
									assign node270 = (inp[11]) ? node278 : node271;
										assign node271 = (inp[8]) ? node273 : 3'b110;
											assign node273 = (inp[5]) ? node275 : 3'b100;
												assign node275 = (inp[10]) ? 3'b110 : 3'b100;
										assign node278 = (inp[8]) ? node280 : 3'b100;
											assign node280 = (inp[5]) ? node284 : node281;
												assign node281 = (inp[10]) ? 3'b110 : 3'b100;
												assign node284 = (inp[10]) ? 3'b100 : 3'b110;
									assign node287 = (inp[8]) ? node295 : node288;
										assign node288 = (inp[10]) ? node292 : node289;
											assign node289 = (inp[11]) ? 3'b011 : 3'b001;
											assign node292 = (inp[11]) ? 3'b110 : 3'b100;
										assign node295 = (inp[10]) ? node301 : node296;
											assign node296 = (inp[11]) ? node298 : 3'b110;
												assign node298 = (inp[5]) ? 3'b100 : 3'b110;
											assign node301 = (inp[11]) ? 3'b001 : 3'b011;
								assign node304 = (inp[11]) ? node320 : node305;
									assign node305 = (inp[8]) ? node311 : node306;
										assign node306 = (inp[5]) ? node308 : 3'b001;
											assign node308 = (inp[2]) ? 3'b001 : 3'b110;
										assign node311 = (inp[2]) ? node315 : node312;
											assign node312 = (inp[5]) ? 3'b110 : 3'b001;
											assign node315 = (inp[5]) ? node317 : 3'b110;
												assign node317 = (inp[10]) ? 3'b001 : 3'b110;
									assign node320 = (inp[5]) ? node328 : node321;
										assign node321 = (inp[2]) ? node323 : 3'b110;
											assign node323 = (inp[10]) ? node325 : 3'b110;
												assign node325 = (inp[8]) ? 3'b001 : 3'b110;
										assign node328 = (inp[2]) ? 3'b110 : 3'b001;
					assign node331 = (inp[1]) ? node333 : 3'b111;
						assign node333 = (inp[7]) ? node375 : node334;
							assign node334 = (inp[4]) ? node366 : node335;
								assign node335 = (inp[10]) ? node343 : node336;
									assign node336 = (inp[5]) ? node340 : node337;
										assign node337 = (inp[11]) ? 3'b011 : 3'b111;
										assign node340 = (inp[11]) ? 3'b111 : 3'b011;
									assign node343 = (inp[2]) ? node359 : node344;
										assign node344 = (inp[8]) ? node352 : node345;
											assign node345 = (inp[11]) ? node349 : node346;
												assign node346 = (inp[5]) ? 3'b011 : 3'b111;
												assign node349 = (inp[5]) ? 3'b111 : 3'b011;
											assign node352 = (inp[5]) ? node356 : node353;
												assign node353 = (inp[11]) ? 3'b011 : 3'b111;
												assign node356 = (inp[11]) ? 3'b111 : 3'b011;
										assign node359 = (inp[5]) ? node363 : node360;
											assign node360 = (inp[11]) ? 3'b011 : 3'b111;
											assign node363 = (inp[11]) ? 3'b111 : 3'b011;
								assign node366 = (inp[2]) ? node368 : 3'b001;
									assign node368 = (inp[8]) ? node372 : node369;
										assign node369 = (inp[10]) ? 3'b001 : 3'b111;
										assign node372 = (inp[10]) ? 3'b111 : 3'b011;
							assign node375 = (inp[2]) ? node385 : node376;
								assign node376 = (inp[4]) ? node378 : 3'b101;
									assign node378 = (inp[5]) ? node382 : node379;
										assign node379 = (inp[11]) ? 3'b011 : 3'b111;
										assign node382 = (inp[11]) ? 3'b111 : 3'b011;
								assign node385 = (inp[4]) ? node387 : 3'b001;
									assign node387 = (inp[11]) ? node395 : node388;
										assign node388 = (inp[8]) ? node390 : 3'b101;
											assign node390 = (inp[10]) ? node392 : 3'b001;
												assign node392 = (inp[5]) ? 3'b101 : 3'b001;
										assign node395 = (inp[8]) ? node397 : 3'b011;
											assign node397 = (inp[10]) ? node401 : node398;
												assign node398 = (inp[5]) ? 3'b101 : 3'b001;
												assign node401 = (inp[5]) ? 3'b011 : 3'b101;
		assign node404 = (inp[3]) ? node584 : node405;
			assign node405 = (inp[6]) ? node543 : node406;
				assign node406 = (inp[9]) ? node450 : node407;
					assign node407 = (inp[4]) ? node409 : 3'b010;
						assign node409 = (inp[7]) ? node413 : node410;
							assign node410 = (inp[1]) ? 3'b000 : 3'b010;
							assign node413 = (inp[1]) ? 3'b010 : node414;
								assign node414 = (inp[2]) ? node436 : node415;
									assign node415 = (inp[11]) ? node421 : node416;
										assign node416 = (inp[10]) ? node418 : 3'b000;
											assign node418 = (inp[5]) ? 3'b010 : 3'b000;
										assign node421 = (inp[8]) ? node429 : node422;
											assign node422 = (inp[10]) ? node426 : node423;
												assign node423 = (inp[5]) ? 3'b010 : 3'b000;
												assign node426 = (inp[5]) ? 3'b000 : 3'b010;
											assign node429 = (inp[10]) ? node433 : node430;
												assign node430 = (inp[5]) ? 3'b010 : 3'b000;
												assign node433 = (inp[5]) ? 3'b000 : 3'b010;
									assign node436 = (inp[11]) ? node442 : node437;
										assign node437 = (inp[10]) ? node439 : 3'b010;
											assign node439 = (inp[5]) ? 3'b000 : 3'b010;
										assign node442 = (inp[5]) ? node446 : node443;
											assign node443 = (inp[10]) ? 3'b000 : 3'b010;
											assign node446 = (inp[10]) ? 3'b010 : 3'b000;
					assign node450 = (inp[4]) ? node484 : node451;
						assign node451 = (inp[2]) ? node461 : node452;
							assign node452 = (inp[7]) ? 3'b000 : node453;
								assign node453 = (inp[11]) ? node457 : node454;
									assign node454 = (inp[5]) ? 3'b010 : 3'b000;
									assign node457 = (inp[5]) ? 3'b000 : 3'b010;
							assign node461 = (inp[7]) ? 3'b010 : node462;
								assign node462 = (inp[10]) ? node476 : node463;
									assign node463 = (inp[8]) ? node469 : node464;
										assign node464 = (inp[5]) ? node466 : 3'b010;
											assign node466 = (inp[11]) ? 3'b000 : 3'b010;
										assign node469 = (inp[5]) ? node473 : node470;
											assign node470 = (inp[11]) ? 3'b010 : 3'b000;
											assign node473 = (inp[11]) ? 3'b000 : 3'b010;
									assign node476 = (inp[5]) ? node480 : node477;
										assign node477 = (inp[11]) ? 3'b010 : 3'b000;
										assign node480 = (inp[11]) ? 3'b000 : 3'b010;
						assign node484 = (inp[2]) ? node494 : node485;
							assign node485 = (inp[7]) ? node487 : 3'b010;
								assign node487 = (inp[5]) ? node491 : node488;
									assign node488 = (inp[11]) ? 3'b010 : 3'b000;
									assign node491 = (inp[11]) ? 3'b000 : 3'b010;
							assign node494 = (inp[7]) ? node502 : node495;
								assign node495 = (inp[8]) ? node499 : node496;
									assign node496 = (inp[10]) ? 3'b010 : 3'b000;
									assign node499 = (inp[10]) ? 3'b000 : 3'b010;
								assign node502 = (inp[1]) ? node526 : node503;
									assign node503 = (inp[5]) ? node517 : node504;
										assign node504 = (inp[10]) ? node510 : node505;
											assign node505 = (inp[8]) ? 3'b010 : node506;
												assign node506 = (inp[11]) ? 3'b010 : 3'b000;
											assign node510 = (inp[11]) ? node514 : node511;
												assign node511 = (inp[8]) ? 3'b010 : 3'b000;
												assign node514 = (inp[8]) ? 3'b000 : 3'b010;
										assign node517 = (inp[11]) ? node523 : node518;
											assign node518 = (inp[10]) ? 3'b000 : node519;
												assign node519 = (inp[8]) ? 3'b010 : 3'b000;
											assign node523 = (inp[8]) ? 3'b000 : 3'b010;
									assign node526 = (inp[11]) ? node534 : node527;
										assign node527 = (inp[8]) ? node529 : 3'b100;
											assign node529 = (inp[5]) ? node531 : 3'b010;
												assign node531 = (inp[10]) ? 3'b100 : 3'b110;
										assign node534 = (inp[8]) ? node536 : 3'b110;
											assign node536 = (inp[5]) ? node540 : node537;
												assign node537 = (inp[10]) ? 3'b100 : 3'b110;
												assign node540 = (inp[10]) ? 3'b010 : 3'b000;
				assign node543 = (inp[4]) ? node545 : 3'b000;
					assign node545 = (inp[9]) ? node547 : 3'b000;
						assign node547 = (inp[1]) ? node581 : node548;
							assign node548 = (inp[11]) ? node564 : node549;
								assign node549 = (inp[5]) ? node555 : node550;
									assign node550 = (inp[8]) ? node552 : 3'b010;
										assign node552 = (inp[2]) ? 3'b110 : 3'b010;
									assign node555 = (inp[2]) ? node559 : node556;
										assign node556 = (inp[10]) ? 3'b100 : 3'b110;
										assign node559 = (inp[10]) ? 3'b010 : node560;
											assign node560 = (inp[8]) ? 3'b110 : 3'b010;
								assign node564 = (inp[2]) ? node572 : node565;
									assign node565 = (inp[5]) ? node569 : node566;
										assign node566 = (inp[10]) ? 3'b100 : 3'b110;
										assign node569 = (inp[10]) ? 3'b010 : 3'b000;
									assign node572 = (inp[8]) ? node574 : 3'b100;
										assign node574 = (inp[5]) ? node578 : node575;
											assign node575 = (inp[10]) ? 3'b000 : 3'b100;
											assign node578 = (inp[10]) ? 3'b100 : 3'b000;
							assign node581 = (inp[7]) ? 3'b000 : 3'b100;
			assign node584 = (inp[9]) ? node722 : node585;
				assign node585 = (inp[1]) ? node653 : node586;
					assign node586 = (inp[6]) ? node624 : node587;
						assign node587 = (inp[4]) ? node589 : 3'b001;
							assign node589 = (inp[7]) ? node621 : node590;
								assign node590 = (inp[2]) ? node604 : node591;
									assign node591 = (inp[11]) ? node595 : node592;
										assign node592 = (inp[8]) ? 3'b011 : 3'b111;
										assign node595 = (inp[8]) ? node597 : 3'b011;
											assign node597 = (inp[10]) ? node601 : node598;
												assign node598 = (inp[5]) ? 3'b111 : 3'b011;
												assign node601 = (inp[5]) ? 3'b011 : 3'b111;
									assign node604 = (inp[11]) ? node612 : node605;
										assign node605 = (inp[8]) ? node607 : 3'b011;
											assign node607 = (inp[10]) ? node609 : 3'b101;
												assign node609 = (inp[5]) ? 3'b011 : 3'b101;
										assign node612 = (inp[8]) ? node614 : 3'b101;
											assign node614 = (inp[10]) ? node618 : node615;
												assign node615 = (inp[5]) ? 3'b011 : 3'b101;
												assign node618 = (inp[5]) ? 3'b101 : 3'b011;
								assign node621 = (inp[2]) ? 3'b001 : 3'b101;
						assign node624 = (inp[4]) ? node626 : 3'b000;
							assign node626 = (inp[7]) ? node628 : 3'b001;
								assign node628 = (inp[11]) ? node640 : node629;
									assign node629 = (inp[2]) ? node635 : node630;
										assign node630 = (inp[10]) ? node632 : 3'b100;
											assign node632 = (inp[5]) ? 3'b010 : 3'b100;
										assign node635 = (inp[10]) ? node637 : 3'b000;
											assign node637 = (inp[5]) ? 3'b100 : 3'b000;
									assign node640 = (inp[2]) ? node646 : node641;
										assign node641 = (inp[10]) ? node643 : 3'b100;
											assign node643 = (inp[8]) ? 3'b010 : 3'b100;
										assign node646 = (inp[10]) ? node650 : node647;
											assign node647 = (inp[5]) ? 3'b110 : 3'b010;
											assign node650 = (inp[5]) ? 3'b010 : 3'b110;
					assign node653 = (inp[4]) ? node655 : 3'b000;
						assign node655 = (inp[7]) ? node685 : node656;
							assign node656 = (inp[6]) ? 3'b100 : node657;
								assign node657 = (inp[2]) ? node669 : node658;
									assign node658 = (inp[11]) ? node664 : node659;
										assign node659 = (inp[8]) ? node661 : 3'b101;
											assign node661 = (inp[5]) ? 3'b101 : 3'b001;
										assign node664 = (inp[8]) ? node666 : 3'b001;
											assign node666 = (inp[10]) ? 3'b001 : 3'b101;
									assign node669 = (inp[11]) ? node675 : node670;
										assign node670 = (inp[8]) ? node672 : 3'b001;
											assign node672 = (inp[10]) ? 3'b001 : 3'b110;
										assign node675 = (inp[8]) ? node677 : 3'b110;
											assign node677 = (inp[10]) ? node681 : node678;
												assign node678 = (inp[5]) ? 3'b001 : 3'b110;
												assign node681 = (inp[5]) ? 3'b110 : 3'b001;
							assign node685 = (inp[6]) ? 3'b000 : node686;
								assign node686 = (inp[2]) ? node704 : node687;
									assign node687 = (inp[10]) ? node697 : node688;
										assign node688 = (inp[8]) ? node692 : node689;
											assign node689 = (inp[11]) ? 3'b110 : 3'b010;
											assign node692 = (inp[5]) ? node694 : 3'b010;
												assign node694 = (inp[11]) ? 3'b010 : 3'b110;
										assign node697 = (inp[5]) ? node701 : node698;
											assign node698 = (inp[11]) ? 3'b110 : 3'b010;
											assign node701 = (inp[11]) ? 3'b010 : 3'b110;
									assign node704 = (inp[11]) ? node712 : node705;
										assign node705 = (inp[8]) ? node707 : 3'b010;
											assign node707 = (inp[10]) ? node709 : 3'b100;
												assign node709 = (inp[5]) ? 3'b010 : 3'b100;
										assign node712 = (inp[8]) ? node714 : 3'b100;
											assign node714 = (inp[5]) ? node718 : node715;
												assign node715 = (inp[10]) ? 3'b010 : 3'b100;
												assign node718 = (inp[10]) ? 3'b100 : 3'b010;
				assign node722 = (inp[6]) ? node832 : node723;
					assign node723 = (inp[1]) ? node725 : 3'b111;
						assign node725 = (inp[4]) ? node781 : node726;
							assign node726 = (inp[11]) ? node756 : node727;
								assign node727 = (inp[8]) ? node739 : node728;
									assign node728 = (inp[2]) ? node734 : node729;
										assign node729 = (inp[5]) ? 3'b010 : node730;
											assign node730 = (inp[7]) ? 3'b110 : 3'b010;
										assign node734 = (inp[10]) ? node736 : 3'b110;
											assign node736 = (inp[7]) ? 3'b110 : 3'b010;
									assign node739 = (inp[10]) ? node747 : node740;
										assign node740 = (inp[2]) ? 3'b001 : node741;
											assign node741 = (inp[7]) ? node743 : 3'b001;
												assign node743 = (inp[5]) ? 3'b001 : 3'b101;
										assign node747 = (inp[5]) ? node753 : node748;
											assign node748 = (inp[2]) ? 3'b001 : node749;
												assign node749 = (inp[7]) ? 3'b101 : 3'b001;
											assign node753 = (inp[2]) ? 3'b110 : 3'b010;
								assign node756 = (inp[8]) ? node768 : node757;
									assign node757 = (inp[5]) ? node759 : 3'b001;
										assign node759 = (inp[2]) ? node763 : node760;
											assign node760 = (inp[7]) ? 3'b101 : 3'b001;
											assign node763 = (inp[10]) ? 3'b001 : node764;
												assign node764 = (inp[7]) ? 3'b001 : 3'b101;
									assign node768 = (inp[10]) ? node774 : node769;
										assign node769 = (inp[5]) ? node771 : 3'b001;
											assign node771 = (inp[7]) ? 3'b110 : 3'b010;
										assign node774 = (inp[5]) ? node778 : node775;
											assign node775 = (inp[2]) ? 3'b110 : 3'b010;
											assign node778 = (inp[2]) ? 3'b001 : 3'b101;
							assign node781 = (inp[7]) ? node807 : node782;
								assign node782 = (inp[11]) ? node790 : node783;
									assign node783 = (inp[8]) ? node785 : 3'b011;
										assign node785 = (inp[5]) ? node787 : 3'b111;
											assign node787 = (inp[10]) ? 3'b011 : 3'b111;
									assign node790 = (inp[8]) ? node792 : 3'b111;
										assign node792 = (inp[2]) ? node800 : node793;
											assign node793 = (inp[10]) ? node797 : node794;
												assign node794 = (inp[5]) ? 3'b011 : 3'b111;
												assign node797 = (inp[5]) ? 3'b111 : 3'b011;
											assign node800 = (inp[10]) ? node804 : node801;
												assign node801 = (inp[5]) ? 3'b011 : 3'b111;
												assign node804 = (inp[5]) ? 3'b111 : 3'b011;
								assign node807 = (inp[2]) ? node823 : node808;
									assign node808 = (inp[8]) ? 3'b001 : node809;
										assign node809 = (inp[10]) ? node815 : node810;
											assign node810 = (inp[5]) ? node812 : 3'b011;
												assign node812 = (inp[11]) ? 3'b011 : 3'b001;
											assign node815 = (inp[5]) ? node819 : node816;
												assign node816 = (inp[11]) ? 3'b001 : 3'b011;
												assign node819 = (inp[11]) ? 3'b011 : 3'b001;
									assign node823 = (inp[8]) ? 3'b101 : node824;
										assign node824 = (inp[5]) ? node828 : node825;
											assign node825 = (inp[11]) ? 3'b101 : 3'b011;
											assign node828 = (inp[11]) ? 3'b011 : 3'b101;
					assign node832 = (inp[1]) ? node896 : node833;
						assign node833 = (inp[7]) ? node859 : node834;
							assign node834 = (inp[4]) ? node850 : node835;
								assign node835 = (inp[2]) ? node843 : node836;
									assign node836 = (inp[11]) ? node840 : node837;
										assign node837 = (inp[5]) ? 3'b001 : 3'b101;
										assign node840 = (inp[5]) ? 3'b101 : 3'b001;
									assign node843 = (inp[5]) ? node847 : node844;
										assign node844 = (inp[11]) ? 3'b001 : 3'b101;
										assign node847 = (inp[11]) ? 3'b101 : 3'b001;
								assign node850 = (inp[2]) ? node852 : 3'b010;
									assign node852 = (inp[10]) ? node856 : node853;
										assign node853 = (inp[8]) ? 3'b001 : 3'b101;
										assign node856 = (inp[8]) ? 3'b101 : 3'b010;
							assign node859 = (inp[4]) ? node863 : node860;
								assign node860 = (inp[2]) ? 3'b010 : 3'b110;
								assign node863 = (inp[2]) ? node879 : node864;
									assign node864 = (inp[8]) ? node872 : node865;
										assign node865 = (inp[11]) ? node869 : node866;
											assign node866 = (inp[5]) ? 3'b001 : 3'b101;
											assign node869 = (inp[5]) ? 3'b101 : 3'b001;
										assign node872 = (inp[11]) ? node876 : node873;
											assign node873 = (inp[5]) ? 3'b001 : 3'b101;
											assign node876 = (inp[5]) ? 3'b101 : 3'b001;
									assign node879 = (inp[11]) ? node887 : node880;
										assign node880 = (inp[8]) ? node882 : 3'b110;
											assign node882 = (inp[5]) ? node884 : 3'b010;
												assign node884 = (inp[10]) ? 3'b110 : 3'b010;
										assign node887 = (inp[8]) ? node889 : 3'b001;
											assign node889 = (inp[10]) ? node893 : node890;
												assign node890 = (inp[5]) ? 3'b110 : 3'b010;
												assign node893 = (inp[5]) ? 3'b001 : 3'b110;
						assign node896 = (inp[7]) ? node918 : node897;
							assign node897 = (inp[4]) ? node905 : node898;
								assign node898 = (inp[11]) ? node902 : node899;
									assign node899 = (inp[5]) ? 3'b010 : 3'b110;
									assign node902 = (inp[5]) ? 3'b110 : 3'b010;
								assign node905 = (inp[2]) ? node911 : node906;
									assign node906 = (inp[8]) ? 3'b000 : node907;
										assign node907 = (inp[10]) ? 3'b001 : 3'b000;
									assign node911 = (inp[10]) ? node915 : node912;
										assign node912 = (inp[8]) ? 3'b010 : 3'b110;
										assign node915 = (inp[8]) ? 3'b110 : 3'b001;
							assign node918 = (inp[4]) ? node922 : node919;
								assign node919 = (inp[2]) ? 3'b000 : 3'b100;
								assign node922 = (inp[2]) ? node954 : node923;
									assign node923 = (inp[10]) ? node939 : node924;
										assign node924 = (inp[8]) ? node932 : node925;
											assign node925 = (inp[5]) ? node929 : node926;
												assign node926 = (inp[11]) ? 3'b010 : 3'b110;
												assign node929 = (inp[11]) ? 3'b110 : 3'b010;
											assign node932 = (inp[11]) ? node936 : node933;
												assign node933 = (inp[5]) ? 3'b010 : 3'b110;
												assign node936 = (inp[5]) ? 3'b110 : 3'b010;
										assign node939 = (inp[8]) ? node947 : node940;
											assign node940 = (inp[11]) ? node944 : node941;
												assign node941 = (inp[5]) ? 3'b010 : 3'b110;
												assign node944 = (inp[5]) ? 3'b110 : 3'b010;
											assign node947 = (inp[11]) ? node951 : node948;
												assign node948 = (inp[5]) ? 3'b010 : 3'b110;
												assign node951 = (inp[5]) ? 3'b110 : 3'b010;
									assign node954 = (inp[11]) ? node962 : node955;
										assign node955 = (inp[8]) ? node957 : 3'b100;
											assign node957 = (inp[5]) ? node959 : 3'b000;
												assign node959 = (inp[10]) ? 3'b100 : 3'b000;
										assign node962 = (inp[8]) ? node964 : 3'b010;
											assign node964 = (inp[10]) ? node968 : node965;
												assign node965 = (inp[5]) ? 3'b100 : 3'b000;
												assign node968 = (inp[5]) ? 3'b010 : 3'b100;

endmodule