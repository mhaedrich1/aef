module dtc_split5_bm61 (
	input  wire [12-1:0] inp,
	output wire [11-1:0] outp
);

	wire [11-1:0] node1;
	wire [11-1:0] node2;
	wire [11-1:0] node3;
	wire [11-1:0] node4;
	wire [11-1:0] node5;
	wire [11-1:0] node6;
	wire [11-1:0] node7;
	wire [11-1:0] node8;
	wire [11-1:0] node9;
	wire [11-1:0] node10;
	wire [11-1:0] node13;
	wire [11-1:0] node14;
	wire [11-1:0] node17;
	wire [11-1:0] node20;
	wire [11-1:0] node22;
	wire [11-1:0] node23;
	wire [11-1:0] node27;
	wire [11-1:0] node28;
	wire [11-1:0] node31;
	wire [11-1:0] node32;
	wire [11-1:0] node35;
	wire [11-1:0] node38;
	wire [11-1:0] node39;
	wire [11-1:0] node40;
	wire [11-1:0] node41;
	wire [11-1:0] node43;
	wire [11-1:0] node47;
	wire [11-1:0] node48;
	wire [11-1:0] node49;
	wire [11-1:0] node54;
	wire [11-1:0] node55;
	wire [11-1:0] node56;
	wire [11-1:0] node59;
	wire [11-1:0] node62;
	wire [11-1:0] node63;
	wire [11-1:0] node65;
	wire [11-1:0] node68;
	wire [11-1:0] node71;
	wire [11-1:0] node72;
	wire [11-1:0] node73;
	wire [11-1:0] node75;
	wire [11-1:0] node76;
	wire [11-1:0] node79;
	wire [11-1:0] node81;
	wire [11-1:0] node84;
	wire [11-1:0] node85;
	wire [11-1:0] node86;
	wire [11-1:0] node89;
	wire [11-1:0] node92;
	wire [11-1:0] node93;
	wire [11-1:0] node96;
	wire [11-1:0] node97;
	wire [11-1:0] node101;
	wire [11-1:0] node102;
	wire [11-1:0] node103;
	wire [11-1:0] node106;
	wire [11-1:0] node108;
	wire [11-1:0] node111;
	wire [11-1:0] node112;
	wire [11-1:0] node113;
	wire [11-1:0] node116;
	wire [11-1:0] node119;
	wire [11-1:0] node121;
	wire [11-1:0] node123;
	wire [11-1:0] node126;
	wire [11-1:0] node127;
	wire [11-1:0] node128;
	wire [11-1:0] node129;
	wire [11-1:0] node130;
	wire [11-1:0] node131;
	wire [11-1:0] node132;
	wire [11-1:0] node135;
	wire [11-1:0] node138;
	wire [11-1:0] node141;
	wire [11-1:0] node142;
	wire [11-1:0] node146;
	wire [11-1:0] node147;
	wire [11-1:0] node148;
	wire [11-1:0] node151;
	wire [11-1:0] node154;
	wire [11-1:0] node155;
	wire [11-1:0] node158;
	wire [11-1:0] node161;
	wire [11-1:0] node162;
	wire [11-1:0] node163;
	wire [11-1:0] node164;
	wire [11-1:0] node165;
	wire [11-1:0] node168;
	wire [11-1:0] node171;
	wire [11-1:0] node173;
	wire [11-1:0] node176;
	wire [11-1:0] node177;
	wire [11-1:0] node180;
	wire [11-1:0] node181;
	wire [11-1:0] node185;
	wire [11-1:0] node186;
	wire [11-1:0] node187;
	wire [11-1:0] node190;
	wire [11-1:0] node191;
	wire [11-1:0] node194;
	wire [11-1:0] node197;
	wire [11-1:0] node198;
	wire [11-1:0] node199;
	wire [11-1:0] node203;
	wire [11-1:0] node205;
	wire [11-1:0] node208;
	wire [11-1:0] node209;
	wire [11-1:0] node210;
	wire [11-1:0] node211;
	wire [11-1:0] node212;
	wire [11-1:0] node216;
	wire [11-1:0] node217;
	wire [11-1:0] node220;
	wire [11-1:0] node221;
	wire [11-1:0] node224;
	wire [11-1:0] node227;
	wire [11-1:0] node228;
	wire [11-1:0] node231;
	wire [11-1:0] node232;
	wire [11-1:0] node233;
	wire [11-1:0] node237;
	wire [11-1:0] node240;
	wire [11-1:0] node241;
	wire [11-1:0] node242;
	wire [11-1:0] node243;
	wire [11-1:0] node246;
	wire [11-1:0] node249;
	wire [11-1:0] node250;
	wire [11-1:0] node253;
	wire [11-1:0] node256;
	wire [11-1:0] node257;
	wire [11-1:0] node258;
	wire [11-1:0] node262;
	wire [11-1:0] node263;
	wire [11-1:0] node264;
	wire [11-1:0] node269;
	wire [11-1:0] node270;
	wire [11-1:0] node271;
	wire [11-1:0] node272;
	wire [11-1:0] node273;
	wire [11-1:0] node274;
	wire [11-1:0] node275;
	wire [11-1:0] node276;
	wire [11-1:0] node280;
	wire [11-1:0] node283;
	wire [11-1:0] node285;
	wire [11-1:0] node288;
	wire [11-1:0] node289;
	wire [11-1:0] node290;
	wire [11-1:0] node291;
	wire [11-1:0] node295;
	wire [11-1:0] node298;
	wire [11-1:0] node299;
	wire [11-1:0] node302;
	wire [11-1:0] node304;
	wire [11-1:0] node307;
	wire [11-1:0] node308;
	wire [11-1:0] node309;
	wire [11-1:0] node310;
	wire [11-1:0] node314;
	wire [11-1:0] node315;
	wire [11-1:0] node319;
	wire [11-1:0] node320;
	wire [11-1:0] node322;
	wire [11-1:0] node323;
	wire [11-1:0] node327;
	wire [11-1:0] node328;
	wire [11-1:0] node329;
	wire [11-1:0] node333;
	wire [11-1:0] node336;
	wire [11-1:0] node337;
	wire [11-1:0] node338;
	wire [11-1:0] node339;
	wire [11-1:0] node340;
	wire [11-1:0] node343;
	wire [11-1:0] node344;
	wire [11-1:0] node348;
	wire [11-1:0] node349;
	wire [11-1:0] node350;
	wire [11-1:0] node354;
	wire [11-1:0] node356;
	wire [11-1:0] node359;
	wire [11-1:0] node360;
	wire [11-1:0] node361;
	wire [11-1:0] node364;
	wire [11-1:0] node367;
	wire [11-1:0] node368;
	wire [11-1:0] node369;
	wire [11-1:0] node372;
	wire [11-1:0] node375;
	wire [11-1:0] node378;
	wire [11-1:0] node379;
	wire [11-1:0] node380;
	wire [11-1:0] node382;
	wire [11-1:0] node384;
	wire [11-1:0] node387;
	wire [11-1:0] node388;
	wire [11-1:0] node390;
	wire [11-1:0] node393;
	wire [11-1:0] node396;
	wire [11-1:0] node397;
	wire [11-1:0] node398;
	wire [11-1:0] node399;
	wire [11-1:0] node402;
	wire [11-1:0] node405;
	wire [11-1:0] node408;
	wire [11-1:0] node409;
	wire [11-1:0] node412;
	wire [11-1:0] node415;
	wire [11-1:0] node416;
	wire [11-1:0] node417;
	wire [11-1:0] node418;
	wire [11-1:0] node419;
	wire [11-1:0] node421;
	wire [11-1:0] node424;
	wire [11-1:0] node425;
	wire [11-1:0] node428;
	wire [11-1:0] node429;
	wire [11-1:0] node432;
	wire [11-1:0] node435;
	wire [11-1:0] node436;
	wire [11-1:0] node438;
	wire [11-1:0] node440;
	wire [11-1:0] node443;
	wire [11-1:0] node444;
	wire [11-1:0] node448;
	wire [11-1:0] node449;
	wire [11-1:0] node450;
	wire [11-1:0] node451;
	wire [11-1:0] node455;
	wire [11-1:0] node456;
	wire [11-1:0] node458;
	wire [11-1:0] node461;
	wire [11-1:0] node462;
	wire [11-1:0] node466;
	wire [11-1:0] node467;
	wire [11-1:0] node469;
	wire [11-1:0] node472;
	wire [11-1:0] node475;
	wire [11-1:0] node476;
	wire [11-1:0] node477;
	wire [11-1:0] node478;
	wire [11-1:0] node479;
	wire [11-1:0] node483;
	wire [11-1:0] node484;
	wire [11-1:0] node485;
	wire [11-1:0] node489;
	wire [11-1:0] node490;
	wire [11-1:0] node494;
	wire [11-1:0] node495;
	wire [11-1:0] node496;
	wire [11-1:0] node497;
	wire [11-1:0] node501;
	wire [11-1:0] node504;
	wire [11-1:0] node505;
	wire [11-1:0] node506;
	wire [11-1:0] node509;
	wire [11-1:0] node512;
	wire [11-1:0] node514;
	wire [11-1:0] node517;
	wire [11-1:0] node518;
	wire [11-1:0] node520;
	wire [11-1:0] node521;
	wire [11-1:0] node523;
	wire [11-1:0] node526;
	wire [11-1:0] node528;
	wire [11-1:0] node531;
	wire [11-1:0] node532;
	wire [11-1:0] node533;
	wire [11-1:0] node536;
	wire [11-1:0] node537;
	wire [11-1:0] node541;
	wire [11-1:0] node544;
	wire [11-1:0] node545;
	wire [11-1:0] node546;
	wire [11-1:0] node547;
	wire [11-1:0] node548;
	wire [11-1:0] node549;
	wire [11-1:0] node550;
	wire [11-1:0] node551;
	wire [11-1:0] node554;
	wire [11-1:0] node555;
	wire [11-1:0] node559;
	wire [11-1:0] node562;
	wire [11-1:0] node563;
	wire [11-1:0] node564;
	wire [11-1:0] node565;
	wire [11-1:0] node568;
	wire [11-1:0] node571;
	wire [11-1:0] node574;
	wire [11-1:0] node577;
	wire [11-1:0] node578;
	wire [11-1:0] node579;
	wire [11-1:0] node580;
	wire [11-1:0] node582;
	wire [11-1:0] node585;
	wire [11-1:0] node589;
	wire [11-1:0] node590;
	wire [11-1:0] node591;
	wire [11-1:0] node594;
	wire [11-1:0] node598;
	wire [11-1:0] node599;
	wire [11-1:0] node600;
	wire [11-1:0] node601;
	wire [11-1:0] node602;
	wire [11-1:0] node606;
	wire [11-1:0] node607;
	wire [11-1:0] node609;
	wire [11-1:0] node613;
	wire [11-1:0] node614;
	wire [11-1:0] node617;
	wire [11-1:0] node618;
	wire [11-1:0] node621;
	wire [11-1:0] node624;
	wire [11-1:0] node625;
	wire [11-1:0] node626;
	wire [11-1:0] node627;
	wire [11-1:0] node631;
	wire [11-1:0] node634;
	wire [11-1:0] node635;
	wire [11-1:0] node636;
	wire [11-1:0] node640;
	wire [11-1:0] node641;
	wire [11-1:0] node642;
	wire [11-1:0] node645;
	wire [11-1:0] node648;
	wire [11-1:0] node650;
	wire [11-1:0] node653;
	wire [11-1:0] node654;
	wire [11-1:0] node655;
	wire [11-1:0] node656;
	wire [11-1:0] node657;
	wire [11-1:0] node658;
	wire [11-1:0] node659;
	wire [11-1:0] node662;
	wire [11-1:0] node665;
	wire [11-1:0] node668;
	wire [11-1:0] node671;
	wire [11-1:0] node672;
	wire [11-1:0] node674;
	wire [11-1:0] node677;
	wire [11-1:0] node679;
	wire [11-1:0] node682;
	wire [11-1:0] node683;
	wire [11-1:0] node684;
	wire [11-1:0] node685;
	wire [11-1:0] node689;
	wire [11-1:0] node690;
	wire [11-1:0] node692;
	wire [11-1:0] node695;
	wire [11-1:0] node698;
	wire [11-1:0] node699;
	wire [11-1:0] node700;
	wire [11-1:0] node702;
	wire [11-1:0] node705;
	wire [11-1:0] node706;
	wire [11-1:0] node710;
	wire [11-1:0] node713;
	wire [11-1:0] node714;
	wire [11-1:0] node715;
	wire [11-1:0] node716;
	wire [11-1:0] node719;
	wire [11-1:0] node721;
	wire [11-1:0] node723;
	wire [11-1:0] node726;
	wire [11-1:0] node727;
	wire [11-1:0] node728;
	wire [11-1:0] node729;
	wire [11-1:0] node732;
	wire [11-1:0] node735;
	wire [11-1:0] node736;
	wire [11-1:0] node740;
	wire [11-1:0] node741;
	wire [11-1:0] node743;
	wire [11-1:0] node747;
	wire [11-1:0] node748;
	wire [11-1:0] node749;
	wire [11-1:0] node752;
	wire [11-1:0] node753;
	wire [11-1:0] node755;
	wire [11-1:0] node758;
	wire [11-1:0] node760;
	wire [11-1:0] node763;
	wire [11-1:0] node765;
	wire [11-1:0] node767;
	wire [11-1:0] node770;
	wire [11-1:0] node771;
	wire [11-1:0] node772;
	wire [11-1:0] node773;
	wire [11-1:0] node774;
	wire [11-1:0] node775;
	wire [11-1:0] node778;
	wire [11-1:0] node779;
	wire [11-1:0] node782;
	wire [11-1:0] node785;
	wire [11-1:0] node786;
	wire [11-1:0] node788;
	wire [11-1:0] node790;
	wire [11-1:0] node793;
	wire [11-1:0] node794;
	wire [11-1:0] node797;
	wire [11-1:0] node798;
	wire [11-1:0] node802;
	wire [11-1:0] node803;
	wire [11-1:0] node804;
	wire [11-1:0] node805;
	wire [11-1:0] node808;
	wire [11-1:0] node811;
	wire [11-1:0] node814;
	wire [11-1:0] node815;
	wire [11-1:0] node816;
	wire [11-1:0] node820;
	wire [11-1:0] node821;
	wire [11-1:0] node825;
	wire [11-1:0] node826;
	wire [11-1:0] node827;
	wire [11-1:0] node828;
	wire [11-1:0] node829;
	wire [11-1:0] node832;
	wire [11-1:0] node835;
	wire [11-1:0] node836;
	wire [11-1:0] node838;
	wire [11-1:0] node841;
	wire [11-1:0] node844;
	wire [11-1:0] node845;
	wire [11-1:0] node846;
	wire [11-1:0] node847;
	wire [11-1:0] node851;
	wire [11-1:0] node854;
	wire [11-1:0] node855;
	wire [11-1:0] node858;
	wire [11-1:0] node861;
	wire [11-1:0] node862;
	wire [11-1:0] node863;
	wire [11-1:0] node864;
	wire [11-1:0] node866;
	wire [11-1:0] node870;
	wire [11-1:0] node871;
	wire [11-1:0] node874;
	wire [11-1:0] node877;
	wire [11-1:0] node878;
	wire [11-1:0] node880;
	wire [11-1:0] node883;
	wire [11-1:0] node885;
	wire [11-1:0] node887;
	wire [11-1:0] node890;
	wire [11-1:0] node891;
	wire [11-1:0] node892;
	wire [11-1:0] node893;
	wire [11-1:0] node894;
	wire [11-1:0] node896;
	wire [11-1:0] node899;
	wire [11-1:0] node900;
	wire [11-1:0] node903;
	wire [11-1:0] node905;
	wire [11-1:0] node908;
	wire [11-1:0] node909;
	wire [11-1:0] node911;
	wire [11-1:0] node912;
	wire [11-1:0] node916;
	wire [11-1:0] node918;
	wire [11-1:0] node921;
	wire [11-1:0] node922;
	wire [11-1:0] node923;
	wire [11-1:0] node924;
	wire [11-1:0] node927;
	wire [11-1:0] node930;
	wire [11-1:0] node931;
	wire [11-1:0] node934;
	wire [11-1:0] node937;
	wire [11-1:0] node938;
	wire [11-1:0] node940;
	wire [11-1:0] node943;
	wire [11-1:0] node946;
	wire [11-1:0] node947;
	wire [11-1:0] node948;
	wire [11-1:0] node949;
	wire [11-1:0] node950;
	wire [11-1:0] node954;
	wire [11-1:0] node955;
	wire [11-1:0] node959;
	wire [11-1:0] node960;
	wire [11-1:0] node961;
	wire [11-1:0] node964;
	wire [11-1:0] node967;
	wire [11-1:0] node969;
	wire [11-1:0] node972;
	wire [11-1:0] node973;
	wire [11-1:0] node974;
	wire [11-1:0] node975;
	wire [11-1:0] node979;
	wire [11-1:0] node981;
	wire [11-1:0] node984;
	wire [11-1:0] node985;
	wire [11-1:0] node986;
	wire [11-1:0] node988;
	wire [11-1:0] node991;
	wire [11-1:0] node994;
	wire [11-1:0] node997;
	wire [11-1:0] node998;
	wire [11-1:0] node999;
	wire [11-1:0] node1000;
	wire [11-1:0] node1001;
	wire [11-1:0] node1002;
	wire [11-1:0] node1003;
	wire [11-1:0] node1004;
	wire [11-1:0] node1005;
	wire [11-1:0] node1008;
	wire [11-1:0] node1011;
	wire [11-1:0] node1012;
	wire [11-1:0] node1015;
	wire [11-1:0] node1018;
	wire [11-1:0] node1019;
	wire [11-1:0] node1020;
	wire [11-1:0] node1023;
	wire [11-1:0] node1026;
	wire [11-1:0] node1027;
	wire [11-1:0] node1030;
	wire [11-1:0] node1033;
	wire [11-1:0] node1034;
	wire [11-1:0] node1035;
	wire [11-1:0] node1038;
	wire [11-1:0] node1039;
	wire [11-1:0] node1043;
	wire [11-1:0] node1044;
	wire [11-1:0] node1045;
	wire [11-1:0] node1047;
	wire [11-1:0] node1050;
	wire [11-1:0] node1051;
	wire [11-1:0] node1055;
	wire [11-1:0] node1056;
	wire [11-1:0] node1060;
	wire [11-1:0] node1061;
	wire [11-1:0] node1062;
	wire [11-1:0] node1063;
	wire [11-1:0] node1065;
	wire [11-1:0] node1067;
	wire [11-1:0] node1070;
	wire [11-1:0] node1073;
	wire [11-1:0] node1074;
	wire [11-1:0] node1075;
	wire [11-1:0] node1078;
	wire [11-1:0] node1081;
	wire [11-1:0] node1082;
	wire [11-1:0] node1085;
	wire [11-1:0] node1088;
	wire [11-1:0] node1089;
	wire [11-1:0] node1090;
	wire [11-1:0] node1091;
	wire [11-1:0] node1094;
	wire [11-1:0] node1097;
	wire [11-1:0] node1099;
	wire [11-1:0] node1101;
	wire [11-1:0] node1104;
	wire [11-1:0] node1105;
	wire [11-1:0] node1107;
	wire [11-1:0] node1108;
	wire [11-1:0] node1112;
	wire [11-1:0] node1113;
	wire [11-1:0] node1115;
	wire [11-1:0] node1118;
	wire [11-1:0] node1119;
	wire [11-1:0] node1123;
	wire [11-1:0] node1124;
	wire [11-1:0] node1125;
	wire [11-1:0] node1126;
	wire [11-1:0] node1127;
	wire [11-1:0] node1128;
	wire [11-1:0] node1130;
	wire [11-1:0] node1133;
	wire [11-1:0] node1134;
	wire [11-1:0] node1138;
	wire [11-1:0] node1139;
	wire [11-1:0] node1142;
	wire [11-1:0] node1145;
	wire [11-1:0] node1146;
	wire [11-1:0] node1147;
	wire [11-1:0] node1150;
	wire [11-1:0] node1153;
	wire [11-1:0] node1154;
	wire [11-1:0] node1155;
	wire [11-1:0] node1159;
	wire [11-1:0] node1162;
	wire [11-1:0] node1163;
	wire [11-1:0] node1164;
	wire [11-1:0] node1166;
	wire [11-1:0] node1169;
	wire [11-1:0] node1170;
	wire [11-1:0] node1173;
	wire [11-1:0] node1176;
	wire [11-1:0] node1177;
	wire [11-1:0] node1178;
	wire [11-1:0] node1180;
	wire [11-1:0] node1183;
	wire [11-1:0] node1186;
	wire [11-1:0] node1187;
	wire [11-1:0] node1189;
	wire [11-1:0] node1192;
	wire [11-1:0] node1193;
	wire [11-1:0] node1196;
	wire [11-1:0] node1199;
	wire [11-1:0] node1200;
	wire [11-1:0] node1201;
	wire [11-1:0] node1202;
	wire [11-1:0] node1203;
	wire [11-1:0] node1204;
	wire [11-1:0] node1207;
	wire [11-1:0] node1210;
	wire [11-1:0] node1212;
	wire [11-1:0] node1215;
	wire [11-1:0] node1216;
	wire [11-1:0] node1219;
	wire [11-1:0] node1222;
	wire [11-1:0] node1223;
	wire [11-1:0] node1224;
	wire [11-1:0] node1227;
	wire [11-1:0] node1230;
	wire [11-1:0] node1231;
	wire [11-1:0] node1234;
	wire [11-1:0] node1237;
	wire [11-1:0] node1238;
	wire [11-1:0] node1239;
	wire [11-1:0] node1241;
	wire [11-1:0] node1244;
	wire [11-1:0] node1246;
	wire [11-1:0] node1249;
	wire [11-1:0] node1250;
	wire [11-1:0] node1251;
	wire [11-1:0] node1254;
	wire [11-1:0] node1257;
	wire [11-1:0] node1258;
	wire [11-1:0] node1259;
	wire [11-1:0] node1263;
	wire [11-1:0] node1266;
	wire [11-1:0] node1267;
	wire [11-1:0] node1268;
	wire [11-1:0] node1269;
	wire [11-1:0] node1270;
	wire [11-1:0] node1271;
	wire [11-1:0] node1272;
	wire [11-1:0] node1275;
	wire [11-1:0] node1276;
	wire [11-1:0] node1279;
	wire [11-1:0] node1282;
	wire [11-1:0] node1283;
	wire [11-1:0] node1285;
	wire [11-1:0] node1288;
	wire [11-1:0] node1289;
	wire [11-1:0] node1293;
	wire [11-1:0] node1294;
	wire [11-1:0] node1295;
	wire [11-1:0] node1299;
	wire [11-1:0] node1301;
	wire [11-1:0] node1304;
	wire [11-1:0] node1305;
	wire [11-1:0] node1306;
	wire [11-1:0] node1307;
	wire [11-1:0] node1310;
	wire [11-1:0] node1313;
	wire [11-1:0] node1315;
	wire [11-1:0] node1318;
	wire [11-1:0] node1319;
	wire [11-1:0] node1321;
	wire [11-1:0] node1324;
	wire [11-1:0] node1325;
	wire [11-1:0] node1326;
	wire [11-1:0] node1330;
	wire [11-1:0] node1331;
	wire [11-1:0] node1335;
	wire [11-1:0] node1336;
	wire [11-1:0] node1337;
	wire [11-1:0] node1338;
	wire [11-1:0] node1339;
	wire [11-1:0] node1342;
	wire [11-1:0] node1345;
	wire [11-1:0] node1348;
	wire [11-1:0] node1349;
	wire [11-1:0] node1350;
	wire [11-1:0] node1351;
	wire [11-1:0] node1355;
	wire [11-1:0] node1358;
	wire [11-1:0] node1359;
	wire [11-1:0] node1360;
	wire [11-1:0] node1364;
	wire [11-1:0] node1367;
	wire [11-1:0] node1368;
	wire [11-1:0] node1369;
	wire [11-1:0] node1370;
	wire [11-1:0] node1374;
	wire [11-1:0] node1375;
	wire [11-1:0] node1379;
	wire [11-1:0] node1380;
	wire [11-1:0] node1381;
	wire [11-1:0] node1384;
	wire [11-1:0] node1387;
	wire [11-1:0] node1388;
	wire [11-1:0] node1389;
	wire [11-1:0] node1393;
	wire [11-1:0] node1396;
	wire [11-1:0] node1397;
	wire [11-1:0] node1398;
	wire [11-1:0] node1399;
	wire [11-1:0] node1400;
	wire [11-1:0] node1401;
	wire [11-1:0] node1404;
	wire [11-1:0] node1405;
	wire [11-1:0] node1409;
	wire [11-1:0] node1412;
	wire [11-1:0] node1413;
	wire [11-1:0] node1414;
	wire [11-1:0] node1418;
	wire [11-1:0] node1419;
	wire [11-1:0] node1420;
	wire [11-1:0] node1424;
	wire [11-1:0] node1426;
	wire [11-1:0] node1429;
	wire [11-1:0] node1430;
	wire [11-1:0] node1431;
	wire [11-1:0] node1434;
	wire [11-1:0] node1435;
	wire [11-1:0] node1437;
	wire [11-1:0] node1441;
	wire [11-1:0] node1442;
	wire [11-1:0] node1444;
	wire [11-1:0] node1447;
	wire [11-1:0] node1449;
	wire [11-1:0] node1450;
	wire [11-1:0] node1454;
	wire [11-1:0] node1455;
	wire [11-1:0] node1456;
	wire [11-1:0] node1458;
	wire [11-1:0] node1459;
	wire [11-1:0] node1463;
	wire [11-1:0] node1464;
	wire [11-1:0] node1465;
	wire [11-1:0] node1468;
	wire [11-1:0] node1471;
	wire [11-1:0] node1474;
	wire [11-1:0] node1475;
	wire [11-1:0] node1476;
	wire [11-1:0] node1477;
	wire [11-1:0] node1481;
	wire [11-1:0] node1484;
	wire [11-1:0] node1486;
	wire [11-1:0] node1487;
	wire [11-1:0] node1491;
	wire [11-1:0] node1492;
	wire [11-1:0] node1493;
	wire [11-1:0] node1494;
	wire [11-1:0] node1495;
	wire [11-1:0] node1496;
	wire [11-1:0] node1497;
	wire [11-1:0] node1498;
	wire [11-1:0] node1499;
	wire [11-1:0] node1502;
	wire [11-1:0] node1505;
	wire [11-1:0] node1508;
	wire [11-1:0] node1509;
	wire [11-1:0] node1512;
	wire [11-1:0] node1515;
	wire [11-1:0] node1516;
	wire [11-1:0] node1517;
	wire [11-1:0] node1518;
	wire [11-1:0] node1522;
	wire [11-1:0] node1525;
	wire [11-1:0] node1527;
	wire [11-1:0] node1529;
	wire [11-1:0] node1532;
	wire [11-1:0] node1533;
	wire [11-1:0] node1534;
	wire [11-1:0] node1535;
	wire [11-1:0] node1538;
	wire [11-1:0] node1541;
	wire [11-1:0] node1542;
	wire [11-1:0] node1545;
	wire [11-1:0] node1547;
	wire [11-1:0] node1550;
	wire [11-1:0] node1551;
	wire [11-1:0] node1552;
	wire [11-1:0] node1554;
	wire [11-1:0] node1557;
	wire [11-1:0] node1559;
	wire [11-1:0] node1562;
	wire [11-1:0] node1563;
	wire [11-1:0] node1564;
	wire [11-1:0] node1567;
	wire [11-1:0] node1570;
	wire [11-1:0] node1572;
	wire [11-1:0] node1575;
	wire [11-1:0] node1576;
	wire [11-1:0] node1577;
	wire [11-1:0] node1578;
	wire [11-1:0] node1579;
	wire [11-1:0] node1582;
	wire [11-1:0] node1583;
	wire [11-1:0] node1586;
	wire [11-1:0] node1589;
	wire [11-1:0] node1590;
	wire [11-1:0] node1591;
	wire [11-1:0] node1595;
	wire [11-1:0] node1597;
	wire [11-1:0] node1600;
	wire [11-1:0] node1601;
	wire [11-1:0] node1604;
	wire [11-1:0] node1605;
	wire [11-1:0] node1607;
	wire [11-1:0] node1610;
	wire [11-1:0] node1613;
	wire [11-1:0] node1614;
	wire [11-1:0] node1615;
	wire [11-1:0] node1616;
	wire [11-1:0] node1619;
	wire [11-1:0] node1622;
	wire [11-1:0] node1623;
	wire [11-1:0] node1624;
	wire [11-1:0] node1628;
	wire [11-1:0] node1629;
	wire [11-1:0] node1633;
	wire [11-1:0] node1634;
	wire [11-1:0] node1635;
	wire [11-1:0] node1638;
	wire [11-1:0] node1639;
	wire [11-1:0] node1643;
	wire [11-1:0] node1644;
	wire [11-1:0] node1646;
	wire [11-1:0] node1649;
	wire [11-1:0] node1650;
	wire [11-1:0] node1654;
	wire [11-1:0] node1655;
	wire [11-1:0] node1656;
	wire [11-1:0] node1657;
	wire [11-1:0] node1658;
	wire [11-1:0] node1659;
	wire [11-1:0] node1660;
	wire [11-1:0] node1665;
	wire [11-1:0] node1666;
	wire [11-1:0] node1669;
	wire [11-1:0] node1672;
	wire [11-1:0] node1673;
	wire [11-1:0] node1675;
	wire [11-1:0] node1678;
	wire [11-1:0] node1679;
	wire [11-1:0] node1682;
	wire [11-1:0] node1684;
	wire [11-1:0] node1687;
	wire [11-1:0] node1688;
	wire [11-1:0] node1689;
	wire [11-1:0] node1691;
	wire [11-1:0] node1694;
	wire [11-1:0] node1695;
	wire [11-1:0] node1698;
	wire [11-1:0] node1700;
	wire [11-1:0] node1703;
	wire [11-1:0] node1704;
	wire [11-1:0] node1706;
	wire [11-1:0] node1709;
	wire [11-1:0] node1710;
	wire [11-1:0] node1713;
	wire [11-1:0] node1714;
	wire [11-1:0] node1717;
	wire [11-1:0] node1720;
	wire [11-1:0] node1721;
	wire [11-1:0] node1722;
	wire [11-1:0] node1723;
	wire [11-1:0] node1725;
	wire [11-1:0] node1728;
	wire [11-1:0] node1729;
	wire [11-1:0] node1730;
	wire [11-1:0] node1733;
	wire [11-1:0] node1736;
	wire [11-1:0] node1739;
	wire [11-1:0] node1740;
	wire [11-1:0] node1741;
	wire [11-1:0] node1744;
	wire [11-1:0] node1745;
	wire [11-1:0] node1749;
	wire [11-1:0] node1750;
	wire [11-1:0] node1751;
	wire [11-1:0] node1755;
	wire [11-1:0] node1758;
	wire [11-1:0] node1759;
	wire [11-1:0] node1760;
	wire [11-1:0] node1761;
	wire [11-1:0] node1762;
	wire [11-1:0] node1766;
	wire [11-1:0] node1769;
	wire [11-1:0] node1771;
	wire [11-1:0] node1772;
	wire [11-1:0] node1776;
	wire [11-1:0] node1777;
	wire [11-1:0] node1778;
	wire [11-1:0] node1781;
	wire [11-1:0] node1783;
	wire [11-1:0] node1786;
	wire [11-1:0] node1788;
	wire [11-1:0] node1791;
	wire [11-1:0] node1792;
	wire [11-1:0] node1793;
	wire [11-1:0] node1794;
	wire [11-1:0] node1795;
	wire [11-1:0] node1796;
	wire [11-1:0] node1797;
	wire [11-1:0] node1800;
	wire [11-1:0] node1802;
	wire [11-1:0] node1805;
	wire [11-1:0] node1808;
	wire [11-1:0] node1809;
	wire [11-1:0] node1810;
	wire [11-1:0] node1811;
	wire [11-1:0] node1814;
	wire [11-1:0] node1817;
	wire [11-1:0] node1820;
	wire [11-1:0] node1823;
	wire [11-1:0] node1824;
	wire [11-1:0] node1825;
	wire [11-1:0] node1826;
	wire [11-1:0] node1830;
	wire [11-1:0] node1831;
	wire [11-1:0] node1835;
	wire [11-1:0] node1836;
	wire [11-1:0] node1837;
	wire [11-1:0] node1838;
	wire [11-1:0] node1843;
	wire [11-1:0] node1845;
	wire [11-1:0] node1848;
	wire [11-1:0] node1849;
	wire [11-1:0] node1850;
	wire [11-1:0] node1851;
	wire [11-1:0] node1854;
	wire [11-1:0] node1857;
	wire [11-1:0] node1858;
	wire [11-1:0] node1859;
	wire [11-1:0] node1862;
	wire [11-1:0] node1865;
	wire [11-1:0] node1868;
	wire [11-1:0] node1869;
	wire [11-1:0] node1870;
	wire [11-1:0] node1871;
	wire [11-1:0] node1874;
	wire [11-1:0] node1877;
	wire [11-1:0] node1878;
	wire [11-1:0] node1881;
	wire [11-1:0] node1884;
	wire [11-1:0] node1885;
	wire [11-1:0] node1886;
	wire [11-1:0] node1890;
	wire [11-1:0] node1891;
	wire [11-1:0] node1893;
	wire [11-1:0] node1897;
	wire [11-1:0] node1898;
	wire [11-1:0] node1899;
	wire [11-1:0] node1900;
	wire [11-1:0] node1901;
	wire [11-1:0] node1902;
	wire [11-1:0] node1905;
	wire [11-1:0] node1906;
	wire [11-1:0] node1909;
	wire [11-1:0] node1912;
	wire [11-1:0] node1913;
	wire [11-1:0] node1916;
	wire [11-1:0] node1919;
	wire [11-1:0] node1920;
	wire [11-1:0] node1921;
	wire [11-1:0] node1922;
	wire [11-1:0] node1926;
	wire [11-1:0] node1929;
	wire [11-1:0] node1930;
	wire [11-1:0] node1933;
	wire [11-1:0] node1935;
	wire [11-1:0] node1938;
	wire [11-1:0] node1939;
	wire [11-1:0] node1940;
	wire [11-1:0] node1941;
	wire [11-1:0] node1944;
	wire [11-1:0] node1945;
	wire [11-1:0] node1949;
	wire [11-1:0] node1951;
	wire [11-1:0] node1954;
	wire [11-1:0] node1955;
	wire [11-1:0] node1956;
	wire [11-1:0] node1959;
	wire [11-1:0] node1961;
	wire [11-1:0] node1964;
	wire [11-1:0] node1967;
	wire [11-1:0] node1968;
	wire [11-1:0] node1969;
	wire [11-1:0] node1970;
	wire [11-1:0] node1973;
	wire [11-1:0] node1975;
	wire [11-1:0] node1977;
	wire [11-1:0] node1980;
	wire [11-1:0] node1981;
	wire [11-1:0] node1982;
	wire [11-1:0] node1985;
	wire [11-1:0] node1989;
	wire [11-1:0] node1990;
	wire [11-1:0] node1991;
	wire [11-1:0] node1994;
	wire [11-1:0] node1997;
	wire [11-1:0] node1998;
	wire [11-1:0] node1999;
	wire [11-1:0] node2002;
	wire [11-1:0] node2005;
	wire [11-1:0] node2007;
	wire [11-1:0] node2010;
	wire [11-1:0] node2011;
	wire [11-1:0] node2012;
	wire [11-1:0] node2013;
	wire [11-1:0] node2014;
	wire [11-1:0] node2015;
	wire [11-1:0] node2016;
	wire [11-1:0] node2017;
	wire [11-1:0] node2018;
	wire [11-1:0] node2020;
	wire [11-1:0] node2023;
	wire [11-1:0] node2024;
	wire [11-1:0] node2027;
	wire [11-1:0] node2028;
	wire [11-1:0] node2031;
	wire [11-1:0] node2034;
	wire [11-1:0] node2035;
	wire [11-1:0] node2037;
	wire [11-1:0] node2040;
	wire [11-1:0] node2041;
	wire [11-1:0] node2043;
	wire [11-1:0] node2047;
	wire [11-1:0] node2048;
	wire [11-1:0] node2049;
	wire [11-1:0] node2052;
	wire [11-1:0] node2053;
	wire [11-1:0] node2054;
	wire [11-1:0] node2059;
	wire [11-1:0] node2060;
	wire [11-1:0] node2062;
	wire [11-1:0] node2065;
	wire [11-1:0] node2066;
	wire [11-1:0] node2069;
	wire [11-1:0] node2071;
	wire [11-1:0] node2074;
	wire [11-1:0] node2075;
	wire [11-1:0] node2076;
	wire [11-1:0] node2077;
	wire [11-1:0] node2079;
	wire [11-1:0] node2082;
	wire [11-1:0] node2085;
	wire [11-1:0] node2086;
	wire [11-1:0] node2087;
	wire [11-1:0] node2091;
	wire [11-1:0] node2093;
	wire [11-1:0] node2096;
	wire [11-1:0] node2097;
	wire [11-1:0] node2098;
	wire [11-1:0] node2101;
	wire [11-1:0] node2103;
	wire [11-1:0] node2106;
	wire [11-1:0] node2107;
	wire [11-1:0] node2108;
	wire [11-1:0] node2110;
	wire [11-1:0] node2114;
	wire [11-1:0] node2115;
	wire [11-1:0] node2117;
	wire [11-1:0] node2120;
	wire [11-1:0] node2123;
	wire [11-1:0] node2124;
	wire [11-1:0] node2125;
	wire [11-1:0] node2126;
	wire [11-1:0] node2127;
	wire [11-1:0] node2128;
	wire [11-1:0] node2129;
	wire [11-1:0] node2134;
	wire [11-1:0] node2135;
	wire [11-1:0] node2138;
	wire [11-1:0] node2141;
	wire [11-1:0] node2142;
	wire [11-1:0] node2143;
	wire [11-1:0] node2146;
	wire [11-1:0] node2147;
	wire [11-1:0] node2151;
	wire [11-1:0] node2152;
	wire [11-1:0] node2156;
	wire [11-1:0] node2157;
	wire [11-1:0] node2158;
	wire [11-1:0] node2159;
	wire [11-1:0] node2160;
	wire [11-1:0] node2165;
	wire [11-1:0] node2166;
	wire [11-1:0] node2169;
	wire [11-1:0] node2170;
	wire [11-1:0] node2174;
	wire [11-1:0] node2175;
	wire [11-1:0] node2176;
	wire [11-1:0] node2178;
	wire [11-1:0] node2181;
	wire [11-1:0] node2182;
	wire [11-1:0] node2186;
	wire [11-1:0] node2187;
	wire [11-1:0] node2189;
	wire [11-1:0] node2192;
	wire [11-1:0] node2195;
	wire [11-1:0] node2196;
	wire [11-1:0] node2197;
	wire [11-1:0] node2198;
	wire [11-1:0] node2200;
	wire [11-1:0] node2203;
	wire [11-1:0] node2204;
	wire [11-1:0] node2205;
	wire [11-1:0] node2210;
	wire [11-1:0] node2211;
	wire [11-1:0] node2212;
	wire [11-1:0] node2214;
	wire [11-1:0] node2218;
	wire [11-1:0] node2220;
	wire [11-1:0] node2221;
	wire [11-1:0] node2225;
	wire [11-1:0] node2226;
	wire [11-1:0] node2227;
	wire [11-1:0] node2230;
	wire [11-1:0] node2231;
	wire [11-1:0] node2234;
	wire [11-1:0] node2235;
	wire [11-1:0] node2238;
	wire [11-1:0] node2241;
	wire [11-1:0] node2242;
	wire [11-1:0] node2243;
	wire [11-1:0] node2246;
	wire [11-1:0] node2247;
	wire [11-1:0] node2250;
	wire [11-1:0] node2253;
	wire [11-1:0] node2254;
	wire [11-1:0] node2256;
	wire [11-1:0] node2259;
	wire [11-1:0] node2262;
	wire [11-1:0] node2263;
	wire [11-1:0] node2264;
	wire [11-1:0] node2265;
	wire [11-1:0] node2266;
	wire [11-1:0] node2267;
	wire [11-1:0] node2268;
	wire [11-1:0] node2271;
	wire [11-1:0] node2272;
	wire [11-1:0] node2276;
	wire [11-1:0] node2279;
	wire [11-1:0] node2280;
	wire [11-1:0] node2282;
	wire [11-1:0] node2285;
	wire [11-1:0] node2286;
	wire [11-1:0] node2289;
	wire [11-1:0] node2290;
	wire [11-1:0] node2293;
	wire [11-1:0] node2296;
	wire [11-1:0] node2297;
	wire [11-1:0] node2298;
	wire [11-1:0] node2299;
	wire [11-1:0] node2302;
	wire [11-1:0] node2303;
	wire [11-1:0] node2307;
	wire [11-1:0] node2308;
	wire [11-1:0] node2312;
	wire [11-1:0] node2313;
	wire [11-1:0] node2314;
	wire [11-1:0] node2317;
	wire [11-1:0] node2320;
	wire [11-1:0] node2322;
	wire [11-1:0] node2325;
	wire [11-1:0] node2326;
	wire [11-1:0] node2327;
	wire [11-1:0] node2328;
	wire [11-1:0] node2331;
	wire [11-1:0] node2332;
	wire [11-1:0] node2333;
	wire [11-1:0] node2337;
	wire [11-1:0] node2339;
	wire [11-1:0] node2342;
	wire [11-1:0] node2343;
	wire [11-1:0] node2345;
	wire [11-1:0] node2348;
	wire [11-1:0] node2349;
	wire [11-1:0] node2352;
	wire [11-1:0] node2354;
	wire [11-1:0] node2357;
	wire [11-1:0] node2358;
	wire [11-1:0] node2359;
	wire [11-1:0] node2360;
	wire [11-1:0] node2364;
	wire [11-1:0] node2365;
	wire [11-1:0] node2369;
	wire [11-1:0] node2370;
	wire [11-1:0] node2373;
	wire [11-1:0] node2374;
	wire [11-1:0] node2377;
	wire [11-1:0] node2380;
	wire [11-1:0] node2381;
	wire [11-1:0] node2382;
	wire [11-1:0] node2383;
	wire [11-1:0] node2384;
	wire [11-1:0] node2385;
	wire [11-1:0] node2386;
	wire [11-1:0] node2391;
	wire [11-1:0] node2392;
	wire [11-1:0] node2395;
	wire [11-1:0] node2398;
	wire [11-1:0] node2399;
	wire [11-1:0] node2400;
	wire [11-1:0] node2403;
	wire [11-1:0] node2406;
	wire [11-1:0] node2407;
	wire [11-1:0] node2409;
	wire [11-1:0] node2412;
	wire [11-1:0] node2413;
	wire [11-1:0] node2416;
	wire [11-1:0] node2419;
	wire [11-1:0] node2420;
	wire [11-1:0] node2421;
	wire [11-1:0] node2423;
	wire [11-1:0] node2424;
	wire [11-1:0] node2427;
	wire [11-1:0] node2430;
	wire [11-1:0] node2431;
	wire [11-1:0] node2434;
	wire [11-1:0] node2436;
	wire [11-1:0] node2439;
	wire [11-1:0] node2440;
	wire [11-1:0] node2441;
	wire [11-1:0] node2443;
	wire [11-1:0] node2446;
	wire [11-1:0] node2447;
	wire [11-1:0] node2450;
	wire [11-1:0] node2453;
	wire [11-1:0] node2454;
	wire [11-1:0] node2456;
	wire [11-1:0] node2459;
	wire [11-1:0] node2462;
	wire [11-1:0] node2463;
	wire [11-1:0] node2464;
	wire [11-1:0] node2465;
	wire [11-1:0] node2466;
	wire [11-1:0] node2467;
	wire [11-1:0] node2470;
	wire [11-1:0] node2473;
	wire [11-1:0] node2474;
	wire [11-1:0] node2478;
	wire [11-1:0] node2479;
	wire [11-1:0] node2482;
	wire [11-1:0] node2485;
	wire [11-1:0] node2486;
	wire [11-1:0] node2487;
	wire [11-1:0] node2488;
	wire [11-1:0] node2493;
	wire [11-1:0] node2494;
	wire [11-1:0] node2497;
	wire [11-1:0] node2498;
	wire [11-1:0] node2501;
	wire [11-1:0] node2504;
	wire [11-1:0] node2505;
	wire [11-1:0] node2506;
	wire [11-1:0] node2509;
	wire [11-1:0] node2511;
	wire [11-1:0] node2513;
	wire [11-1:0] node2516;
	wire [11-1:0] node2517;
	wire [11-1:0] node2518;
	wire [11-1:0] node2521;
	wire [11-1:0] node2524;
	wire [11-1:0] node2525;
	wire [11-1:0] node2529;
	wire [11-1:0] node2530;
	wire [11-1:0] node2531;
	wire [11-1:0] node2532;
	wire [11-1:0] node2533;
	wire [11-1:0] node2534;
	wire [11-1:0] node2535;
	wire [11-1:0] node2536;
	wire [11-1:0] node2537;
	wire [11-1:0] node2540;
	wire [11-1:0] node2543;
	wire [11-1:0] node2546;
	wire [11-1:0] node2547;
	wire [11-1:0] node2551;
	wire [11-1:0] node2552;
	wire [11-1:0] node2553;
	wire [11-1:0] node2556;
	wire [11-1:0] node2557;
	wire [11-1:0] node2561;
	wire [11-1:0] node2562;
	wire [11-1:0] node2565;
	wire [11-1:0] node2568;
	wire [11-1:0] node2569;
	wire [11-1:0] node2570;
	wire [11-1:0] node2571;
	wire [11-1:0] node2574;
	wire [11-1:0] node2577;
	wire [11-1:0] node2579;
	wire [11-1:0] node2580;
	wire [11-1:0] node2583;
	wire [11-1:0] node2586;
	wire [11-1:0] node2587;
	wire [11-1:0] node2589;
	wire [11-1:0] node2592;
	wire [11-1:0] node2593;
	wire [11-1:0] node2595;
	wire [11-1:0] node2598;
	wire [11-1:0] node2601;
	wire [11-1:0] node2602;
	wire [11-1:0] node2603;
	wire [11-1:0] node2604;
	wire [11-1:0] node2605;
	wire [11-1:0] node2608;
	wire [11-1:0] node2609;
	wire [11-1:0] node2612;
	wire [11-1:0] node2615;
	wire [11-1:0] node2616;
	wire [11-1:0] node2618;
	wire [11-1:0] node2621;
	wire [11-1:0] node2622;
	wire [11-1:0] node2625;
	wire [11-1:0] node2628;
	wire [11-1:0] node2629;
	wire [11-1:0] node2632;
	wire [11-1:0] node2634;
	wire [11-1:0] node2636;
	wire [11-1:0] node2639;
	wire [11-1:0] node2640;
	wire [11-1:0] node2641;
	wire [11-1:0] node2642;
	wire [11-1:0] node2645;
	wire [11-1:0] node2648;
	wire [11-1:0] node2649;
	wire [11-1:0] node2653;
	wire [11-1:0] node2654;
	wire [11-1:0] node2656;
	wire [11-1:0] node2659;
	wire [11-1:0] node2661;
	wire [11-1:0] node2662;
	wire [11-1:0] node2665;
	wire [11-1:0] node2668;
	wire [11-1:0] node2669;
	wire [11-1:0] node2670;
	wire [11-1:0] node2671;
	wire [11-1:0] node2672;
	wire [11-1:0] node2674;
	wire [11-1:0] node2676;
	wire [11-1:0] node2679;
	wire [11-1:0] node2680;
	wire [11-1:0] node2684;
	wire [11-1:0] node2685;
	wire [11-1:0] node2688;
	wire [11-1:0] node2689;
	wire [11-1:0] node2690;
	wire [11-1:0] node2694;
	wire [11-1:0] node2695;
	wire [11-1:0] node2699;
	wire [11-1:0] node2700;
	wire [11-1:0] node2701;
	wire [11-1:0] node2703;
	wire [11-1:0] node2706;
	wire [11-1:0] node2707;
	wire [11-1:0] node2711;
	wire [11-1:0] node2712;
	wire [11-1:0] node2713;
	wire [11-1:0] node2715;
	wire [11-1:0] node2719;
	wire [11-1:0] node2721;
	wire [11-1:0] node2724;
	wire [11-1:0] node2725;
	wire [11-1:0] node2726;
	wire [11-1:0] node2727;
	wire [11-1:0] node2728;
	wire [11-1:0] node2731;
	wire [11-1:0] node2734;
	wire [11-1:0] node2735;
	wire [11-1:0] node2737;
	wire [11-1:0] node2740;
	wire [11-1:0] node2743;
	wire [11-1:0] node2744;
	wire [11-1:0] node2747;
	wire [11-1:0] node2749;
	wire [11-1:0] node2751;
	wire [11-1:0] node2754;
	wire [11-1:0] node2755;
	wire [11-1:0] node2756;
	wire [11-1:0] node2757;
	wire [11-1:0] node2758;
	wire [11-1:0] node2763;
	wire [11-1:0] node2766;
	wire [11-1:0] node2767;
	wire [11-1:0] node2770;
	wire [11-1:0] node2773;
	wire [11-1:0] node2774;
	wire [11-1:0] node2775;
	wire [11-1:0] node2776;
	wire [11-1:0] node2777;
	wire [11-1:0] node2778;
	wire [11-1:0] node2779;
	wire [11-1:0] node2780;
	wire [11-1:0] node2783;
	wire [11-1:0] node2787;
	wire [11-1:0] node2788;
	wire [11-1:0] node2791;
	wire [11-1:0] node2793;
	wire [11-1:0] node2796;
	wire [11-1:0] node2797;
	wire [11-1:0] node2800;
	wire [11-1:0] node2801;
	wire [11-1:0] node2805;
	wire [11-1:0] node2806;
	wire [11-1:0] node2807;
	wire [11-1:0] node2809;
	wire [11-1:0] node2810;
	wire [11-1:0] node2813;
	wire [11-1:0] node2816;
	wire [11-1:0] node2817;
	wire [11-1:0] node2818;
	wire [11-1:0] node2821;
	wire [11-1:0] node2825;
	wire [11-1:0] node2826;
	wire [11-1:0] node2829;
	wire [11-1:0] node2830;
	wire [11-1:0] node2833;
	wire [11-1:0] node2835;
	wire [11-1:0] node2838;
	wire [11-1:0] node2839;
	wire [11-1:0] node2840;
	wire [11-1:0] node2841;
	wire [11-1:0] node2844;
	wire [11-1:0] node2845;
	wire [11-1:0] node2848;
	wire [11-1:0] node2851;
	wire [11-1:0] node2852;
	wire [11-1:0] node2853;
	wire [11-1:0] node2857;
	wire [11-1:0] node2858;
	wire [11-1:0] node2862;
	wire [11-1:0] node2863;
	wire [11-1:0] node2864;
	wire [11-1:0] node2866;
	wire [11-1:0] node2867;
	wire [11-1:0] node2871;
	wire [11-1:0] node2872;
	wire [11-1:0] node2874;
	wire [11-1:0] node2878;
	wire [11-1:0] node2879;
	wire [11-1:0] node2880;
	wire [11-1:0] node2883;
	wire [11-1:0] node2886;
	wire [11-1:0] node2887;
	wire [11-1:0] node2891;
	wire [11-1:0] node2892;
	wire [11-1:0] node2893;
	wire [11-1:0] node2894;
	wire [11-1:0] node2895;
	wire [11-1:0] node2896;
	wire [11-1:0] node2897;
	wire [11-1:0] node2900;
	wire [11-1:0] node2903;
	wire [11-1:0] node2904;
	wire [11-1:0] node2908;
	wire [11-1:0] node2909;
	wire [11-1:0] node2912;
	wire [11-1:0] node2915;
	wire [11-1:0] node2916;
	wire [11-1:0] node2917;
	wire [11-1:0] node2920;
	wire [11-1:0] node2921;
	wire [11-1:0] node2925;
	wire [11-1:0] node2926;
	wire [11-1:0] node2929;
	wire [11-1:0] node2930;
	wire [11-1:0] node2933;
	wire [11-1:0] node2936;
	wire [11-1:0] node2937;
	wire [11-1:0] node2938;
	wire [11-1:0] node2939;
	wire [11-1:0] node2942;
	wire [11-1:0] node2945;
	wire [11-1:0] node2946;
	wire [11-1:0] node2948;
	wire [11-1:0] node2951;
	wire [11-1:0] node2952;
	wire [11-1:0] node2956;
	wire [11-1:0] node2957;
	wire [11-1:0] node2958;
	wire [11-1:0] node2960;
	wire [11-1:0] node2964;
	wire [11-1:0] node2966;
	wire [11-1:0] node2967;
	wire [11-1:0] node2971;
	wire [11-1:0] node2972;
	wire [11-1:0] node2973;
	wire [11-1:0] node2974;
	wire [11-1:0] node2975;
	wire [11-1:0] node2978;
	wire [11-1:0] node2981;
	wire [11-1:0] node2982;
	wire [11-1:0] node2985;
	wire [11-1:0] node2986;
	wire [11-1:0] node2990;
	wire [11-1:0] node2991;
	wire [11-1:0] node2992;
	wire [11-1:0] node2995;
	wire [11-1:0] node2998;
	wire [11-1:0] node3000;
	wire [11-1:0] node3003;
	wire [11-1:0] node3004;
	wire [11-1:0] node3005;
	wire [11-1:0] node3007;
	wire [11-1:0] node3008;
	wire [11-1:0] node3012;
	wire [11-1:0] node3014;
	wire [11-1:0] node3015;
	wire [11-1:0] node3019;
	wire [11-1:0] node3020;
	wire [11-1:0] node3021;
	wire [11-1:0] node3025;
	wire [11-1:0] node3026;
	wire [11-1:0] node3027;
	wire [11-1:0] node3031;
	wire [11-1:0] node3034;
	wire [11-1:0] node3035;
	wire [11-1:0] node3036;
	wire [11-1:0] node3037;
	wire [11-1:0] node3038;
	wire [11-1:0] node3039;
	wire [11-1:0] node3040;
	wire [11-1:0] node3041;
	wire [11-1:0] node3042;
	wire [11-1:0] node3044;
	wire [11-1:0] node3047;
	wire [11-1:0] node3048;
	wire [11-1:0] node3052;
	wire [11-1:0] node3053;
	wire [11-1:0] node3056;
	wire [11-1:0] node3059;
	wire [11-1:0] node3060;
	wire [11-1:0] node3061;
	wire [11-1:0] node3065;
	wire [11-1:0] node3066;
	wire [11-1:0] node3070;
	wire [11-1:0] node3071;
	wire [11-1:0] node3072;
	wire [11-1:0] node3073;
	wire [11-1:0] node3075;
	wire [11-1:0] node3079;
	wire [11-1:0] node3080;
	wire [11-1:0] node3084;
	wire [11-1:0] node3085;
	wire [11-1:0] node3086;
	wire [11-1:0] node3087;
	wire [11-1:0] node3092;
	wire [11-1:0] node3094;
	wire [11-1:0] node3095;
	wire [11-1:0] node3099;
	wire [11-1:0] node3100;
	wire [11-1:0] node3101;
	wire [11-1:0] node3102;
	wire [11-1:0] node3103;
	wire [11-1:0] node3107;
	wire [11-1:0] node3110;
	wire [11-1:0] node3111;
	wire [11-1:0] node3112;
	wire [11-1:0] node3116;
	wire [11-1:0] node3117;
	wire [11-1:0] node3121;
	wire [11-1:0] node3122;
	wire [11-1:0] node3123;
	wire [11-1:0] node3124;
	wire [11-1:0] node3125;
	wire [11-1:0] node3129;
	wire [11-1:0] node3132;
	wire [11-1:0] node3133;
	wire [11-1:0] node3136;
	wire [11-1:0] node3139;
	wire [11-1:0] node3140;
	wire [11-1:0] node3141;
	wire [11-1:0] node3142;
	wire [11-1:0] node3146;
	wire [11-1:0] node3148;
	wire [11-1:0] node3151;
	wire [11-1:0] node3152;
	wire [11-1:0] node3154;
	wire [11-1:0] node3157;
	wire [11-1:0] node3160;
	wire [11-1:0] node3161;
	wire [11-1:0] node3162;
	wire [11-1:0] node3163;
	wire [11-1:0] node3164;
	wire [11-1:0] node3165;
	wire [11-1:0] node3169;
	wire [11-1:0] node3171;
	wire [11-1:0] node3174;
	wire [11-1:0] node3175;
	wire [11-1:0] node3176;
	wire [11-1:0] node3179;
	wire [11-1:0] node3182;
	wire [11-1:0] node3185;
	wire [11-1:0] node3186;
	wire [11-1:0] node3187;
	wire [11-1:0] node3188;
	wire [11-1:0] node3191;
	wire [11-1:0] node3194;
	wire [11-1:0] node3195;
	wire [11-1:0] node3196;
	wire [11-1:0] node3199;
	wire [11-1:0] node3203;
	wire [11-1:0] node3204;
	wire [11-1:0] node3206;
	wire [11-1:0] node3209;
	wire [11-1:0] node3210;
	wire [11-1:0] node3212;
	wire [11-1:0] node3215;
	wire [11-1:0] node3218;
	wire [11-1:0] node3219;
	wire [11-1:0] node3220;
	wire [11-1:0] node3221;
	wire [11-1:0] node3222;
	wire [11-1:0] node3226;
	wire [11-1:0] node3227;
	wire [11-1:0] node3230;
	wire [11-1:0] node3233;
	wire [11-1:0] node3234;
	wire [11-1:0] node3236;
	wire [11-1:0] node3239;
	wire [11-1:0] node3241;
	wire [11-1:0] node3242;
	wire [11-1:0] node3246;
	wire [11-1:0] node3247;
	wire [11-1:0] node3248;
	wire [11-1:0] node3250;
	wire [11-1:0] node3253;
	wire [11-1:0] node3256;
	wire [11-1:0] node3257;
	wire [11-1:0] node3258;
	wire [11-1:0] node3261;
	wire [11-1:0] node3262;
	wire [11-1:0] node3265;
	wire [11-1:0] node3268;
	wire [11-1:0] node3271;
	wire [11-1:0] node3272;
	wire [11-1:0] node3273;
	wire [11-1:0] node3274;
	wire [11-1:0] node3275;
	wire [11-1:0] node3277;
	wire [11-1:0] node3278;
	wire [11-1:0] node3281;
	wire [11-1:0] node3282;
	wire [11-1:0] node3286;
	wire [11-1:0] node3287;
	wire [11-1:0] node3289;
	wire [11-1:0] node3292;
	wire [11-1:0] node3293;
	wire [11-1:0] node3295;
	wire [11-1:0] node3298;
	wire [11-1:0] node3300;
	wire [11-1:0] node3303;
	wire [11-1:0] node3304;
	wire [11-1:0] node3306;
	wire [11-1:0] node3307;
	wire [11-1:0] node3310;
	wire [11-1:0] node3313;
	wire [11-1:0] node3314;
	wire [11-1:0] node3315;
	wire [11-1:0] node3317;
	wire [11-1:0] node3320;
	wire [11-1:0] node3321;
	wire [11-1:0] node3324;
	wire [11-1:0] node3327;
	wire [11-1:0] node3329;
	wire [11-1:0] node3330;
	wire [11-1:0] node3334;
	wire [11-1:0] node3335;
	wire [11-1:0] node3336;
	wire [11-1:0] node3337;
	wire [11-1:0] node3338;
	wire [11-1:0] node3341;
	wire [11-1:0] node3344;
	wire [11-1:0] node3345;
	wire [11-1:0] node3348;
	wire [11-1:0] node3351;
	wire [11-1:0] node3352;
	wire [11-1:0] node3353;
	wire [11-1:0] node3354;
	wire [11-1:0] node3357;
	wire [11-1:0] node3361;
	wire [11-1:0] node3362;
	wire [11-1:0] node3364;
	wire [11-1:0] node3367;
	wire [11-1:0] node3370;
	wire [11-1:0] node3371;
	wire [11-1:0] node3372;
	wire [11-1:0] node3374;
	wire [11-1:0] node3377;
	wire [11-1:0] node3379;
	wire [11-1:0] node3382;
	wire [11-1:0] node3383;
	wire [11-1:0] node3385;
	wire [11-1:0] node3387;
	wire [11-1:0] node3390;
	wire [11-1:0] node3391;
	wire [11-1:0] node3395;
	wire [11-1:0] node3396;
	wire [11-1:0] node3397;
	wire [11-1:0] node3398;
	wire [11-1:0] node3400;
	wire [11-1:0] node3401;
	wire [11-1:0] node3405;
	wire [11-1:0] node3406;
	wire [11-1:0] node3407;
	wire [11-1:0] node3411;
	wire [11-1:0] node3413;
	wire [11-1:0] node3415;
	wire [11-1:0] node3418;
	wire [11-1:0] node3419;
	wire [11-1:0] node3420;
	wire [11-1:0] node3423;
	wire [11-1:0] node3426;
	wire [11-1:0] node3427;
	wire [11-1:0] node3428;
	wire [11-1:0] node3430;
	wire [11-1:0] node3433;
	wire [11-1:0] node3436;
	wire [11-1:0] node3439;
	wire [11-1:0] node3440;
	wire [11-1:0] node3441;
	wire [11-1:0] node3442;
	wire [11-1:0] node3443;
	wire [11-1:0] node3446;
	wire [11-1:0] node3448;
	wire [11-1:0] node3451;
	wire [11-1:0] node3452;
	wire [11-1:0] node3453;
	wire [11-1:0] node3457;
	wire [11-1:0] node3460;
	wire [11-1:0] node3461;
	wire [11-1:0] node3464;
	wire [11-1:0] node3465;
	wire [11-1:0] node3468;
	wire [11-1:0] node3471;
	wire [11-1:0] node3472;
	wire [11-1:0] node3473;
	wire [11-1:0] node3474;
	wire [11-1:0] node3479;
	wire [11-1:0] node3480;
	wire [11-1:0] node3481;
	wire [11-1:0] node3485;
	wire [11-1:0] node3487;
	wire [11-1:0] node3488;
	wire [11-1:0] node3492;
	wire [11-1:0] node3493;
	wire [11-1:0] node3494;
	wire [11-1:0] node3495;
	wire [11-1:0] node3496;
	wire [11-1:0] node3497;
	wire [11-1:0] node3498;
	wire [11-1:0] node3499;
	wire [11-1:0] node3500;
	wire [11-1:0] node3505;
	wire [11-1:0] node3506;
	wire [11-1:0] node3509;
	wire [11-1:0] node3510;
	wire [11-1:0] node3514;
	wire [11-1:0] node3515;
	wire [11-1:0] node3516;
	wire [11-1:0] node3519;
	wire [11-1:0] node3522;
	wire [11-1:0] node3523;
	wire [11-1:0] node3524;
	wire [11-1:0] node3527;
	wire [11-1:0] node3530;
	wire [11-1:0] node3533;
	wire [11-1:0] node3534;
	wire [11-1:0] node3535;
	wire [11-1:0] node3538;
	wire [11-1:0] node3539;
	wire [11-1:0] node3541;
	wire [11-1:0] node3544;
	wire [11-1:0] node3547;
	wire [11-1:0] node3548;
	wire [11-1:0] node3550;
	wire [11-1:0] node3552;
	wire [11-1:0] node3555;
	wire [11-1:0] node3556;
	wire [11-1:0] node3557;
	wire [11-1:0] node3561;
	wire [11-1:0] node3564;
	wire [11-1:0] node3565;
	wire [11-1:0] node3566;
	wire [11-1:0] node3567;
	wire [11-1:0] node3568;
	wire [11-1:0] node3571;
	wire [11-1:0] node3572;
	wire [11-1:0] node3576;
	wire [11-1:0] node3579;
	wire [11-1:0] node3580;
	wire [11-1:0] node3581;
	wire [11-1:0] node3585;
	wire [11-1:0] node3586;
	wire [11-1:0] node3587;
	wire [11-1:0] node3590;
	wire [11-1:0] node3593;
	wire [11-1:0] node3596;
	wire [11-1:0] node3597;
	wire [11-1:0] node3598;
	wire [11-1:0] node3600;
	wire [11-1:0] node3603;
	wire [11-1:0] node3605;
	wire [11-1:0] node3608;
	wire [11-1:0] node3609;
	wire [11-1:0] node3610;
	wire [11-1:0] node3614;
	wire [11-1:0] node3615;
	wire [11-1:0] node3618;
	wire [11-1:0] node3621;
	wire [11-1:0] node3622;
	wire [11-1:0] node3623;
	wire [11-1:0] node3624;
	wire [11-1:0] node3625;
	wire [11-1:0] node3626;
	wire [11-1:0] node3627;
	wire [11-1:0] node3631;
	wire [11-1:0] node3632;
	wire [11-1:0] node3636;
	wire [11-1:0] node3637;
	wire [11-1:0] node3640;
	wire [11-1:0] node3643;
	wire [11-1:0] node3644;
	wire [11-1:0] node3646;
	wire [11-1:0] node3649;
	wire [11-1:0] node3650;
	wire [11-1:0] node3651;
	wire [11-1:0] node3655;
	wire [11-1:0] node3658;
	wire [11-1:0] node3659;
	wire [11-1:0] node3660;
	wire [11-1:0] node3661;
	wire [11-1:0] node3662;
	wire [11-1:0] node3666;
	wire [11-1:0] node3669;
	wire [11-1:0] node3671;
	wire [11-1:0] node3674;
	wire [11-1:0] node3676;
	wire [11-1:0] node3677;
	wire [11-1:0] node3678;
	wire [11-1:0] node3682;
	wire [11-1:0] node3684;
	wire [11-1:0] node3687;
	wire [11-1:0] node3688;
	wire [11-1:0] node3689;
	wire [11-1:0] node3690;
	wire [11-1:0] node3692;
	wire [11-1:0] node3695;
	wire [11-1:0] node3697;
	wire [11-1:0] node3698;
	wire [11-1:0] node3701;
	wire [11-1:0] node3704;
	wire [11-1:0] node3705;
	wire [11-1:0] node3707;
	wire [11-1:0] node3710;
	wire [11-1:0] node3711;
	wire [11-1:0] node3714;
	wire [11-1:0] node3717;
	wire [11-1:0] node3718;
	wire [11-1:0] node3719;
	wire [11-1:0] node3721;
	wire [11-1:0] node3722;
	wire [11-1:0] node3726;
	wire [11-1:0] node3727;
	wire [11-1:0] node3728;
	wire [11-1:0] node3732;
	wire [11-1:0] node3733;
	wire [11-1:0] node3737;
	wire [11-1:0] node3738;
	wire [11-1:0] node3739;
	wire [11-1:0] node3740;
	wire [11-1:0] node3744;
	wire [11-1:0] node3745;
	wire [11-1:0] node3749;
	wire [11-1:0] node3752;
	wire [11-1:0] node3753;
	wire [11-1:0] node3754;
	wire [11-1:0] node3755;
	wire [11-1:0] node3756;
	wire [11-1:0] node3757;
	wire [11-1:0] node3758;
	wire [11-1:0] node3761;
	wire [11-1:0] node3763;
	wire [11-1:0] node3766;
	wire [11-1:0] node3767;
	wire [11-1:0] node3770;
	wire [11-1:0] node3771;
	wire [11-1:0] node3775;
	wire [11-1:0] node3777;
	wire [11-1:0] node3778;
	wire [11-1:0] node3779;
	wire [11-1:0] node3783;
	wire [11-1:0] node3786;
	wire [11-1:0] node3787;
	wire [11-1:0] node3788;
	wire [11-1:0] node3789;
	wire [11-1:0] node3790;
	wire [11-1:0] node3794;
	wire [11-1:0] node3795;
	wire [11-1:0] node3798;
	wire [11-1:0] node3801;
	wire [11-1:0] node3802;
	wire [11-1:0] node3806;
	wire [11-1:0] node3807;
	wire [11-1:0] node3808;
	wire [11-1:0] node3811;
	wire [11-1:0] node3814;
	wire [11-1:0] node3816;
	wire [11-1:0] node3819;
	wire [11-1:0] node3820;
	wire [11-1:0] node3821;
	wire [11-1:0] node3822;
	wire [11-1:0] node3823;
	wire [11-1:0] node3825;
	wire [11-1:0] node3829;
	wire [11-1:0] node3831;
	wire [11-1:0] node3832;
	wire [11-1:0] node3835;
	wire [11-1:0] node3838;
	wire [11-1:0] node3839;
	wire [11-1:0] node3841;
	wire [11-1:0] node3844;
	wire [11-1:0] node3845;
	wire [11-1:0] node3846;
	wire [11-1:0] node3850;
	wire [11-1:0] node3852;
	wire [11-1:0] node3855;
	wire [11-1:0] node3856;
	wire [11-1:0] node3857;
	wire [11-1:0] node3858;
	wire [11-1:0] node3859;
	wire [11-1:0] node3862;
	wire [11-1:0] node3865;
	wire [11-1:0] node3866;
	wire [11-1:0] node3870;
	wire [11-1:0] node3872;
	wire [11-1:0] node3875;
	wire [11-1:0] node3876;
	wire [11-1:0] node3877;
	wire [11-1:0] node3879;
	wire [11-1:0] node3883;
	wire [11-1:0] node3884;
	wire [11-1:0] node3887;
	wire [11-1:0] node3890;
	wire [11-1:0] node3891;
	wire [11-1:0] node3892;
	wire [11-1:0] node3893;
	wire [11-1:0] node3894;
	wire [11-1:0] node3895;
	wire [11-1:0] node3898;
	wire [11-1:0] node3901;
	wire [11-1:0] node3902;
	wire [11-1:0] node3905;
	wire [11-1:0] node3908;
	wire [11-1:0] node3909;
	wire [11-1:0] node3910;
	wire [11-1:0] node3914;
	wire [11-1:0] node3915;
	wire [11-1:0] node3918;
	wire [11-1:0] node3921;
	wire [11-1:0] node3922;
	wire [11-1:0] node3923;
	wire [11-1:0] node3925;
	wire [11-1:0] node3928;
	wire [11-1:0] node3929;
	wire [11-1:0] node3930;
	wire [11-1:0] node3933;
	wire [11-1:0] node3937;
	wire [11-1:0] node3938;
	wire [11-1:0] node3940;
	wire [11-1:0] node3943;
	wire [11-1:0] node3946;
	wire [11-1:0] node3947;
	wire [11-1:0] node3948;
	wire [11-1:0] node3949;
	wire [11-1:0] node3950;
	wire [11-1:0] node3953;
	wire [11-1:0] node3956;
	wire [11-1:0] node3957;
	wire [11-1:0] node3960;
	wire [11-1:0] node3963;
	wire [11-1:0] node3964;
	wire [11-1:0] node3965;
	wire [11-1:0] node3968;
	wire [11-1:0] node3971;
	wire [11-1:0] node3972;
	wire [11-1:0] node3976;
	wire [11-1:0] node3977;
	wire [11-1:0] node3978;
	wire [11-1:0] node3979;
	wire [11-1:0] node3982;
	wire [11-1:0] node3985;
	wire [11-1:0] node3986;
	wire [11-1:0] node3989;
	wire [11-1:0] node3990;
	wire [11-1:0] node3994;
	wire [11-1:0] node3995;
	wire [11-1:0] node3997;
	wire [11-1:0] node4000;
	wire [11-1:0] node4001;

	assign outp = (inp[1]) ? node2010 : node1;
		assign node1 = (inp[7]) ? node997 : node2;
			assign node2 = (inp[2]) ? node544 : node3;
				assign node3 = (inp[0]) ? node269 : node4;
					assign node4 = (inp[4]) ? node126 : node5;
						assign node5 = (inp[9]) ? node71 : node6;
							assign node6 = (inp[10]) ? node38 : node7;
								assign node7 = (inp[3]) ? node27 : node8;
									assign node8 = (inp[5]) ? node20 : node9;
										assign node9 = (inp[6]) ? node13 : node10;
											assign node10 = (inp[11]) ? 11'b01000001001 : 11'b01000001010;
											assign node13 = (inp[8]) ? node17 : node14;
												assign node14 = (inp[11]) ? 11'b01010000010 : 11'b01001100010;
												assign node17 = (inp[11]) ? 11'b01011101000 : 11'b01000101010;
										assign node20 = (inp[11]) ? node22 : 11'b01000111011;
											assign node22 = (inp[6]) ? 11'b01011011001 : node23;
												assign node23 = (inp[8]) ? 11'b01001011010 : 11'b01000011000;
									assign node27 = (inp[11]) ? node31 : node28;
										assign node28 = (inp[6]) ? 11'b11111001010 : 11'b11101101011;
										assign node31 = (inp[5]) ? node35 : node32;
											assign node32 = (inp[8]) ? 11'b11101111000 : 11'b11000010010;
											assign node35 = (inp[8]) ? 11'b11010001010 : 11'b11101101000;
								assign node38 = (inp[3]) ? node54 : node39;
									assign node39 = (inp[5]) ? node47 : node40;
										assign node40 = (inp[6]) ? 11'b11110101000 : node41;
											assign node41 = (inp[8]) ? node43 : 11'b11000101011;
												assign node43 = (inp[11]) ? 11'b11111101001 : 11'b11001101011;
										assign node47 = (inp[6]) ? 11'b11101011001 : node48;
											assign node48 = (inp[11]) ? 11'b11101111000 : node49;
												assign node49 = (inp[8]) ? 11'b11101111010 : 11'b11100111010;
									assign node54 = (inp[11]) ? node62 : node55;
										assign node55 = (inp[5]) ? node59 : node56;
											assign node56 = (inp[6]) ? 11'b01010100110 : 11'b01000101111;
											assign node59 = (inp[6]) ? 11'b01110011101 : 11'b01100111110;
										assign node62 = (inp[5]) ? node68 : node63;
											assign node63 = (inp[8]) ? node65 : 11'b01001111101;
												assign node65 = (inp[6]) ? 11'b01010111110 : 11'b01011111101;
											assign node68 = (inp[8]) ? 11'b01001101110 : 11'b01010101100;
							assign node71 = (inp[6]) ? node101 : node72;
								assign node72 = (inp[5]) ? node84 : node73;
									assign node73 = (inp[10]) ? node75 : 11'b11001101111;
										assign node75 = (inp[3]) ? node79 : node76;
											assign node76 = (inp[11]) ? 11'b11100111111 : 11'b11000111111;
											assign node79 = (inp[8]) ? node81 : 11'b01010111111;
												assign node81 = (inp[11]) ? 11'b01101111101 : 11'b01110111111;
									assign node84 = (inp[3]) ? node92 : node85;
										assign node85 = (inp[10]) ? node89 : node86;
											assign node86 = (inp[8]) ? 11'b01001101010 : 11'b01110101000;
											assign node89 = (inp[11]) ? 11'b11110101110 : 11'b11100101110;
										assign node92 = (inp[10]) ? node96 : node93;
											assign node93 = (inp[11]) ? 11'b11100111110 : 11'b11001111110;
											assign node96 = (inp[8]) ? 11'b01101101100 : node97;
												assign node97 = (inp[11]) ? 11'b01000101100 : 11'b01010101110;
								assign node101 = (inp[5]) ? node111 : node102;
									assign node102 = (inp[8]) ? node106 : node103;
										assign node103 = (inp[3]) ? 11'b11011100100 : 11'b01111111001;
										assign node106 = (inp[10]) ? node108 : 11'b11111001110;
											assign node108 = (inp[11]) ? 11'b11011011100 : 11'b11001011110;
									assign node111 = (inp[8]) ? node119 : node112;
										assign node112 = (inp[3]) ? node116 : node113;
											assign node113 = (inp[11]) ? 11'b01111001011 : 11'b01010011001;
											assign node116 = (inp[11]) ? 11'b11010011111 : 11'b11001111111;
										assign node119 = (inp[10]) ? node121 : 11'b11100111111;
											assign node121 = (inp[11]) ? node123 : 11'b11010101111;
												assign node123 = (inp[3]) ? 11'b01111101111 : 11'b11111101111;
						assign node126 = (inp[5]) ? node208 : node127;
							assign node127 = (inp[6]) ? node161 : node128;
								assign node128 = (inp[10]) ? node146 : node129;
									assign node129 = (inp[3]) ? node141 : node130;
										assign node130 = (inp[11]) ? node138 : node131;
											assign node131 = (inp[8]) ? node135 : node132;
												assign node132 = (inp[9]) ? 11'b01101001111 : 11'b01001001111;
												assign node135 = (inp[9]) ? 11'b01110001111 : 11'b01100101111;
											assign node138 = (inp[8]) ? 11'b01000011111 : 11'b01011011111;
										assign node141 = (inp[9]) ? 11'b11011011011 : node142;
											assign node142 = (inp[11]) ? 11'b11010101101 : 11'b11001001111;
									assign node146 = (inp[3]) ? node154 : node147;
										assign node147 = (inp[9]) ? node151 : node148;
											assign node148 = (inp[8]) ? 11'b11111011101 : 11'b11110011111;
											assign node151 = (inp[8]) ? 11'b11111011011 : 11'b11110011011;
										assign node154 = (inp[8]) ? node158 : node155;
											assign node155 = (inp[9]) ? 11'b01100011011 : 11'b01110011011;
											assign node158 = (inp[11]) ? 11'b01111011011 : 11'b01101011001;
								assign node161 = (inp[11]) ? node185 : node162;
									assign node162 = (inp[8]) ? node176 : node163;
										assign node163 = (inp[3]) ? node171 : node164;
											assign node164 = (inp[9]) ? node168 : node165;
												assign node165 = (inp[10]) ? 11'b11001010110 : 11'b01000100110;
												assign node168 = (inp[10]) ? 11'b11101000000 : 11'b01100000100;
											assign node171 = (inp[9]) ? node173 : 11'b01110000010;
												assign node173 = (inp[10]) ? 11'b01111010000 : 11'b11110010000;
										assign node176 = (inp[9]) ? node180 : node177;
											assign node177 = (inp[10]) ? 11'b11110011100 : 11'b11000001100;
											assign node180 = (inp[10]) ? 11'b11000101010 : node181;
												assign node181 = (inp[3]) ? 11'b11010111010 : 11'b01111101100;
									assign node185 = (inp[10]) ? node197 : node186;
										assign node186 = (inp[9]) ? node190 : node187;
											assign node187 = (inp[8]) ? 11'b11011001110 : 11'b11100101111;
											assign node190 = (inp[8]) ? node194 : node191;
												assign node191 = (inp[3]) ? 11'b11011011001 : 11'b01001011101;
												assign node194 = (inp[3]) ? 11'b11000011000 : 11'b01010011100;
										assign node197 = (inp[3]) ? node203 : node198;
											assign node198 = (inp[9]) ? 11'b11111111001 : node199;
												assign node199 = (inp[8]) ? 11'b11101011110 : 11'b11110111111;
											assign node203 = (inp[9]) ? node205 : 11'b01110011010;
												assign node205 = (inp[8]) ? 11'b01111111011 : 11'b01110011011;
							assign node208 = (inp[6]) ? node240 : node209;
								assign node209 = (inp[9]) ? node227 : node210;
									assign node210 = (inp[10]) ? node216 : node211;
										assign node211 = (inp[11]) ? 11'b11101111100 : node212;
											assign node212 = (inp[3]) ? 11'b11010111100 : 11'b01111111100;
										assign node216 = (inp[11]) ? node220 : node217;
											assign node217 = (inp[8]) ? 11'b01001011000 : 11'b01010011010;
											assign node220 = (inp[8]) ? node224 : node221;
												assign node221 = (inp[3]) ? 11'b01100001000 : 11'b11001001100;
												assign node224 = (inp[3]) ? 11'b01110101000 : 11'b11110101100;
									assign node227 = (inp[3]) ? node231 : node228;
										assign node228 = (inp[10]) ? 11'b11011001000 : 11'b01010001100;
										assign node231 = (inp[10]) ? node237 : node232;
											assign node232 = (inp[8]) ? 11'b11110001000 : node233;
												assign node233 = (inp[11]) ? 11'b11111001000 : 11'b11001001000;
											assign node237 = (inp[11]) ? 11'b01110001000 : 11'b01100001000;
								assign node240 = (inp[8]) ? node256 : node241;
									assign node241 = (inp[11]) ? node249 : node242;
										assign node242 = (inp[3]) ? node246 : node243;
											assign node243 = (inp[10]) ? 11'b11001011011 : 11'b01100111111;
											assign node246 = (inp[9]) ? 11'b11010101011 : 11'b01011111001;
										assign node249 = (inp[3]) ? node253 : node250;
											assign node250 = (inp[10]) ? 11'b11010101110 : 11'b01001111100;
											assign node253 = (inp[9]) ? 11'b11101101000 : 11'b01100101010;
									assign node256 = (inp[11]) ? node262 : node257;
										assign node257 = (inp[10]) ? 11'b11101011001 : node258;
											assign node258 = (inp[3]) ? 11'b11011011101 : 11'b01111011101;
										assign node262 = (inp[9]) ? 11'b01101001111 : node263;
											assign node263 = (inp[10]) ? 11'b11110101101 : node264;
												assign node264 = (inp[3]) ? 11'b11100111101 : 11'b01101111101;
					assign node269 = (inp[3]) ? node415 : node270;
						assign node270 = (inp[4]) ? node336 : node271;
							assign node271 = (inp[11]) ? node307 : node272;
								assign node272 = (inp[6]) ? node288 : node273;
									assign node273 = (inp[8]) ? node283 : node274;
										assign node274 = (inp[10]) ? node280 : node275;
											assign node275 = (inp[5]) ? 11'b01001101000 : node276;
												assign node276 = (inp[9]) ? 11'b01001101101 : 11'b01001101001;
											assign node280 = (inp[5]) ? 11'b01100101100 : 11'b01000101101;
										assign node283 = (inp[5]) ? node285 : 11'b01111111001;
											assign node285 = (inp[9]) ? 11'b01001111010 : 11'b01011101100;
									assign node288 = (inp[5]) ? node298 : node289;
										assign node289 = (inp[8]) ? node295 : node290;
											assign node290 = (inp[9]) ? 11'b01011100110 : node291;
												assign node291 = (inp[10]) ? 11'b01010100100 : 11'b01011100000;
											assign node295 = (inp[10]) ? 11'b01111001100 : 11'b01100001110;
										assign node298 = (inp[9]) ? node302 : node299;
											assign node299 = (inp[10]) ? 11'b01001101111 : 11'b01110101001;
											assign node302 = (inp[10]) ? node304 : 11'b01011101111;
												assign node304 = (inp[8]) ? 11'b01010111001 : 11'b01111111001;
								assign node307 = (inp[5]) ? node319 : node308;
									assign node308 = (inp[8]) ? node314 : node309;
										assign node309 = (inp[9]) ? 11'b01010101001 : node310;
											assign node310 = (inp[10]) ? 11'b01011111101 : 11'b01001111001;
										assign node314 = (inp[9]) ? 11'b01101101011 : node315;
											assign node315 = (inp[10]) ? 11'b01111111111 : 11'b01111111010;
									assign node319 = (inp[6]) ? node327 : node320;
										assign node320 = (inp[10]) ? node322 : 11'b01101011000;
											assign node322 = (inp[9]) ? 11'b01010101000 : node323;
												assign node323 = (inp[8]) ? 11'b01110011100 : 11'b01010111110;
										assign node327 = (inp[10]) ? node333 : node328;
											assign node328 = (inp[9]) ? 11'b01101011101 : node329;
												assign node329 = (inp[8]) ? 11'b01110011001 : 11'b01010011011;
											assign node333 = (inp[8]) ? 11'b01101111111 : 11'b01000011101;
							assign node336 = (inp[5]) ? node378 : node337;
								assign node337 = (inp[6]) ? node359 : node338;
									assign node338 = (inp[11]) ? node348 : node339;
										assign node339 = (inp[10]) ? node343 : node340;
											assign node340 = (inp[9]) ? 11'b01010011101 : 11'b01001001001;
											assign node343 = (inp[8]) ? 11'b01001011011 : node344;
												assign node344 = (inp[9]) ? 11'b01100011001 : 11'b01000011101;
										assign node348 = (inp[10]) ? node354 : node349;
											assign node349 = (inp[8]) ? 11'b01110111011 : node350;
												assign node350 = (inp[9]) ? 11'b01011001101 : 11'b01011011001;
											assign node354 = (inp[8]) ? node356 : 11'b01110001101;
												assign node356 = (inp[9]) ? 11'b01011001001 : 11'b01001001101;
									assign node359 = (inp[11]) ? node367 : node360;
										assign node360 = (inp[9]) ? node364 : node361;
											assign node361 = (inp[8]) ? 11'b01110001000 : 11'b01010100000;
											assign node364 = (inp[10]) ? 11'b01010111000 : 11'b01001111100;
										assign node367 = (inp[8]) ? node375 : node368;
											assign node368 = (inp[10]) ? node372 : node369;
												assign node369 = (inp[9]) ? 11'b01001001111 : 11'b01001111001;
												assign node372 = (inp[9]) ? 11'b01100001001 : 11'b01100101111;
											assign node375 = (inp[10]) ? 11'b01011001100 : 11'b01100011000;
								assign node378 = (inp[8]) ? node396 : node379;
									assign node379 = (inp[10]) ? node387 : node380;
										assign node380 = (inp[11]) ? node382 : 11'b01111011100;
											assign node382 = (inp[9]) ? node384 : 11'b01101011010;
												assign node384 = (inp[6]) ? 11'b01101101110 : 11'b01111001110;
										assign node387 = (inp[6]) ? node393 : node388;
											assign node388 = (inp[9]) ? node390 : 11'b01100001110;
												assign node390 = (inp[11]) ? 11'b01110001010 : 11'b01100011010;
											assign node393 = (inp[9]) ? 11'b01100101010 : 11'b01110101100;
									assign node396 = (inp[6]) ? node408 : node397;
										assign node397 = (inp[11]) ? node405 : node398;
											assign node398 = (inp[10]) ? node402 : node399;
												assign node399 = (inp[9]) ? 11'b01010011110 : 11'b01010101010;
												assign node402 = (inp[9]) ? 11'b01000011000 : 11'b01101011110;
											assign node405 = (inp[10]) ? 11'b01010101110 : 11'b01001001110;
										assign node408 = (inp[10]) ? node412 : node409;
											assign node409 = (inp[11]) ? 11'b01011001101 : 11'b01001011111;
											assign node412 = (inp[9]) ? 11'b01010011011 : 11'b01110011101;
						assign node415 = (inp[10]) ? node475 : node416;
							assign node416 = (inp[4]) ? node448 : node417;
								assign node417 = (inp[9]) ? node435 : node418;
									assign node418 = (inp[5]) ? node424 : node419;
										assign node419 = (inp[6]) ? node421 : 11'b01001101001;
											assign node421 = (inp[8]) ? 11'b01010101010 : 11'b01000000000;
										assign node424 = (inp[8]) ? node428 : node425;
											assign node425 = (inp[6]) ? 11'b01100001011 : 11'b01101101010;
											assign node428 = (inp[11]) ? node432 : node429;
												assign node429 = (inp[6]) ? 11'b01100101011 : 11'b01100001001;
												assign node432 = (inp[6]) ? 11'b01111101001 : 11'b01110001000;
									assign node435 = (inp[5]) ? node443 : node436;
										assign node436 = (inp[6]) ? node438 : 11'b01011111001;
											assign node438 = (inp[8]) ? node440 : 11'b01001110010;
												assign node440 = (inp[11]) ? 11'b01101011010 : 11'b01011011010;
										assign node443 = (inp[11]) ? 11'b01010011001 : node444;
											assign node444 = (inp[8]) ? 11'b01100111001 : 11'b01101111000;
								assign node448 = (inp[9]) ? node466 : node449;
									assign node449 = (inp[5]) ? node455 : node450;
										assign node450 = (inp[6]) ? 11'b01000011010 : node451;
											assign node451 = (inp[11]) ? 11'b01111011011 : 11'b01001011001;
										assign node455 = (inp[11]) ? node461 : node456;
											assign node456 = (inp[6]) ? node458 : 11'b01111011000;
												assign node458 = (inp[8]) ? 11'b01110011011 : 11'b01111111011;
											assign node461 = (inp[8]) ? 11'b01010111010 : node462;
												assign node462 = (inp[6]) ? 11'b01001111000 : 11'b01001011010;
									assign node466 = (inp[5]) ? node472 : node467;
										assign node467 = (inp[6]) ? node469 : 11'b01111001001;
											assign node469 = (inp[8]) ? 11'b01110101000 : 11'b01110001011;
										assign node472 = (inp[6]) ? 11'b01011001011 : 11'b01010001010;
							assign node475 = (inp[9]) ? node517 : node476;
								assign node476 = (inp[5]) ? node494 : node477;
									assign node477 = (inp[6]) ? node483 : node478;
										assign node478 = (inp[4]) ? 11'b01110001001 : node479;
											assign node479 = (inp[8]) ? 11'b01110101011 : 11'b01100101001;
										assign node483 = (inp[8]) ? node489 : node484;
											assign node484 = (inp[11]) ? 11'b01011001011 : node485;
												assign node485 = (inp[4]) ? 11'b01100000010 : 11'b01000100010;
											assign node489 = (inp[4]) ? 11'b01111101010 : node490;
												assign node490 = (inp[11]) ? 11'b01110101000 : 11'b01010001010;
									assign node494 = (inp[6]) ? node504 : node495;
										assign node495 = (inp[4]) ? node501 : node496;
											assign node496 = (inp[11]) ? 11'b01101101000 : node497;
												assign node497 = (inp[8]) ? 11'b01011101000 : 11'b01000101000;
											assign node501 = (inp[11]) ? 11'b01001001010 : 11'b01101001010;
										assign node504 = (inp[4]) ? node512 : node505;
											assign node505 = (inp[8]) ? node509 : node506;
												assign node506 = (inp[11]) ? 11'b01111001001 : 11'b01000001011;
												assign node509 = (inp[11]) ? 11'b01100101011 : 11'b01011101011;
											assign node512 = (inp[8]) ? node514 : 11'b01010101000;
												assign node514 = (inp[11]) ? 11'b01001001001 : 11'b01100001001;
								assign node517 = (inp[5]) ? node531 : node518;
									assign node518 = (inp[6]) ? node520 : 11'b01000101001;
										assign node520 = (inp[11]) ? node526 : node521;
											assign node521 = (inp[8]) ? node523 : 11'b01001000000;
												assign node523 = (inp[4]) ? 11'b01001101010 : 11'b01001001000;
											assign node526 = (inp[4]) ? node528 : 11'b01011101001;
												assign node528 = (inp[8]) ? 11'b01001101001 : 11'b01000001001;
									assign node531 = (inp[11]) ? node541 : node532;
										assign node532 = (inp[6]) ? node536 : node533;
											assign node533 = (inp[8]) ? 11'b01011101010 : 11'b01010101000;
											assign node536 = (inp[4]) ? 11'b01001001011 : node537;
												assign node537 = (inp[8]) ? 11'b01011001011 : 11'b01010101001;
										assign node541 = (inp[6]) ? 11'b01001101010 : 11'b01000101010;
				assign node544 = (inp[0]) ? node770 : node545;
					assign node545 = (inp[8]) ? node653 : node546;
						assign node546 = (inp[11]) ? node598 : node547;
							assign node547 = (inp[5]) ? node577 : node548;
								assign node548 = (inp[10]) ? node562 : node549;
									assign node549 = (inp[4]) ? node559 : node550;
										assign node550 = (inp[3]) ? node554 : node551;
											assign node551 = (inp[9]) ? 11'b01100001001 : 11'b01101001011;
											assign node554 = (inp[9]) ? 11'b11101101110 : node555;
												assign node555 = (inp[6]) ? 11'b11101001011 : 11'b11101001010;
										assign node559 = (inp[6]) ? 11'b11100101100 : 11'b01100100101;
									assign node562 = (inp[4]) ? node574 : node563;
										assign node563 = (inp[9]) ? node571 : node564;
											assign node564 = (inp[3]) ? node568 : node565;
												assign node565 = (inp[6]) ? 11'b11110001011 : 11'b11110001010;
												assign node568 = (inp[6]) ? 11'b01110001101 : 11'b01110001110;
											assign node571 = (inp[3]) ? 11'b01110111110 : 11'b11110110111;
										assign node574 = (inp[6]) ? 11'b01011101010 : 11'b01000100001;
								assign node577 = (inp[6]) ? node589 : node578;
									assign node578 = (inp[4]) ? 11'b01111110100 : node579;
										assign node579 = (inp[9]) ? node585 : node580;
											assign node580 = (inp[10]) ? node582 : 11'b01100010011;
												assign node582 = (inp[3]) ? 11'b01001010101 : 11'b11011010011;
											assign node585 = (inp[10]) ? 11'b11000000101 : 11'b11110010101;
									assign node589 = (inp[9]) ? 11'b01100001100 : node590;
										assign node590 = (inp[10]) ? node594 : node591;
											assign node591 = (inp[4]) ? 11'b01111011100 : 11'b01100111010;
											assign node594 = (inp[4]) ? 11'b01100011000 : 11'b01011011100;
							assign node598 = (inp[5]) ? node624 : node599;
								assign node599 = (inp[6]) ? node613 : node600;
									assign node600 = (inp[9]) ? node606 : node601;
										assign node601 = (inp[10]) ? 11'b01100010111 : node602;
											assign node602 = (inp[3]) ? 11'b11111010011 : 11'b01100000011;
										assign node606 = (inp[3]) ? 11'b11011100111 : node607;
											assign node607 = (inp[10]) ? node609 : 11'b01010010011;
												assign node609 = (inp[4]) ? 11'b11011010011 : 11'b11001110101;
									assign node613 = (inp[4]) ? node617 : node614;
										assign node614 = (inp[3]) ? 11'b11011001110 : 11'b01011011000;
										assign node617 = (inp[9]) ? node621 : node618;
											assign node618 = (inp[3]) ? 11'b11011101100 : 11'b11011111110;
											assign node621 = (inp[3]) ? 11'b11110111000 : 11'b01100111100;
								assign node624 = (inp[6]) ? node634 : node625;
									assign node625 = (inp[4]) ? node631 : node626;
										assign node626 = (inp[9]) ? 11'b01110000110 : node627;
											assign node627 = (inp[3]) ? 11'b11011000000 : 11'b01101010000;
										assign node631 = (inp[10]) ? 11'b11101100000 : 11'b11001100000;
									assign node634 = (inp[4]) ? node640 : node635;
										assign node635 = (inp[10]) ? 11'b01101100111 : node636;
											assign node636 = (inp[3]) ? 11'b11010100001 : 11'b01110110001;
										assign node640 = (inp[10]) ? node648 : node641;
											assign node641 = (inp[3]) ? node645 : node642;
												assign node642 = (inp[9]) ? 11'b01111000111 : 11'b01101010111;
												assign node645 = (inp[9]) ? 11'b11011000011 : 11'b11001010101;
											assign node648 = (inp[3]) ? node650 : 11'b11100000101;
												assign node650 = (inp[9]) ? 11'b01010000001 : 11'b01000000011;
						assign node653 = (inp[5]) ? node713 : node654;
							assign node654 = (inp[10]) ? node682 : node655;
								assign node655 = (inp[3]) ? node671 : node656;
									assign node656 = (inp[4]) ? node668 : node657;
										assign node657 = (inp[11]) ? node665 : node658;
											assign node658 = (inp[9]) ? node662 : node659;
												assign node659 = (inp[6]) ? 11'b01100000011 : 11'b01100100010;
												assign node662 = (inp[6]) ? 11'b01110100001 : 11'b01110000010;
											assign node665 = (inp[6]) ? 11'b01110000001 : 11'b01101100001;
										assign node668 = (inp[6]) ? 11'b01011100101 : 11'b01000000100;
									assign node671 = (inp[4]) ? node677 : node672;
										assign node672 = (inp[11]) ? node674 : 11'b11000000100;
											assign node674 = (inp[6]) ? 11'b11000000101 : 11'b11010000111;
										assign node677 = (inp[11]) ? node679 : 11'b11100110011;
											assign node679 = (inp[6]) ? 11'b11110100100 : 11'b11101000101;
								assign node682 = (inp[3]) ? node698 : node683;
									assign node683 = (inp[6]) ? node689 : node684;
										assign node684 = (inp[11]) ? 11'b11000100001 : node685;
											assign node685 = (inp[9]) ? 11'b11111100011 : 11'b11111000010;
										assign node689 = (inp[4]) ? node695 : node690;
											assign node690 = (inp[9]) ? node692 : 11'b11101100001;
												assign node692 = (inp[11]) ? 11'b11101110110 : 11'b11111110111;
											assign node695 = (inp[11]) ? 11'b11010110000 : 11'b11000110111;
									assign node698 = (inp[4]) ? node710 : node699;
										assign node699 = (inp[11]) ? node705 : node700;
											assign node700 = (inp[9]) ? node702 : 11'b01000000110;
												assign node702 = (inp[6]) ? 11'b01011110101 : 11'b01011010100;
											assign node705 = (inp[6]) ? 11'b01100010111 : node706;
												assign node706 = (inp[9]) ? 11'b01001010111 : 11'b01111010101;
										assign node710 = (inp[9]) ? 11'b01010110011 : 11'b01101100011;
							assign node713 = (inp[10]) ? node747 : node714;
								assign node714 = (inp[3]) ? node726 : node715;
									assign node715 = (inp[4]) ? node719 : node716;
										assign node716 = (inp[9]) ? 11'b01110100010 : 11'b01100110010;
										assign node719 = (inp[6]) ? node721 : 11'b01010010101;
											assign node721 = (inp[11]) ? node723 : 11'b01011110110;
												assign node723 = (inp[9]) ? 11'b01011000110 : 11'b01010010110;
									assign node726 = (inp[9]) ? node740 : node727;
										assign node727 = (inp[4]) ? node735 : node728;
											assign node728 = (inp[11]) ? node732 : node729;
												assign node729 = (inp[6]) ? 11'b11101010000 : 11'b11111110011;
												assign node732 = (inp[6]) ? 11'b11111100010 : 11'b11110100010;
											assign node735 = (inp[11]) ? 11'b11010010110 : node736;
												assign node736 = (inp[6]) ? 11'b11110010110 : 11'b11101010111;
										assign node740 = (inp[4]) ? 11'b11010100010 : node741;
											assign node741 = (inp[11]) ? node743 : 11'b11100010100;
												assign node743 = (inp[6]) ? 11'b11011010110 : 11'b11010110100;
								assign node747 = (inp[3]) ? node763 : node748;
									assign node748 = (inp[4]) ? node752 : node749;
										assign node749 = (inp[9]) ? 11'b11101000100 : 11'b11001110001;
										assign node752 = (inp[9]) ? node758 : node753;
											assign node753 = (inp[6]) ? node755 : 11'b11111000111;
												assign node755 = (inp[11]) ? 11'b11010000100 : 11'b11110000100;
											assign node758 = (inp[11]) ? node760 : 11'b11010110000;
												assign node760 = (inp[6]) ? 11'b11010000000 : 11'b11000000000;
									assign node763 = (inp[11]) ? node765 : 11'b01000010110;
										assign node765 = (inp[4]) ? node767 : 11'b01011000100;
											assign node767 = (inp[6]) ? 11'b01011000000 : 11'b01011000010;
					assign node770 = (inp[3]) ? node890 : node771;
						assign node771 = (inp[5]) ? node825 : node772;
							assign node772 = (inp[4]) ? node802 : node773;
								assign node773 = (inp[10]) ? node785 : node774;
									assign node774 = (inp[8]) ? node778 : node775;
										assign node775 = (inp[6]) ? 11'b01101011100 : 11'b01110010101;
										assign node778 = (inp[11]) ? node782 : node779;
											assign node779 = (inp[9]) ? 11'b01100100101 : 11'b01110000001;
											assign node782 = (inp[9]) ? 11'b01010010111 : 11'b01110110011;
									assign node785 = (inp[9]) ? node793 : node786;
										assign node786 = (inp[11]) ? node788 : 11'b01101000100;
											assign node788 = (inp[8]) ? node790 : 11'b01001010101;
												assign node790 = (inp[6]) ? 11'b01111010101 : 11'b01101010111;
										assign node793 = (inp[8]) ? node797 : node794;
											assign node794 = (inp[11]) ? 11'b01001100011 : 11'b01010110001;
											assign node797 = (inp[11]) ? 11'b01111100000 : node798;
												assign node798 = (inp[6]) ? 11'b01101110011 : 11'b01111010010;
								assign node802 = (inp[6]) ? node814 : node803;
									assign node803 = (inp[10]) ? node811 : node804;
										assign node804 = (inp[9]) ? node808 : node805;
											assign node805 = (inp[11]) ? 11'b01010110011 : 11'b01001100011;
											assign node808 = (inp[11]) ? 11'b01000100101 : 11'b01000110101;
										assign node811 = (inp[8]) ? 11'b01010100001 : 11'b01110010011;
									assign node814 = (inp[8]) ? node820 : node815;
										assign node815 = (inp[10]) ? 11'b01001111100 : node816;
											assign node816 = (inp[9]) ? 11'b01010101110 : 11'b01010101010;
										assign node820 = (inp[11]) ? 11'b01100110010 : node821;
											assign node821 = (inp[9]) ? 11'b01011010111 : 11'b01110110101;
							assign node825 = (inp[8]) ? node861 : node826;
								assign node826 = (inp[6]) ? node844 : node827;
									assign node827 = (inp[4]) ? node835 : node828;
										assign node828 = (inp[9]) ? node832 : node829;
											assign node829 = (inp[10]) ? 11'b01000010110 : 11'b01011010010;
											assign node832 = (inp[11]) ? 11'b01110000000 : 11'b01101110010;
										assign node835 = (inp[10]) ? node841 : node836;
											assign node836 = (inp[9]) ? node838 : 11'b01110100010;
												assign node838 = (inp[11]) ? 11'b01111100110 : 11'b01101110100;
											assign node841 = (inp[9]) ? 11'b01110100010 : 11'b01100100110;
									assign node844 = (inp[11]) ? node854 : node845;
										assign node845 = (inp[9]) ? node851 : node846;
											assign node846 = (inp[10]) ? 11'b01101001110 : node847;
												assign node847 = (inp[4]) ? 11'b01101001000 : 11'b01010101000;
											assign node851 = (inp[4]) ? 11'b01111110111 : 11'b01110011010;
										assign node854 = (inp[10]) ? node858 : node855;
											assign node855 = (inp[4]) ? 11'b01111010001 : 11'b01000110011;
											assign node858 = (inp[4]) ? 11'b01100000011 : 11'b01100100001;
								assign node861 = (inp[6]) ? node877 : node862;
									assign node862 = (inp[11]) ? node870 : node863;
										assign node863 = (inp[4]) ? 11'b01010010111 : node864;
											assign node864 = (inp[9]) ? node866 : 11'b01000100111;
												assign node866 = (inp[10]) ? 11'b01001010001 : 11'b01101000111;
										assign node870 = (inp[4]) ? node874 : node871;
											assign node871 = (inp[10]) ? 11'b01111110100 : 11'b01010110110;
											assign node874 = (inp[10]) ? 11'b01010000100 : 11'b01011010000;
									assign node877 = (inp[10]) ? node883 : node878;
										assign node878 = (inp[9]) ? node880 : 11'b01101110000;
											assign node880 = (inp[11]) ? 11'b01001000100 : 11'b01001110100;
										assign node883 = (inp[9]) ? node885 : 11'b01010000110;
											assign node885 = (inp[11]) ? node887 : 11'b01000110010;
												assign node887 = (inp[4]) ? 11'b01000000010 : 11'b01001000010;
						assign node890 = (inp[4]) ? node946 : node891;
							assign node891 = (inp[9]) ? node921 : node892;
								assign node892 = (inp[8]) ? node908 : node893;
									assign node893 = (inp[5]) ? node899 : node894;
										assign node894 = (inp[10]) ? node896 : 11'b01010001000;
											assign node896 = (inp[6]) ? 11'b01101001010 : 11'b01000001000;
										assign node899 = (inp[10]) ? node903 : node900;
											assign node900 = (inp[6]) ? 11'b01110101010 : 11'b01110000010;
											assign node903 = (inp[11]) ? node905 : 11'b01001000011;
												assign node905 = (inp[6]) ? 11'b01111100001 : 11'b01111000010;
									assign node908 = (inp[11]) ? node916 : node909;
										assign node909 = (inp[10]) ? node911 : 11'b01111000010;
											assign node911 = (inp[6]) ? 11'b01010000000 : node912;
												assign node912 = (inp[5]) ? 11'b01010100011 : 11'b01010000000;
										assign node916 = (inp[10]) ? node918 : 11'b01000100011;
											assign node918 = (inp[6]) ? 11'b01110000001 : 11'b01111000011;
								assign node921 = (inp[10]) ? node937 : node922;
									assign node922 = (inp[8]) ? node930 : node923;
										assign node923 = (inp[5]) ? node927 : node924;
											assign node924 = (inp[11]) ? 11'b01111011000 : 11'b01011111000;
											assign node927 = (inp[11]) ? 11'b01000110011 : 11'b01110011000;
										assign node930 = (inp[5]) ? node934 : node931;
											assign node931 = (inp[11]) ? 11'b01110010001 : 11'b01001010010;
											assign node934 = (inp[11]) ? 11'b01001010010 : 11'b01111010010;
									assign node937 = (inp[11]) ? node943 : node938;
										assign node938 = (inp[5]) ? node940 : 11'b01000000010;
											assign node940 = (inp[6]) ? 11'b01011001010 : 11'b01011100010;
										assign node943 = (inp[6]) ? 11'b01011100000 : 11'b01011000001;
							assign node946 = (inp[10]) ? node972 : node947;
								assign node947 = (inp[9]) ? node959 : node948;
									assign node948 = (inp[8]) ? node954 : node949;
										assign node949 = (inp[6]) ? 11'b01101111000 : node950;
											assign node950 = (inp[11]) ? 11'b01101110011 : 11'b01011110011;
										assign node954 = (inp[6]) ? 11'b01100010010 : node955;
											assign node955 = (inp[11]) ? 11'b01100010011 : 11'b01101010001;
									assign node959 = (inp[5]) ? node967 : node960;
										assign node960 = (inp[11]) ? node964 : node961;
											assign node961 = (inp[8]) ? 11'b01100100001 : 11'b01111000011;
											assign node964 = (inp[8]) ? 11'b01101100001 : 11'b01100100001;
										assign node967 = (inp[8]) ? node969 : 11'b01001000011;
											assign node969 = (inp[11]) ? 11'b01000000010 : 11'b01001100010;
								assign node972 = (inp[8]) ? node984 : node973;
									assign node973 = (inp[9]) ? node979 : node974;
										assign node974 = (inp[6]) ? 11'b01010101000 : node975;
											assign node975 = (inp[5]) ? 11'b01010100010 : 11'b01010100011;
										assign node979 = (inp[5]) ? node981 : 11'b01000000001;
											assign node981 = (inp[11]) ? 11'b01000000001 : 11'b01000100011;
									assign node984 = (inp[11]) ? node994 : node985;
										assign node985 = (inp[9]) ? node991 : node986;
											assign node986 = (inp[5]) ? node988 : 11'b01111000011;
												assign node988 = (inp[6]) ? 11'b01101100000 : 11'b01100000011;
											assign node991 = (inp[6]) ? 11'b01000000011 : 11'b01001100011;
										assign node994 = (inp[6]) ? 11'b01001100000 : 11'b01001100011;
			assign node997 = (inp[6]) ? node1491 : node998;
				assign node998 = (inp[2]) ? node1266 : node999;
					assign node999 = (inp[8]) ? node1123 : node1000;
						assign node1000 = (inp[5]) ? node1060 : node1001;
							assign node1001 = (inp[0]) ? node1033 : node1002;
								assign node1002 = (inp[11]) ? node1018 : node1003;
									assign node1003 = (inp[10]) ? node1011 : node1004;
										assign node1004 = (inp[9]) ? node1008 : node1005;
											assign node1005 = (inp[4]) ? 11'b11010100111 : 11'b11011100011;
											assign node1008 = (inp[4]) ? 11'b01111000111 : 11'b01010100011;
										assign node1011 = (inp[3]) ? node1015 : node1012;
											assign node1012 = (inp[9]) ? 11'b11011110101 : 11'b11011100001;
											assign node1015 = (inp[9]) ? 11'b01011110101 : 11'b01010100101;
									assign node1018 = (inp[4]) ? node1026 : node1019;
										assign node1019 = (inp[3]) ? node1023 : node1020;
											assign node1020 = (inp[10]) ? 11'b11111110101 : 11'b01110010011;
											assign node1023 = (inp[10]) ? 11'b01001110111 : 11'b11111100111;
										assign node1026 = (inp[10]) ? node1030 : node1027;
											assign node1027 = (inp[9]) ? 11'b01001110111 : 11'b11100100101;
											assign node1030 = (inp[3]) ? 11'b01101110011 : 11'b11100110001;
								assign node1033 = (inp[4]) ? node1043 : node1034;
									assign node1034 = (inp[3]) ? node1038 : node1035;
										assign node1035 = (inp[9]) ? 11'b01000100101 : 11'b01001100001;
										assign node1038 = (inp[9]) ? 11'b01101110011 : node1039;
											assign node1039 = (inp[11]) ? 11'b01001000011 : 11'b01001100011;
									assign node1043 = (inp[11]) ? node1055 : node1044;
										assign node1044 = (inp[3]) ? node1050 : node1045;
											assign node1045 = (inp[10]) ? node1047 : 11'b01101010101;
												assign node1047 = (inp[9]) ? 11'b01100010011 : 11'b01001010111;
											assign node1050 = (inp[10]) ? 11'b01101000001 : node1051;
												assign node1051 = (inp[9]) ? 11'b01100000011 : 11'b01000110011;
										assign node1055 = (inp[9]) ? 11'b01110100011 : node1056;
											assign node1056 = (inp[3]) ? 11'b01110110011 : 11'b01010110001;
							assign node1060 = (inp[0]) ? node1088 : node1061;
								assign node1061 = (inp[9]) ? node1073 : node1062;
									assign node1062 = (inp[11]) ? node1070 : node1063;
										assign node1063 = (inp[4]) ? node1065 : 11'b01011010011;
											assign node1065 = (inp[10]) ? node1067 : 11'b11100010101;
												assign node1067 = (inp[3]) ? 11'b01001110010 : 11'b11000000111;
										assign node1070 = (inp[4]) ? 11'b11110010110 : 11'b11111100000;
									assign node1073 = (inp[11]) ? node1081 : node1074;
										assign node1074 = (inp[10]) ? node1078 : node1075;
											assign node1075 = (inp[3]) ? 11'b11011100000 : 11'b01101110100;
											assign node1078 = (inp[3]) ? 11'b01110100010 : 11'b11010110010;
										assign node1081 = (inp[4]) ? node1085 : node1082;
											assign node1082 = (inp[3]) ? 11'b11000110110 : 11'b01100100000;
											assign node1085 = (inp[10]) ? 11'b01100000000 : 11'b11101000010;
								assign node1088 = (inp[3]) ? node1104 : node1089;
									assign node1089 = (inp[11]) ? node1097 : node1090;
										assign node1090 = (inp[10]) ? node1094 : node1091;
											assign node1091 = (inp[9]) ? 11'b01000000111 : 11'b01110000011;
											assign node1094 = (inp[9]) ? 11'b01100110000 : 11'b01010010101;
										assign node1097 = (inp[4]) ? node1099 : 11'b01110110110;
											assign node1099 = (inp[10]) ? node1101 : 11'b01101010000;
												assign node1101 = (inp[9]) ? 11'b01110000010 : 11'b01100000110;
									assign node1104 = (inp[11]) ? node1112 : node1105;
										assign node1105 = (inp[10]) ? node1107 : 11'b01101010011;
											assign node1107 = (inp[4]) ? 11'b01000100010 : node1108;
												assign node1108 = (inp[9]) ? 11'b01011000001 : 11'b01000000001;
										assign node1112 = (inp[10]) ? node1118 : node1113;
											assign node1113 = (inp[9]) ? node1115 : 11'b01000010000;
												assign node1115 = (inp[4]) ? 11'b01011000000 : 11'b01010110000;
											assign node1118 = (inp[9]) ? 11'b01001000010 : node1119;
												assign node1119 = (inp[4]) ? 11'b01011000010 : 11'b01110100010;
						assign node1123 = (inp[5]) ? node1199 : node1124;
							assign node1124 = (inp[11]) ? node1162 : node1125;
								assign node1125 = (inp[0]) ? node1145 : node1126;
									assign node1126 = (inp[10]) ? node1138 : node1127;
										assign node1127 = (inp[9]) ? node1133 : node1128;
											assign node1128 = (inp[3]) ? node1130 : 11'b01010000010;
												assign node1130 = (inp[4]) ? 11'b11011100100 : 11'b11111100010;
											assign node1133 = (inp[3]) ? 11'b11100100100 : node1134;
												assign node1134 = (inp[4]) ? 11'b01100100100 : 11'b01000100010;
										assign node1138 = (inp[9]) ? node1142 : node1139;
											assign node1139 = (inp[3]) ? 11'b01000100010 : 11'b11110110100;
											assign node1142 = (inp[3]) ? 11'b01110010010 : 11'b11011000010;
									assign node1145 = (inp[3]) ? node1153 : node1146;
										assign node1146 = (inp[4]) ? node1150 : node1147;
											assign node1147 = (inp[10]) ? 11'b01101100110 : 11'b01110100100;
											assign node1150 = (inp[9]) ? 11'b01001010000 : 11'b01100110100;
										assign node1153 = (inp[4]) ? node1159 : node1154;
											assign node1154 = (inp[9]) ? 11'b01010110010 : node1155;
												assign node1155 = (inp[10]) ? 11'b01011100000 : 11'b01001100010;
											assign node1159 = (inp[10]) ? 11'b01110100000 : 11'b01111000010;
								assign node1162 = (inp[4]) ? node1176 : node1163;
									assign node1163 = (inp[3]) ? node1169 : node1164;
										assign node1164 = (inp[0]) ? node1166 : 11'b11101000010;
											assign node1166 = (inp[10]) ? 11'b01100000010 : 11'b01100010010;
										assign node1169 = (inp[10]) ? node1173 : node1170;
											assign node1170 = (inp[0]) ? 11'b01100010000 : 11'b11110010000;
											assign node1173 = (inp[9]) ? 11'b01110010100 : 11'b01111000010;
									assign node1176 = (inp[0]) ? node1186 : node1177;
										assign node1177 = (inp[10]) ? node1183 : node1178;
											assign node1178 = (inp[9]) ? node1180 : 11'b10001101111;
												assign node1180 = (inp[3]) ? 11'b10000111001 : 11'b00010111111;
											assign node1183 = (inp[9]) ? 11'b10101111001 : 11'b10101111101;
										assign node1186 = (inp[10]) ? node1192 : node1187;
											assign node1187 = (inp[3]) ? node1189 : 11'b00100101101;
												assign node1189 = (inp[9]) ? 11'b00111101011 : 11'b00111111001;
											assign node1192 = (inp[9]) ? node1196 : node1193;
												assign node1193 = (inp[3]) ? 11'b00000101001 : 11'b00000101111;
												assign node1196 = (inp[3]) ? 11'b00001101001 : 11'b00011101011;
							assign node1199 = (inp[0]) ? node1237 : node1200;
								assign node1200 = (inp[9]) ? node1222 : node1201;
									assign node1201 = (inp[4]) ? node1215 : node1202;
										assign node1202 = (inp[10]) ? node1210 : node1203;
											assign node1203 = (inp[3]) ? node1207 : node1204;
												assign node1204 = (inp[11]) ? 11'b00011111011 : 11'b00010111011;
												assign node1207 = (inp[11]) ? 11'b10001101001 : 11'b10010111001;
											assign node1210 = (inp[3]) ? node1212 : 11'b10110111001;
												assign node1212 = (inp[11]) ? 11'b00010101111 : 11'b00101011111;
										assign node1215 = (inp[3]) ? node1219 : node1216;
											assign node1216 = (inp[11]) ? 11'b10101001111 : 11'b10011001111;
											assign node1219 = (inp[10]) ? 11'b00011011001 : 11'b10001011111;
									assign node1222 = (inp[3]) ? node1230 : node1223;
										assign node1223 = (inp[10]) ? node1227 : node1224;
											assign node1224 = (inp[4]) ? 11'b00111001101 : 11'b00001011001;
											assign node1227 = (inp[11]) ? 11'b10100001001 : 11'b10100011001;
										assign node1230 = (inp[4]) ? node1234 : node1231;
											assign node1231 = (inp[11]) ? 11'b00100101111 : 11'b00110001111;
											assign node1234 = (inp[10]) ? 11'b00100001001 : 11'b10110001011;
								assign node1237 = (inp[9]) ? node1249 : node1238;
									assign node1238 = (inp[11]) ? node1244 : node1239;
										assign node1239 = (inp[10]) ? node1241 : 11'b00100101011;
											assign node1241 = (inp[4]) ? 11'b00100001011 : 11'b00010101101;
										assign node1244 = (inp[4]) ? node1246 : 11'b00110101011;
											assign node1246 = (inp[3]) ? 11'b00010111001 : 11'b00000111011;
									assign node1249 = (inp[11]) ? node1257 : node1250;
										assign node1250 = (inp[10]) ? node1254 : node1251;
											assign node1251 = (inp[4]) ? 11'b00010001001 : 11'b00101011001;
											assign node1254 = (inp[4]) ? 11'b00001111011 : 11'b00000011001;
										assign node1257 = (inp[4]) ? node1263 : node1258;
											assign node1258 = (inp[10]) ? 11'b00011101001 : node1259;
												assign node1259 = (inp[3]) ? 11'b00011111011 : 11'b00001111111;
											assign node1263 = (inp[10]) ? 11'b00010001011 : 11'b00001001101;
					assign node1266 = (inp[0]) ? node1396 : node1267;
						assign node1267 = (inp[4]) ? node1335 : node1268;
							assign node1268 = (inp[9]) ? node1304 : node1269;
								assign node1269 = (inp[10]) ? node1293 : node1270;
									assign node1270 = (inp[3]) ? node1282 : node1271;
										assign node1271 = (inp[5]) ? node1275 : node1272;
											assign node1272 = (inp[8]) ? 11'b00111101001 : 11'b00110101010;
											assign node1275 = (inp[11]) ? node1279 : node1276;
												assign node1276 = (inp[8]) ? 11'b00111011011 : 11'b00110111010;
												assign node1279 = (inp[8]) ? 11'b00110111010 : 11'b00111011000;
										assign node1282 = (inp[11]) ? node1288 : node1283;
											assign node1283 = (inp[5]) ? node1285 : 11'b10111001011;
												assign node1285 = (inp[8]) ? 11'b10101011001 : 11'b10110111000;
											assign node1288 = (inp[5]) ? 11'b10001001010 : node1289;
												assign node1289 = (inp[8]) ? 11'b10000111011 : 11'b10100111000;
									assign node1293 = (inp[3]) ? node1299 : node1294;
										assign node1294 = (inp[5]) ? 11'b10110111000 : node1295;
											assign node1295 = (inp[8]) ? 11'b10101001001 : 11'b10101001000;
										assign node1299 = (inp[11]) ? node1301 : 11'b00001011101;
											assign node1301 = (inp[8]) ? 11'b00101001110 : 11'b00110001100;
								assign node1304 = (inp[10]) ? node1318 : node1305;
									assign node1305 = (inp[11]) ? node1313 : node1306;
										assign node1306 = (inp[3]) ? node1310 : node1307;
											assign node1307 = (inp[5]) ? 11'b00100011001 : 11'b00110001011;
											assign node1310 = (inp[5]) ? 11'b10110011111 : 11'b10110001101;
										assign node1313 = (inp[5]) ? node1315 : 11'b10000001100;
											assign node1315 = (inp[8]) ? 11'b10001011110 : 11'b10111111111;
									assign node1318 = (inp[3]) ? node1324 : node1319;
										assign node1319 = (inp[11]) ? node1321 : 11'b10101111110;
											assign node1321 = (inp[8]) ? 11'b10101111101 : 11'b10001101101;
										assign node1324 = (inp[8]) ? node1330 : node1325;
											assign node1325 = (inp[5]) ? 11'b00110101100 : node1326;
												assign node1326 = (inp[11]) ? 11'b00111011110 : 11'b00101111110;
											assign node1330 = (inp[5]) ? 11'b00000001100 : node1331;
												assign node1331 = (inp[11]) ? 11'b00010111111 : 11'b00000011101;
							assign node1335 = (inp[9]) ? node1367 : node1336;
								assign node1336 = (inp[3]) ? node1348 : node1337;
									assign node1337 = (inp[5]) ? node1345 : node1338;
										assign node1338 = (inp[11]) ? node1342 : node1339;
											assign node1339 = (inp[10]) ? 11'b10011011101 : 11'b00011001101;
											assign node1342 = (inp[8]) ? 11'b10001011111 : 11'b10010011110;
										assign node1345 = (inp[11]) ? 11'b00010011110 : 11'b10100101110;
									assign node1348 = (inp[10]) ? node1358 : node1349;
										assign node1349 = (inp[5]) ? node1355 : node1350;
											assign node1350 = (inp[8]) ? 11'b10110101101 : node1351;
												assign node1351 = (inp[11]) ? 11'b10011001110 : 11'b10110101100;
											assign node1355 = (inp[11]) ? 11'b10000111101 : 11'b10011011110;
										assign node1358 = (inp[11]) ? node1364 : node1359;
											assign node1359 = (inp[5]) ? 11'b00110111010 : node1360;
												assign node1360 = (inp[8]) ? 11'b00110001001 : 11'b00010101000;
											assign node1364 = (inp[8]) ? 11'b00011011001 : 11'b00011101011;
								assign node1367 = (inp[10]) ? node1379 : node1368;
									assign node1368 = (inp[3]) ? node1374 : node1369;
										assign node1369 = (inp[8]) ? 11'b00000001111 : node1370;
											assign node1370 = (inp[5]) ? 11'b00010011110 : 11'b00100011110;
										assign node1374 = (inp[11]) ? 11'b10000001010 : node1375;
											assign node1375 = (inp[5]) ? 11'b10011101010 : 11'b10001111010;
									assign node1379 = (inp[3]) ? node1387 : node1380;
										assign node1380 = (inp[5]) ? node1384 : node1381;
											assign node1381 = (inp[11]) ? 11'b10001111000 : 11'b10001101000;
											assign node1384 = (inp[8]) ? 11'b10001111000 : 11'b10100011010;
										assign node1387 = (inp[5]) ? node1393 : node1388;
											assign node1388 = (inp[11]) ? 11'b00001111010 : node1389;
												assign node1389 = (inp[8]) ? 11'b00011111011 : 11'b00010111000;
											assign node1393 = (inp[8]) ? 11'b00000001000 : 11'b00000101001;
						assign node1396 = (inp[9]) ? node1454 : node1397;
							assign node1397 = (inp[3]) ? node1429 : node1398;
								assign node1398 = (inp[10]) ? node1412 : node1399;
									assign node1399 = (inp[11]) ? node1409 : node1400;
										assign node1400 = (inp[8]) ? node1404 : node1401;
											assign node1401 = (inp[5]) ? 11'b00110101000 : 11'b00001001001;
											assign node1404 = (inp[5]) ? 11'b00101001011 : node1405;
												assign node1405 = (inp[4]) ? 11'b00101001001 : 11'b00100101001;
										assign node1409 = (inp[8]) ? 11'b00110111011 : 11'b00100111011;
									assign node1412 = (inp[5]) ? node1418 : node1413;
										assign node1413 = (inp[11]) ? 11'b00100111111 : node1414;
											assign node1414 = (inp[4]) ? 11'b00100011111 : 11'b00101001101;
										assign node1418 = (inp[8]) ? node1424 : node1419;
											assign node1419 = (inp[11]) ? 11'b00100101101 : node1420;
												assign node1420 = (inp[4]) ? 11'b00011011110 : 11'b00110101100;
											assign node1424 = (inp[4]) ? node1426 : 11'b00001001101;
												assign node1426 = (inp[11]) ? 11'b00011001100 : 11'b00110111100;
								assign node1429 = (inp[4]) ? node1441 : node1430;
									assign node1430 = (inp[11]) ? node1434 : node1431;
										assign node1431 = (inp[8]) ? 11'b00111001011 : 11'b00011001011;
										assign node1434 = (inp[8]) ? 11'b00100101010 : node1435;
											assign node1435 = (inp[5]) ? node1437 : 11'b00101001000;
												assign node1437 = (inp[10]) ? 11'b00110001010 : 11'b00111001000;
									assign node1441 = (inp[8]) ? node1447 : node1442;
										assign node1442 = (inp[5]) ? node1444 : 11'b00010001010;
											assign node1444 = (inp[10]) ? 11'b00011101011 : 11'b00010111011;
										assign node1447 = (inp[5]) ? node1449 : 11'b00011011001;
											assign node1449 = (inp[11]) ? 11'b00001011010 : node1450;
												assign node1450 = (inp[10]) ? 11'b00100101010 : 11'b00100111010;
							assign node1454 = (inp[3]) ? node1474 : node1455;
								assign node1455 = (inp[10]) ? node1463 : node1456;
									assign node1456 = (inp[5]) ? node1458 : 11'b00000001111;
										assign node1458 = (inp[8]) ? 11'b00010001110 : node1459;
											assign node1459 = (inp[4]) ? 11'b00111101111 : 11'b00011101110;
									assign node1463 = (inp[11]) ? node1471 : node1464;
										assign node1464 = (inp[8]) ? node1468 : node1465;
											assign node1465 = (inp[5]) ? 11'b00110011000 : 11'b00011111000;
											assign node1468 = (inp[4]) ? 11'b00011111010 : 11'b00001111010;
										assign node1471 = (inp[5]) ? 11'b00010001010 : 11'b00010001011;
								assign node1474 = (inp[5]) ? node1484 : node1475;
									assign node1475 = (inp[10]) ? node1481 : node1476;
										assign node1476 = (inp[4]) ? 11'b00111101000 : node1477;
											assign node1477 = (inp[8]) ? 11'b00111111011 : 11'b00011111010;
										assign node1481 = (inp[4]) ? 11'b00000001001 : 11'b00001001011;
									assign node1484 = (inp[8]) ? node1486 : 11'b00001101001;
										assign node1486 = (inp[11]) ? 11'b00000001000 : node1487;
											assign node1487 = (inp[4]) ? 11'b00001101000 : 11'b00011101000;
				assign node1491 = (inp[8]) ? node1791 : node1492;
					assign node1492 = (inp[5]) ? node1654 : node1493;
						assign node1493 = (inp[2]) ? node1575 : node1494;
							assign node1494 = (inp[4]) ? node1532 : node1495;
								assign node1495 = (inp[11]) ? node1515 : node1496;
									assign node1496 = (inp[3]) ? node1508 : node1497;
										assign node1497 = (inp[9]) ? node1505 : node1498;
											assign node1498 = (inp[10]) ? node1502 : node1499;
												assign node1499 = (inp[0]) ? 11'b00011101000 : 11'b00011101010;
												assign node1502 = (inp[0]) ? 11'b00011101100 : 11'b10011101000;
											assign node1505 = (inp[10]) ? 11'b00011111010 : 11'b00010101110;
										assign node1508 = (inp[0]) ? node1512 : node1509;
											assign node1509 = (inp[9]) ? 11'b10000101110 : 11'b10001101000;
											assign node1512 = (inp[9]) ? 11'b00000111000 : 11'b00000101010;
									assign node1515 = (inp[3]) ? node1525 : node1516;
										assign node1516 = (inp[0]) ? node1522 : node1517;
											assign node1517 = (inp[9]) ? 11'b10101011100 : node1518;
												assign node1518 = (inp[10]) ? 11'b10000001010 : 11'b00000001010;
											assign node1522 = (inp[9]) ? 11'b00000001010 : 11'b00010011100;
										assign node1525 = (inp[10]) ? node1527 : 11'b10010011000;
											assign node1527 = (inp[9]) ? node1529 : 11'b00011011110;
												assign node1529 = (inp[0]) ? 11'b00010001000 : 11'b00010011100;
								assign node1532 = (inp[11]) ? node1550 : node1533;
									assign node1533 = (inp[3]) ? node1541 : node1534;
										assign node1534 = (inp[9]) ? node1538 : node1535;
											assign node1535 = (inp[0]) ? 11'b00011101000 : 11'b00011101110;
											assign node1538 = (inp[0]) ? 11'b00111011110 : 11'b00110101100;
										assign node1541 = (inp[9]) ? node1545 : node1542;
											assign node1542 = (inp[10]) ? 11'b00100101010 : 11'b00000111010;
											assign node1545 = (inp[0]) ? node1547 : 11'b00101011000;
												assign node1547 = (inp[10]) ? 11'b00001001000 : 11'b00101001000;
									assign node1550 = (inp[0]) ? node1562 : node1551;
										assign node1551 = (inp[3]) ? node1557 : node1552;
											assign node1552 = (inp[9]) ? node1554 : 11'b10101110111;
												assign node1554 = (inp[10]) ? 11'b10110110001 : 11'b00011110101;
											assign node1557 = (inp[10]) ? node1559 : 11'b10000110011;
												assign node1559 = (inp[9]) ? 11'b00100110011 : 11'b00111110011;
										assign node1562 = (inp[9]) ? node1570 : node1563;
											assign node1563 = (inp[10]) ? node1567 : node1564;
												assign node1564 = (inp[3]) ? 11'b00111110011 : 11'b00000011010;
												assign node1567 = (inp[3]) ? 11'b00011100011 : 11'b00101100101;
											assign node1570 = (inp[10]) ? node1572 : 11'b00110100001;
												assign node1572 = (inp[3]) ? 11'b00000100001 : 11'b00100100011;
							assign node1575 = (inp[0]) ? node1613 : node1576;
								assign node1576 = (inp[10]) ? node1600 : node1577;
									assign node1577 = (inp[3]) ? node1589 : node1578;
										assign node1578 = (inp[9]) ? node1582 : node1579;
											assign node1579 = (inp[11]) ? 11'b00101100011 : 11'b00111000010;
											assign node1582 = (inp[4]) ? node1586 : node1583;
												assign node1583 = (inp[11]) ? 11'b00000110011 : 11'b00110000000;
												assign node1586 = (inp[11]) ? 11'b00110010101 : 11'b00000100101;
										assign node1589 = (inp[11]) ? node1595 : node1590;
											assign node1590 = (inp[4]) ? 11'b10111100111 : node1591;
												assign node1591 = (inp[9]) ? 11'b10110000110 : 11'b10111000000;
											assign node1595 = (inp[4]) ? node1597 : 11'b10111110001;
												assign node1597 = (inp[9]) ? 11'b10101010011 : 11'b10000000111;
									assign node1600 = (inp[4]) ? node1604 : node1601;
										assign node1601 = (inp[9]) ? 11'b00101110111 : 11'b00100110101;
										assign node1604 = (inp[3]) ? node1610 : node1605;
											assign node1605 = (inp[9]) ? node1607 : 11'b10101110101;
												assign node1607 = (inp[11]) ? 11'b10001010001 : 11'b10011100011;
											assign node1610 = (inp[9]) ? 11'b00001110001 : 11'b00000100011;
								assign node1613 = (inp[3]) ? node1633 : node1614;
									assign node1614 = (inp[4]) ? node1622 : node1615;
										assign node1615 = (inp[11]) ? node1619 : node1616;
											assign node1616 = (inp[10]) ? 11'b00000010000 : 11'b00010000100;
											assign node1619 = (inp[10]) ? 11'b00010110101 : 11'b00100110101;
										assign node1622 = (inp[11]) ? node1628 : node1623;
											assign node1623 = (inp[10]) ? 11'b00000110111 : node1624;
												assign node1624 = (inp[9]) ? 11'b00110110111 : 11'b00011100011;
											assign node1628 = (inp[10]) ? 11'b00110000111 : node1629;
												assign node1629 = (inp[9]) ? 11'b00011000111 : 11'b00001010001;
									assign node1633 = (inp[4]) ? node1643 : node1634;
										assign node1634 = (inp[11]) ? node1638 : node1635;
											assign node1635 = (inp[10]) ? 11'b00000000010 : 11'b00011000010;
											assign node1638 = (inp[9]) ? 11'b00111010011 : node1639;
												assign node1639 = (inp[10]) ? 11'b00100100011 : 11'b00010100011;
										assign node1643 = (inp[11]) ? node1649 : node1644;
											assign node1644 = (inp[9]) ? node1646 : 11'b00011110001;
												assign node1646 = (inp[10]) ? 11'b00001100001 : 11'b00110100001;
											assign node1649 = (inp[10]) ? 11'b00010000001 : node1650;
												assign node1650 = (inp[9]) ? 11'b00101000001 : 11'b00100010011;
						assign node1654 = (inp[9]) ? node1720 : node1655;
							assign node1655 = (inp[0]) ? node1687 : node1656;
								assign node1656 = (inp[2]) ? node1672 : node1657;
									assign node1657 = (inp[10]) ? node1665 : node1658;
										assign node1658 = (inp[4]) ? 11'b10111010101 : node1659;
											assign node1659 = (inp[11]) ? 11'b00001010001 : node1660;
												assign node1660 = (inp[3]) ? 11'b10001110001 : 11'b00011110011;
										assign node1665 = (inp[3]) ? node1669 : node1666;
											assign node1666 = (inp[4]) ? 11'b10000100101 : 11'b10100010001;
											assign node1669 = (inp[11]) ? 11'b00111100011 : 11'b00000010001;
									assign node1672 = (inp[3]) ? node1678 : node1673;
										assign node1673 = (inp[10]) ? node1675 : 11'b00110010011;
											assign node1675 = (inp[11]) ? 11'b10010110001 : 11'b10010010011;
										assign node1678 = (inp[11]) ? node1682 : node1679;
											assign node1679 = (inp[4]) ? 11'b10000110101 : 11'b00000010101;
											assign node1682 = (inp[10]) ? node1684 : 11'b10010010101;
												assign node1684 = (inp[4]) ? 11'b00011000001 : 11'b00111000111;
								assign node1687 = (inp[3]) ? node1703 : node1688;
									assign node1688 = (inp[10]) ? node1694 : node1689;
										assign node1689 = (inp[4]) ? node1691 : 11'b00010010011;
											assign node1691 = (inp[2]) ? 11'b00100100001 : 11'b00110110001;
										assign node1694 = (inp[11]) ? node1698 : node1695;
											assign node1695 = (inp[2]) ? 11'b00100000111 : 11'b00000010111;
											assign node1698 = (inp[4]) ? node1700 : 11'b00011010111;
												assign node1700 = (inp[2]) ? 11'b00111000111 : 11'b00111100111;
									assign node1703 = (inp[4]) ? node1709 : node1704;
										assign node1704 = (inp[2]) ? node1706 : 11'b00110000001;
											assign node1706 = (inp[10]) ? 11'b00000000001 : 11'b00110000001;
										assign node1709 = (inp[11]) ? node1713 : node1710;
											assign node1710 = (inp[10]) ? 11'b00110000011 : 11'b00111010001;
											assign node1713 = (inp[10]) ? node1717 : node1714;
												assign node1714 = (inp[2]) ? 11'b00010010001 : 11'b00000110011;
												assign node1717 = (inp[2]) ? 11'b00011000001 : 11'b00011100001;
							assign node1720 = (inp[0]) ? node1758 : node1721;
								assign node1721 = (inp[4]) ? node1739 : node1722;
									assign node1722 = (inp[11]) ? node1728 : node1723;
										assign node1723 = (inp[3]) ? node1725 : 11'b10100100101;
											assign node1725 = (inp[10]) ? 11'b00111100101 : 11'b10111110101;
										assign node1728 = (inp[2]) ? node1736 : node1729;
											assign node1729 = (inp[3]) ? node1733 : node1730;
												assign node1730 = (inp[10]) ? 11'b10111100111 : 11'b00101100011;
												assign node1733 = (inp[10]) ? 11'b00001100101 : 11'b10001110101;
											assign node1736 = (inp[3]) ? 11'b00100000111 : 11'b10001000101;
									assign node1739 = (inp[3]) ? node1749 : node1740;
										assign node1740 = (inp[10]) ? node1744 : node1741;
											assign node1741 = (inp[2]) ? 11'b00011110101 : 11'b00001100101;
											assign node1744 = (inp[11]) ? 11'b10100000011 : node1745;
												assign node1745 = (inp[2]) ? 11'b10101110001 : 11'b10011010001;
										assign node1749 = (inp[10]) ? node1755 : node1750;
											assign node1750 = (inp[2]) ? 11'b10111100011 : node1751;
												assign node1751 = (inp[11]) ? 11'b10111100001 : 11'b10000000001;
											assign node1755 = (inp[11]) ? 11'b00100100001 : 11'b00101000011;
								assign node1758 = (inp[11]) ? node1776 : node1759;
									assign node1759 = (inp[3]) ? node1769 : node1760;
										assign node1760 = (inp[10]) ? node1766 : node1761;
											assign node1761 = (inp[4]) ? 11'b00111110101 : node1762;
												assign node1762 = (inp[2]) ? 11'b00001100111 : 11'b00010100101;
											assign node1766 = (inp[4]) ? 11'b00101110001 : 11'b00111110001;
										assign node1769 = (inp[2]) ? node1771 : 11'b00100110011;
											assign node1771 = (inp[10]) ? 11'b00010100011 : node1772;
												assign node1772 = (inp[4]) ? 11'b00011100011 : 11'b00111110011;
									assign node1776 = (inp[3]) ? node1786 : node1777;
										assign node1777 = (inp[10]) ? node1781 : node1778;
											assign node1778 = (inp[2]) ? 11'b00101000111 : 11'b00101100111;
											assign node1781 = (inp[4]) ? node1783 : 11'b00101100001;
												assign node1783 = (inp[2]) ? 11'b00100000011 : 11'b00100100011;
										assign node1786 = (inp[2]) ? node1788 : 11'b00011100001;
											assign node1788 = (inp[10]) ? 11'b00000000001 : 11'b00001010001;
					assign node1791 = (inp[0]) ? node1897 : node1792;
						assign node1792 = (inp[2]) ? node1848 : node1793;
							assign node1793 = (inp[11]) ? node1823 : node1794;
								assign node1794 = (inp[5]) ? node1808 : node1795;
									assign node1795 = (inp[9]) ? node1805 : node1796;
										assign node1796 = (inp[4]) ? node1800 : node1797;
											assign node1797 = (inp[10]) ? 11'b00111000111 : 11'b10100100001;
											assign node1800 = (inp[3]) ? node1802 : 11'b00111000111;
												assign node1802 = (inp[10]) ? 11'b00011000001 : 11'b10011000101;
										assign node1805 = (inp[4]) ? 11'b00100000111 : 11'b00001000001;
									assign node1808 = (inp[10]) ? node1820 : node1809;
										assign node1809 = (inp[9]) ? node1817 : node1810;
											assign node1810 = (inp[4]) ? node1814 : node1811;
												assign node1811 = (inp[3]) ? 11'b10010010000 : 11'b00010010010;
												assign node1814 = (inp[3]) ? 11'b10000010110 : 11'b00100010100;
											assign node1817 = (inp[4]) ? 11'b10111100000 : 11'b10001010100;
										assign node1820 = (inp[4]) ? 11'b00011110010 : 11'b00110000110;
								assign node1823 = (inp[5]) ? node1835 : node1824;
									assign node1824 = (inp[10]) ? node1830 : node1825;
										assign node1825 = (inp[9]) ? 11'b10011010010 : node1826;
											assign node1826 = (inp[4]) ? 11'b10001100100 : 11'b10111110010;
										assign node1830 = (inp[4]) ? 11'b00101010010 : node1831;
											assign node1831 = (inp[9]) ? 11'b10001110110 : 11'b00000110110;
									assign node1835 = (inp[9]) ? node1843 : node1836;
										assign node1836 = (inp[4]) ? 11'b00110110100 : node1837;
											assign node1837 = (inp[3]) ? 11'b10010100000 : node1838;
												assign node1838 = (inp[10]) ? 11'b10011110010 : 11'b00000110010;
										assign node1843 = (inp[3]) ? node1845 : 11'b10100000010;
											assign node1845 = (inp[10]) ? 11'b00100100110 : 11'b10110110110;
							assign node1848 = (inp[11]) ? node1868 : node1849;
								assign node1849 = (inp[9]) ? node1857 : node1850;
									assign node1850 = (inp[5]) ? node1854 : node1851;
										assign node1851 = (inp[4]) ? 11'b00111100010 : 11'b00011100100;
										assign node1854 = (inp[4]) ? 11'b00101110000 : 11'b10111110000;
									assign node1857 = (inp[5]) ? node1865 : node1858;
										assign node1858 = (inp[3]) ? node1862 : node1859;
											assign node1859 = (inp[10]) ? 11'b10100110110 : 11'b00011100100;
											assign node1862 = (inp[10]) ? 11'b00000110010 : 11'b10100110010;
										assign node1865 = (inp[10]) ? 11'b00000100000 : 11'b10000100000;
								assign node1868 = (inp[9]) ? node1884 : node1869;
									assign node1869 = (inp[4]) ? node1877 : node1870;
										assign node1870 = (inp[3]) ? node1874 : node1871;
											assign node1871 = (inp[10]) ? 11'b10001000000 : 11'b00100100000;
											assign node1874 = (inp[10]) ? 11'b00101000100 : 11'b10101000000;
										assign node1877 = (inp[5]) ? node1881 : node1878;
											assign node1878 = (inp[10]) ? 11'b10001010100 : 11'b00010000100;
											assign node1881 = (inp[3]) ? 11'b10001010100 : 11'b00001010110;
									assign node1884 = (inp[5]) ? node1890 : node1885;
										assign node1885 = (inp[4]) ? 11'b10100010010 : node1886;
											assign node1886 = (inp[10]) ? 11'b00010010110 : 11'b00011010000;
										assign node1890 = (inp[4]) ? 11'b10000000000 : node1891;
											assign node1891 = (inp[10]) ? node1893 : 11'b10000010100;
												assign node1893 = (inp[3]) ? 11'b00000000100 : 11'b10000000110;
						assign node1897 = (inp[3]) ? node1967 : node1898;
							assign node1898 = (inp[11]) ? node1938 : node1899;
								assign node1899 = (inp[2]) ? node1919 : node1900;
									assign node1900 = (inp[5]) ? node1912 : node1901;
										assign node1901 = (inp[9]) ? node1905 : node1902;
											assign node1902 = (inp[10]) ? 11'b00111010101 : 11'b00111000011;
											assign node1905 = (inp[10]) ? node1909 : node1906;
												assign node1906 = (inp[4]) ? 11'b00000010101 : 11'b00101000101;
												assign node1909 = (inp[4]) ? 11'b00010010001 : 11'b00100010011;
										assign node1912 = (inp[9]) ? node1916 : node1913;
											assign node1913 = (inp[10]) ? 11'b00000000110 : 11'b00000000000;
											assign node1916 = (inp[10]) ? 11'b00011010000 : 11'b00101000100;
									assign node1919 = (inp[9]) ? node1929 : node1920;
										assign node1920 = (inp[5]) ? node1926 : node1921;
											assign node1921 = (inp[10]) ? 11'b00111100100 : node1922;
												assign node1922 = (inp[4]) ? 11'b00110100000 : 11'b00110000001;
											assign node1926 = (inp[4]) ? 11'b00011100010 : 11'b00111100010;
										assign node1929 = (inp[10]) ? node1933 : node1930;
											assign node1930 = (inp[4]) ? 11'b00011110100 : 11'b00101100100;
											assign node1933 = (inp[4]) ? node1935 : 11'b00100110000;
												assign node1935 = (inp[5]) ? 11'b00000110010 : 11'b00000110000;
								assign node1938 = (inp[4]) ? node1954 : node1939;
									assign node1939 = (inp[2]) ? node1949 : node1940;
										assign node1940 = (inp[9]) ? node1944 : node1941;
											assign node1941 = (inp[5]) ? 11'b00101110100 : 11'b00100110110;
											assign node1944 = (inp[10]) ? 11'b00111100000 : node1945;
												assign node1945 = (inp[5]) ? 11'b00011110100 : 11'b00010110110;
										assign node1949 = (inp[9]) ? node1951 : 11'b00101010010;
											assign node1951 = (inp[5]) ? 11'b00000010110 : 11'b00010010110;
									assign node1954 = (inp[5]) ? node1964 : node1955;
										assign node1955 = (inp[10]) ? node1959 : node1956;
											assign node1956 = (inp[9]) ? 11'b00111000110 : 11'b00101010010;
											assign node1959 = (inp[9]) ? node1961 : 11'b00001000110;
												assign node1961 = (inp[2]) ? 11'b00000000010 : 11'b00001000010;
										assign node1964 = (inp[2]) ? 11'b00000000110 : 11'b00010000110;
							assign node1967 = (inp[10]) ? node1989 : node1968;
								assign node1968 = (inp[5]) ? node1980 : node1969;
									assign node1969 = (inp[11]) ? node1973 : node1970;
										assign node1970 = (inp[2]) ? 11'b00000110010 : 11'b00010010001;
										assign node1973 = (inp[9]) ? node1975 : 11'b00110110010;
											assign node1975 = (inp[4]) ? node1977 : 11'b00100110000;
												assign node1977 = (inp[2]) ? 11'b00100000000 : 11'b00111000000;
									assign node1980 = (inp[4]) ? 11'b00000100000 : node1981;
										assign node1981 = (inp[2]) ? node1985 : node1982;
											assign node1982 = (inp[11]) ? 11'b00111100010 : 11'b00100000000;
											assign node1985 = (inp[11]) ? 11'b00101000000 : 11'b00111100000;
								assign node1989 = (inp[9]) ? node1997 : node1990;
									assign node1990 = (inp[11]) ? node1994 : node1991;
										assign node1991 = (inp[5]) ? 11'b00011000010 : 11'b00110000011;
										assign node1994 = (inp[4]) ? 11'b00001000000 : 11'b00101000000;
									assign node1997 = (inp[5]) ? node2005 : node1998;
										assign node1998 = (inp[11]) ? node2002 : node1999;
											assign node1999 = (inp[2]) ? 11'b00000100010 : 11'b00001100010;
											assign node2002 = (inp[2]) ? 11'b00010000000 : 11'b00011100010;
										assign node2005 = (inp[4]) ? node2007 : 11'b00000100010;
											assign node2007 = (inp[11]) ? 11'b00000000000 : 11'b00000100000;
		assign node2010 = (inp[7]) ? node3034 : node2011;
			assign node2011 = (inp[6]) ? node2529 : node2012;
				assign node2012 = (inp[8]) ? node2262 : node2013;
					assign node2013 = (inp[0]) ? node2123 : node2014;
						assign node2014 = (inp[4]) ? node2074 : node2015;
							assign node2015 = (inp[9]) ? node2047 : node2016;
								assign node2016 = (inp[3]) ? node2034 : node2017;
									assign node2017 = (inp[5]) ? node2023 : node2018;
										assign node2018 = (inp[10]) ? node2020 : 11'b00100101011;
											assign node2020 = (inp[11]) ? 11'b10001001011 : 11'b10001101011;
										assign node2023 = (inp[10]) ? node2027 : node2024;
											assign node2024 = (inp[11]) ? 11'b00000111001 : 11'b00000011001;
											assign node2027 = (inp[2]) ? node2031 : node2028;
												assign node2028 = (inp[11]) ? 11'b10101011001 : 11'b10101111001;
												assign node2031 = (inp[11]) ? 11'b10001111011 : 11'b10010011001;
									assign node2034 = (inp[10]) ? node2040 : node2035;
										assign node2035 = (inp[5]) ? node2037 : 11'b10101001000;
											assign node2037 = (inp[2]) ? 11'b10100011011 : 11'b10001111011;
										assign node2040 = (inp[2]) ? 11'b00101111111 : node2041;
											assign node2041 = (inp[11]) ? node2043 : 11'b00101111111;
												assign node2043 = (inp[5]) ? 11'b00011001111 : 11'b00001011101;
								assign node2047 = (inp[2]) ? node2059 : node2048;
									assign node2048 = (inp[3]) ? node2052 : node2049;
										assign node2049 = (inp[11]) ? 11'b10100011111 : 11'b10100101101;
										assign node2052 = (inp[11]) ? 11'b00000001101 : node2053;
											assign node2053 = (inp[5]) ? 11'b10000111111 : node2054;
												assign node2054 = (inp[10]) ? 11'b00000111101 : 11'b10000101101;
									assign node2059 = (inp[11]) ? node2065 : node2060;
										assign node2060 = (inp[3]) ? node2062 : 11'b00101001000;
											assign node2062 = (inp[5]) ? 11'b00101001101 : 11'b00110011110;
										assign node2065 = (inp[3]) ? node2069 : node2066;
											assign node2066 = (inp[5]) ? 11'b10010101111 : 11'b00011111001;
											assign node2069 = (inp[10]) ? node2071 : 11'b10100111101;
												assign node2071 = (inp[5]) ? 11'b00110101101 : 11'b00100111111;
							assign node2074 = (inp[3]) ? node2096 : node2075;
								assign node2075 = (inp[10]) ? node2085 : node2076;
									assign node2076 = (inp[2]) ? node2082 : node2077;
										assign node2077 = (inp[11]) ? node2079 : 11'b00010111101;
											assign node2079 = (inp[5]) ? 11'b00011001111 : 11'b00010011111;
										assign node2082 = (inp[5]) ? 11'b00111101101 : 11'b00111011111;
									assign node2085 = (inp[9]) ? node2091 : node2086;
										assign node2086 = (inp[2]) ? 11'b10111101101 : node2087;
											assign node2087 = (inp[5]) ? 11'b10001001111 : 11'b10111011111;
										assign node2091 = (inp[5]) ? node2093 : 11'b10010101011;
											assign node2093 = (inp[11]) ? 11'b10010001011 : 11'b10110011001;
								assign node2096 = (inp[10]) ? node2106 : node2097;
									assign node2097 = (inp[9]) ? node2101 : node2098;
										assign node2098 = (inp[5]) ? 11'b10001011101 : 11'b10101101111;
										assign node2101 = (inp[11]) ? node2103 : 11'b10000101011;
											assign node2103 = (inp[2]) ? 11'b10001101001 : 11'b10111001001;
									assign node2106 = (inp[2]) ? node2114 : node2107;
										assign node2107 = (inp[5]) ? 11'b00011111011 : node2108;
											assign node2108 = (inp[11]) ? node2110 : 11'b00100111001;
												assign node2110 = (inp[9]) ? 11'b00110011001 : 11'b00111011001;
										assign node2114 = (inp[5]) ? node2120 : node2115;
											assign node2115 = (inp[11]) ? node2117 : 11'b00000111001;
												assign node2117 = (inp[9]) ? 11'b00011011001 : 11'b00010111001;
											assign node2120 = (inp[11]) ? 11'b00010101001 : 11'b00110011001;
						assign node2123 = (inp[3]) ? node2195 : node2124;
							assign node2124 = (inp[5]) ? node2156 : node2125;
								assign node2125 = (inp[2]) ? node2141 : node2126;
									assign node2126 = (inp[11]) ? node2134 : node2127;
										assign node2127 = (inp[9]) ? 11'b00000111011 : node2128;
											assign node2128 = (inp[4]) ? 11'b00001111111 : node2129;
												assign node2129 = (inp[10]) ? 11'b00001101111 : 11'b00001101011;
										assign node2134 = (inp[9]) ? node2138 : node2135;
											assign node2135 = (inp[4]) ? 11'b00111001111 : 11'b00001011111;
											assign node2138 = (inp[4]) ? 11'b00010001111 : 11'b00010001011;
									assign node2141 = (inp[4]) ? node2151 : node2142;
										assign node2142 = (inp[11]) ? node2146 : node2143;
											assign node2143 = (inp[10]) ? 11'b00010011010 : 11'b00000001110;
											assign node2146 = (inp[10]) ? 11'b00001101001 : node2147;
												assign node2147 = (inp[9]) ? 11'b00111111111 : 11'b00010111011;
										assign node2151 = (inp[11]) ? 11'b00010111001 : node2152;
											assign node2152 = (inp[9]) ? 11'b00101111101 : 11'b00011111101;
								assign node2156 = (inp[11]) ? node2174 : node2157;
									assign node2157 = (inp[9]) ? node2165 : node2158;
										assign node2158 = (inp[4]) ? 11'b00111001001 : node2159;
											assign node2159 = (inp[10]) ? 11'b00110001111 : node2160;
												assign node2160 = (inp[2]) ? 11'b00000001011 : 11'b00001101011;
										assign node2165 = (inp[10]) ? node2169 : node2166;
											assign node2166 = (inp[2]) ? 11'b00100011111 : 11'b00110111111;
											assign node2169 = (inp[2]) ? 11'b00101011001 : node2170;
												assign node2170 = (inp[4]) ? 11'b00100111001 : 11'b00100111011;
									assign node2174 = (inp[9]) ? node2186 : node2175;
										assign node2175 = (inp[4]) ? node2181 : node2176;
											assign node2176 = (inp[10]) ? node2178 : 11'b00011111001;
												assign node2178 = (inp[2]) ? 11'b00001111101 : 11'b00011011101;
											assign node2181 = (inp[10]) ? 11'b00101101101 : node2182;
												assign node2182 = (inp[2]) ? 11'b00101111011 : 11'b00100011001;
										assign node2186 = (inp[10]) ? node2192 : node2187;
											assign node2187 = (inp[2]) ? node2189 : 11'b00111011101;
												assign node2189 = (inp[4]) ? 11'b00111101101 : 11'b00110111101;
											assign node2192 = (inp[2]) ? 11'b00110101001 : 11'b00110001001;
							assign node2195 = (inp[9]) ? node2225 : node2196;
								assign node2196 = (inp[10]) ? node2210 : node2197;
									assign node2197 = (inp[4]) ? node2203 : node2198;
										assign node2198 = (inp[5]) ? node2200 : 11'b00001001001;
											assign node2200 = (inp[11]) ? 11'b00111101011 : 11'b00101101001;
										assign node2203 = (inp[2]) ? 11'b00011111001 : node2204;
											assign node2204 = (inp[11]) ? 11'b00111011001 : node2205;
												assign node2205 = (inp[5]) ? 11'b00111111001 : 11'b00001111001;
									assign node2210 = (inp[5]) ? node2218 : node2211;
										assign node2211 = (inp[11]) ? 11'b00011001001 : node2212;
											assign node2212 = (inp[4]) ? node2214 : 11'b00001001000;
												assign node2214 = (inp[2]) ? 11'b00101101011 : 11'b00101101001;
										assign node2218 = (inp[2]) ? node2220 : 11'b00011001011;
											assign node2220 = (inp[4]) ? 11'b00110001001 : node2221;
												assign node2221 = (inp[11]) ? 11'b00110101011 : 11'b00000001011;
								assign node2225 = (inp[4]) ? node2241 : node2226;
									assign node2226 = (inp[10]) ? node2230 : node2227;
										assign node2227 = (inp[2]) ? 11'b00010011000 : 11'b00010011011;
										assign node2230 = (inp[2]) ? node2234 : node2231;
											assign node2231 = (inp[11]) ? 11'b00010001001 : 11'b00010101001;
											assign node2234 = (inp[11]) ? node2238 : node2235;
												assign node2235 = (inp[5]) ? 11'b00011001011 : 11'b00000001010;
												assign node2238 = (inp[5]) ? 11'b00000101001 : 11'b00010101011;
									assign node2241 = (inp[5]) ? node2253 : node2242;
										assign node2242 = (inp[11]) ? node2246 : node2243;
											assign node2243 = (inp[10]) ? 11'b00000101001 : 11'b00100101001;
											assign node2246 = (inp[2]) ? node2250 : node2247;
												assign node2247 = (inp[10]) ? 11'b00000001001 : 11'b00110001001;
												assign node2250 = (inp[10]) ? 11'b00001001001 : 11'b00101001001;
										assign node2253 = (inp[10]) ? node2259 : node2254;
											assign node2254 = (inp[11]) ? node2256 : 11'b00010001001;
												assign node2256 = (inp[2]) ? 11'b00000101011 : 11'b00010001011;
											assign node2259 = (inp[11]) ? 11'b00000001001 : 11'b00000101011;
					assign node2262 = (inp[0]) ? node2380 : node2263;
						assign node2263 = (inp[2]) ? node2325 : node2264;
							assign node2264 = (inp[11]) ? node2296 : node2265;
								assign node2265 = (inp[4]) ? node2279 : node2266;
									assign node2266 = (inp[9]) ? node2276 : node2267;
										assign node2267 = (inp[5]) ? node2271 : node2268;
											assign node2268 = (inp[3]) ? 11'b10100001001 : 11'b00000001011;
											assign node2271 = (inp[3]) ? 11'b10000011010 : node2272;
												assign node2272 = (inp[10]) ? 11'b10100011000 : 11'b00001011000;
										assign node2276 = (inp[3]) ? 11'b10001111110 : 11'b10001101100;
									assign node2279 = (inp[3]) ? node2285 : node2280;
										assign node2280 = (inp[5]) ? node2282 : 11'b00100101100;
											assign node2282 = (inp[9]) ? 11'b00100111110 : 11'b00111111100;
										assign node2285 = (inp[10]) ? node2289 : node2286;
											assign node2286 = (inp[5]) ? 11'b10110101000 : 11'b10000101110;
											assign node2289 = (inp[9]) ? node2293 : node2290;
												assign node2290 = (inp[5]) ? 11'b00000111000 : 11'b00011101010;
												assign node2293 = (inp[5]) ? 11'b00101101000 : 11'b00100111010;
								assign node2296 = (inp[4]) ? node2312 : node2297;
									assign node2297 = (inp[9]) ? node2307 : node2298;
										assign node2298 = (inp[5]) ? node2302 : node2299;
											assign node2299 = (inp[3]) ? 11'b10100111010 : 11'b10110101000;
											assign node2302 = (inp[3]) ? 11'b00000101110 : node2303;
												assign node2303 = (inp[10]) ? 11'b10010111010 : 11'b00001111010;
										assign node2307 = (inp[5]) ? 11'b10110101100 : node2308;
											assign node2308 = (inp[10]) ? 11'b00101011100 : 11'b00111011000;
									assign node2312 = (inp[10]) ? node2320 : node2313;
										assign node2313 = (inp[3]) ? node2317 : node2314;
											assign node2314 = (inp[9]) ? 11'b00001011110 : 11'b00101011100;
											assign node2317 = (inp[5]) ? 11'b10101011110 : 11'b10010001100;
										assign node2320 = (inp[9]) ? node2322 : 11'b00100011000;
											assign node2322 = (inp[3]) ? 11'b00111011000 : 11'b10111011010;
							assign node2325 = (inp[5]) ? node2357 : node2326;
								assign node2326 = (inp[11]) ? node2342 : node2327;
									assign node2327 = (inp[9]) ? node2331 : node2328;
										assign node2328 = (inp[4]) ? 11'b10110001101 : 11'b00100101011;
										assign node2331 = (inp[10]) ? node2337 : node2332;
											assign node2332 = (inp[3]) ? 11'b10001001111 : node2333;
												assign node2333 = (inp[4]) ? 11'b00011001111 : 11'b00111001001;
											assign node2337 = (inp[3]) ? node2339 : 11'b10101011101;
												assign node2339 = (inp[4]) ? 11'b00001011011 : 11'b00010011111;
									assign node2342 = (inp[4]) ? node2348 : node2343;
										assign node2343 = (inp[3]) ? node2345 : 11'b10111111110;
											assign node2345 = (inp[9]) ? 11'b10010001101 : 11'b00110011101;
										assign node2348 = (inp[10]) ? node2352 : node2349;
											assign node2349 = (inp[9]) ? 11'b10110111000 : 11'b10101101110;
											assign node2352 = (inp[3]) ? node2354 : 11'b10000111010;
												assign node2354 = (inp[9]) ? 11'b00010111000 : 11'b00001111000;
								assign node2357 = (inp[3]) ? node2369 : node2358;
									assign node2358 = (inp[10]) ? node2364 : node2359;
										assign node2359 = (inp[11]) ? 11'b00100011010 : node2360;
											assign node2360 = (inp[9]) ? 11'b00111111000 : 11'b00100111000;
										assign node2364 = (inp[11]) ? 11'b10001001110 : node2365;
											assign node2365 = (inp[9]) ? 11'b10110101110 : 11'b10110101100;
									assign node2369 = (inp[11]) ? node2373 : node2370;
										assign node2370 = (inp[9]) ? 11'b10001001000 : 11'b00101011010;
										assign node2373 = (inp[9]) ? node2377 : node2374;
											assign node2374 = (inp[4]) ? 11'b10011011100 : 11'b10110001000;
											assign node2377 = (inp[4]) ? 11'b00010001000 : 11'b00011001100;
						assign node2380 = (inp[3]) ? node2462 : node2381;
							assign node2381 = (inp[5]) ? node2419 : node2382;
								assign node2382 = (inp[11]) ? node2398 : node2383;
									assign node2383 = (inp[2]) ? node2391 : node2384;
										assign node2384 = (inp[9]) ? 11'b00110111010 : node2385;
											assign node2385 = (inp[10]) ? 11'b00101101110 : node2386;
												assign node2386 = (inp[4]) ? 11'b00100101010 : 11'b00100001011;
										assign node2391 = (inp[4]) ? node2395 : node2392;
											assign node2392 = (inp[9]) ? 11'b00111001111 : 11'b00101001111;
											assign node2395 = (inp[10]) ? 11'b00100011111 : 11'b00001011111;
									assign node2398 = (inp[4]) ? node2406 : node2399;
										assign node2399 = (inp[9]) ? node2403 : node2400;
											assign node2400 = (inp[10]) ? 11'b00100011101 : 11'b00111011001;
											assign node2403 = (inp[2]) ? 11'b00000011111 : 11'b00001011100;
										assign node2406 = (inp[2]) ? node2412 : node2407;
											assign node2407 = (inp[9]) ? node2409 : 11'b00000001110;
												assign node2409 = (inp[10]) ? 11'b00011001010 : 11'b00101001110;
											assign node2412 = (inp[9]) ? node2416 : node2413;
												assign node2413 = (inp[10]) ? 11'b00011101100 : 11'b00111111010;
												assign node2416 = (inp[10]) ? 11'b00010101010 : 11'b00110101100;
								assign node2419 = (inp[11]) ? node2439 : node2420;
									assign node2420 = (inp[4]) ? node2430 : node2421;
										assign node2421 = (inp[2]) ? node2423 : 11'b00010001110;
											assign node2423 = (inp[10]) ? node2427 : node2424;
												assign node2424 = (inp[9]) ? 11'b00101101100 : 11'b00101101010;
												assign node2427 = (inp[9]) ? 11'b00000111010 : 11'b00001101100;
										assign node2430 = (inp[9]) ? node2434 : node2431;
											assign node2431 = (inp[10]) ? 11'b00111011110 : 11'b00000101010;
											assign node2434 = (inp[2]) ? node2436 : 11'b00001111010;
												assign node2436 = (inp[10]) ? 11'b00011011000 : 11'b00011011100;
									assign node2439 = (inp[4]) ? node2453 : node2440;
										assign node2440 = (inp[9]) ? node2446 : node2441;
											assign node2441 = (inp[10]) ? node2443 : 11'b00101111010;
												assign node2443 = (inp[2]) ? 11'b00110011110 : 11'b00110111110;
											assign node2446 = (inp[10]) ? node2450 : node2447;
												assign node2447 = (inp[2]) ? 11'b00010011100 : 11'b00000111110;
												assign node2450 = (inp[2]) ? 11'b00011001000 : 11'b00011001010;
										assign node2453 = (inp[9]) ? node2459 : node2454;
											assign node2454 = (inp[10]) ? node2456 : 11'b00011011010;
												assign node2456 = (inp[2]) ? 11'b00010001110 : 11'b00011001100;
											assign node2459 = (inp[10]) ? 11'b00010001000 : 11'b00010001100;
							assign node2462 = (inp[10]) ? node2504 : node2463;
								assign node2463 = (inp[2]) ? node2485 : node2464;
									assign node2464 = (inp[9]) ? node2478 : node2465;
										assign node2465 = (inp[11]) ? node2473 : node2466;
											assign node2466 = (inp[4]) ? node2470 : node2467;
												assign node2467 = (inp[5]) ? 11'b00100001000 : 11'b00000001001;
												assign node2470 = (inp[5]) ? 11'b00110111010 : 11'b00000111000;
											assign node2473 = (inp[4]) ? 11'b00011011010 : node2474;
												assign node2474 = (inp[5]) ? 11'b00111101000 : 11'b00010101010;
										assign node2478 = (inp[4]) ? node2482 : node2479;
											assign node2479 = (inp[5]) ? 11'b00010111000 : 11'b00011111000;
											assign node2482 = (inp[5]) ? 11'b00011101010 : 11'b00111101000;
									assign node2485 = (inp[11]) ? node2493 : node2486;
										assign node2486 = (inp[5]) ? 11'b00110111010 : node2487;
											assign node2487 = (inp[9]) ? 11'b00101001001 : node2488;
												assign node2488 = (inp[4]) ? 11'b00010011011 : 11'b00010101001;
										assign node2493 = (inp[5]) ? node2497 : node2494;
											assign node2494 = (inp[9]) ? 11'b00100101000 : 11'b00101111010;
											assign node2497 = (inp[9]) ? node2501 : node2498;
												assign node2498 = (inp[4]) ? 11'b00001011000 : 11'b00100001000;
												assign node2501 = (inp[4]) ? 11'b00000001010 : 11'b00001011010;
								assign node2504 = (inp[11]) ? node2516 : node2505;
									assign node2505 = (inp[2]) ? node2509 : node2506;
										assign node2506 = (inp[4]) ? 11'b00111101000 : 11'b00011101000;
										assign node2509 = (inp[4]) ? node2511 : 11'b00011101010;
											assign node2511 = (inp[5]) ? node2513 : 11'b00001001011;
												assign node2513 = (inp[9]) ? 11'b00001001000 : 11'b00101001010;
									assign node2516 = (inp[4]) ? node2524 : node2517;
										assign node2517 = (inp[9]) ? node2521 : node2518;
											assign node2518 = (inp[5]) ? 11'b00100001010 : 11'b00110001011;
											assign node2521 = (inp[5]) ? 11'b00001001000 : 11'b00010001010;
										assign node2524 = (inp[5]) ? 11'b00000001000 : node2525;
											assign node2525 = (inp[9]) ? 11'b00001001000 : 11'b00000001000;
				assign node2529 = (inp[2]) ? node2773 : node2530;
					assign node2530 = (inp[8]) ? node2668 : node2531;
						assign node2531 = (inp[5]) ? node2601 : node2532;
							assign node2532 = (inp[11]) ? node2568 : node2533;
								assign node2533 = (inp[9]) ? node2551 : node2534;
									assign node2534 = (inp[4]) ? node2546 : node2535;
										assign node2535 = (inp[0]) ? node2543 : node2536;
											assign node2536 = (inp[3]) ? node2540 : node2537;
												assign node2537 = (inp[10]) ? 11'b10001101000 : 11'b00001101010;
												assign node2540 = (inp[10]) ? 11'b00011101110 : 11'b10011101000;
											assign node2543 = (inp[3]) ? 11'b00001101010 : 11'b00011101110;
										assign node2546 = (inp[0]) ? 11'b00000111000 : node2547;
											assign node2547 = (inp[3]) ? 11'b10010101100 : 11'b00000101110;
									assign node2551 = (inp[4]) ? node2561 : node2552;
										assign node2552 = (inp[10]) ? node2556 : node2553;
											assign node2553 = (inp[3]) ? 11'b00000111010 : 11'b00001101000;
											assign node2556 = (inp[0]) ? 11'b00010111000 : node2557;
												assign node2557 = (inp[3]) ? 11'b00010111100 : 11'b10000111110;
										assign node2561 = (inp[3]) ? node2565 : node2562;
											assign node2562 = (inp[0]) ? 11'b00111111100 : 11'b00101101100;
											assign node2565 = (inp[0]) ? 11'b00101101010 : 11'b10111111010;
								assign node2568 = (inp[0]) ? node2586 : node2569;
									assign node2569 = (inp[4]) ? node2577 : node2570;
										assign node2570 = (inp[9]) ? node2574 : node2571;
											assign node2571 = (inp[3]) ? 11'b00000111110 : 11'b10010101000;
											assign node2574 = (inp[3]) ? 11'b00001011100 : 11'b10111011110;
										assign node2577 = (inp[9]) ? node2579 : 11'b10111011100;
											assign node2579 = (inp[3]) ? node2583 : node2580;
												assign node2580 = (inp[10]) ? 11'b10100011010 : 11'b00000011110;
												assign node2583 = (inp[10]) ? 11'b00110011000 : 11'b10010011000;
									assign node2586 = (inp[10]) ? node2592 : node2587;
										assign node2587 = (inp[3]) ? node2589 : 11'b00001011010;
											assign node2589 = (inp[9]) ? 11'b00101011010 : 11'b00111011000;
										assign node2592 = (inp[9]) ? node2598 : node2593;
											assign node2593 = (inp[3]) ? node2595 : 11'b00010111110;
												assign node2595 = (inp[4]) ? 11'b00010001010 : 11'b00100101010;
											assign node2598 = (inp[4]) ? 11'b00100001010 : 11'b00001001010;
							assign node2601 = (inp[11]) ? node2639 : node2602;
								assign node2602 = (inp[9]) ? node2628 : node2603;
									assign node2603 = (inp[0]) ? node2615 : node2604;
										assign node2604 = (inp[4]) ? node2608 : node2605;
											assign node2605 = (inp[3]) ? 11'b10011011010 : 11'b00000011000;
											assign node2608 = (inp[3]) ? node2612 : node2609;
												assign node2609 = (inp[10]) ? 11'b10000001110 : 11'b00010011100;
												assign node2612 = (inp[10]) ? 11'b00010011000 : 11'b10100011110;
										assign node2615 = (inp[3]) ? node2621 : node2616;
											assign node2616 = (inp[4]) ? node2618 : 11'b00111001100;
												assign node2618 = (inp[10]) ? 11'b00000011100 : 11'b00100001000;
											assign node2621 = (inp[4]) ? node2625 : node2622;
												assign node2622 = (inp[10]) ? 11'b00001001010 : 11'b00101001010;
												assign node2625 = (inp[10]) ? 11'b00111100011 : 11'b00110011010;
									assign node2628 = (inp[3]) ? node2632 : node2629;
										assign node2629 = (inp[10]) ? 11'b00111110011 : 11'b00101110111;
										assign node2632 = (inp[4]) ? node2634 : 11'b00101011000;
											assign node2634 = (inp[0]) ? node2636 : 11'b10011100001;
												assign node2636 = (inp[10]) ? 11'b00001100011 : 11'b00001100001;
								assign node2639 = (inp[0]) ? node2653 : node2640;
									assign node2640 = (inp[4]) ? node2648 : node2641;
										assign node2641 = (inp[3]) ? node2645 : node2642;
											assign node2642 = (inp[10]) ? 11'b10110110011 : 11'b00011110001;
											assign node2645 = (inp[10]) ? 11'b00011100111 : 11'b10010110111;
										assign node2648 = (inp[3]) ? 11'b10100100011 : node2649;
											assign node2649 = (inp[9]) ? 11'b00011100101 : 11'b10011100111;
									assign node2653 = (inp[3]) ? node2659 : node2654;
										assign node2654 = (inp[9]) ? node2656 : 11'b00000110111;
											assign node2656 = (inp[4]) ? 11'b00101100101 : 11'b00100100001;
										assign node2659 = (inp[9]) ? node2661 : 11'b00001110001;
											assign node2661 = (inp[10]) ? node2665 : node2662;
												assign node2662 = (inp[4]) ? 11'b00010100011 : 11'b00010110001;
												assign node2665 = (inp[4]) ? 11'b00000100001 : 11'b00001100011;
						assign node2668 = (inp[0]) ? node2724 : node2669;
							assign node2669 = (inp[5]) ? node2699 : node2670;
								assign node2670 = (inp[10]) ? node2684 : node2671;
									assign node2671 = (inp[3]) ? node2679 : node2672;
										assign node2672 = (inp[4]) ? node2674 : 11'b00011000001;
											assign node2674 = (inp[11]) ? node2676 : 11'b00110000111;
												assign node2676 = (inp[9]) ? 11'b00011110101 : 11'b00110000111;
										assign node2679 = (inp[9]) ? 11'b10110000111 : node2680;
											assign node2680 = (inp[11]) ? 11'b10101010001 : 11'b10110100001;
									assign node2684 = (inp[3]) ? node2688 : node2685;
										assign node2685 = (inp[4]) ? 11'b10110010101 : 11'b10001010111;
										assign node2688 = (inp[4]) ? node2694 : node2689;
											assign node2689 = (inp[11]) ? 11'b00011010101 : node2690;
												assign node2690 = (inp[9]) ? 11'b00111010101 : 11'b00101000111;
											assign node2694 = (inp[11]) ? 11'b00111110011 : node2695;
												assign node2695 = (inp[9]) ? 11'b00111010011 : 11'b00000000001;
								assign node2699 = (inp[9]) ? node2711 : node2700;
									assign node2700 = (inp[4]) ? node2706 : node2701;
										assign node2701 = (inp[3]) ? node2703 : 11'b00010110011;
											assign node2703 = (inp[11]) ? 11'b10000100011 : 11'b10000110011;
										assign node2706 = (inp[10]) ? 11'b10001100111 : node2707;
											assign node2707 = (inp[3]) ? 11'b10011110101 : 11'b00111110101;
									assign node2711 = (inp[4]) ? node2719 : node2712;
										assign node2712 = (inp[11]) ? 11'b10101010101 : node2713;
											assign node2713 = (inp[10]) ? node2715 : 11'b10010110101;
												assign node2715 = (inp[3]) ? 11'b00101100111 : 11'b10010100101;
										assign node2719 = (inp[3]) ? node2721 : 11'b10100110011;
											assign node2721 = (inp[10]) ? 11'b00110100001 : 11'b10100100011;
							assign node2724 = (inp[9]) ? node2754 : node2725;
								assign node2725 = (inp[10]) ? node2743 : node2726;
									assign node2726 = (inp[4]) ? node2734 : node2727;
										assign node2727 = (inp[11]) ? node2731 : node2728;
											assign node2728 = (inp[3]) ? 11'b00100100011 : 11'b00110100011;
											assign node2731 = (inp[3]) ? 11'b00110100001 : 11'b00110110011;
										assign node2734 = (inp[11]) ? node2740 : node2735;
											assign node2735 = (inp[5]) ? node2737 : 11'b00110000011;
												assign node2737 = (inp[3]) ? 11'b00111110011 : 11'b00001100001;
											assign node2740 = (inp[5]) ? 11'b00010010011 : 11'b00100010011;
									assign node2743 = (inp[3]) ? node2747 : node2744;
										assign node2744 = (inp[5]) ? 11'b00111110111 : 11'b00011100111;
										assign node2747 = (inp[5]) ? node2749 : 11'b00110000011;
											assign node2749 = (inp[4]) ? node2751 : 11'b00101000011;
												assign node2751 = (inp[11]) ? 11'b00000000001 : 11'b00101100001;
								assign node2754 = (inp[10]) ? node2766 : node2755;
									assign node2755 = (inp[3]) ? node2763 : node2756;
										assign node2756 = (inp[11]) ? 11'b00011010101 : node2757;
											assign node2757 = (inp[4]) ? 11'b00001110101 : node2758;
												assign node2758 = (inp[5]) ? 11'b00100100111 : 11'b00101000101;
										assign node2763 = (inp[5]) ? 11'b00010000011 : 11'b00011010011;
									assign node2766 = (inp[11]) ? node2770 : node2767;
										assign node2767 = (inp[4]) ? 11'b00010110001 : 11'b00011110011;
										assign node2770 = (inp[3]) ? 11'b00001100001 : 11'b00001100011;
					assign node2773 = (inp[5]) ? node2891 : node2774;
						assign node2774 = (inp[11]) ? node2838 : node2775;
							assign node2775 = (inp[8]) ? node2805 : node2776;
								assign node2776 = (inp[9]) ? node2796 : node2777;
									assign node2777 = (inp[4]) ? node2787 : node2778;
										assign node2778 = (inp[0]) ? 11'b00001000101 : node2779;
											assign node2779 = (inp[10]) ? node2783 : node2780;
												assign node2780 = (inp[3]) ? 11'b10101000011 : 11'b00101000011;
												assign node2783 = (inp[3]) ? 11'b00111000111 : 11'b10111000001;
										assign node2787 = (inp[3]) ? node2791 : node2788;
											assign node2788 = (inp[0]) ? 11'b00000010111 : 11'b00100000101;
											assign node2791 = (inp[10]) ? node2793 : 11'b00010010011;
												assign node2793 = (inp[0]) ? 11'b00100000001 : 11'b00010000001;
									assign node2796 = (inp[4]) ? node2800 : node2797;
										assign node2797 = (inp[3]) ? 11'b00011010001 : 11'b00011000101;
										assign node2800 = (inp[10]) ? 11'b00101110000 : node2801;
											assign node2801 = (inp[3]) ? 11'b00111100010 : 11'b00111110110;
								assign node2805 = (inp[0]) ? node2825 : node2806;
									assign node2806 = (inp[9]) ? node2816 : node2807;
										assign node2807 = (inp[4]) ? node2809 : 11'b00000000100;
											assign node2809 = (inp[3]) ? node2813 : node2810;
												assign node2810 = (inp[10]) ? 11'b10001110100 : 11'b00011100110;
												assign node2813 = (inp[10]) ? 11'b00100100010 : 11'b10101100100;
										assign node2816 = (inp[4]) ? 11'b10110100010 : node2817;
											assign node2817 = (inp[10]) ? node2821 : node2818;
												assign node2818 = (inp[3]) ? 11'b10011100100 : 11'b00111100010;
												assign node2821 = (inp[3]) ? 11'b00011110110 : 11'b10111110100;
									assign node2825 = (inp[3]) ? node2829 : node2826;
										assign node2826 = (inp[4]) ? 11'b00111100000 : 11'b00110000010;
										assign node2829 = (inp[10]) ? node2833 : node2830;
											assign node2830 = (inp[4]) ? 11'b00011110000 : 11'b00001110000;
											assign node2833 = (inp[9]) ? node2835 : 11'b00011100010;
												assign node2835 = (inp[4]) ? 11'b00000100010 : 11'b00001100010;
							assign node2838 = (inp[0]) ? node2862 : node2839;
								assign node2839 = (inp[4]) ? node2851 : node2840;
									assign node2840 = (inp[9]) ? node2844 : node2841;
										assign node2841 = (inp[10]) ? 11'b00110110110 : 11'b10101110010;
										assign node2844 = (inp[10]) ? node2848 : node2845;
											assign node2845 = (inp[3]) ? 11'b10010100100 : 11'b00010110010;
											assign node2848 = (inp[3]) ? 11'b00100110110 : 11'b10000110100;
									assign node2851 = (inp[9]) ? node2857 : node2852;
										assign node2852 = (inp[10]) ? 11'b00010110000 : node2853;
											assign node2853 = (inp[8]) ? 11'b00001100100 : 11'b00110100100;
										assign node2857 = (inp[8]) ? 11'b10110110010 : node2858;
											assign node2858 = (inp[3]) ? 11'b00011110000 : 11'b10011110010;
								assign node2862 = (inp[10]) ? node2878 : node2863;
									assign node2863 = (inp[9]) ? node2871 : node2864;
										assign node2864 = (inp[4]) ? node2866 : 11'b00000100000;
											assign node2866 = (inp[8]) ? 11'b00100110010 : node2867;
												assign node2867 = (inp[3]) ? 11'b00100110000 : 11'b00000110000;
										assign node2871 = (inp[4]) ? 11'b00100100010 : node2872;
											assign node2872 = (inp[8]) ? node2874 : 11'b00100110110;
												assign node2874 = (inp[3]) ? 11'b00111110010 : 11'b00011110100;
									assign node2878 = (inp[3]) ? node2886 : node2879;
										assign node2879 = (inp[9]) ? node2883 : node2880;
											assign node2880 = (inp[4]) ? 11'b00111100110 : 11'b00111110110;
											assign node2883 = (inp[4]) ? 11'b00000100010 : 11'b00111100010;
										assign node2886 = (inp[8]) ? 11'b00000100000 : node2887;
											assign node2887 = (inp[9]) ? 11'b00001100000 : 11'b00011100000;
						assign node2891 = (inp[0]) ? node2971 : node2892;
							assign node2892 = (inp[4]) ? node2936 : node2893;
								assign node2893 = (inp[11]) ? node2915 : node2894;
									assign node2894 = (inp[9]) ? node2908 : node2895;
										assign node2895 = (inp[10]) ? node2903 : node2896;
											assign node2896 = (inp[3]) ? node2900 : node2897;
												assign node2897 = (inp[8]) ? 11'b00100110000 : 11'b00101110000;
												assign node2900 = (inp[8]) ? 11'b10101010010 : 11'b10100110010;
											assign node2903 = (inp[3]) ? 11'b00001010100 : node2904;
												assign node2904 = (inp[8]) ? 11'b10001010010 : 11'b10000110010;
										assign node2908 = (inp[8]) ? node2912 : node2909;
											assign node2909 = (inp[10]) ? 11'b00100100100 : 11'b10100110110;
											assign node2912 = (inp[10]) ? 11'b10101000110 : 11'b10101010110;
									assign node2915 = (inp[9]) ? node2925 : node2916;
										assign node2916 = (inp[8]) ? node2920 : node2917;
											assign node2917 = (inp[3]) ? 11'b00100000110 : 11'b10000010010;
											assign node2920 = (inp[3]) ? 11'b00111000100 : node2921;
												assign node2921 = (inp[10]) ? 11'b10111010000 : 11'b00111010010;
										assign node2925 = (inp[10]) ? node2929 : node2926;
											assign node2926 = (inp[8]) ? 11'b10011010110 : 11'b00000000000;
											assign node2929 = (inp[3]) ? node2933 : node2930;
												assign node2930 = (inp[8]) ? 11'b10011000100 : 11'b10011000110;
												assign node2933 = (inp[8]) ? 11'b00011000100 : 11'b00111000100;
								assign node2936 = (inp[9]) ? node2956 : node2937;
									assign node2937 = (inp[8]) ? node2945 : node2938;
										assign node2938 = (inp[3]) ? node2942 : node2939;
											assign node2939 = (inp[11]) ? 11'b00101010100 : 11'b10111000100;
											assign node2942 = (inp[10]) ? 11'b00101010010 : 11'b10011010100;
										assign node2945 = (inp[10]) ? node2951 : node2946;
											assign node2946 = (inp[3]) ? node2948 : 11'b00001010100;
												assign node2948 = (inp[11]) ? 11'b10010010110 : 11'b10110010110;
											assign node2951 = (inp[3]) ? 11'b00010000000 : node2952;
												assign node2952 = (inp[11]) ? 11'b10010000100 : 11'b10110000100;
									assign node2956 = (inp[10]) ? node2964 : node2957;
										assign node2957 = (inp[3]) ? 11'b10010000010 : node2958;
											assign node2958 = (inp[8]) ? node2960 : 11'b00001010110;
												assign node2960 = (inp[11]) ? 11'b00010000110 : 11'b00010010110;
										assign node2964 = (inp[3]) ? node2966 : 11'b10110000000;
											assign node2966 = (inp[11]) ? 11'b00010000000 : node2967;
												assign node2967 = (inp[8]) ? 11'b00010000000 : 11'b00010000010;
							assign node2971 = (inp[10]) ? node3003 : node2972;
								assign node2972 = (inp[3]) ? node2990 : node2973;
									assign node2973 = (inp[9]) ? node2981 : node2974;
										assign node2974 = (inp[11]) ? node2978 : node2975;
											assign node2975 = (inp[8]) ? 11'b00111000010 : 11'b00010100010;
											assign node2978 = (inp[4]) ? 11'b00000010010 : 11'b00000010000;
										assign node2981 = (inp[4]) ? node2985 : node2982;
											assign node2982 = (inp[8]) ? 11'b00111000110 : 11'b00000100110;
											assign node2985 = (inp[8]) ? 11'b00000010110 : node2986;
												assign node2986 = (inp[11]) ? 11'b00100000110 : 11'b00111010100;
									assign node2990 = (inp[8]) ? node2998 : node2991;
										assign node2991 = (inp[11]) ? node2995 : node2992;
											assign node2992 = (inp[9]) ? 11'b00011000000 : 11'b00101010000;
											assign node2995 = (inp[9]) ? 11'b00001010010 : 11'b00011010010;
										assign node2998 = (inp[11]) ? node3000 : 11'b00100010010;
											assign node3000 = (inp[4]) ? 11'b00000010010 : 11'b00001010010;
								assign node3003 = (inp[3]) ? node3019 : node3004;
									assign node3004 = (inp[9]) ? node3012 : node3005;
										assign node3005 = (inp[4]) ? node3007 : 11'b00010010110;
											assign node3007 = (inp[8]) ? 11'b00000000100 : node3008;
												assign node3008 = (inp[11]) ? 11'b00111000100 : 11'b00001010100;
										assign node3012 = (inp[8]) ? node3014 : 11'b00110110000;
											assign node3014 = (inp[4]) ? 11'b00000010000 : node3015;
												assign node3015 = (inp[11]) ? 11'b00001000000 : 11'b00011010000;
									assign node3019 = (inp[11]) ? node3025 : node3020;
										assign node3020 = (inp[4]) ? 11'b00111000010 : node3021;
											assign node3021 = (inp[9]) ? 11'b00011000010 : 11'b00000100000;
										assign node3025 = (inp[9]) ? node3031 : node3026;
											assign node3026 = (inp[4]) ? 11'b00011000000 : node3027;
												assign node3027 = (inp[8]) ? 11'b00101000000 : 11'b00110000000;
											assign node3031 = (inp[4]) ? 11'b00000000000 : 11'b00001000000;
			assign node3034 = (inp[6]) ? node3492 : node3035;
				assign node3035 = (inp[2]) ? node3271 : node3036;
					assign node3036 = (inp[5]) ? node3160 : node3037;
						assign node3037 = (inp[0]) ? node3099 : node3038;
							assign node3038 = (inp[11]) ? node3070 : node3039;
								assign node3039 = (inp[10]) ? node3059 : node3040;
									assign node3040 = (inp[3]) ? node3052 : node3041;
										assign node3041 = (inp[4]) ? node3047 : node3042;
											assign node3042 = (inp[8]) ? node3044 : 11'b00011100011;
												assign node3044 = (inp[9]) ? 11'b00000000001 : 11'b00010000011;
											assign node3047 = (inp[8]) ? 11'b00111100101 : node3048;
												assign node3048 = (inp[9]) ? 11'b00110100111 : 11'b00010100111;
										assign node3052 = (inp[9]) ? node3056 : node3053;
											assign node3053 = (inp[8]) ? 11'b10011100111 : 11'b10010100111;
											assign node3056 = (inp[8]) ? 11'b10101100111 : 11'b10011100111;
									assign node3059 = (inp[8]) ? node3065 : node3060;
										assign node3060 = (inp[3]) ? 11'b00110110001 : node3061;
											assign node3061 = (inp[9]) ? 11'b10011110101 : 11'b10010110101;
										assign node3065 = (inp[3]) ? 11'b00001100011 : node3066;
											assign node3066 = (inp[9]) ? 11'b10010100011 : 11'b10010000001;
								assign node3070 = (inp[9]) ? node3084 : node3071;
									assign node3071 = (inp[4]) ? node3079 : node3072;
										assign node3072 = (inp[3]) ? 11'b00000110111 : node3073;
											assign node3073 = (inp[8]) ? node3075 : 11'b10011100001;
												assign node3075 = (inp[10]) ? 11'b10100100001 : 11'b00010100001;
										assign node3079 = (inp[10]) ? 11'b00111110001 : node3080;
											assign node3080 = (inp[3]) ? 11'b10001100111 : 11'b00101100111;
									assign node3084 = (inp[10]) ? node3092 : node3085;
										assign node3085 = (inp[3]) ? 11'b10000110011 : node3086;
											assign node3086 = (inp[4]) ? 11'b00011110111 : node3087;
												assign node3087 = (inp[8]) ? 11'b00100110011 : 11'b00111110011;
										assign node3092 = (inp[4]) ? node3094 : 11'b10111110101;
											assign node3094 = (inp[3]) ? 11'b00100110001 : node3095;
												assign node3095 = (inp[8]) ? 11'b10101110011 : 11'b10100110011;
							assign node3099 = (inp[10]) ? node3121 : node3100;
								assign node3100 = (inp[11]) ? node3110 : node3101;
									assign node3101 = (inp[4]) ? node3107 : node3102;
										assign node3102 = (inp[9]) ? 11'b00011110011 : node3103;
											assign node3103 = (inp[3]) ? 11'b00000000011 : 11'b00100000011;
										assign node3107 = (inp[8]) ? 11'b00101100001 : 11'b00100100011;
									assign node3110 = (inp[4]) ? node3116 : node3111;
										assign node3111 = (inp[8]) ? 11'b00100110001 : node3112;
											assign node3112 = (inp[9]) ? 11'b00101110011 : 11'b00001100011;
										assign node3116 = (inp[9]) ? 11'b00010100111 : node3117;
											assign node3117 = (inp[8]) ? 11'b00111110011 : 11'b00110110011;
								assign node3121 = (inp[11]) ? node3139 : node3122;
									assign node3122 = (inp[3]) ? node3132 : node3123;
										assign node3123 = (inp[9]) ? node3129 : node3124;
											assign node3124 = (inp[8]) ? 11'b00101110111 : node3125;
												assign node3125 = (inp[4]) ? 11'b00000110101 : 11'b00001100101;
											assign node3129 = (inp[8]) ? 11'b00000110011 : 11'b00100110001;
										assign node3132 = (inp[9]) ? node3136 : node3133;
											assign node3133 = (inp[8]) ? 11'b00111100001 : 11'b00100100001;
											assign node3136 = (inp[8]) ? 11'b00000100011 : 11'b00001100001;
									assign node3139 = (inp[4]) ? node3151 : node3140;
										assign node3140 = (inp[8]) ? node3146 : node3141;
											assign node3141 = (inp[9]) ? 11'b00011100001 : node3142;
												assign node3142 = (inp[3]) ? 11'b00101100001 : 11'b00001110101;
											assign node3146 = (inp[3]) ? node3148 : 11'b00100100001;
												assign node3148 = (inp[9]) ? 11'b00011100011 : 11'b00110100011;
										assign node3151 = (inp[8]) ? node3157 : node3152;
											assign node3152 = (inp[3]) ? node3154 : 11'b00110100001;
												assign node3154 = (inp[9]) ? 11'b00000100001 : 11'b00010100001;
											assign node3157 = (inp[3]) ? 11'b00001100001 : 11'b00011100001;
						assign node3160 = (inp[0]) ? node3218 : node3161;
							assign node3161 = (inp[9]) ? node3185 : node3162;
								assign node3162 = (inp[4]) ? node3174 : node3163;
									assign node3163 = (inp[8]) ? node3169 : node3164;
										assign node3164 = (inp[10]) ? 11'b10111010011 : node3165;
											assign node3165 = (inp[3]) ? 11'b10011010011 : 11'b00010010001;
										assign node3169 = (inp[3]) ? node3171 : 11'b10001010011;
											assign node3171 = (inp[10]) ? 11'b00011000101 : 11'b10001000011;
									assign node3174 = (inp[10]) ? node3182 : node3175;
										assign node3175 = (inp[3]) ? node3179 : node3176;
											assign node3176 = (inp[8]) ? 11'b00110010101 : 11'b00011010111;
											assign node3179 = (inp[11]) ? 11'b10110010101 : 11'b10101010101;
										assign node3182 = (inp[11]) ? 11'b00100000011 : 11'b00000010011;
								assign node3185 = (inp[3]) ? node3203 : node3186;
									assign node3186 = (inp[4]) ? node3194 : node3187;
										assign node3187 = (inp[11]) ? node3191 : node3188;
											assign node3188 = (inp[8]) ? 11'b00000110001 : 11'b00011010001;
											assign node3191 = (inp[8]) ? 11'b00011000001 : 11'b00101000011;
										assign node3194 = (inp[10]) ? 11'b10100000001 : node3195;
											assign node3195 = (inp[11]) ? node3199 : node3196;
												assign node3196 = (inp[8]) ? 11'b00111010111 : 11'b00100010101;
												assign node3199 = (inp[8]) ? 11'b00110000111 : 11'b00000000111;
									assign node3203 = (inp[4]) ? node3209 : node3204;
										assign node3204 = (inp[10]) ? node3206 : 11'b10110010111;
											assign node3206 = (inp[11]) ? 11'b00100000111 : 11'b00110100111;
										assign node3209 = (inp[10]) ? node3215 : node3210;
											assign node3210 = (inp[11]) ? node3212 : 11'b10101000011;
												assign node3212 = (inp[8]) ? 11'b10110000001 : 11'b10100000011;
											assign node3215 = (inp[8]) ? 11'b00111000001 : 11'b00110000011;
							assign node3218 = (inp[3]) ? node3246 : node3219;
								assign node3219 = (inp[8]) ? node3233 : node3220;
									assign node3220 = (inp[11]) ? node3226 : node3221;
										assign node3221 = (inp[10]) ? 11'b00101010011 : node3222;
											assign node3222 = (inp[9]) ? 11'b00001000101 : 11'b00000100001;
										assign node3226 = (inp[4]) ? node3230 : node3227;
											assign node3227 = (inp[10]) ? 11'b00111000011 : 11'b00111010101;
											assign node3230 = (inp[10]) ? 11'b00110000001 : 11'b00110000111;
									assign node3233 = (inp[4]) ? node3239 : node3234;
										assign node3234 = (inp[10]) ? node3236 : 11'b00110100101;
											assign node3236 = (inp[9]) ? 11'b00000110011 : 11'b00010100111;
										assign node3239 = (inp[11]) ? node3241 : 11'b00001010001;
											assign node3241 = (inp[10]) ? 11'b00010000111 : node3242;
												assign node3242 = (inp[9]) ? 11'b00000000111 : 11'b00000010001;
								assign node3246 = (inp[9]) ? node3256 : node3247;
									assign node3247 = (inp[4]) ? node3253 : node3248;
										assign node3248 = (inp[10]) ? node3250 : 11'b00111000011;
											assign node3250 = (inp[8]) ? 11'b00101000001 : 11'b00111000011;
										assign node3253 = (inp[11]) ? 11'b00001010001 : 11'b00101000011;
									assign node3256 = (inp[4]) ? node3268 : node3257;
										assign node3257 = (inp[10]) ? node3261 : node3258;
											assign node3258 = (inp[11]) ? 11'b00010010011 : 11'b00100110001;
											assign node3261 = (inp[11]) ? node3265 : node3262;
												assign node3262 = (inp[8]) ? 11'b00010100011 : 11'b00011000001;
												assign node3265 = (inp[8]) ? 11'b00000000011 : 11'b00001000011;
										assign node3268 = (inp[11]) ? 11'b00010000001 : 11'b00011000001;
					assign node3271 = (inp[8]) ? node3395 : node3272;
						assign node3272 = (inp[5]) ? node3334 : node3273;
							assign node3273 = (inp[11]) ? node3303 : node3274;
								assign node3274 = (inp[4]) ? node3286 : node3275;
									assign node3275 = (inp[0]) ? node3277 : 11'b10111000011;
										assign node3277 = (inp[9]) ? node3281 : node3278;
											assign node3278 = (inp[10]) ? 11'b00001000001 : 11'b00011000011;
											assign node3281 = (inp[10]) ? 11'b00011010011 : node3282;
												assign node3282 = (inp[3]) ? 11'b00011010011 : 11'b00001000101;
									assign node3286 = (inp[9]) ? node3292 : node3287;
										assign node3287 = (inp[10]) ? node3289 : 11'b10111000101;
											assign node3289 = (inp[0]) ? 11'b00010010111 : 11'b00010000011;
										assign node3292 = (inp[0]) ? node3298 : node3293;
											assign node3293 = (inp[3]) ? node3295 : 11'b10000000001;
												assign node3295 = (inp[10]) ? 11'b00010010001 : 11'b10000010011;
											assign node3298 = (inp[3]) ? node3300 : 11'b00100010111;
												assign node3300 = (inp[10]) ? 11'b00000000001 : 11'b00110000001;
								assign node3303 = (inp[4]) ? node3313 : node3304;
									assign node3304 = (inp[0]) ? node3306 : 11'b10100010011;
										assign node3306 = (inp[3]) ? node3310 : node3307;
											assign node3307 = (inp[10]) ? 11'b00000010111 : 11'b00010010011;
											assign node3310 = (inp[10]) ? 11'b00100000001 : 11'b00010000011;
									assign node3313 = (inp[0]) ? node3327 : node3314;
										assign node3314 = (inp[9]) ? node3320 : node3315;
											assign node3315 = (inp[10]) ? node3317 : 11'b10011100100;
												assign node3317 = (inp[3]) ? 11'b00001110000 : 11'b10011110100;
											assign node3320 = (inp[10]) ? node3324 : node3321;
												assign node3321 = (inp[3]) ? 11'b10111110010 : 11'b00101110110;
												assign node3324 = (inp[3]) ? 11'b00001110000 : 11'b10001110010;
										assign node3327 = (inp[10]) ? node3329 : 11'b00001100110;
											assign node3329 = (inp[3]) ? 11'b00011100010 : node3330;
												assign node3330 = (inp[9]) ? 11'b00111100000 : 11'b00101100100;
							assign node3334 = (inp[10]) ? node3370 : node3335;
								assign node3335 = (inp[9]) ? node3351 : node3336;
									assign node3336 = (inp[3]) ? node3344 : node3337;
										assign node3337 = (inp[0]) ? node3341 : node3338;
											assign node3338 = (inp[11]) ? 11'b00111110100 : 11'b00111110000;
											assign node3341 = (inp[4]) ? 11'b00101110000 : 11'b00011110000;
										assign node3344 = (inp[4]) ? node3348 : node3345;
											assign node3345 = (inp[0]) ? 11'b00111100000 : 11'b10001100000;
											assign node3348 = (inp[0]) ? 11'b00010110010 : 11'b10010110110;
									assign node3351 = (inp[11]) ? node3361 : node3352;
										assign node3352 = (inp[4]) ? 11'b00100110100 : node3353;
											assign node3353 = (inp[3]) ? node3357 : node3354;
												assign node3354 = (inp[0]) ? 11'b00010100100 : 11'b00110110000;
												assign node3357 = (inp[0]) ? 11'b00110110000 : 11'b10100110100;
										assign node3361 = (inp[3]) ? node3367 : node3362;
											assign node3362 = (inp[4]) ? node3364 : 11'b00001100010;
												assign node3364 = (inp[0]) ? 11'b00110100100 : 11'b00100100110;
											assign node3367 = (inp[4]) ? 11'b10010100000 : 11'b10111110110;
								assign node3370 = (inp[9]) ? node3382 : node3371;
									assign node3371 = (inp[3]) ? node3377 : node3372;
										assign node3372 = (inp[0]) ? node3374 : 11'b10100100110;
											assign node3374 = (inp[4]) ? 11'b00010110100 : 11'b00110100110;
										assign node3377 = (inp[0]) ? node3379 : 11'b00010110110;
											assign node3379 = (inp[4]) ? 11'b00010100010 : 11'b00000100010;
									assign node3382 = (inp[11]) ? node3390 : node3383;
										assign node3383 = (inp[3]) ? node3385 : 11'b10101110010;
											assign node3385 = (inp[4]) ? node3387 : 11'b00110100110;
												assign node3387 = (inp[0]) ? 11'b00001100010 : 11'b00011100010;
										assign node3390 = (inp[4]) ? 11'b00000100000 : node3391;
											assign node3391 = (inp[0]) ? 11'b00001100000 : 11'b00101100100;
						assign node3395 = (inp[11]) ? node3439 : node3396;
							assign node3396 = (inp[0]) ? node3418 : node3397;
								assign node3397 = (inp[9]) ? node3405 : node3398;
									assign node3398 = (inp[4]) ? node3400 : 11'b10000100010;
										assign node3400 = (inp[5]) ? 11'b10101000110 : node3401;
											assign node3401 = (inp[10]) ? 11'b10011010100 : 11'b00011000110;
									assign node3405 = (inp[4]) ? node3411 : node3406;
										assign node3406 = (inp[3]) ? 11'b10111010100 : node3407;
											assign node3407 = (inp[5]) ? 11'b00101010010 : 11'b10111010110;
										assign node3411 = (inp[5]) ? node3413 : 11'b10111010010;
											assign node3413 = (inp[3]) ? node3415 : 11'b10001010000;
												assign node3415 = (inp[10]) ? 11'b00011000000 : 11'b10011000000;
								assign node3418 = (inp[10]) ? node3426 : node3419;
									assign node3419 = (inp[5]) ? node3423 : node3420;
										assign node3420 = (inp[3]) ? 11'b00010100010 : 11'b00100100010;
										assign node3423 = (inp[9]) ? 11'b00111010000 : 11'b00111000010;
									assign node3426 = (inp[3]) ? node3436 : node3427;
										assign node3427 = (inp[9]) ? node3433 : node3428;
											assign node3428 = (inp[4]) ? node3430 : 11'b00001000110;
												assign node3430 = (inp[5]) ? 11'b00111010110 : 11'b00101010100;
											assign node3433 = (inp[5]) ? 11'b00011010000 : 11'b00111010010;
										assign node3436 = (inp[5]) ? 11'b00101000010 : 11'b00001000010;
							assign node3439 = (inp[3]) ? node3471 : node3440;
								assign node3440 = (inp[5]) ? node3460 : node3441;
									assign node3441 = (inp[9]) ? node3451 : node3442;
										assign node3442 = (inp[0]) ? node3446 : node3443;
											assign node3443 = (inp[10]) ? 11'b10011000000 : 11'b00111000000;
											assign node3446 = (inp[4]) ? node3448 : 11'b00101010100;
												assign node3448 = (inp[10]) ? 11'b00010000110 : 11'b00110010000;
										assign node3451 = (inp[10]) ? node3457 : node3452;
											assign node3452 = (inp[4]) ? 11'b00110010110 : node3453;
												assign node3453 = (inp[0]) ? 11'b00000010110 : 11'b00010010010;
											assign node3457 = (inp[0]) ? 11'b00100000010 : 11'b10100010110;
									assign node3460 = (inp[9]) ? node3464 : node3461;
										assign node3461 = (inp[0]) ? 11'b00110010110 : 11'b10010000110;
										assign node3464 = (inp[0]) ? node3468 : node3465;
											assign node3465 = (inp[10]) ? 11'b10010000000 : 11'b00110000000;
											assign node3468 = (inp[4]) ? 11'b00010000100 : 11'b00010000000;
								assign node3471 = (inp[10]) ? node3479 : node3472;
									assign node3472 = (inp[0]) ? 11'b00110010010 : node3473;
										assign node3473 = (inp[4]) ? 11'b10110000100 : node3474;
											assign node3474 = (inp[9]) ? 11'b10000000110 : 11'b10001010000;
									assign node3479 = (inp[9]) ? node3485 : node3480;
										assign node3480 = (inp[4]) ? 11'b00000000010 : node3481;
											assign node3481 = (inp[0]) ? 11'b00100000010 : 11'b00100000110;
										assign node3485 = (inp[5]) ? node3487 : 11'b00000010000;
											assign node3487 = (inp[4]) ? 11'b00000000000 : node3488;
												assign node3488 = (inp[0]) ? 11'b00000000000 : 11'b00000000100;
				assign node3492 = (inp[2]) ? node3752 : node3493;
					assign node3493 = (inp[8]) ? node3621 : node3494;
						assign node3494 = (inp[11]) ? node3564 : node3495;
							assign node3495 = (inp[3]) ? node3533 : node3496;
								assign node3496 = (inp[9]) ? node3514 : node3497;
									assign node3497 = (inp[10]) ? node3505 : node3498;
										assign node3498 = (inp[5]) ? 11'b00001110100 : node3499;
											assign node3499 = (inp[0]) ? 11'b00011100010 : node3500;
												assign node3500 = (inp[4]) ? 11'b00011100110 : 11'b00011100010;
										assign node3505 = (inp[4]) ? node3509 : node3506;
											assign node3506 = (inp[0]) ? 11'b00111100110 : 11'b10111110010;
											assign node3509 = (inp[5]) ? 11'b10011100100 : node3510;
												assign node3510 = (inp[0]) ? 11'b00011110110 : 11'b10011110110;
									assign node3514 = (inp[5]) ? node3522 : node3515;
										assign node3515 = (inp[10]) ? node3519 : node3516;
											assign node3516 = (inp[0]) ? 11'b00111110100 : 11'b00111100100;
											assign node3519 = (inp[0]) ? 11'b00011110000 : 11'b10011110100;
										assign node3522 = (inp[10]) ? node3530 : node3523;
											assign node3523 = (inp[4]) ? node3527 : node3524;
												assign node3524 = (inp[0]) ? 11'b00011100110 : 11'b00001110010;
												assign node3527 = (inp[0]) ? 11'b00101110110 : 11'b00111110110;
											assign node3530 = (inp[4]) ? 11'b00111110010 : 11'b00111110000;
								assign node3533 = (inp[4]) ? node3547 : node3534;
									assign node3534 = (inp[9]) ? node3538 : node3535;
										assign node3535 = (inp[10]) ? 11'b00101110110 : 11'b10000110000;
										assign node3538 = (inp[5]) ? node3544 : node3539;
											assign node3539 = (inp[0]) ? node3541 : 11'b00001110100;
												assign node3541 = (inp[10]) ? 11'b00001100000 : 11'b00001110000;
											assign node3544 = (inp[0]) ? 11'b00011100000 : 11'b00011100100;
									assign node3547 = (inp[9]) ? node3555 : node3548;
										assign node3548 = (inp[10]) ? node3550 : 11'b00001110010;
											assign node3550 = (inp[5]) ? node3552 : 11'b00101100010;
												assign node3552 = (inp[0]) ? 11'b00111100010 : 11'b00001110000;
										assign node3555 = (inp[0]) ? node3561 : node3556;
											assign node3556 = (inp[5]) ? 11'b00101100010 : node3557;
												assign node3557 = (inp[10]) ? 11'b00101110000 : 11'b10101110000;
											assign node3561 = (inp[10]) ? 11'b00001100000 : 11'b00101100000;
							assign node3564 = (inp[0]) ? node3596 : node3565;
								assign node3565 = (inp[5]) ? node3579 : node3566;
									assign node3566 = (inp[10]) ? node3576 : node3567;
										assign node3567 = (inp[3]) ? node3571 : node3568;
											assign node3568 = (inp[9]) ? 11'b00010110110 : 11'b00000100100;
											assign node3571 = (inp[9]) ? 11'b10110100100 : node3572;
												assign node3572 = (inp[4]) ? 11'b10110100110 : 11'b10010110010;
										assign node3576 = (inp[3]) ? 11'b00110110010 : 11'b10110110000;
									assign node3579 = (inp[9]) ? node3585 : node3580;
										assign node3580 = (inp[4]) ? 11'b10100110110 : node3581;
											assign node3581 = (inp[10]) ? 11'b10101110000 : 11'b10111100000;
										assign node3585 = (inp[4]) ? node3593 : node3586;
											assign node3586 = (inp[10]) ? node3590 : node3587;
												assign node3587 = (inp[3]) ? 11'b10001110100 : 11'b00101100000;
												assign node3590 = (inp[3]) ? 11'b00000100110 : 11'b10110100110;
											assign node3593 = (inp[10]) ? 11'b00100100000 : 11'b10110100000;
								assign node3596 = (inp[3]) ? node3608 : node3597;
									assign node3597 = (inp[4]) ? node3603 : node3598;
										assign node3598 = (inp[9]) ? node3600 : 11'b00001110100;
											assign node3600 = (inp[10]) ? 11'b00100100010 : 11'b00101110100;
										assign node3603 = (inp[10]) ? node3605 : 11'b00000100110;
											assign node3605 = (inp[9]) ? 11'b00100100000 : 11'b00110100100;
									assign node3608 = (inp[9]) ? node3614 : node3609;
										assign node3609 = (inp[4]) ? 11'b00000110010 : node3610;
											assign node3610 = (inp[5]) ? 11'b00101100000 : 11'b00100100010;
										assign node3614 = (inp[10]) ? node3618 : node3615;
											assign node3615 = (inp[4]) ? 11'b00110100000 : 11'b00010110010;
											assign node3618 = (inp[5]) ? 11'b00000100000 : 11'b00010100000;
						assign node3621 = (inp[5]) ? node3687 : node3622;
							assign node3622 = (inp[11]) ? node3658 : node3623;
								assign node3623 = (inp[0]) ? node3643 : node3624;
									assign node3624 = (inp[4]) ? node3636 : node3625;
										assign node3625 = (inp[3]) ? node3631 : node3626;
											assign node3626 = (inp[10]) ? 11'b10000100010 : node3627;
												assign node3627 = (inp[9]) ? 11'b00000100010 : 11'b00010100010;
											assign node3631 = (inp[9]) ? 11'b00100110100 : node3632;
												assign node3632 = (inp[10]) ? 11'b00110100110 : 11'b10100100010;
										assign node3636 = (inp[9]) ? node3640 : node3637;
											assign node3637 = (inp[3]) ? 11'b10010100100 : 11'b10100110100;
											assign node3640 = (inp[3]) ? 11'b10001010010 : 11'b00101000110;
									assign node3643 = (inp[3]) ? node3649 : node3644;
										assign node3644 = (inp[4]) ? node3646 : 11'b00100110000;
											assign node3646 = (inp[9]) ? 11'b00011010010 : 11'b00110100000;
										assign node3649 = (inp[10]) ? node3655 : node3650;
											assign node3650 = (inp[9]) ? 11'b00010110000 : node3651;
												assign node3651 = (inp[4]) ? 11'b00000110000 : 11'b00000100010;
											assign node3655 = (inp[4]) ? 11'b00001000010 : 11'b00000100000;
								assign node3658 = (inp[0]) ? node3674 : node3659;
									assign node3659 = (inp[10]) ? node3669 : node3660;
										assign node3660 = (inp[3]) ? node3666 : node3661;
											assign node3661 = (inp[9]) ? 11'b00111010000 : node3662;
												assign node3662 = (inp[4]) ? 11'b00101000110 : 11'b00001000010;
											assign node3666 = (inp[9]) ? 11'b10101000100 : 11'b10111010000;
										assign node3669 = (inp[4]) ? node3671 : 11'b00111010110;
											assign node3671 = (inp[9]) ? 11'b00101010000 : 11'b00101010010;
									assign node3674 = (inp[3]) ? node3676 : 11'b00101010100;
										assign node3676 = (inp[9]) ? node3682 : node3677;
											assign node3677 = (inp[4]) ? 11'b00111010010 : node3678;
												assign node3678 = (inp[10]) ? 11'b00111000000 : 11'b00011000000;
											assign node3682 = (inp[4]) ? node3684 : 11'b00011000010;
												assign node3684 = (inp[10]) ? 11'b00001000000 : 11'b00111000000;
							assign node3687 = (inp[4]) ? node3717 : node3688;
								assign node3688 = (inp[3]) ? node3704 : node3689;
									assign node3689 = (inp[9]) ? node3695 : node3690;
										assign node3690 = (inp[11]) ? node3692 : 11'b00001000100;
											assign node3692 = (inp[10]) ? 11'b00100010110 : 11'b00000010000;
										assign node3695 = (inp[11]) ? node3697 : 11'b00010010010;
											assign node3697 = (inp[0]) ? node3701 : node3698;
												assign node3698 = (inp[10]) ? 11'b10100000110 : 11'b00000000010;
												assign node3701 = (inp[10]) ? 11'b00000000010 : 11'b00010010110;
									assign node3704 = (inp[0]) ? node3710 : node3705;
										assign node3705 = (inp[9]) ? node3707 : 11'b10010000010;
											assign node3707 = (inp[11]) ? 11'b00100000110 : 11'b00110000110;
										assign node3710 = (inp[11]) ? node3714 : node3711;
											assign node3711 = (inp[10]) ? 11'b00010000010 : 11'b00100010010;
											assign node3714 = (inp[10]) ? 11'b00100000010 : 11'b00110000010;
								assign node3717 = (inp[0]) ? node3737 : node3718;
									assign node3718 = (inp[10]) ? node3726 : node3719;
										assign node3719 = (inp[11]) ? node3721 : 11'b10000010110;
											assign node3721 = (inp[9]) ? 11'b00110000100 : node3722;
												assign node3722 = (inp[3]) ? 11'b10110010100 : 11'b00110010100;
										assign node3726 = (inp[3]) ? node3732 : node3727;
											assign node3727 = (inp[9]) ? 11'b10110010000 : node3728;
												assign node3728 = (inp[11]) ? 11'b10100000100 : 11'b10010000100;
											assign node3732 = (inp[9]) ? 11'b00100000000 : node3733;
												assign node3733 = (inp[11]) ? 11'b00100000000 : 11'b00010010000;
									assign node3737 = (inp[3]) ? node3749 : node3738;
										assign node3738 = (inp[10]) ? node3744 : node3739;
											assign node3739 = (inp[11]) ? 11'b00010010000 : node3740;
												assign node3740 = (inp[9]) ? 11'b00000010100 : 11'b00000000010;
											assign node3744 = (inp[11]) ? 11'b00000000100 : node3745;
												assign node3745 = (inp[9]) ? 11'b00010010000 : 11'b00110010100;
										assign node3749 = (inp[10]) ? 11'b00000000000 : 11'b00010000000;
					assign node3752 = (inp[8]) ? node3890 : node3753;
						assign node3753 = (inp[5]) ? node3819 : node3754;
							assign node3754 = (inp[4]) ? node3786 : node3755;
								assign node3755 = (inp[0]) ? node3775 : node3756;
									assign node3756 = (inp[9]) ? node3766 : node3757;
										assign node3757 = (inp[11]) ? node3761 : node3758;
											assign node3758 = (inp[3]) ? 11'b10111000010 : 11'b00111000010;
											assign node3761 = (inp[3]) ? node3763 : 11'b10111000010;
												assign node3763 = (inp[10]) ? 11'b00101010110 : 11'b10111010010;
										assign node3766 = (inp[11]) ? node3770 : node3767;
											assign node3767 = (inp[3]) ? 11'b00101010110 : 11'b00111000010;
											assign node3770 = (inp[10]) ? 11'b10011010110 : node3771;
												assign node3771 = (inp[3]) ? 11'b10001000110 : 11'b00001010010;
									assign node3775 = (inp[10]) ? node3777 : 11'b00011000010;
										assign node3777 = (inp[11]) ? node3783 : node3778;
											assign node3778 = (inp[9]) ? 11'b00001010010 : node3779;
												assign node3779 = (inp[3]) ? 11'b00001000010 : 11'b00001000110;
											assign node3783 = (inp[9]) ? 11'b00011000010 : 11'b00011010110;
								assign node3786 = (inp[10]) ? node3806 : node3787;
									assign node3787 = (inp[11]) ? node3801 : node3788;
										assign node3788 = (inp[0]) ? node3794 : node3789;
											assign node3789 = (inp[9]) ? 11'b10011010000 : node3790;
												assign node3790 = (inp[3]) ? 11'b10111000100 : 11'b00111000100;
											assign node3794 = (inp[9]) ? node3798 : node3795;
												assign node3795 = (inp[3]) ? 11'b00011010000 : 11'b00011000000;
												assign node3798 = (inp[3]) ? 11'b00111000000 : 11'b00111010100;
										assign node3801 = (inp[9]) ? 11'b00011000100 : node3802;
											assign node3802 = (inp[3]) ? 11'b00101010010 : 11'b00001010010;
									assign node3806 = (inp[3]) ? node3814 : node3807;
										assign node3807 = (inp[0]) ? node3811 : node3808;
											assign node3808 = (inp[9]) ? 11'b10011000000 : 11'b10001010110;
											assign node3811 = (inp[9]) ? 11'b00101010000 : 11'b00001010100;
										assign node3814 = (inp[0]) ? node3816 : 11'b00001010000;
											assign node3816 = (inp[9]) ? 11'b00001000000 : 11'b00101000000;
							assign node3819 = (inp[11]) ? node3855 : node3820;
								assign node3820 = (inp[4]) ? node3838 : node3821;
									assign node3821 = (inp[9]) ? node3829 : node3822;
										assign node3822 = (inp[0]) ? 11'b00101000100 : node3823;
											assign node3823 = (inp[10]) ? node3825 : 11'b10111010000;
												assign node3825 = (inp[3]) ? 11'b00001010100 : 11'b10011010000;
										assign node3829 = (inp[10]) ? node3831 : 11'b00101010000;
											assign node3831 = (inp[0]) ? node3835 : node3832;
												assign node3832 = (inp[3]) ? 11'b00110000110 : 11'b10010000110;
												assign node3835 = (inp[3]) ? 11'b00010000010 : 11'b00110010010;
									assign node3838 = (inp[0]) ? node3844 : node3839;
										assign node3839 = (inp[10]) ? node3841 : 11'b10000010110;
											assign node3841 = (inp[3]) ? 11'b00110010010 : 11'b10100010010;
										assign node3844 = (inp[9]) ? node3850 : node3845;
											assign node3845 = (inp[10]) ? 11'b00110000010 : node3846;
												assign node3846 = (inp[3]) ? 11'b00100010010 : 11'b00100000010;
											assign node3850 = (inp[10]) ? node3852 : 11'b00110010110;
												assign node3852 = (inp[3]) ? 11'b00000000010 : 11'b00100010010;
								assign node3855 = (inp[9]) ? node3875 : node3856;
									assign node3856 = (inp[10]) ? node3870 : node3857;
										assign node3857 = (inp[4]) ? node3865 : node3858;
											assign node3858 = (inp[3]) ? node3862 : node3859;
												assign node3859 = (inp[0]) ? 11'b00000010010 : 11'b00100010010;
												assign node3862 = (inp[0]) ? 11'b00110000000 : 11'b10000000010;
											assign node3865 = (inp[3]) ? 11'b10010010100 : node3866;
												assign node3866 = (inp[0]) ? 11'b00110010000 : 11'b00110010100;
										assign node3870 = (inp[0]) ? node3872 : 11'b00110000100;
											assign node3872 = (inp[3]) ? 11'b00010000000 : 11'b00110000100;
									assign node3875 = (inp[0]) ? node3883 : node3876;
										assign node3876 = (inp[3]) ? 11'b00100000100 : node3877;
											assign node3877 = (inp[10]) ? node3879 : 11'b00100000100;
												assign node3879 = (inp[4]) ? 11'b10100000000 : 11'b10000000100;
										assign node3883 = (inp[3]) ? node3887 : node3884;
											assign node3884 = (inp[4]) ? 11'b00100000000 : 11'b00100010100;
											assign node3887 = (inp[10]) ? 11'b00000000000 : 11'b00000010000;
						assign node3890 = (inp[0]) ? node3946 : node3891;
							assign node3891 = (inp[4]) ? node3921 : node3892;
								assign node3892 = (inp[5]) ? node3908 : node3893;
									assign node3893 = (inp[9]) ? node3901 : node3894;
										assign node3894 = (inp[11]) ? node3898 : node3895;
											assign node3895 = (inp[3]) ? 11'b00010000110 : 11'b10110000010;
											assign node3898 = (inp[3]) ? 11'b10000010010 : 11'b10000000010;
										assign node3901 = (inp[11]) ? node3905 : node3902;
											assign node3902 = (inp[10]) ? 11'b00000010110 : 11'b10000000110;
											assign node3905 = (inp[10]) ? 11'b00010010100 : 11'b00010010000;
									assign node3908 = (inp[10]) ? node3914 : node3909;
										assign node3909 = (inp[9]) ? 11'b10110010100 : node3910;
											assign node3910 = (inp[3]) ? 11'b10110010000 : 11'b00110010000;
										assign node3914 = (inp[3]) ? node3918 : node3915;
											assign node3915 = (inp[11]) ? 11'b10000000100 : 11'b10110000100;
											assign node3918 = (inp[11]) ? 11'b00000000100 : 11'b00010000100;
								assign node3921 = (inp[10]) ? node3937 : node3922;
									assign node3922 = (inp[3]) ? node3928 : node3923;
										assign node3923 = (inp[9]) ? node3925 : 11'b00010000100;
											assign node3925 = (inp[11]) ? 11'b00100010100 : 11'b00000010100;
										assign node3928 = (inp[9]) ? 11'b10000000000 : node3929;
											assign node3929 = (inp[5]) ? node3933 : node3930;
												assign node3930 = (inp[11]) ? 11'b10100000100 : 11'b10110000110;
												assign node3933 = (inp[11]) ? 11'b10000010100 : 11'b10100010100;
									assign node3937 = (inp[3]) ? node3943 : node3938;
										assign node3938 = (inp[11]) ? node3940 : 11'b10000010000;
											assign node3940 = (inp[5]) ? 11'b10000000000 : 11'b10000010000;
										assign node3943 = (inp[5]) ? 11'b00000000000 : 11'b00000010000;
							assign node3946 = (inp[5]) ? node3976 : node3947;
								assign node3947 = (inp[11]) ? node3963 : node3948;
									assign node3948 = (inp[3]) ? node3956 : node3949;
										assign node3949 = (inp[4]) ? node3953 : node3950;
											assign node3950 = (inp[10]) ? 11'b00110000110 : 11'b00100000110;
											assign node3953 = (inp[9]) ? 11'b00010010110 : 11'b00110010110;
										assign node3956 = (inp[9]) ? node3960 : node3957;
											assign node3957 = (inp[4]) ? 11'b00010010010 : 11'b00010000010;
											assign node3960 = (inp[10]) ? 11'b00000000010 : 11'b00000010010;
									assign node3963 = (inp[10]) ? node3971 : node3964;
										assign node3964 = (inp[9]) ? node3968 : node3965;
											assign node3965 = (inp[4]) ? 11'b00100010000 : 11'b00100010010;
											assign node3968 = (inp[3]) ? 11'b00110010000 : 11'b00010010100;
										assign node3971 = (inp[4]) ? 11'b00000000000 : node3972;
											assign node3972 = (inp[3]) ? 11'b00010000000 : 11'b00110000000;
								assign node3976 = (inp[11]) ? node3994 : node3977;
									assign node3977 = (inp[4]) ? node3985 : node3978;
										assign node3978 = (inp[10]) ? node3982 : node3979;
											assign node3979 = (inp[3]) ? 11'b00110010000 : 11'b00110000100;
											assign node3982 = (inp[9]) ? 11'b00010010000 : 11'b00010000000;
										assign node3985 = (inp[3]) ? node3989 : node3986;
											assign node3986 = (inp[10]) ? 11'b00100010100 : 11'b00000010100;
											assign node3989 = (inp[9]) ? 11'b00000000000 : node3990;
												assign node3990 = (inp[10]) ? 11'b00100000000 : 11'b00100010000;
									assign node3994 = (inp[9]) ? node4000 : node3995;
										assign node3995 = (inp[3]) ? node3997 : 11'b00000000100;
											assign node3997 = (inp[4]) ? 11'b00000000000 : 11'b00100000000;
										assign node4000 = (inp[10]) ? 11'b00000000000 : node4001;
											assign node4001 = (inp[4]) ? 11'b00000000000 : 11'b00000010000;

endmodule