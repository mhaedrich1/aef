module dtc_split125_bm88 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node80;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node111;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node194;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node206;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node264;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node283;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node289;
	wire [3-1:0] node293;
	wire [3-1:0] node295;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node319;
	wire [3-1:0] node322;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node334;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node381;

	assign outp = (inp[6]) ? node128 : node1;
		assign node1 = (inp[9]) ? node91 : node2;
			assign node2 = (inp[3]) ? node60 : node3;
				assign node3 = (inp[0]) ? node27 : node4;
					assign node4 = (inp[5]) ? node14 : node5;
						assign node5 = (inp[2]) ? 3'b000 : node6;
							assign node6 = (inp[11]) ? node8 : 3'b000;
								assign node8 = (inp[4]) ? 3'b000 : node9;
									assign node9 = (inp[8]) ? 3'b000 : 3'b010;
						assign node14 = (inp[10]) ? node20 : node15;
							assign node15 = (inp[11]) ? 3'b000 : node16;
								assign node16 = (inp[8]) ? 3'b000 : 3'b010;
							assign node20 = (inp[1]) ? node22 : 3'b110;
								assign node22 = (inp[7]) ? node24 : 3'b010;
									assign node24 = (inp[4]) ? 3'b000 : 3'b010;
					assign node27 = (inp[11]) ? node43 : node28;
						assign node28 = (inp[10]) ? node38 : node29;
							assign node29 = (inp[7]) ? node31 : 3'b110;
								assign node31 = (inp[4]) ? 3'b111 : node32;
									assign node32 = (inp[1]) ? 3'b001 : node33;
										assign node33 = (inp[2]) ? 3'b001 : 3'b010;
							assign node38 = (inp[5]) ? node40 : 3'b000;
								assign node40 = (inp[8]) ? 3'b000 : 3'b100;
						assign node43 = (inp[4]) ? node55 : node44;
							assign node44 = (inp[5]) ? node50 : node45;
								assign node45 = (inp[1]) ? 3'b110 : node46;
									assign node46 = (inp[10]) ? 3'b100 : 3'b010;
								assign node50 = (inp[1]) ? 3'b100 : node51;
									assign node51 = (inp[10]) ? 3'b000 : 3'b100;
							assign node55 = (inp[10]) ? 3'b000 : node56;
								assign node56 = (inp[7]) ? 3'b000 : 3'b100;
				assign node60 = (inp[7]) ? node70 : node61;
					assign node61 = (inp[10]) ? 3'b000 : node62;
						assign node62 = (inp[11]) ? 3'b000 : node63;
							assign node63 = (inp[2]) ? 3'b000 : node64;
								assign node64 = (inp[1]) ? 3'b000 : 3'b100;
					assign node70 = (inp[8]) ? node84 : node71;
						assign node71 = (inp[4]) ? 3'b000 : node72;
							assign node72 = (inp[1]) ? node80 : node73;
								assign node73 = (inp[0]) ? 3'b000 : node74;
									assign node74 = (inp[10]) ? 3'b000 : node75;
										assign node75 = (inp[5]) ? 3'b010 : 3'b000;
								assign node80 = (inp[5]) ? 3'b100 : 3'b010;
						assign node84 = (inp[0]) ? node86 : 3'b100;
							assign node86 = (inp[2]) ? 3'b000 : node87;
								assign node87 = (inp[10]) ? 3'b100 : 3'b000;
			assign node91 = (inp[8]) ? node93 : 3'b000;
				assign node93 = (inp[7]) ? node101 : node94;
					assign node94 = (inp[1]) ? node96 : 3'b000;
						assign node96 = (inp[10]) ? 3'b000 : node97;
							assign node97 = (inp[11]) ? 3'b000 : 3'b100;
					assign node101 = (inp[11]) ? node121 : node102;
						assign node102 = (inp[3]) ? node114 : node103;
							assign node103 = (inp[0]) ? node105 : 3'b000;
								assign node105 = (inp[1]) ? node111 : node106;
									assign node106 = (inp[10]) ? 3'b110 : node107;
										assign node107 = (inp[5]) ? 3'b010 : 3'b110;
									assign node111 = (inp[4]) ? 3'b000 : 3'b100;
							assign node114 = (inp[10]) ? 3'b000 : node115;
								assign node115 = (inp[0]) ? node117 : 3'b000;
									assign node117 = (inp[4]) ? 3'b000 : 3'b010;
						assign node121 = (inp[10]) ? 3'b000 : node122;
							assign node122 = (inp[0]) ? 3'b000 : node123;
								assign node123 = (inp[3]) ? 3'b100 : 3'b000;
		assign node128 = (inp[3]) ? node238 : node129;
			assign node129 = (inp[0]) ? node161 : node130;
				assign node130 = (inp[7]) ? node140 : node131;
					assign node131 = (inp[8]) ? 3'b001 : node132;
						assign node132 = (inp[5]) ? node134 : 3'b001;
							assign node134 = (inp[9]) ? 3'b000 : node135;
								assign node135 = (inp[11]) ? 3'b000 : 3'b001;
					assign node140 = (inp[5]) ? node152 : node141;
						assign node141 = (inp[11]) ? node143 : 3'b111;
							assign node143 = (inp[1]) ? 3'b011 : node144;
								assign node144 = (inp[8]) ? node148 : node145;
									assign node145 = (inp[2]) ? 3'b111 : 3'b101;
									assign node148 = (inp[2]) ? 3'b011 : 3'b111;
						assign node152 = (inp[8]) ? node154 : 3'b000;
							assign node154 = (inp[2]) ? node156 : 3'b011;
								assign node156 = (inp[1]) ? node158 : 3'b011;
									assign node158 = (inp[4]) ? 3'b101 : 3'b111;
				assign node161 = (inp[7]) ? node199 : node162;
					assign node162 = (inp[10]) ? node188 : node163;
						assign node163 = (inp[5]) ? node175 : node164;
							assign node164 = (inp[8]) ? node172 : node165;
								assign node165 = (inp[4]) ? node169 : node166;
									assign node166 = (inp[11]) ? 3'b111 : 3'b011;
									assign node169 = (inp[11]) ? 3'b011 : 3'b001;
								assign node172 = (inp[9]) ? 3'b111 : 3'b101;
							assign node175 = (inp[4]) ? node179 : node176;
								assign node176 = (inp[11]) ? 3'b111 : 3'b101;
								assign node179 = (inp[1]) ? node185 : node180;
									assign node180 = (inp[8]) ? 3'b011 : node181;
										assign node181 = (inp[9]) ? 3'b110 : 3'b010;
									assign node185 = (inp[2]) ? 3'b110 : 3'b100;
						assign node188 = (inp[4]) ? node194 : node189;
							assign node189 = (inp[11]) ? 3'b010 : node190;
								assign node190 = (inp[1]) ? 3'b110 : 3'b100;
							assign node194 = (inp[8]) ? node196 : 3'b110;
								assign node196 = (inp[11]) ? 3'b100 : 3'b110;
					assign node199 = (inp[4]) ? node219 : node200;
						assign node200 = (inp[10]) ? node210 : node201;
							assign node201 = (inp[5]) ? node203 : 3'b011;
								assign node203 = (inp[1]) ? 3'b111 : node204;
									assign node204 = (inp[8]) ? node206 : 3'b111;
										assign node206 = (inp[9]) ? 3'b011 : 3'b111;
							assign node210 = (inp[2]) ? 3'b101 : node211;
								assign node211 = (inp[9]) ? 3'b110 : node212;
									assign node212 = (inp[5]) ? node214 : 3'b101;
										assign node214 = (inp[1]) ? 3'b011 : 3'b111;
						assign node219 = (inp[1]) ? node225 : node220;
							assign node220 = (inp[8]) ? node222 : 3'b001;
								assign node222 = (inp[9]) ? 3'b001 : 3'b011;
							assign node225 = (inp[8]) ? node229 : node226;
								assign node226 = (inp[10]) ? 3'b100 : 3'b101;
								assign node229 = (inp[10]) ? node233 : node230;
									assign node230 = (inp[9]) ? 3'b001 : 3'b011;
									assign node233 = (inp[9]) ? 3'b110 : node234;
										assign node234 = (inp[2]) ? 3'b101 : 3'b001;
			assign node238 = (inp[7]) ? node302 : node239;
				assign node239 = (inp[0]) ? node275 : node240;
					assign node240 = (inp[10]) ? node260 : node241;
						assign node241 = (inp[1]) ? node245 : node242;
							assign node242 = (inp[4]) ? 3'b010 : 3'b000;
							assign node245 = (inp[4]) ? node257 : node246;
								assign node246 = (inp[9]) ? node254 : node247;
									assign node247 = (inp[5]) ? node249 : 3'b110;
										assign node249 = (inp[8]) ? node251 : 3'b010;
											assign node251 = (inp[2]) ? 3'b110 : 3'b010;
									assign node254 = (inp[11]) ? 3'b010 : 3'b000;
								assign node257 = (inp[9]) ? 3'b010 : 3'b000;
						assign node260 = (inp[8]) ? node268 : node261;
							assign node261 = (inp[11]) ? 3'b100 : node262;
								assign node262 = (inp[5]) ? node264 : 3'b010;
									assign node264 = (inp[9]) ? 3'b100 : 3'b110;
							assign node268 = (inp[11]) ? node272 : node269;
								assign node269 = (inp[5]) ? 3'b010 : 3'b000;
								assign node272 = (inp[5]) ? 3'b100 : 3'b000;
					assign node275 = (inp[9]) ? node293 : node276;
						assign node276 = (inp[10]) ? node286 : node277;
							assign node277 = (inp[2]) ? node283 : node278;
								assign node278 = (inp[5]) ? 3'b010 : node279;
									assign node279 = (inp[4]) ? 3'b010 : 3'b100;
								assign node283 = (inp[8]) ? 3'b100 : 3'b110;
							assign node286 = (inp[11]) ? 3'b000 : node287;
								assign node287 = (inp[1]) ? node289 : 3'b100;
									assign node289 = (inp[4]) ? 3'b000 : 3'b100;
						assign node293 = (inp[2]) ? node295 : 3'b000;
							assign node295 = (inp[11]) ? node297 : 3'b100;
								assign node297 = (inp[10]) ? 3'b000 : node298;
									assign node298 = (inp[5]) ? 3'b000 : 3'b100;
				assign node302 = (inp[10]) ? node342 : node303;
					assign node303 = (inp[4]) ? node327 : node304;
						assign node304 = (inp[8]) ? node312 : node305;
							assign node305 = (inp[5]) ? node309 : node306;
								assign node306 = (inp[11]) ? 3'b001 : 3'b101;
								assign node309 = (inp[0]) ? 3'b000 : 3'b110;
							assign node312 = (inp[5]) ? node322 : node313;
								assign node313 = (inp[1]) ? node319 : node314;
									assign node314 = (inp[0]) ? 3'b011 : node315;
										assign node315 = (inp[11]) ? 3'b101 : 3'b011;
									assign node319 = (inp[2]) ? 3'b111 : 3'b101;
								assign node322 = (inp[1]) ? node324 : 3'b101;
									assign node324 = (inp[9]) ? 3'b001 : 3'b011;
						assign node327 = (inp[0]) ? node339 : node328;
							assign node328 = (inp[9]) ? node334 : node329;
								assign node329 = (inp[1]) ? 3'b001 : node330;
									assign node330 = (inp[11]) ? 3'b101 : 3'b000;
								assign node334 = (inp[5]) ? node336 : 3'b000;
									assign node336 = (inp[1]) ? 3'b010 : 3'b110;
							assign node339 = (inp[2]) ? 3'b100 : 3'b110;
					assign node342 = (inp[0]) ? node364 : node343;
						assign node343 = (inp[11]) ? node353 : node344;
							assign node344 = (inp[5]) ? node348 : node345;
								assign node345 = (inp[9]) ? 3'b110 : 3'b101;
								assign node348 = (inp[2]) ? 3'b001 : node349;
									assign node349 = (inp[4]) ? 3'b001 : 3'b011;
							assign node353 = (inp[9]) ? node359 : node354;
								assign node354 = (inp[8]) ? 3'b101 : node355;
									assign node355 = (inp[4]) ? 3'b110 : 3'b101;
								assign node359 = (inp[1]) ? 3'b110 : node360;
									assign node360 = (inp[2]) ? 3'b110 : 3'b010;
						assign node364 = (inp[9]) ? node378 : node365;
							assign node365 = (inp[4]) ? node373 : node366;
								assign node366 = (inp[1]) ? 3'b110 : node367;
									assign node367 = (inp[5]) ? 3'b010 : node368;
										assign node368 = (inp[8]) ? 3'b101 : 3'b001;
								assign node373 = (inp[11]) ? 3'b010 : node374;
									assign node374 = (inp[2]) ? 3'b010 : 3'b110;
							assign node378 = (inp[1]) ? 3'b000 : node379;
								assign node379 = (inp[11]) ? node381 : 3'b010;
									assign node381 = (inp[8]) ? 3'b110 : 3'b010;

endmodule