module dtc_split125_bm93 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node47;
	wire [3-1:0] node49;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node92;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node101;

	assign outp = (inp[0]) ? node24 : node1;
		assign node1 = (inp[7]) ? 3'b000 : node2;
			assign node2 = (inp[3]) ? node4 : 3'b000;
				assign node4 = (inp[6]) ? 3'b000 : node5;
					assign node5 = (inp[5]) ? node11 : node6;
						assign node6 = (inp[8]) ? 3'b000 : node7;
							assign node7 = (inp[4]) ? 3'b100 : 3'b000;
						assign node11 = (inp[8]) ? node17 : node12;
							assign node12 = (inp[4]) ? node14 : 3'b010;
								assign node14 = (inp[11]) ? 3'b100 : 3'b010;
							assign node17 = (inp[2]) ? 3'b100 : node18;
								assign node18 = (inp[4]) ? 3'b000 : 3'b100;
		assign node24 = (inp[3]) ? node70 : node25;
			assign node25 = (inp[5]) ? node35 : node26;
				assign node26 = (inp[8]) ? 3'b000 : node27;
					assign node27 = (inp[7]) ? 3'b000 : node28;
						assign node28 = (inp[6]) ? 3'b000 : node29;
							assign node29 = (inp[4]) ? 3'b110 : 3'b000;
				assign node35 = (inp[7]) ? node53 : node36;
					assign node36 = (inp[6]) ? 3'b100 : node37;
						assign node37 = (inp[8]) ? node47 : node38;
							assign node38 = (inp[2]) ? 3'b100 : node39;
								assign node39 = (inp[9]) ? 3'b000 : node40;
									assign node40 = (inp[11]) ? 3'b000 : node41;
										assign node41 = (inp[10]) ? 3'b100 : 3'b110;
							assign node47 = (inp[4]) ? node49 : 3'b110;
								assign node49 = (inp[10]) ? 3'b110 : 3'b100;
					assign node53 = (inp[2]) ? node55 : 3'b000;
						assign node55 = (inp[1]) ? node57 : 3'b000;
							assign node57 = (inp[11]) ? node65 : node58;
								assign node58 = (inp[4]) ? node60 : 3'b100;
									assign node60 = (inp[8]) ? 3'b100 : node61;
										assign node61 = (inp[10]) ? 3'b100 : 3'b000;
								assign node65 = (inp[8]) ? 3'b000 : node66;
									assign node66 = (inp[6]) ? 3'b000 : 3'b100;
			assign node70 = (inp[7]) ? node92 : node71;
				assign node71 = (inp[5]) ? node81 : node72;
					assign node72 = (inp[4]) ? node74 : 3'b011;
						assign node74 = (inp[10]) ? node76 : 3'b011;
							assign node76 = (inp[6]) ? 3'b011 : node77;
								assign node77 = (inp[8]) ? 3'b011 : 3'b111;
					assign node81 = (inp[6]) ? 3'b110 : node82;
						assign node82 = (inp[2]) ? 3'b111 : node83;
							assign node83 = (inp[9]) ? 3'b011 : node84;
								assign node84 = (inp[11]) ? node86 : 3'b111;
									assign node86 = (inp[1]) ? 3'b111 : 3'b011;
				assign node92 = (inp[5]) ? node94 : 3'b000;
					assign node94 = (inp[6]) ? 3'b000 : node95;
						assign node95 = (inp[8]) ? node101 : node96;
							assign node96 = (inp[9]) ? node98 : 3'b011;
								assign node98 = (inp[1]) ? 3'b111 : 3'b011;
							assign node101 = (inp[11]) ? 3'b011 : 3'b001;

endmodule