module dtc_split875_bm78 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node195;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node204;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node227;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node278;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node285;
	wire [3-1:0] node287;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node343;
	wire [3-1:0] node346;
	wire [3-1:0] node348;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node362;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node383;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node399;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node405;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node412;
	wire [3-1:0] node414;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node423;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node436;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node445;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node456;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node478;
	wire [3-1:0] node481;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node497;
	wire [3-1:0] node499;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node506;
	wire [3-1:0] node509;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node514;
	wire [3-1:0] node516;
	wire [3-1:0] node519;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node536;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node545;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node553;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node575;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node605;
	wire [3-1:0] node607;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node612;
	wire [3-1:0] node613;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node644;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node654;
	wire [3-1:0] node657;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node669;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node683;
	wire [3-1:0] node687;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node695;
	wire [3-1:0] node696;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node708;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node714;
	wire [3-1:0] node717;
	wire [3-1:0] node719;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node728;
	wire [3-1:0] node731;
	wire [3-1:0] node733;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node741;
	wire [3-1:0] node745;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node752;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node770;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node791;
	wire [3-1:0] node793;
	wire [3-1:0] node796;
	wire [3-1:0] node798;
	wire [3-1:0] node800;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node819;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node827;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node834;
	wire [3-1:0] node836;
	wire [3-1:0] node839;
	wire [3-1:0] node841;
	wire [3-1:0] node843;
	wire [3-1:0] node845;
	wire [3-1:0] node848;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node855;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node861;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node868;
	wire [3-1:0] node872;
	wire [3-1:0] node874;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node887;
	wire [3-1:0] node889;
	wire [3-1:0] node891;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node897;
	wire [3-1:0] node900;
	wire [3-1:0] node903;
	wire [3-1:0] node905;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node913;
	wire [3-1:0] node916;
	wire [3-1:0] node918;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node925;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node940;
	wire [3-1:0] node942;
	wire [3-1:0] node943;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node951;
	wire [3-1:0] node953;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node967;
	wire [3-1:0] node969;
	wire [3-1:0] node971;
	wire [3-1:0] node973;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node982;
	wire [3-1:0] node984;
	wire [3-1:0] node986;
	wire [3-1:0] node989;
	wire [3-1:0] node990;
	wire [3-1:0] node993;
	wire [3-1:0] node994;
	wire [3-1:0] node998;
	wire [3-1:0] node1000;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1017;
	wire [3-1:0] node1018;
	wire [3-1:0] node1019;
	wire [3-1:0] node1020;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1027;
	wire [3-1:0] node1030;
	wire [3-1:0] node1033;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1045;
	wire [3-1:0] node1046;
	wire [3-1:0] node1050;
	wire [3-1:0] node1051;
	wire [3-1:0] node1052;
	wire [3-1:0] node1056;
	wire [3-1:0] node1057;
	wire [3-1:0] node1062;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1065;
	wire [3-1:0] node1066;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1074;
	wire [3-1:0] node1077;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1083;
	wire [3-1:0] node1084;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1090;
	wire [3-1:0] node1092;
	wire [3-1:0] node1095;
	wire [3-1:0] node1097;
	wire [3-1:0] node1100;
	wire [3-1:0] node1101;
	wire [3-1:0] node1103;
	wire [3-1:0] node1106;
	wire [3-1:0] node1108;
	wire [3-1:0] node1111;
	wire [3-1:0] node1112;
	wire [3-1:0] node1116;
	wire [3-1:0] node1117;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1121;
	wire [3-1:0] node1123;
	wire [3-1:0] node1125;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1132;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1136;
	wire [3-1:0] node1137;
	wire [3-1:0] node1138;
	wire [3-1:0] node1140;
	wire [3-1:0] node1143;
	wire [3-1:0] node1145;
	wire [3-1:0] node1151;
	wire [3-1:0] node1152;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1155;
	wire [3-1:0] node1156;
	wire [3-1:0] node1158;
	wire [3-1:0] node1160;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1168;
	wire [3-1:0] node1169;
	wire [3-1:0] node1170;
	wire [3-1:0] node1173;
	wire [3-1:0] node1175;
	wire [3-1:0] node1178;
	wire [3-1:0] node1180;
	wire [3-1:0] node1182;
	wire [3-1:0] node1185;
	wire [3-1:0] node1187;
	wire [3-1:0] node1189;
	wire [3-1:0] node1192;
	wire [3-1:0] node1193;
	wire [3-1:0] node1194;
	wire [3-1:0] node1195;
	wire [3-1:0] node1196;
	wire [3-1:0] node1199;
	wire [3-1:0] node1202;
	wire [3-1:0] node1203;
	wire [3-1:0] node1206;
	wire [3-1:0] node1209;
	wire [3-1:0] node1210;
	wire [3-1:0] node1211;
	wire [3-1:0] node1212;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;
	wire [3-1:0] node1220;
	wire [3-1:0] node1223;
	wire [3-1:0] node1224;
	wire [3-1:0] node1226;
	wire [3-1:0] node1229;
	wire [3-1:0] node1231;
	wire [3-1:0] node1234;
	wire [3-1:0] node1235;
	wire [3-1:0] node1236;
	wire [3-1:0] node1238;
	wire [3-1:0] node1239;
	wire [3-1:0] node1243;
	wire [3-1:0] node1244;
	wire [3-1:0] node1245;
	wire [3-1:0] node1249;
	wire [3-1:0] node1252;
	wire [3-1:0] node1253;
	wire [3-1:0] node1256;
	wire [3-1:0] node1258;
	wire [3-1:0] node1261;
	wire [3-1:0] node1262;
	wire [3-1:0] node1263;
	wire [3-1:0] node1264;
	wire [3-1:0] node1265;
	wire [3-1:0] node1266;
	wire [3-1:0] node1269;
	wire [3-1:0] node1271;
	wire [3-1:0] node1274;
	wire [3-1:0] node1275;
	wire [3-1:0] node1278;
	wire [3-1:0] node1280;
	wire [3-1:0] node1283;
	wire [3-1:0] node1284;
	wire [3-1:0] node1285;
	wire [3-1:0] node1288;
	wire [3-1:0] node1291;
	wire [3-1:0] node1293;
	wire [3-1:0] node1294;
	wire [3-1:0] node1298;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1301;
	wire [3-1:0] node1304;
	wire [3-1:0] node1305;
	wire [3-1:0] node1309;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1315;
	wire [3-1:0] node1316;
	wire [3-1:0] node1320;
	wire [3-1:0] node1321;
	wire [3-1:0] node1322;
	wire [3-1:0] node1326;
	wire [3-1:0] node1327;
	wire [3-1:0] node1328;
	wire [3-1:0] node1332;
	wire [3-1:0] node1335;
	wire [3-1:0] node1336;
	wire [3-1:0] node1337;
	wire [3-1:0] node1338;
	wire [3-1:0] node1339;
	wire [3-1:0] node1344;
	wire [3-1:0] node1345;
	wire [3-1:0] node1346;
	wire [3-1:0] node1349;
	wire [3-1:0] node1351;
	wire [3-1:0] node1354;
	wire [3-1:0] node1355;
	wire [3-1:0] node1360;
	wire [3-1:0] node1362;
	wire [3-1:0] node1364;
	wire [3-1:0] node1365;
	wire [3-1:0] node1366;
	wire [3-1:0] node1367;
	wire [3-1:0] node1369;
	wire [3-1:0] node1371;
	wire [3-1:0] node1374;
	wire [3-1:0] node1375;
	wire [3-1:0] node1378;
	wire [3-1:0] node1380;
	wire [3-1:0] node1384;
	wire [3-1:0] node1385;
	wire [3-1:0] node1386;
	wire [3-1:0] node1387;
	wire [3-1:0] node1389;
	wire [3-1:0] node1391;
	wire [3-1:0] node1394;
	wire [3-1:0] node1395;
	wire [3-1:0] node1396;
	wire [3-1:0] node1400;
	wire [3-1:0] node1402;
	wire [3-1:0] node1405;
	wire [3-1:0] node1407;
	wire [3-1:0] node1410;
	wire [3-1:0] node1412;
	wire [3-1:0] node1413;
	wire [3-1:0] node1415;
	wire [3-1:0] node1418;
	wire [3-1:0] node1419;

	assign outp = (inp[3]) ? node1116 : node1;
		assign node1 = (inp[4]) ? node759 : node2;
			assign node2 = (inp[0]) ? node526 : node3;
				assign node3 = (inp[6]) ? node315 : node4;
					assign node4 = (inp[9]) ? node146 : node5;
						assign node5 = (inp[1]) ? node73 : node6;
							assign node6 = (inp[5]) ? node50 : node7;
								assign node7 = (inp[7]) ? node27 : node8;
									assign node8 = (inp[2]) ? node16 : node9;
										assign node9 = (inp[8]) ? node11 : 3'b000;
											assign node11 = (inp[11]) ? 3'b000 : node12;
												assign node12 = (inp[10]) ? 3'b000 : 3'b100;
										assign node16 = (inp[10]) ? node22 : node17;
											assign node17 = (inp[11]) ? node19 : 3'b000;
												assign node19 = (inp[8]) ? 3'b100 : 3'b000;
											assign node22 = (inp[8]) ? node24 : 3'b100;
												assign node24 = (inp[11]) ? 3'b000 : 3'b100;
									assign node27 = (inp[11]) ? node39 : node28;
										assign node28 = (inp[10]) ? node34 : node29;
											assign node29 = (inp[2]) ? 3'b000 : node30;
												assign node30 = (inp[8]) ? 3'b100 : 3'b000;
											assign node34 = (inp[8]) ? node36 : 3'b100;
												assign node36 = (inp[2]) ? 3'b100 : 3'b010;
										assign node39 = (inp[2]) ? node45 : node40;
											assign node40 = (inp[10]) ? node42 : 3'b100;
												assign node42 = (inp[8]) ? 3'b010 : 3'b100;
											assign node45 = (inp[10]) ? node47 : 3'b010;
												assign node47 = (inp[8]) ? 3'b110 : 3'b010;
								assign node50 = (inp[11]) ? node62 : node51;
									assign node51 = (inp[7]) ? 3'b000 : node52;
										assign node52 = (inp[10]) ? node54 : 3'b000;
											assign node54 = (inp[8]) ? node58 : node55;
												assign node55 = (inp[2]) ? 3'b100 : 3'b000;
												assign node58 = (inp[2]) ? 3'b000 : 3'b100;
									assign node62 = (inp[2]) ? node68 : node63;
										assign node63 = (inp[10]) ? node65 : 3'b000;
											assign node65 = (inp[7]) ? 3'b000 : 3'b100;
										assign node68 = (inp[10]) ? node70 : 3'b100;
											assign node70 = (inp[7]) ? 3'b100 : 3'b000;
							assign node73 = (inp[5]) ? node115 : node74;
								assign node74 = (inp[2]) ? node98 : node75;
									assign node75 = (inp[10]) ? node87 : node76;
										assign node76 = (inp[7]) ? node82 : node77;
											assign node77 = (inp[8]) ? node79 : 3'b100;
												assign node79 = (inp[11]) ? 3'b000 : 3'b100;
											assign node82 = (inp[8]) ? node84 : 3'b010;
												assign node84 = (inp[11]) ? 3'b000 : 3'b010;
										assign node87 = (inp[7]) ? node93 : node88;
											assign node88 = (inp[11]) ? node90 : 3'b010;
												assign node90 = (inp[8]) ? 3'b110 : 3'b010;
											assign node93 = (inp[8]) ? node95 : 3'b110;
												assign node95 = (inp[11]) ? 3'b001 : 3'b011;
									assign node98 = (inp[7]) ? node110 : node99;
										assign node99 = (inp[8]) ? node103 : node100;
											assign node100 = (inp[10]) ? 3'b110 : 3'b010;
											assign node103 = (inp[11]) ? node107 : node104;
												assign node104 = (inp[10]) ? 3'b110 : 3'b010;
												assign node107 = (inp[10]) ? 3'b001 : 3'b101;
										assign node110 = (inp[10]) ? 3'b101 : node111;
											assign node111 = (inp[8]) ? 3'b111 : 3'b110;
								assign node115 = (inp[10]) ? node131 : node116;
									assign node116 = (inp[2]) ? node122 : node117;
										assign node117 = (inp[7]) ? node119 : 3'b000;
											assign node119 = (inp[11]) ? 3'b100 : 3'b000;
										assign node122 = (inp[11]) ? node128 : node123;
											assign node123 = (inp[8]) ? 3'b100 : node124;
												assign node124 = (inp[7]) ? 3'b100 : 3'b000;
											assign node128 = (inp[7]) ? 3'b010 : 3'b100;
									assign node131 = (inp[7]) ? node141 : node132;
										assign node132 = (inp[2]) ? node138 : node133;
											assign node133 = (inp[11]) ? 3'b100 : node134;
												assign node134 = (inp[8]) ? 3'b100 : 3'b000;
											assign node138 = (inp[11]) ? 3'b010 : 3'b000;
										assign node141 = (inp[2]) ? node143 : 3'b010;
											assign node143 = (inp[11]) ? 3'b110 : 3'b100;
						assign node146 = (inp[1]) ? node230 : node147;
							assign node147 = (inp[5]) ? node187 : node148;
								assign node148 = (inp[10]) ? node168 : node149;
									assign node149 = (inp[2]) ? node159 : node150;
										assign node150 = (inp[7]) ? 3'b010 : node151;
											assign node151 = (inp[11]) ? node155 : node152;
												assign node152 = (inp[8]) ? 3'b110 : 3'b010;
												assign node155 = (inp[8]) ? 3'b010 : 3'b110;
										assign node159 = (inp[7]) ? node163 : node160;
											assign node160 = (inp[8]) ? 3'b110 : 3'b010;
											assign node163 = (inp[11]) ? node165 : 3'b110;
												assign node165 = (inp[8]) ? 3'b111 : 3'b110;
									assign node168 = (inp[2]) ? node176 : node169;
										assign node169 = (inp[8]) ? node173 : node170;
											assign node170 = (inp[7]) ? 3'b110 : 3'b010;
											assign node173 = (inp[7]) ? 3'b001 : 3'b110;
										assign node176 = (inp[7]) ? node182 : node177;
											assign node177 = (inp[8]) ? node179 : 3'b110;
												assign node179 = (inp[11]) ? 3'b001 : 3'b110;
											assign node182 = (inp[11]) ? 3'b101 : node183;
												assign node183 = (inp[8]) ? 3'b101 : 3'b001;
								assign node187 = (inp[10]) ? node209 : node188;
									assign node188 = (inp[8]) ? node200 : node189;
										assign node189 = (inp[2]) ? node195 : node190;
											assign node190 = (inp[11]) ? 3'b100 : node191;
												assign node191 = (inp[7]) ? 3'b000 : 3'b010;
											assign node195 = (inp[11]) ? node197 : 3'b100;
												assign node197 = (inp[7]) ? 3'b010 : 3'b100;
										assign node200 = (inp[2]) ? node204 : node201;
											assign node201 = (inp[7]) ? 3'b100 : 3'b000;
											assign node204 = (inp[7]) ? node206 : 3'b100;
												assign node206 = (inp[11]) ? 3'b010 : 3'b000;
									assign node209 = (inp[11]) ? node223 : node210;
										assign node210 = (inp[2]) ? node216 : node211;
											assign node211 = (inp[7]) ? 3'b110 : node212;
												assign node212 = (inp[8]) ? 3'b100 : 3'b000;
											assign node216 = (inp[8]) ? node220 : node217;
												assign node217 = (inp[7]) ? 3'b000 : 3'b100;
												assign node220 = (inp[7]) ? 3'b100 : 3'b010;
										assign node223 = (inp[7]) ? node227 : node224;
											assign node224 = (inp[2]) ? 3'b010 : 3'b100;
											assign node227 = (inp[2]) ? 3'b110 : 3'b010;
							assign node230 = (inp[5]) ? node266 : node231;
								assign node231 = (inp[10]) ? node243 : node232;
									assign node232 = (inp[2]) ? node238 : node233;
										assign node233 = (inp[7]) ? node235 : 3'b110;
											assign node235 = (inp[8]) ? 3'b101 : 3'b001;
										assign node238 = (inp[7]) ? 3'b011 : node239;
											assign node239 = (inp[8]) ? 3'b101 : 3'b001;
									assign node243 = (inp[2]) ? node255 : node244;
										assign node244 = (inp[7]) ? node250 : node245;
											assign node245 = (inp[11]) ? 3'b101 : node246;
												assign node246 = (inp[8]) ? 3'b101 : 3'b001;
											assign node250 = (inp[11]) ? 3'b011 : node251;
												assign node251 = (inp[8]) ? 3'b011 : 3'b101;
										assign node255 = (inp[7]) ? node261 : node256;
											assign node256 = (inp[11]) ? 3'b011 : node257;
												assign node257 = (inp[8]) ? 3'b011 : 3'b101;
											assign node261 = (inp[11]) ? 3'b111 : node262;
												assign node262 = (inp[8]) ? 3'b111 : 3'b011;
								assign node266 = (inp[10]) ? node290 : node267;
									assign node267 = (inp[11]) ? node281 : node268;
										assign node268 = (inp[8]) ? node276 : node269;
											assign node269 = (inp[7]) ? node273 : node270;
												assign node270 = (inp[2]) ? 3'b010 : 3'b100;
												assign node273 = (inp[2]) ? 3'b100 : 3'b010;
											assign node276 = (inp[2]) ? node278 : 3'b110;
												assign node278 = (inp[7]) ? 3'b100 : 3'b110;
										assign node281 = (inp[7]) ? node285 : node282;
											assign node282 = (inp[2]) ? 3'b110 : 3'b010;
											assign node285 = (inp[2]) ? node287 : 3'b110;
												assign node287 = (inp[8]) ? 3'b011 : 3'b001;
									assign node290 = (inp[7]) ? node304 : node291;
										assign node291 = (inp[2]) ? node297 : node292;
											assign node292 = (inp[11]) ? 3'b110 : node293;
												assign node293 = (inp[8]) ? 3'b110 : 3'b010;
											assign node297 = (inp[8]) ? node301 : node298;
												assign node298 = (inp[11]) ? 3'b001 : 3'b110;
												assign node301 = (inp[11]) ? 3'b101 : 3'b001;
										assign node304 = (inp[11]) ? node308 : node305;
											assign node305 = (inp[2]) ? 3'b101 : 3'b100;
											assign node308 = (inp[2]) ? node312 : node309;
												assign node309 = (inp[8]) ? 3'b101 : 3'b001;
												assign node312 = (inp[8]) ? 3'b011 : 3'b101;
					assign node315 = (inp[9]) ? node389 : node316;
						assign node316 = (inp[1]) ? node378 : node317;
							assign node317 = (inp[5]) ? node333 : node318;
								assign node318 = (inp[2]) ? 3'b011 : node319;
									assign node319 = (inp[10]) ? 3'b011 : node320;
										assign node320 = (inp[7]) ? node326 : node321;
											assign node321 = (inp[8]) ? 3'b010 : node322;
												assign node322 = (inp[11]) ? 3'b010 : 3'b011;
											assign node326 = (inp[8]) ? 3'b011 : node327;
												assign node327 = (inp[11]) ? 3'b011 : 3'b010;
								assign node333 = (inp[7]) ? node351 : node334;
									assign node334 = (inp[10]) ? node340 : node335;
										assign node335 = (inp[2]) ? 3'b011 : node336;
											assign node336 = (inp[8]) ? 3'b010 : 3'b011;
										assign node340 = (inp[2]) ? node346 : node341;
											assign node341 = (inp[8]) ? node343 : 3'b011;
												assign node343 = (inp[11]) ? 3'b010 : 3'b011;
											assign node346 = (inp[8]) ? node348 : 3'b010;
												assign node348 = (inp[11]) ? 3'b011 : 3'b010;
									assign node351 = (inp[11]) ? node365 : node352;
										assign node352 = (inp[10]) ? node358 : node353;
											assign node353 = (inp[2]) ? 3'b010 : node354;
												assign node354 = (inp[8]) ? 3'b010 : 3'b011;
											assign node358 = (inp[8]) ? node362 : node359;
												assign node359 = (inp[2]) ? 3'b011 : 3'b010;
												assign node362 = (inp[2]) ? 3'b010 : 3'b011;
										assign node365 = (inp[2]) ? node373 : node366;
											assign node366 = (inp[8]) ? node370 : node367;
												assign node367 = (inp[10]) ? 3'b010 : 3'b011;
												assign node370 = (inp[10]) ? 3'b011 : 3'b010;
											assign node373 = (inp[8]) ? 3'b011 : node374;
												assign node374 = (inp[10]) ? 3'b011 : 3'b010;
							assign node378 = (inp[2]) ? 3'b011 : node379;
								assign node379 = (inp[7]) ? 3'b011 : node380;
									assign node380 = (inp[10]) ? 3'b011 : node381;
										assign node381 = (inp[5]) ? node383 : 3'b011;
											assign node383 = (inp[8]) ? 3'b011 : 3'b010;
						assign node389 = (inp[7]) ? node473 : node390;
							assign node390 = (inp[5]) ? node426 : node391;
								assign node391 = (inp[11]) ? node409 : node392;
									assign node392 = (inp[8]) ? node402 : node393;
										assign node393 = (inp[2]) ? node399 : node394;
											assign node394 = (inp[10]) ? 3'b011 : node395;
												assign node395 = (inp[1]) ? 3'b101 : 3'b001;
											assign node399 = (inp[10]) ? 3'b111 : 3'b011;
										assign node402 = (inp[2]) ? 3'b111 : node403;
											assign node403 = (inp[10]) ? node405 : 3'b011;
												assign node405 = (inp[1]) ? 3'b111 : 3'b011;
									assign node409 = (inp[8]) ? node417 : node410;
										assign node410 = (inp[2]) ? node412 : 3'b111;
											assign node412 = (inp[10]) ? node414 : 3'b111;
												assign node414 = (inp[1]) ? 3'b111 : 3'b011;
										assign node417 = (inp[10]) ? node421 : node418;
											assign node418 = (inp[2]) ? 3'b111 : 3'b011;
											assign node421 = (inp[2]) ? node423 : 3'b111;
												assign node423 = (inp[1]) ? 3'b111 : 3'b011;
								assign node426 = (inp[10]) ? node450 : node427;
									assign node427 = (inp[2]) ? node439 : node428;
										assign node428 = (inp[8]) ? node432 : node429;
											assign node429 = (inp[11]) ? 3'b011 : 3'b111;
											assign node432 = (inp[11]) ? node436 : node433;
												assign node433 = (inp[1]) ? 3'b001 : 3'b101;
												assign node436 = (inp[1]) ? 3'b101 : 3'b001;
										assign node439 = (inp[8]) ? node445 : node440;
											assign node440 = (inp[1]) ? 3'b101 : node441;
												assign node441 = (inp[11]) ? 3'b101 : 3'b001;
											assign node445 = (inp[11]) ? node447 : 3'b101;
												assign node447 = (inp[1]) ? 3'b011 : 3'b111;
									assign node450 = (inp[11]) ? node464 : node451;
										assign node451 = (inp[2]) ? node459 : node452;
											assign node452 = (inp[8]) ? node456 : node453;
												assign node453 = (inp[1]) ? 3'b101 : 3'b001;
												assign node456 = (inp[1]) ? 3'b111 : 3'b011;
											assign node459 = (inp[8]) ? 3'b001 : node460;
												assign node460 = (inp[1]) ? 3'b011 : 3'b111;
										assign node464 = (inp[8]) ? node468 : node465;
											assign node465 = (inp[2]) ? 3'b011 : 3'b101;
											assign node468 = (inp[2]) ? 3'b111 : node469;
												assign node469 = (inp[1]) ? 3'b011 : 3'b111;
							assign node473 = (inp[5]) ? node493 : node474;
								assign node474 = (inp[1]) ? node484 : node475;
									assign node475 = (inp[2]) ? node481 : node476;
										assign node476 = (inp[11]) ? node478 : 3'b011;
											assign node478 = (inp[10]) ? 3'b011 : 3'b111;
										assign node481 = (inp[11]) ? 3'b011 : 3'b111;
									assign node484 = (inp[8]) ? 3'b111 : node485;
										assign node485 = (inp[10]) ? 3'b111 : node486;
											assign node486 = (inp[2]) ? 3'b111 : node487;
												assign node487 = (inp[11]) ? 3'b111 : 3'b011;
								assign node493 = (inp[2]) ? node509 : node494;
									assign node494 = (inp[11]) ? node502 : node495;
										assign node495 = (inp[1]) ? node497 : 3'b011;
											assign node497 = (inp[8]) ? node499 : 3'b011;
												assign node499 = (inp[10]) ? 3'b111 : 3'b011;
										assign node502 = (inp[10]) ? node504 : 3'b111;
											assign node504 = (inp[1]) ? node506 : 3'b011;
												assign node506 = (inp[8]) ? 3'b111 : 3'b011;
									assign node509 = (inp[10]) ? node519 : node510;
										assign node510 = (inp[11]) ? node514 : node511;
											assign node511 = (inp[1]) ? 3'b011 : 3'b111;
											assign node514 = (inp[8]) ? node516 : 3'b011;
												assign node516 = (inp[1]) ? 3'b111 : 3'b011;
										assign node519 = (inp[8]) ? node521 : 3'b111;
											assign node521 = (inp[11]) ? 3'b111 : node522;
												assign node522 = (inp[1]) ? 3'b011 : 3'b111;
				assign node526 = (inp[6]) ? 3'b111 : node527;
					assign node527 = (inp[1]) ? node677 : node528;
						assign node528 = (inp[9]) ? node610 : node529;
							assign node529 = (inp[7]) ? node569 : node530;
								assign node530 = (inp[5]) ? node548 : node531;
									assign node531 = (inp[11]) ? node539 : node532;
										assign node532 = (inp[10]) ? node536 : node533;
											assign node533 = (inp[2]) ? 3'b011 : 3'b010;
											assign node536 = (inp[2]) ? 3'b101 : 3'b001;
										assign node539 = (inp[10]) ? node545 : node540;
											assign node540 = (inp[2]) ? 3'b101 : node541;
												assign node541 = (inp[8]) ? 3'b111 : 3'b110;
											assign node545 = (inp[2]) ? 3'b011 : 3'b101;
									assign node548 = (inp[2]) ? node556 : node549;
										assign node549 = (inp[11]) ? node553 : node550;
											assign node550 = (inp[10]) ? 3'b010 : 3'b110;
											assign node553 = (inp[10]) ? 3'b110 : 3'b010;
										assign node556 = (inp[10]) ? node562 : node557;
											assign node557 = (inp[8]) ? 3'b110 : node558;
												assign node558 = (inp[11]) ? 3'b110 : 3'b010;
											assign node562 = (inp[11]) ? node566 : node563;
												assign node563 = (inp[8]) ? 3'b010 : 3'b110;
												assign node566 = (inp[8]) ? 3'b101 : 3'b001;
								assign node569 = (inp[2]) ? node589 : node570;
									assign node570 = (inp[10]) ? node578 : node571;
										assign node571 = (inp[5]) ? node575 : node572;
											assign node572 = (inp[11]) ? 3'b101 : 3'b001;
											assign node575 = (inp[11]) ? 3'b111 : 3'b011;
										assign node578 = (inp[5]) ? node584 : node579;
											assign node579 = (inp[11]) ? 3'b011 : node580;
												assign node580 = (inp[8]) ? 3'b011 : 3'b001;
											assign node584 = (inp[11]) ? 3'b001 : node585;
												assign node585 = (inp[8]) ? 3'b001 : 3'b011;
									assign node589 = (inp[11]) ? node599 : node590;
										assign node590 = (inp[5]) ? node594 : node591;
											assign node591 = (inp[10]) ? 3'b111 : 3'b101;
											assign node594 = (inp[8]) ? 3'b101 : node595;
												assign node595 = (inp[10]) ? 3'b101 : 3'b111;
										assign node599 = (inp[10]) ? node605 : node600;
											assign node600 = (inp[8]) ? 3'b011 : node601;
												assign node601 = (inp[5]) ? 3'b001 : 3'b011;
											assign node605 = (inp[5]) ? node607 : 3'b111;
												assign node607 = (inp[8]) ? 3'b111 : 3'b101;
							assign node610 = (inp[5]) ? node638 : node611;
								assign node611 = (inp[2]) ? node631 : node612;
									assign node612 = (inp[10]) ? node624 : node613;
										assign node613 = (inp[7]) ? node619 : node614;
											assign node614 = (inp[11]) ? 3'b011 : node615;
												assign node615 = (inp[8]) ? 3'b011 : 3'b101;
											assign node619 = (inp[11]) ? 3'b111 : node620;
												assign node620 = (inp[8]) ? 3'b111 : 3'b011;
										assign node624 = (inp[8]) ? 3'b111 : node625;
											assign node625 = (inp[11]) ? 3'b111 : node626;
												assign node626 = (inp[7]) ? 3'b111 : 3'b011;
									assign node631 = (inp[11]) ? 3'b111 : node632;
										assign node632 = (inp[8]) ? 3'b111 : node633;
											assign node633 = (inp[7]) ? 3'b111 : 3'b011;
								assign node638 = (inp[2]) ? node660 : node639;
									assign node639 = (inp[8]) ? node647 : node640;
										assign node640 = (inp[10]) ? node644 : node641;
											assign node641 = (inp[7]) ? 3'b101 : 3'b110;
											assign node644 = (inp[7]) ? 3'b011 : 3'b101;
										assign node647 = (inp[10]) ? node653 : node648;
											assign node648 = (inp[11]) ? node650 : 3'b001;
												assign node650 = (inp[7]) ? 3'b011 : 3'b101;
											assign node653 = (inp[11]) ? node657 : node654;
												assign node654 = (inp[7]) ? 3'b111 : 3'b101;
												assign node657 = (inp[7]) ? 3'b111 : 3'b011;
									assign node660 = (inp[11]) ? node666 : node661;
										assign node661 = (inp[7]) ? 3'b011 : node662;
											assign node662 = (inp[10]) ? 3'b011 : 3'b101;
										assign node666 = (inp[7]) ? node672 : node667;
											assign node667 = (inp[10]) ? node669 : 3'b011;
												assign node669 = (inp[8]) ? 3'b111 : 3'b011;
											assign node672 = (inp[10]) ? 3'b111 : node673;
												assign node673 = (inp[8]) ? 3'b111 : 3'b011;
						assign node677 = (inp[9]) ? node745 : node678;
							assign node678 = (inp[5]) ? node700 : node679;
								assign node679 = (inp[2]) ? node695 : node680;
									assign node680 = (inp[10]) ? node690 : node681;
										assign node681 = (inp[7]) ? node687 : node682;
											assign node682 = (inp[11]) ? 3'b011 : node683;
												assign node683 = (inp[8]) ? 3'b011 : 3'b111;
											assign node687 = (inp[11]) ? 3'b111 : 3'b011;
										assign node690 = (inp[8]) ? 3'b111 : node691;
											assign node691 = (inp[11]) ? 3'b111 : 3'b011;
									assign node695 = (inp[11]) ? 3'b111 : node696;
										assign node696 = (inp[7]) ? 3'b111 : 3'b011;
								assign node700 = (inp[7]) ? node722 : node701;
									assign node701 = (inp[10]) ? node711 : node702;
										assign node702 = (inp[11]) ? node704 : 3'b101;
											assign node704 = (inp[8]) ? node708 : node705;
												assign node705 = (inp[2]) ? 3'b101 : 3'b001;
												assign node708 = (inp[2]) ? 3'b001 : 3'b111;
										assign node711 = (inp[2]) ? node717 : node712;
											assign node712 = (inp[11]) ? node714 : 3'b101;
												assign node714 = (inp[8]) ? 3'b011 : 3'b101;
											assign node717 = (inp[11]) ? node719 : 3'b011;
												assign node719 = (inp[8]) ? 3'b111 : 3'b011;
									assign node722 = (inp[11]) ? node736 : node723;
										assign node723 = (inp[2]) ? node731 : node724;
											assign node724 = (inp[8]) ? node728 : node725;
												assign node725 = (inp[10]) ? 3'b011 : 3'b111;
												assign node728 = (inp[10]) ? 3'b111 : 3'b011;
											assign node731 = (inp[10]) ? node733 : 3'b011;
												assign node733 = (inp[8]) ? 3'b011 : 3'b111;
										assign node736 = (inp[10]) ? 3'b111 : node737;
											assign node737 = (inp[8]) ? node741 : node738;
												assign node738 = (inp[2]) ? 3'b011 : 3'b111;
												assign node741 = (inp[2]) ? 3'b111 : 3'b011;
							assign node745 = (inp[7]) ? 3'b111 : node746;
								assign node746 = (inp[10]) ? 3'b111 : node747;
									assign node747 = (inp[5]) ? node749 : 3'b111;
										assign node749 = (inp[2]) ? 3'b111 : node750;
											assign node750 = (inp[11]) ? node752 : 3'b011;
												assign node752 = (inp[8]) ? 3'b111 : 3'b011;
			assign node759 = (inp[0]) ? node881 : node760;
				assign node760 = (inp[9]) ? node762 : 3'b000;
					assign node762 = (inp[6]) ? node848 : node763;
						assign node763 = (inp[7]) ? node803 : node764;
							assign node764 = (inp[1]) ? node774 : node765;
								assign node765 = (inp[2]) ? node767 : 3'b000;
									assign node767 = (inp[5]) ? 3'b000 : node768;
										assign node768 = (inp[10]) ? node770 : 3'b000;
											assign node770 = (inp[8]) ? 3'b100 : 3'b000;
								assign node774 = (inp[5]) ? node796 : node775;
									assign node775 = (inp[10]) ? node787 : node776;
										assign node776 = (inp[11]) ? node782 : node777;
											assign node777 = (inp[8]) ? 3'b100 : node778;
												assign node778 = (inp[2]) ? 3'b100 : 3'b000;
											assign node782 = (inp[2]) ? 3'b010 : node783;
												assign node783 = (inp[8]) ? 3'b100 : 3'b000;
										assign node787 = (inp[8]) ? node791 : node788;
											assign node788 = (inp[2]) ? 3'b010 : 3'b100;
											assign node791 = (inp[2]) ? node793 : 3'b010;
												assign node793 = (inp[11]) ? 3'b110 : 3'b010;
									assign node796 = (inp[10]) ? node798 : 3'b000;
										assign node798 = (inp[11]) ? node800 : 3'b000;
											assign node800 = (inp[2]) ? 3'b100 : 3'b000;
							assign node803 = (inp[5]) ? node839 : node804;
								assign node804 = (inp[10]) ? node822 : node805;
									assign node805 = (inp[2]) ? node809 : node806;
										assign node806 = (inp[8]) ? 3'b000 : 3'b100;
										assign node809 = (inp[1]) ? node815 : node810;
											assign node810 = (inp[11]) ? 3'b100 : node811;
												assign node811 = (inp[8]) ? 3'b100 : 3'b000;
											assign node815 = (inp[11]) ? node819 : node816;
												assign node816 = (inp[8]) ? 3'b110 : 3'b010;
												assign node819 = (inp[8]) ? 3'b101 : 3'b110;
									assign node822 = (inp[1]) ? node830 : node823;
										assign node823 = (inp[8]) ? node827 : node824;
											assign node824 = (inp[2]) ? 3'b100 : 3'b000;
											assign node827 = (inp[2]) ? 3'b010 : 3'b100;
										assign node830 = (inp[2]) ? node834 : node831;
											assign node831 = (inp[8]) ? 3'b110 : 3'b010;
											assign node834 = (inp[11]) ? node836 : 3'b010;
												assign node836 = (inp[8]) ? 3'b001 : 3'b110;
								assign node839 = (inp[11]) ? node841 : 3'b100;
									assign node841 = (inp[2]) ? node843 : 3'b100;
										assign node843 = (inp[1]) ? node845 : 3'b000;
											assign node845 = (inp[10]) ? 3'b010 : 3'b000;
						assign node848 = (inp[1]) ? node850 : 3'b000;
							assign node850 = (inp[7]) ? node872 : node851;
								assign node851 = (inp[5]) ? 3'b000 : node852;
									assign node852 = (inp[2]) ? node858 : node853;
										assign node853 = (inp[8]) ? node855 : 3'b000;
											assign node855 = (inp[10]) ? 3'b001 : 3'b000;
										assign node858 = (inp[11]) ? node864 : node859;
											assign node859 = (inp[10]) ? node861 : 3'b000;
												assign node861 = (inp[8]) ? 3'b000 : 3'b001;
											assign node864 = (inp[8]) ? node868 : node865;
												assign node865 = (inp[10]) ? 3'b001 : 3'b000;
												assign node868 = (inp[10]) ? 3'b000 : 3'b001;
								assign node872 = (inp[5]) ? node874 : 3'b001;
									assign node874 = (inp[2]) ? node876 : 3'b000;
										assign node876 = (inp[11]) ? 3'b001 : node877;
											assign node877 = (inp[8]) ? 3'b001 : 3'b000;
				assign node881 = (inp[9]) ? node977 : node882;
					assign node882 = (inp[6]) ? 3'b000 : node883;
						assign node883 = (inp[7]) ? node947 : node884;
							assign node884 = (inp[1]) ? node908 : node885;
								assign node885 = (inp[5]) ? node903 : node886;
									assign node886 = (inp[2]) ? node894 : node887;
										assign node887 = (inp[8]) ? node889 : 3'b100;
											assign node889 = (inp[10]) ? node891 : 3'b000;
												assign node891 = (inp[11]) ? 3'b010 : 3'b110;
										assign node894 = (inp[8]) ? node900 : node895;
											assign node895 = (inp[11]) ? node897 : 3'b010;
												assign node897 = (inp[10]) ? 3'b010 : 3'b110;
											assign node900 = (inp[11]) ? 3'b000 : 3'b010;
									assign node903 = (inp[2]) ? node905 : 3'b000;
										assign node905 = (inp[11]) ? 3'b100 : 3'b000;
								assign node908 = (inp[5]) ? node928 : node909;
									assign node909 = (inp[10]) ? node921 : node910;
										assign node910 = (inp[2]) ? node916 : node911;
											assign node911 = (inp[8]) ? node913 : 3'b010;
												assign node913 = (inp[11]) ? 3'b110 : 3'b010;
											assign node916 = (inp[11]) ? node918 : 3'b110;
												assign node918 = (inp[8]) ? 3'b111 : 3'b110;
										assign node921 = (inp[8]) ? node925 : node922;
											assign node922 = (inp[2]) ? 3'b101 : 3'b110;
											assign node925 = (inp[2]) ? 3'b101 : 3'b001;
									assign node928 = (inp[10]) ? node940 : node929;
										assign node929 = (inp[2]) ? node935 : node930;
											assign node930 = (inp[11]) ? 3'b100 : node931;
												assign node931 = (inp[8]) ? 3'b100 : 3'b000;
											assign node935 = (inp[11]) ? 3'b010 : node936;
												assign node936 = (inp[8]) ? 3'b010 : 3'b100;
										assign node940 = (inp[2]) ? node942 : 3'b010;
											assign node942 = (inp[8]) ? 3'b110 : node943;
												assign node943 = (inp[11]) ? 3'b110 : 3'b010;
							assign node947 = (inp[5]) ? node967 : node948;
								assign node948 = (inp[1]) ? node956 : node949;
									assign node949 = (inp[8]) ? node951 : 3'b110;
										assign node951 = (inp[10]) ? node953 : 3'b110;
											assign node953 = (inp[2]) ? 3'b111 : 3'b110;
									assign node956 = (inp[11]) ? node962 : node957;
										assign node957 = (inp[2]) ? 3'b111 : node958;
											assign node958 = (inp[10]) ? 3'b111 : 3'b110;
										assign node962 = (inp[8]) ? 3'b110 : node963;
											assign node963 = (inp[2]) ? 3'b111 : 3'b110;
								assign node967 = (inp[11]) ? node969 : 3'b110;
									assign node969 = (inp[10]) ? node971 : 3'b110;
										assign node971 = (inp[2]) ? node973 : 3'b110;
											assign node973 = (inp[1]) ? 3'b111 : 3'b110;
					assign node977 = (inp[6]) ? node1111 : node978;
						assign node978 = (inp[1]) ? node1036 : node979;
							assign node979 = (inp[5]) ? node1003 : node980;
								assign node980 = (inp[7]) ? node998 : node981;
									assign node981 = (inp[10]) ? node989 : node982;
										assign node982 = (inp[2]) ? node984 : 3'b010;
											assign node984 = (inp[11]) ? node986 : 3'b110;
												assign node986 = (inp[8]) ? 3'b111 : 3'b110;
										assign node989 = (inp[2]) ? node993 : node990;
											assign node990 = (inp[8]) ? 3'b001 : 3'b110;
											assign node993 = (inp[8]) ? 3'b101 : node994;
												assign node994 = (inp[11]) ? 3'b101 : 3'b001;
									assign node998 = (inp[2]) ? node1000 : 3'b101;
										assign node1000 = (inp[11]) ? 3'b011 : 3'b101;
								assign node1003 = (inp[2]) ? node1017 : node1004;
									assign node1004 = (inp[10]) ? node1012 : node1005;
										assign node1005 = (inp[11]) ? 3'b100 : node1006;
											assign node1006 = (inp[8]) ? 3'b100 : node1007;
												assign node1007 = (inp[7]) ? 3'b100 : 3'b000;
										assign node1012 = (inp[7]) ? 3'b110 : node1013;
											assign node1013 = (inp[11]) ? 3'b010 : 3'b100;
									assign node1017 = (inp[7]) ? node1025 : node1018;
										assign node1018 = (inp[10]) ? 3'b110 : node1019;
											assign node1019 = (inp[8]) ? 3'b010 : node1020;
												assign node1020 = (inp[11]) ? 3'b010 : 3'b100;
										assign node1025 = (inp[11]) ? node1033 : node1026;
											assign node1026 = (inp[8]) ? node1030 : node1027;
												assign node1027 = (inp[10]) ? 3'b110 : 3'b100;
												assign node1030 = (inp[10]) ? 3'b101 : 3'b111;
											assign node1033 = (inp[10]) ? 3'b001 : 3'b011;
							assign node1036 = (inp[5]) ? node1062 : node1037;
								assign node1037 = (inp[7]) ? 3'b111 : node1038;
									assign node1038 = (inp[10]) ? node1050 : node1039;
										assign node1039 = (inp[2]) ? node1045 : node1040;
											assign node1040 = (inp[11]) ? 3'b101 : node1041;
												assign node1041 = (inp[8]) ? 3'b101 : 3'b001;
											assign node1045 = (inp[11]) ? 3'b011 : node1046;
												assign node1046 = (inp[8]) ? 3'b001 : 3'b101;
										assign node1050 = (inp[2]) ? node1056 : node1051;
											assign node1051 = (inp[8]) ? 3'b011 : node1052;
												assign node1052 = (inp[11]) ? 3'b011 : 3'b101;
											assign node1056 = (inp[8]) ? 3'b111 : node1057;
												assign node1057 = (inp[11]) ? 3'b111 : 3'b011;
								assign node1062 = (inp[7]) ? node1088 : node1063;
									assign node1063 = (inp[10]) ? node1077 : node1064;
										assign node1064 = (inp[2]) ? node1070 : node1065;
											assign node1065 = (inp[11]) ? 3'b110 : node1066;
												assign node1066 = (inp[8]) ? 3'b110 : 3'b010;
											assign node1070 = (inp[11]) ? node1074 : node1071;
												assign node1071 = (inp[8]) ? 3'b100 : 3'b110;
												assign node1074 = (inp[8]) ? 3'b011 : 3'b001;
										assign node1077 = (inp[11]) ? node1083 : node1078;
											assign node1078 = (inp[2]) ? 3'b101 : node1079;
												assign node1079 = (inp[8]) ? 3'b001 : 3'b110;
											assign node1083 = (inp[2]) ? 3'b011 : node1084;
												assign node1084 = (inp[8]) ? 3'b101 : 3'b001;
									assign node1088 = (inp[10]) ? node1100 : node1089;
										assign node1089 = (inp[2]) ? node1095 : node1090;
											assign node1090 = (inp[8]) ? node1092 : 3'b001;
												assign node1092 = (inp[11]) ? 3'b011 : 3'b001;
											assign node1095 = (inp[8]) ? node1097 : 3'b001;
												assign node1097 = (inp[11]) ? 3'b101 : 3'b001;
										assign node1100 = (inp[2]) ? node1106 : node1101;
											assign node1101 = (inp[8]) ? node1103 : 3'b101;
												assign node1103 = (inp[11]) ? 3'b011 : 3'b001;
											assign node1106 = (inp[11]) ? node1108 : 3'b011;
												assign node1108 = (inp[8]) ? 3'b111 : 3'b011;
						assign node1111 = (inp[10]) ? 3'b111 : node1112;
							assign node1112 = (inp[7]) ? 3'b111 : 3'b011;
		assign node1116 = (inp[0]) ? node1130 : node1117;
			assign node1117 = (inp[6]) ? 3'b000 : node1118;
				assign node1118 = (inp[4]) ? 3'b000 : node1119;
					assign node1119 = (inp[7]) ? node1121 : 3'b000;
						assign node1121 = (inp[11]) ? node1123 : 3'b000;
							assign node1123 = (inp[8]) ? node1125 : 3'b000;
								assign node1125 = (inp[9]) ? 3'b100 : 3'b000;
			assign node1130 = (inp[4]) ? node1360 : node1131;
				assign node1131 = (inp[9]) ? node1151 : node1132;
					assign node1132 = (inp[6]) ? 3'b000 : node1133;
						assign node1133 = (inp[7]) ? 3'b100 : node1134;
							assign node1134 = (inp[1]) ? node1136 : 3'b000;
								assign node1136 = (inp[5]) ? 3'b000 : node1137;
									assign node1137 = (inp[2]) ? node1143 : node1138;
										assign node1138 = (inp[10]) ? node1140 : 3'b000;
											assign node1140 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1143 = (inp[8]) ? node1145 : 3'b100;
											assign node1145 = (inp[11]) ? 3'b000 : 3'b100;
					assign node1151 = (inp[6]) ? node1261 : node1152;
						assign node1152 = (inp[1]) ? node1192 : node1153;
							assign node1153 = (inp[5]) ? node1185 : node1154;
								assign node1154 = (inp[8]) ? node1168 : node1155;
									assign node1155 = (inp[10]) ? node1163 : node1156;
										assign node1156 = (inp[2]) ? node1158 : 3'b000;
											assign node1158 = (inp[7]) ? node1160 : 3'b000;
												assign node1160 = (inp[11]) ? 3'b010 : 3'b100;
										assign node1163 = (inp[7]) ? 3'b100 : node1164;
											assign node1164 = (inp[2]) ? 3'b100 : 3'b000;
									assign node1168 = (inp[10]) ? node1178 : node1169;
										assign node1169 = (inp[2]) ? node1173 : node1170;
											assign node1170 = (inp[7]) ? 3'b100 : 3'b000;
											assign node1173 = (inp[7]) ? node1175 : 3'b100;
												assign node1175 = (inp[11]) ? 3'b010 : 3'b000;
										assign node1178 = (inp[7]) ? node1180 : 3'b010;
											assign node1180 = (inp[2]) ? node1182 : 3'b010;
												assign node1182 = (inp[11]) ? 3'b110 : 3'b100;
								assign node1185 = (inp[7]) ? node1187 : 3'b000;
									assign node1187 = (inp[2]) ? node1189 : 3'b000;
										assign node1189 = (inp[11]) ? 3'b100 : 3'b000;
							assign node1192 = (inp[5]) ? node1234 : node1193;
								assign node1193 = (inp[8]) ? node1209 : node1194;
									assign node1194 = (inp[10]) ? node1202 : node1195;
										assign node1195 = (inp[2]) ? node1199 : node1196;
											assign node1196 = (inp[7]) ? 3'b010 : 3'b100;
											assign node1199 = (inp[7]) ? 3'b110 : 3'b010;
										assign node1202 = (inp[7]) ? node1206 : node1203;
											assign node1203 = (inp[2]) ? 3'b110 : 3'b010;
											assign node1206 = (inp[2]) ? 3'b101 : 3'b110;
									assign node1209 = (inp[11]) ? node1223 : node1210;
										assign node1210 = (inp[7]) ? node1216 : node1211;
											assign node1211 = (inp[10]) ? 3'b010 : node1212;
												assign node1212 = (inp[2]) ? 3'b010 : 3'b000;
											assign node1216 = (inp[10]) ? node1220 : node1217;
												assign node1217 = (inp[2]) ? 3'b110 : 3'b010;
												assign node1220 = (inp[2]) ? 3'b101 : 3'b011;
										assign node1223 = (inp[2]) ? node1229 : node1224;
											assign node1224 = (inp[7]) ? node1226 : 3'b100;
												assign node1226 = (inp[10]) ? 3'b001 : 3'b000;
											assign node1229 = (inp[7]) ? node1231 : 3'b001;
												assign node1231 = (inp[10]) ? 3'b101 : 3'b111;
								assign node1234 = (inp[7]) ? node1252 : node1235;
									assign node1235 = (inp[10]) ? node1243 : node1236;
										assign node1236 = (inp[2]) ? node1238 : 3'b000;
											assign node1238 = (inp[11]) ? 3'b100 : node1239;
												assign node1239 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1243 = (inp[2]) ? node1249 : node1244;
											assign node1244 = (inp[8]) ? 3'b100 : node1245;
												assign node1245 = (inp[11]) ? 3'b100 : 3'b000;
											assign node1249 = (inp[11]) ? 3'b010 : 3'b100;
									assign node1252 = (inp[2]) ? node1256 : node1253;
										assign node1253 = (inp[10]) ? 3'b010 : 3'b000;
										assign node1256 = (inp[11]) ? node1258 : 3'b100;
											assign node1258 = (inp[10]) ? 3'b110 : 3'b010;
						assign node1261 = (inp[7]) ? node1335 : node1262;
							assign node1262 = (inp[1]) ? node1298 : node1263;
								assign node1263 = (inp[10]) ? node1283 : node1264;
									assign node1264 = (inp[2]) ? node1274 : node1265;
										assign node1265 = (inp[11]) ? node1269 : node1266;
											assign node1266 = (inp[8]) ? 3'b010 : 3'b011;
											assign node1269 = (inp[8]) ? node1271 : 3'b010;
												assign node1271 = (inp[5]) ? 3'b011 : 3'b010;
										assign node1274 = (inp[8]) ? node1278 : node1275;
											assign node1275 = (inp[11]) ? 3'b011 : 3'b010;
											assign node1278 = (inp[11]) ? node1280 : 3'b011;
												assign node1280 = (inp[5]) ? 3'b010 : 3'b011;
									assign node1283 = (inp[11]) ? node1291 : node1284;
										assign node1284 = (inp[2]) ? node1288 : node1285;
											assign node1285 = (inp[5]) ? 3'b011 : 3'b010;
											assign node1288 = (inp[5]) ? 3'b010 : 3'b011;
										assign node1291 = (inp[5]) ? node1293 : 3'b011;
											assign node1293 = (inp[8]) ? 3'b011 : node1294;
												assign node1294 = (inp[2]) ? 3'b010 : 3'b011;
								assign node1298 = (inp[8]) ? node1320 : node1299;
									assign node1299 = (inp[11]) ? node1309 : node1300;
										assign node1300 = (inp[5]) ? node1304 : node1301;
											assign node1301 = (inp[2]) ? 3'b011 : 3'b001;
											assign node1304 = (inp[10]) ? 3'b011 : node1305;
												assign node1305 = (inp[2]) ? 3'b011 : 3'b010;
										assign node1309 = (inp[10]) ? node1315 : node1310;
											assign node1310 = (inp[2]) ? 3'b001 : node1311;
												assign node1311 = (inp[5]) ? 3'b010 : 3'b001;
											assign node1315 = (inp[5]) ? 3'b001 : node1316;
												assign node1316 = (inp[2]) ? 3'b011 : 3'b001;
									assign node1320 = (inp[5]) ? node1326 : node1321;
										assign node1321 = (inp[2]) ? 3'b011 : node1322;
											assign node1322 = (inp[11]) ? 3'b011 : 3'b001;
										assign node1326 = (inp[2]) ? node1332 : node1327;
											assign node1327 = (inp[11]) ? 3'b011 : node1328;
												assign node1328 = (inp[10]) ? 3'b011 : 3'b010;
											assign node1332 = (inp[10]) ? 3'b011 : 3'b001;
							assign node1335 = (inp[1]) ? 3'b101 : node1336;
								assign node1336 = (inp[5]) ? node1344 : node1337;
									assign node1337 = (inp[10]) ? 3'b101 : node1338;
										assign node1338 = (inp[11]) ? 3'b101 : node1339;
											assign node1339 = (inp[2]) ? 3'b101 : 3'b100;
									assign node1344 = (inp[10]) ? node1354 : node1345;
										assign node1345 = (inp[8]) ? node1349 : node1346;
											assign node1346 = (inp[2]) ? 3'b100 : 3'b101;
											assign node1349 = (inp[2]) ? node1351 : 3'b100;
												assign node1351 = (inp[11]) ? 3'b101 : 3'b100;
										assign node1354 = (inp[2]) ? 3'b101 : node1355;
											assign node1355 = (inp[8]) ? 3'b101 : 3'b100;
				assign node1360 = (inp[1]) ? node1362 : 3'b000;
					assign node1362 = (inp[9]) ? node1364 : 3'b000;
						assign node1364 = (inp[6]) ? node1384 : node1365;
							assign node1365 = (inp[5]) ? 3'b000 : node1366;
								assign node1366 = (inp[7]) ? node1374 : node1367;
									assign node1367 = (inp[2]) ? node1369 : 3'b000;
										assign node1369 = (inp[11]) ? node1371 : 3'b000;
											assign node1371 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1374 = (inp[2]) ? node1378 : node1375;
										assign node1375 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1378 = (inp[11]) ? node1380 : 3'b100;
											assign node1380 = (inp[8]) ? 3'b010 : 3'b100;
							assign node1384 = (inp[7]) ? node1410 : node1385;
								assign node1385 = (inp[5]) ? node1405 : node1386;
									assign node1386 = (inp[2]) ? node1394 : node1387;
										assign node1387 = (inp[11]) ? node1389 : 3'b100;
											assign node1389 = (inp[8]) ? node1391 : 3'b100;
												assign node1391 = (inp[10]) ? 3'b010 : 3'b000;
										assign node1394 = (inp[8]) ? node1400 : node1395;
											assign node1395 = (inp[11]) ? 3'b100 : node1396;
												assign node1396 = (inp[10]) ? 3'b010 : 3'b000;
											assign node1400 = (inp[11]) ? node1402 : 3'b000;
												assign node1402 = (inp[10]) ? 3'b000 : 3'b010;
									assign node1405 = (inp[2]) ? node1407 : 3'b000;
										assign node1407 = (inp[11]) ? 3'b100 : 3'b000;
								assign node1410 = (inp[5]) ? node1412 : 3'b110;
									assign node1412 = (inp[2]) ? node1418 : node1413;
										assign node1413 = (inp[11]) ? node1415 : 3'b000;
											assign node1415 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1418 = (inp[11]) ? 3'b010 : node1419;
											assign node1419 = (inp[8]) ? 3'b010 : 3'b100;

endmodule