module dtc_split75_bm39 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node5;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node10;
	wire [14-1:0] node11;
	wire [14-1:0] node12;
	wire [14-1:0] node13;
	wire [14-1:0] node18;
	wire [14-1:0] node19;
	wire [14-1:0] node20;
	wire [14-1:0] node24;
	wire [14-1:0] node25;
	wire [14-1:0] node28;
	wire [14-1:0] node31;
	wire [14-1:0] node32;
	wire [14-1:0] node33;
	wire [14-1:0] node34;
	wire [14-1:0] node37;
	wire [14-1:0] node40;
	wire [14-1:0] node41;
	wire [14-1:0] node44;
	wire [14-1:0] node47;
	wire [14-1:0] node48;
	wire [14-1:0] node50;
	wire [14-1:0] node53;
	wire [14-1:0] node54;
	wire [14-1:0] node57;
	wire [14-1:0] node60;
	wire [14-1:0] node61;
	wire [14-1:0] node62;
	wire [14-1:0] node64;
	wire [14-1:0] node65;
	wire [14-1:0] node68;
	wire [14-1:0] node71;
	wire [14-1:0] node72;
	wire [14-1:0] node73;
	wire [14-1:0] node76;
	wire [14-1:0] node79;
	wire [14-1:0] node80;
	wire [14-1:0] node83;
	wire [14-1:0] node86;
	wire [14-1:0] node87;
	wire [14-1:0] node88;
	wire [14-1:0] node89;
	wire [14-1:0] node92;
	wire [14-1:0] node95;
	wire [14-1:0] node96;
	wire [14-1:0] node99;
	wire [14-1:0] node102;
	wire [14-1:0] node103;
	wire [14-1:0] node104;
	wire [14-1:0] node107;
	wire [14-1:0] node110;
	wire [14-1:0] node111;
	wire [14-1:0] node114;
	wire [14-1:0] node117;
	wire [14-1:0] node118;
	wire [14-1:0] node119;
	wire [14-1:0] node120;
	wire [14-1:0] node121;
	wire [14-1:0] node122;
	wire [14-1:0] node125;
	wire [14-1:0] node128;
	wire [14-1:0] node129;
	wire [14-1:0] node132;
	wire [14-1:0] node135;
	wire [14-1:0] node136;
	wire [14-1:0] node137;
	wire [14-1:0] node140;
	wire [14-1:0] node143;
	wire [14-1:0] node144;
	wire [14-1:0] node147;
	wire [14-1:0] node150;
	wire [14-1:0] node151;
	wire [14-1:0] node152;
	wire [14-1:0] node155;
	wire [14-1:0] node158;
	wire [14-1:0] node159;
	wire [14-1:0] node160;
	wire [14-1:0] node163;
	wire [14-1:0] node166;
	wire [14-1:0] node167;
	wire [14-1:0] node170;
	wire [14-1:0] node173;
	wire [14-1:0] node174;
	wire [14-1:0] node175;
	wire [14-1:0] node177;
	wire [14-1:0] node178;
	wire [14-1:0] node181;
	wire [14-1:0] node184;
	wire [14-1:0] node185;
	wire [14-1:0] node186;
	wire [14-1:0] node189;
	wire [14-1:0] node192;
	wire [14-1:0] node194;
	wire [14-1:0] node195;
	wire [14-1:0] node199;
	wire [14-1:0] node200;
	wire [14-1:0] node201;
	wire [14-1:0] node202;
	wire [14-1:0] node205;
	wire [14-1:0] node209;
	wire [14-1:0] node211;
	wire [14-1:0] node212;
	wire [14-1:0] node215;
	wire [14-1:0] node218;
	wire [14-1:0] node219;
	wire [14-1:0] node220;
	wire [14-1:0] node221;
	wire [14-1:0] node222;
	wire [14-1:0] node224;
	wire [14-1:0] node225;
	wire [14-1:0] node228;
	wire [14-1:0] node231;
	wire [14-1:0] node232;
	wire [14-1:0] node233;
	wire [14-1:0] node236;
	wire [14-1:0] node239;
	wire [14-1:0] node240;
	wire [14-1:0] node243;
	wire [14-1:0] node246;
	wire [14-1:0] node247;
	wire [14-1:0] node248;
	wire [14-1:0] node249;
	wire [14-1:0] node252;
	wire [14-1:0] node255;
	wire [14-1:0] node256;
	wire [14-1:0] node259;
	wire [14-1:0] node262;
	wire [14-1:0] node263;
	wire [14-1:0] node264;
	wire [14-1:0] node267;
	wire [14-1:0] node270;
	wire [14-1:0] node271;
	wire [14-1:0] node274;
	wire [14-1:0] node277;
	wire [14-1:0] node278;
	wire [14-1:0] node279;
	wire [14-1:0] node280;
	wire [14-1:0] node282;
	wire [14-1:0] node285;
	wire [14-1:0] node287;
	wire [14-1:0] node290;
	wire [14-1:0] node291;
	wire [14-1:0] node292;
	wire [14-1:0] node295;
	wire [14-1:0] node298;
	wire [14-1:0] node299;
	wire [14-1:0] node303;
	wire [14-1:0] node305;
	wire [14-1:0] node306;
	wire [14-1:0] node307;
	wire [14-1:0] node311;
	wire [14-1:0] node312;
	wire [14-1:0] node315;
	wire [14-1:0] node318;
	wire [14-1:0] node319;
	wire [14-1:0] node320;
	wire [14-1:0] node322;
	wire [14-1:0] node323;
	wire [14-1:0] node325;
	wire [14-1:0] node328;
	wire [14-1:0] node329;
	wire [14-1:0] node332;
	wire [14-1:0] node335;
	wire [14-1:0] node336;
	wire [14-1:0] node337;
	wire [14-1:0] node338;
	wire [14-1:0] node342;
	wire [14-1:0] node343;
	wire [14-1:0] node346;
	wire [14-1:0] node351;
	wire [14-1:0] node352;
	wire [14-1:0] node353;
	wire [14-1:0] node354;
	wire [14-1:0] node355;
	wire [14-1:0] node356;
	wire [14-1:0] node357;
	wire [14-1:0] node360;
	wire [14-1:0] node361;
	wire [14-1:0] node364;
	wire [14-1:0] node367;
	wire [14-1:0] node368;
	wire [14-1:0] node369;
	wire [14-1:0] node372;
	wire [14-1:0] node375;
	wire [14-1:0] node376;
	wire [14-1:0] node380;
	wire [14-1:0] node381;
	wire [14-1:0] node382;
	wire [14-1:0] node383;
	wire [14-1:0] node386;
	wire [14-1:0] node389;
	wire [14-1:0] node391;
	wire [14-1:0] node394;
	wire [14-1:0] node395;
	wire [14-1:0] node396;
	wire [14-1:0] node399;
	wire [14-1:0] node402;
	wire [14-1:0] node404;
	wire [14-1:0] node407;
	wire [14-1:0] node408;
	wire [14-1:0] node409;
	wire [14-1:0] node410;
	wire [14-1:0] node411;
	wire [14-1:0] node414;
	wire [14-1:0] node417;
	wire [14-1:0] node418;
	wire [14-1:0] node421;
	wire [14-1:0] node424;
	wire [14-1:0] node425;
	wire [14-1:0] node426;
	wire [14-1:0] node429;
	wire [14-1:0] node432;
	wire [14-1:0] node433;
	wire [14-1:0] node436;
	wire [14-1:0] node439;
	wire [14-1:0] node440;
	wire [14-1:0] node441;
	wire [14-1:0] node442;
	wire [14-1:0] node445;
	wire [14-1:0] node448;
	wire [14-1:0] node449;
	wire [14-1:0] node452;
	wire [14-1:0] node455;
	wire [14-1:0] node456;
	wire [14-1:0] node457;
	wire [14-1:0] node461;
	wire [14-1:0] node464;
	wire [14-1:0] node465;
	wire [14-1:0] node466;
	wire [14-1:0] node467;
	wire [14-1:0] node468;
	wire [14-1:0] node469;
	wire [14-1:0] node473;
	wire [14-1:0] node474;
	wire [14-1:0] node477;
	wire [14-1:0] node480;
	wire [14-1:0] node481;
	wire [14-1:0] node482;
	wire [14-1:0] node485;
	wire [14-1:0] node488;
	wire [14-1:0] node489;
	wire [14-1:0] node492;
	wire [14-1:0] node495;
	wire [14-1:0] node496;
	wire [14-1:0] node497;
	wire [14-1:0] node498;
	wire [14-1:0] node501;
	wire [14-1:0] node504;
	wire [14-1:0] node505;
	wire [14-1:0] node509;
	wire [14-1:0] node511;
	wire [14-1:0] node512;
	wire [14-1:0] node515;
	wire [14-1:0] node518;
	wire [14-1:0] node519;
	wire [14-1:0] node520;
	wire [14-1:0] node522;
	wire [14-1:0] node523;
	wire [14-1:0] node526;
	wire [14-1:0] node529;
	wire [14-1:0] node530;
	wire [14-1:0] node531;
	wire [14-1:0] node534;
	wire [14-1:0] node539;
	wire [14-1:0] node540;
	wire [14-1:0] node542;
	wire [14-1:0] node543;
	wire [14-1:0] node545;
	wire [14-1:0] node546;
	wire [14-1:0] node547;
	wire [14-1:0] node554;
	wire [14-1:0] node555;
	wire [14-1:0] node556;
	wire [14-1:0] node557;
	wire [14-1:0] node558;
	wire [14-1:0] node559;
	wire [14-1:0] node560;
	wire [14-1:0] node561;
	wire [14-1:0] node563;
	wire [14-1:0] node566;
	wire [14-1:0] node567;
	wire [14-1:0] node570;
	wire [14-1:0] node573;
	wire [14-1:0] node574;
	wire [14-1:0] node575;
	wire [14-1:0] node578;
	wire [14-1:0] node581;
	wire [14-1:0] node582;
	wire [14-1:0] node586;
	wire [14-1:0] node587;
	wire [14-1:0] node588;
	wire [14-1:0] node590;
	wire [14-1:0] node593;
	wire [14-1:0] node594;
	wire [14-1:0] node598;
	wire [14-1:0] node599;
	wire [14-1:0] node600;
	wire [14-1:0] node603;
	wire [14-1:0] node606;
	wire [14-1:0] node607;
	wire [14-1:0] node611;
	wire [14-1:0] node612;
	wire [14-1:0] node613;
	wire [14-1:0] node614;
	wire [14-1:0] node616;
	wire [14-1:0] node619;
	wire [14-1:0] node620;
	wire [14-1:0] node623;
	wire [14-1:0] node626;
	wire [14-1:0] node627;
	wire [14-1:0] node628;
	wire [14-1:0] node632;
	wire [14-1:0] node633;
	wire [14-1:0] node636;
	wire [14-1:0] node639;
	wire [14-1:0] node640;
	wire [14-1:0] node641;
	wire [14-1:0] node643;
	wire [14-1:0] node647;
	wire [14-1:0] node649;
	wire [14-1:0] node650;
	wire [14-1:0] node653;
	wire [14-1:0] node656;
	wire [14-1:0] node657;
	wire [14-1:0] node658;
	wire [14-1:0] node659;
	wire [14-1:0] node660;
	wire [14-1:0] node661;
	wire [14-1:0] node664;
	wire [14-1:0] node667;
	wire [14-1:0] node668;
	wire [14-1:0] node671;
	wire [14-1:0] node674;
	wire [14-1:0] node675;
	wire [14-1:0] node676;
	wire [14-1:0] node680;
	wire [14-1:0] node681;
	wire [14-1:0] node684;
	wire [14-1:0] node687;
	wire [14-1:0] node688;
	wire [14-1:0] node689;
	wire [14-1:0] node690;
	wire [14-1:0] node693;
	wire [14-1:0] node696;
	wire [14-1:0] node697;
	wire [14-1:0] node700;
	wire [14-1:0] node703;
	wire [14-1:0] node705;
	wire [14-1:0] node706;
	wire [14-1:0] node709;
	wire [14-1:0] node712;
	wire [14-1:0] node713;
	wire [14-1:0] node714;
	wire [14-1:0] node716;
	wire [14-1:0] node717;
	wire [14-1:0] node720;
	wire [14-1:0] node723;
	wire [14-1:0] node724;
	wire [14-1:0] node725;
	wire [14-1:0] node728;
	wire [14-1:0] node733;
	wire [14-1:0] node735;
	wire [14-1:0] node736;
	wire [14-1:0] node737;
	wire [14-1:0] node738;
	wire [14-1:0] node739;
	wire [14-1:0] node740;
	wire [14-1:0] node743;
	wire [14-1:0] node746;
	wire [14-1:0] node747;
	wire [14-1:0] node750;
	wire [14-1:0] node753;
	wire [14-1:0] node754;
	wire [14-1:0] node755;
	wire [14-1:0] node758;
	wire [14-1:0] node761;
	wire [14-1:0] node762;
	wire [14-1:0] node765;
	wire [14-1:0] node768;
	wire [14-1:0] node769;
	wire [14-1:0] node770;
	wire [14-1:0] node771;
	wire [14-1:0] node774;
	wire [14-1:0] node777;
	wire [14-1:0] node778;
	wire [14-1:0] node781;
	wire [14-1:0] node784;
	wire [14-1:0] node785;
	wire [14-1:0] node786;
	wire [14-1:0] node789;
	wire [14-1:0] node794;
	wire [14-1:0] node795;
	wire [14-1:0] node796;
	wire [14-1:0] node797;
	wire [14-1:0] node798;
	wire [14-1:0] node799;
	wire [14-1:0] node801;
	wire [14-1:0] node802;
	wire [14-1:0] node806;
	wire [14-1:0] node807;
	wire [14-1:0] node808;
	wire [14-1:0] node817;
	wire [14-1:0] node818;
	wire [14-1:0] node819;
	wire [14-1:0] node820;
	wire [14-1:0] node821;
	wire [14-1:0] node822;
	wire [14-1:0] node823;
	wire [14-1:0] node825;
	wire [14-1:0] node826;
	wire [14-1:0] node827;
	wire [14-1:0] node830;
	wire [14-1:0] node833;
	wire [14-1:0] node834;
	wire [14-1:0] node837;
	wire [14-1:0] node840;
	wire [14-1:0] node841;
	wire [14-1:0] node842;
	wire [14-1:0] node843;
	wire [14-1:0] node847;
	wire [14-1:0] node848;
	wire [14-1:0] node851;
	wire [14-1:0] node854;
	wire [14-1:0] node855;
	wire [14-1:0] node856;
	wire [14-1:0] node859;
	wire [14-1:0] node862;
	wire [14-1:0] node863;
	wire [14-1:0] node866;
	wire [14-1:0] node869;
	wire [14-1:0] node870;
	wire [14-1:0] node871;
	wire [14-1:0] node872;
	wire [14-1:0] node873;
	wire [14-1:0] node876;
	wire [14-1:0] node879;
	wire [14-1:0] node882;
	wire [14-1:0] node883;
	wire [14-1:0] node884;
	wire [14-1:0] node887;
	wire [14-1:0] node890;
	wire [14-1:0] node891;
	wire [14-1:0] node894;
	wire [14-1:0] node897;
	wire [14-1:0] node898;
	wire [14-1:0] node899;
	wire [14-1:0] node901;
	wire [14-1:0] node904;
	wire [14-1:0] node905;
	wire [14-1:0] node908;
	wire [14-1:0] node911;
	wire [14-1:0] node912;
	wire [14-1:0] node913;
	wire [14-1:0] node916;
	wire [14-1:0] node919;
	wire [14-1:0] node920;
	wire [14-1:0] node923;
	wire [14-1:0] node926;
	wire [14-1:0] node927;
	wire [14-1:0] node928;
	wire [14-1:0] node929;
	wire [14-1:0] node930;
	wire [14-1:0] node932;
	wire [14-1:0] node935;
	wire [14-1:0] node936;
	wire [14-1:0] node939;
	wire [14-1:0] node942;
	wire [14-1:0] node943;
	wire [14-1:0] node944;
	wire [14-1:0] node947;
	wire [14-1:0] node950;
	wire [14-1:0] node951;
	wire [14-1:0] node954;
	wire [14-1:0] node957;
	wire [14-1:0] node958;
	wire [14-1:0] node959;
	wire [14-1:0] node960;
	wire [14-1:0] node963;
	wire [14-1:0] node966;
	wire [14-1:0] node967;
	wire [14-1:0] node970;
	wire [14-1:0] node973;
	wire [14-1:0] node974;
	wire [14-1:0] node975;
	wire [14-1:0] node979;
	wire [14-1:0] node980;
	wire [14-1:0] node983;
	wire [14-1:0] node987;
	wire [14-1:0] node988;
	wire [14-1:0] node989;
	wire [14-1:0] node990;
	wire [14-1:0] node991;
	wire [14-1:0] node992;
	wire [14-1:0] node993;
	wire [14-1:0] node996;
	wire [14-1:0] node999;
	wire [14-1:0] node1000;
	wire [14-1:0] node1004;
	wire [14-1:0] node1005;
	wire [14-1:0] node1007;
	wire [14-1:0] node1010;
	wire [14-1:0] node1011;
	wire [14-1:0] node1014;
	wire [14-1:0] node1017;
	wire [14-1:0] node1018;
	wire [14-1:0] node1019;
	wire [14-1:0] node1020;
	wire [14-1:0] node1023;
	wire [14-1:0] node1026;
	wire [14-1:0] node1027;
	wire [14-1:0] node1030;
	wire [14-1:0] node1033;
	wire [14-1:0] node1034;
	wire [14-1:0] node1036;
	wire [14-1:0] node1039;
	wire [14-1:0] node1040;
	wire [14-1:0] node1043;
	wire [14-1:0] node1047;
	wire [14-1:0] node1048;
	wire [14-1:0] node1050;
	wire [14-1:0] node1051;
	wire [14-1:0] node1052;
	wire [14-1:0] node1053;
	wire [14-1:0] node1056;
	wire [14-1:0] node1059;
	wire [14-1:0] node1060;
	wire [14-1:0] node1063;
	wire [14-1:0] node1068;
	wire [14-1:0] node1069;
	wire [14-1:0] node1070;
	wire [14-1:0] node1071;
	wire [14-1:0] node1072;
	wire [14-1:0] node1073;
	wire [14-1:0] node1075;
	wire [14-1:0] node1076;
	wire [14-1:0] node1079;
	wire [14-1:0] node1082;
	wire [14-1:0] node1083;
	wire [14-1:0] node1085;
	wire [14-1:0] node1091;
	wire [14-1:0] node1092;
	wire [14-1:0] node1093;
	wire [14-1:0] node1094;
	wire [14-1:0] node1095;
	wire [14-1:0] node1097;
	wire [14-1:0] node1100;
	wire [14-1:0] node1101;
	wire [14-1:0] node1104;
	wire [14-1:0] node1107;
	wire [14-1:0] node1108;
	wire [14-1:0] node1109;
	wire [14-1:0] node1112;
	wire [14-1:0] node1115;
	wire [14-1:0] node1116;
	wire [14-1:0] node1119;
	wire [14-1:0] node1122;
	wire [14-1:0] node1123;
	wire [14-1:0] node1124;
	wire [14-1:0] node1125;
	wire [14-1:0] node1128;
	wire [14-1:0] node1131;
	wire [14-1:0] node1132;
	wire [14-1:0] node1135;
	wire [14-1:0] node1139;
	wire [14-1:0] node1140;
	wire [14-1:0] node1141;
	wire [14-1:0] node1142;
	wire [14-1:0] node1143;
	wire [14-1:0] node1146;
	wire [14-1:0] node1149;
	wire [14-1:0] node1150;
	wire [14-1:0] node1153;
	wire [14-1:0] node1156;
	wire [14-1:0] node1157;
	wire [14-1:0] node1159;
	wire [14-1:0] node1164;
	wire [14-1:0] node1165;
	wire [14-1:0] node1167;
	wire [14-1:0] node1168;
	wire [14-1:0] node1169;
	wire [14-1:0] node1171;
	wire [14-1:0] node1178;
	wire [14-1:0] node1179;
	wire [14-1:0] node1180;
	wire [14-1:0] node1181;
	wire [14-1:0] node1182;
	wire [14-1:0] node1183;
	wire [14-1:0] node1184;
	wire [14-1:0] node1185;
	wire [14-1:0] node1186;
	wire [14-1:0] node1187;
	wire [14-1:0] node1188;
	wire [14-1:0] node1189;
	wire [14-1:0] node1194;
	wire [14-1:0] node1195;
	wire [14-1:0] node1196;
	wire [14-1:0] node1197;
	wire [14-1:0] node1200;
	wire [14-1:0] node1203;
	wire [14-1:0] node1206;
	wire [14-1:0] node1207;
	wire [14-1:0] node1208;
	wire [14-1:0] node1211;
	wire [14-1:0] node1214;
	wire [14-1:0] node1215;
	wire [14-1:0] node1218;
	wire [14-1:0] node1221;
	wire [14-1:0] node1222;
	wire [14-1:0] node1223;
	wire [14-1:0] node1224;
	wire [14-1:0] node1226;
	wire [14-1:0] node1229;
	wire [14-1:0] node1232;
	wire [14-1:0] node1233;
	wire [14-1:0] node1235;
	wire [14-1:0] node1238;
	wire [14-1:0] node1239;
	wire [14-1:0] node1243;
	wire [14-1:0] node1244;
	wire [14-1:0] node1245;
	wire [14-1:0] node1247;
	wire [14-1:0] node1250;
	wire [14-1:0] node1252;
	wire [14-1:0] node1255;
	wire [14-1:0] node1256;
	wire [14-1:0] node1258;
	wire [14-1:0] node1261;
	wire [14-1:0] node1262;
	wire [14-1:0] node1265;
	wire [14-1:0] node1268;
	wire [14-1:0] node1269;
	wire [14-1:0] node1270;
	wire [14-1:0] node1271;
	wire [14-1:0] node1272;
	wire [14-1:0] node1274;
	wire [14-1:0] node1277;
	wire [14-1:0] node1278;
	wire [14-1:0] node1281;
	wire [14-1:0] node1284;
	wire [14-1:0] node1285;
	wire [14-1:0] node1286;
	wire [14-1:0] node1291;
	wire [14-1:0] node1292;
	wire [14-1:0] node1293;
	wire [14-1:0] node1294;
	wire [14-1:0] node1297;
	wire [14-1:0] node1300;
	wire [14-1:0] node1301;
	wire [14-1:0] node1305;
	wire [14-1:0] node1306;
	wire [14-1:0] node1308;
	wire [14-1:0] node1311;
	wire [14-1:0] node1313;
	wire [14-1:0] node1316;
	wire [14-1:0] node1317;
	wire [14-1:0] node1318;
	wire [14-1:0] node1320;
	wire [14-1:0] node1321;
	wire [14-1:0] node1324;
	wire [14-1:0] node1327;
	wire [14-1:0] node1328;
	wire [14-1:0] node1331;
	wire [14-1:0] node1333;
	wire [14-1:0] node1336;
	wire [14-1:0] node1337;
	wire [14-1:0] node1338;
	wire [14-1:0] node1339;
	wire [14-1:0] node1342;
	wire [14-1:0] node1345;
	wire [14-1:0] node1347;
	wire [14-1:0] node1350;
	wire [14-1:0] node1351;
	wire [14-1:0] node1354;
	wire [14-1:0] node1355;
	wire [14-1:0] node1359;
	wire [14-1:0] node1360;
	wire [14-1:0] node1361;
	wire [14-1:0] node1362;
	wire [14-1:0] node1363;
	wire [14-1:0] node1364;
	wire [14-1:0] node1367;
	wire [14-1:0] node1370;
	wire [14-1:0] node1371;
	wire [14-1:0] node1373;
	wire [14-1:0] node1376;
	wire [14-1:0] node1378;
	wire [14-1:0] node1381;
	wire [14-1:0] node1382;
	wire [14-1:0] node1383;
	wire [14-1:0] node1385;
	wire [14-1:0] node1388;
	wire [14-1:0] node1389;
	wire [14-1:0] node1393;
	wire [14-1:0] node1394;
	wire [14-1:0] node1395;
	wire [14-1:0] node1398;
	wire [14-1:0] node1401;
	wire [14-1:0] node1403;
	wire [14-1:0] node1408;
	wire [14-1:0] node1409;
	wire [14-1:0] node1410;
	wire [14-1:0] node1411;
	wire [14-1:0] node1412;
	wire [14-1:0] node1413;
	wire [14-1:0] node1418;
	wire [14-1:0] node1419;
	wire [14-1:0] node1420;
	wire [14-1:0] node1423;
	wire [14-1:0] node1426;
	wire [14-1:0] node1427;
	wire [14-1:0] node1430;
	wire [14-1:0] node1433;
	wire [14-1:0] node1434;
	wire [14-1:0] node1435;
	wire [14-1:0] node1437;
	wire [14-1:0] node1440;
	wire [14-1:0] node1441;
	wire [14-1:0] node1444;
	wire [14-1:0] node1447;
	wire [14-1:0] node1448;
	wire [14-1:0] node1449;
	wire [14-1:0] node1452;
	wire [14-1:0] node1455;
	wire [14-1:0] node1456;
	wire [14-1:0] node1459;
	wire [14-1:0] node1462;
	wire [14-1:0] node1463;
	wire [14-1:0] node1464;
	wire [14-1:0] node1466;
	wire [14-1:0] node1467;
	wire [14-1:0] node1470;
	wire [14-1:0] node1473;
	wire [14-1:0] node1474;
	wire [14-1:0] node1475;
	wire [14-1:0] node1478;
	wire [14-1:0] node1481;
	wire [14-1:0] node1482;
	wire [14-1:0] node1485;
	wire [14-1:0] node1488;
	wire [14-1:0] node1489;
	wire [14-1:0] node1490;
	wire [14-1:0] node1491;
	wire [14-1:0] node1494;
	wire [14-1:0] node1497;
	wire [14-1:0] node1498;
	wire [14-1:0] node1501;
	wire [14-1:0] node1504;
	wire [14-1:0] node1505;
	wire [14-1:0] node1506;
	wire [14-1:0] node1509;
	wire [14-1:0] node1512;
	wire [14-1:0] node1513;
	wire [14-1:0] node1516;
	wire [14-1:0] node1519;
	wire [14-1:0] node1520;
	wire [14-1:0] node1521;
	wire [14-1:0] node1522;
	wire [14-1:0] node1523;
	wire [14-1:0] node1524;
	wire [14-1:0] node1525;
	wire [14-1:0] node1527;
	wire [14-1:0] node1528;
	wire [14-1:0] node1531;
	wire [14-1:0] node1534;
	wire [14-1:0] node1535;
	wire [14-1:0] node1536;
	wire [14-1:0] node1539;
	wire [14-1:0] node1542;
	wire [14-1:0] node1543;
	wire [14-1:0] node1547;
	wire [14-1:0] node1548;
	wire [14-1:0] node1549;
	wire [14-1:0] node1551;
	wire [14-1:0] node1554;
	wire [14-1:0] node1555;
	wire [14-1:0] node1558;
	wire [14-1:0] node1561;
	wire [14-1:0] node1562;
	wire [14-1:0] node1563;
	wire [14-1:0] node1566;
	wire [14-1:0] node1569;
	wire [14-1:0] node1571;
	wire [14-1:0] node1574;
	wire [14-1:0] node1575;
	wire [14-1:0] node1576;
	wire [14-1:0] node1577;
	wire [14-1:0] node1579;
	wire [14-1:0] node1582;
	wire [14-1:0] node1585;
	wire [14-1:0] node1586;
	wire [14-1:0] node1587;
	wire [14-1:0] node1591;
	wire [14-1:0] node1595;
	wire [14-1:0] node1596;
	wire [14-1:0] node1597;
	wire [14-1:0] node1599;
	wire [14-1:0] node1602;
	wire [14-1:0] node1603;
	wire [14-1:0] node1606;
	wire [14-1:0] node1609;
	wire [14-1:0] node1610;
	wire [14-1:0] node1611;
	wire [14-1:0] node1614;
	wire [14-1:0] node1617;
	wire [14-1:0] node1618;
	wire [14-1:0] node1621;
	wire [14-1:0] node1624;
	wire [14-1:0] node1625;
	wire [14-1:0] node1626;
	wire [14-1:0] node1627;
	wire [14-1:0] node1628;
	wire [14-1:0] node1629;
	wire [14-1:0] node1631;
	wire [14-1:0] node1634;
	wire [14-1:0] node1636;
	wire [14-1:0] node1639;
	wire [14-1:0] node1640;
	wire [14-1:0] node1641;
	wire [14-1:0] node1644;
	wire [14-1:0] node1647;
	wire [14-1:0] node1649;
	wire [14-1:0] node1652;
	wire [14-1:0] node1653;
	wire [14-1:0] node1654;
	wire [14-1:0] node1656;
	wire [14-1:0] node1659;
	wire [14-1:0] node1660;
	wire [14-1:0] node1663;
	wire [14-1:0] node1666;
	wire [14-1:0] node1667;
	wire [14-1:0] node1668;
	wire [14-1:0] node1672;
	wire [14-1:0] node1673;
	wire [14-1:0] node1676;
	wire [14-1:0] node1681;
	wire [14-1:0] node1682;
	wire [14-1:0] node1683;
	wire [14-1:0] node1684;
	wire [14-1:0] node1685;
	wire [14-1:0] node1686;
	wire [14-1:0] node1687;
	wire [14-1:0] node1690;
	wire [14-1:0] node1693;
	wire [14-1:0] node1694;
	wire [14-1:0] node1696;
	wire [14-1:0] node1699;
	wire [14-1:0] node1701;
	wire [14-1:0] node1704;
	wire [14-1:0] node1705;
	wire [14-1:0] node1706;
	wire [14-1:0] node1709;
	wire [14-1:0] node1711;
	wire [14-1:0] node1714;
	wire [14-1:0] node1715;
	wire [14-1:0] node1716;
	wire [14-1:0] node1719;
	wire [14-1:0] node1722;
	wire [14-1:0] node1725;
	wire [14-1:0] node1727;
	wire [14-1:0] node1728;
	wire [14-1:0] node1730;
	wire [14-1:0] node1732;
	wire [14-1:0] node1735;
	wire [14-1:0] node1736;
	wire [14-1:0] node1737;
	wire [14-1:0] node1741;
	wire [14-1:0] node1744;
	wire [14-1:0] node1746;
	wire [14-1:0] node1747;
	wire [14-1:0] node1748;
	wire [14-1:0] node1749;
	wire [14-1:0] node1752;
	wire [14-1:0] node1755;
	wire [14-1:0] node1756;
	wire [14-1:0] node1759;
	wire [14-1:0] node1763;
	wire [14-1:0] node1765;
	wire [14-1:0] node1766;
	wire [14-1:0] node1768;
	wire [14-1:0] node1769;
	wire [14-1:0] node1770;
	wire [14-1:0] node1773;
	wire [14-1:0] node1776;
	wire [14-1:0] node1777;
	wire [14-1:0] node1780;
	wire [14-1:0] node1784;
	wire [14-1:0] node1785;
	wire [14-1:0] node1786;
	wire [14-1:0] node1787;
	wire [14-1:0] node1788;
	wire [14-1:0] node1789;
	wire [14-1:0] node1790;
	wire [14-1:0] node1791;
	wire [14-1:0] node1793;
	wire [14-1:0] node1794;
	wire [14-1:0] node1797;
	wire [14-1:0] node1800;
	wire [14-1:0] node1801;
	wire [14-1:0] node1804;
	wire [14-1:0] node1806;
	wire [14-1:0] node1809;
	wire [14-1:0] node1810;
	wire [14-1:0] node1811;
	wire [14-1:0] node1812;
	wire [14-1:0] node1816;
	wire [14-1:0] node1817;
	wire [14-1:0] node1821;
	wire [14-1:0] node1822;
	wire [14-1:0] node1824;
	wire [14-1:0] node1827;
	wire [14-1:0] node1828;
	wire [14-1:0] node1832;
	wire [14-1:0] node1833;
	wire [14-1:0] node1834;
	wire [14-1:0] node1835;
	wire [14-1:0] node1837;
	wire [14-1:0] node1840;
	wire [14-1:0] node1843;
	wire [14-1:0] node1844;
	wire [14-1:0] node1845;
	wire [14-1:0] node1849;
	wire [14-1:0] node1850;
	wire [14-1:0] node1853;
	wire [14-1:0] node1856;
	wire [14-1:0] node1857;
	wire [14-1:0] node1858;
	wire [14-1:0] node1859;
	wire [14-1:0] node1864;
	wire [14-1:0] node1865;
	wire [14-1:0] node1867;
	wire [14-1:0] node1870;
	wire [14-1:0] node1871;
	wire [14-1:0] node1874;
	wire [14-1:0] node1877;
	wire [14-1:0] node1878;
	wire [14-1:0] node1879;
	wire [14-1:0] node1880;
	wire [14-1:0] node1882;
	wire [14-1:0] node1884;
	wire [14-1:0] node1887;
	wire [14-1:0] node1888;
	wire [14-1:0] node1890;
	wire [14-1:0] node1893;
	wire [14-1:0] node1894;
	wire [14-1:0] node1897;
	wire [14-1:0] node1900;
	wire [14-1:0] node1901;
	wire [14-1:0] node1902;
	wire [14-1:0] node1903;
	wire [14-1:0] node1906;
	wire [14-1:0] node1909;
	wire [14-1:0] node1911;
	wire [14-1:0] node1914;
	wire [14-1:0] node1915;
	wire [14-1:0] node1918;
	wire [14-1:0] node1919;
	wire [14-1:0] node1922;
	wire [14-1:0] node1926;
	wire [14-1:0] node1927;
	wire [14-1:0] node1928;
	wire [14-1:0] node1930;
	wire [14-1:0] node1931;
	wire [14-1:0] node1934;
	wire [14-1:0] node1937;
	wire [14-1:0] node1938;
	wire [14-1:0] node1939;
	wire [14-1:0] node1942;
	wire [14-1:0] node1945;
	wire [14-1:0] node1946;
	wire [14-1:0] node1949;
	wire [14-1:0] node1952;
	wire [14-1:0] node1953;
	wire [14-1:0] node1954;
	wire [14-1:0] node1955;
	wire [14-1:0] node1958;
	wire [14-1:0] node1961;
	wire [14-1:0] node1962;
	wire [14-1:0] node1965;
	wire [14-1:0] node1968;
	wire [14-1:0] node1969;
	wire [14-1:0] node1970;
	wire [14-1:0] node1973;
	wire [14-1:0] node1976;
	wire [14-1:0] node1977;
	wire [14-1:0] node1980;
	wire [14-1:0] node1983;
	wire [14-1:0] node1984;
	wire [14-1:0] node1985;
	wire [14-1:0] node1986;
	wire [14-1:0] node1987;
	wire [14-1:0] node1988;
	wire [14-1:0] node1990;
	wire [14-1:0] node1991;
	wire [14-1:0] node1994;
	wire [14-1:0] node1997;
	wire [14-1:0] node1998;
	wire [14-1:0] node1999;
	wire [14-1:0] node2002;
	wire [14-1:0] node2005;
	wire [14-1:0] node2008;
	wire [14-1:0] node2009;
	wire [14-1:0] node2010;
	wire [14-1:0] node2012;
	wire [14-1:0] node2015;
	wire [14-1:0] node2018;
	wire [14-1:0] node2019;
	wire [14-1:0] node2020;
	wire [14-1:0] node2023;
	wire [14-1:0] node2026;
	wire [14-1:0] node2027;
	wire [14-1:0] node2030;
	wire [14-1:0] node2033;
	wire [14-1:0] node2034;
	wire [14-1:0] node2035;
	wire [14-1:0] node2036;
	wire [14-1:0] node2039;
	wire [14-1:0] node2041;
	wire [14-1:0] node2044;
	wire [14-1:0] node2045;
	wire [14-1:0] node2048;
	wire [14-1:0] node2049;
	wire [14-1:0] node2052;
	wire [14-1:0] node2055;
	wire [14-1:0] node2056;
	wire [14-1:0] node2057;
	wire [14-1:0] node2058;
	wire [14-1:0] node2061;
	wire [14-1:0] node2064;
	wire [14-1:0] node2065;
	wire [14-1:0] node2069;
	wire [14-1:0] node2070;
	wire [14-1:0] node2072;
	wire [14-1:0] node2075;
	wire [14-1:0] node2076;
	wire [14-1:0] node2079;
	wire [14-1:0] node2082;
	wire [14-1:0] node2084;
	wire [14-1:0] node2085;
	wire [14-1:0] node2086;
	wire [14-1:0] node2087;
	wire [14-1:0] node2088;
	wire [14-1:0] node2091;
	wire [14-1:0] node2094;
	wire [14-1:0] node2095;
	wire [14-1:0] node2099;
	wire [14-1:0] node2100;
	wire [14-1:0] node2101;
	wire [14-1:0] node2105;
	wire [14-1:0] node2106;
	wire [14-1:0] node2111;
	wire [14-1:0] node2113;
	wire [14-1:0] node2114;
	wire [14-1:0] node2115;
	wire [14-1:0] node2117;
	wire [14-1:0] node2122;
	wire [14-1:0] node2123;
	wire [14-1:0] node2124;
	wire [14-1:0] node2125;
	wire [14-1:0] node2126;
	wire [14-1:0] node2128;
	wire [14-1:0] node2129;
	wire [14-1:0] node2130;
	wire [14-1:0] node2132;
	wire [14-1:0] node2135;
	wire [14-1:0] node2138;
	wire [14-1:0] node2139;
	wire [14-1:0] node2140;
	wire [14-1:0] node2143;
	wire [14-1:0] node2146;
	wire [14-1:0] node2147;
	wire [14-1:0] node2151;
	wire [14-1:0] node2152;
	wire [14-1:0] node2153;
	wire [14-1:0] node2154;
	wire [14-1:0] node2156;
	wire [14-1:0] node2159;
	wire [14-1:0] node2160;
	wire [14-1:0] node2164;
	wire [14-1:0] node2165;
	wire [14-1:0] node2167;
	wire [14-1:0] node2170;
	wire [14-1:0] node2171;
	wire [14-1:0] node2174;
	wire [14-1:0] node2178;
	wire [14-1:0] node2179;
	wire [14-1:0] node2180;
	wire [14-1:0] node2182;
	wire [14-1:0] node2185;
	wire [14-1:0] node2186;
	wire [14-1:0] node2189;
	wire [14-1:0] node2192;
	wire [14-1:0] node2193;
	wire [14-1:0] node2194;
	wire [14-1:0] node2197;
	wire [14-1:0] node2200;
	wire [14-1:0] node2201;
	wire [14-1:0] node2204;
	wire [14-1:0] node2207;
	wire [14-1:0] node2208;
	wire [14-1:0] node2209;
	wire [14-1:0] node2210;
	wire [14-1:0] node2211;
	wire [14-1:0] node2212;
	wire [14-1:0] node2214;
	wire [14-1:0] node2217;
	wire [14-1:0] node2218;
	wire [14-1:0] node2222;
	wire [14-1:0] node2223;
	wire [14-1:0] node2226;
	wire [14-1:0] node2227;
	wire [14-1:0] node2231;
	wire [14-1:0] node2232;
	wire [14-1:0] node2233;
	wire [14-1:0] node2234;
	wire [14-1:0] node2237;
	wire [14-1:0] node2240;
	wire [14-1:0] node2242;
	wire [14-1:0] node2245;
	wire [14-1:0] node2246;
	wire [14-1:0] node2249;
	wire [14-1:0] node2250;
	wire [14-1:0] node2253;
	wire [14-1:0] node2258;
	wire [14-1:0] node2259;
	wire [14-1:0] node2261;
	wire [14-1:0] node2263;
	wire [14-1:0] node2265;
	wire [14-1:0] node2267;
	wire [14-1:0] node2268;
	wire [14-1:0] node2273;
	wire [14-1:0] node2274;
	wire [14-1:0] node2275;
	wire [14-1:0] node2276;
	wire [14-1:0] node2277;
	wire [14-1:0] node2278;
	wire [14-1:0] node2279;
	wire [14-1:0] node2280;
	wire [14-1:0] node2281;
	wire [14-1:0] node2283;
	wire [14-1:0] node2285;
	wire [14-1:0] node2288;
	wire [14-1:0] node2289;
	wire [14-1:0] node2290;
	wire [14-1:0] node2293;
	wire [14-1:0] node2296;
	wire [14-1:0] node2297;
	wire [14-1:0] node2300;
	wire [14-1:0] node2303;
	wire [14-1:0] node2304;
	wire [14-1:0] node2305;
	wire [14-1:0] node2306;
	wire [14-1:0] node2309;
	wire [14-1:0] node2312;
	wire [14-1:0] node2313;
	wire [14-1:0] node2317;
	wire [14-1:0] node2318;
	wire [14-1:0] node2319;
	wire [14-1:0] node2322;
	wire [14-1:0] node2325;
	wire [14-1:0] node2327;
	wire [14-1:0] node2330;
	wire [14-1:0] node2331;
	wire [14-1:0] node2332;
	wire [14-1:0] node2333;
	wire [14-1:0] node2335;
	wire [14-1:0] node2339;
	wire [14-1:0] node2340;
	wire [14-1:0] node2341;
	wire [14-1:0] node2345;
	wire [14-1:0] node2346;
	wire [14-1:0] node2350;
	wire [14-1:0] node2351;
	wire [14-1:0] node2352;
	wire [14-1:0] node2356;
	wire [14-1:0] node2358;
	wire [14-1:0] node2359;
	wire [14-1:0] node2362;
	wire [14-1:0] node2365;
	wire [14-1:0] node2366;
	wire [14-1:0] node2367;
	wire [14-1:0] node2368;
	wire [14-1:0] node2369;
	wire [14-1:0] node2370;
	wire [14-1:0] node2374;
	wire [14-1:0] node2375;
	wire [14-1:0] node2378;
	wire [14-1:0] node2381;
	wire [14-1:0] node2382;
	wire [14-1:0] node2383;
	wire [14-1:0] node2387;
	wire [14-1:0] node2388;
	wire [14-1:0] node2391;
	wire [14-1:0] node2394;
	wire [14-1:0] node2395;
	wire [14-1:0] node2396;
	wire [14-1:0] node2399;
	wire [14-1:0] node2401;
	wire [14-1:0] node2404;
	wire [14-1:0] node2406;
	wire [14-1:0] node2408;
	wire [14-1:0] node2411;
	wire [14-1:0] node2412;
	wire [14-1:0] node2413;
	wire [14-1:0] node2415;
	wire [14-1:0] node2416;
	wire [14-1:0] node2420;
	wire [14-1:0] node2421;
	wire [14-1:0] node2422;
	wire [14-1:0] node2425;
	wire [14-1:0] node2430;
	wire [14-1:0] node2431;
	wire [14-1:0] node2432;
	wire [14-1:0] node2433;
	wire [14-1:0] node2434;
	wire [14-1:0] node2435;
	wire [14-1:0] node2436;
	wire [14-1:0] node2440;
	wire [14-1:0] node2443;
	wire [14-1:0] node2444;
	wire [14-1:0] node2445;
	wire [14-1:0] node2449;
	wire [14-1:0] node2450;
	wire [14-1:0] node2454;
	wire [14-1:0] node2455;
	wire [14-1:0] node2456;
	wire [14-1:0] node2459;
	wire [14-1:0] node2460;
	wire [14-1:0] node2463;
	wire [14-1:0] node2466;
	wire [14-1:0] node2467;
	wire [14-1:0] node2468;
	wire [14-1:0] node2471;
	wire [14-1:0] node2474;
	wire [14-1:0] node2476;
	wire [14-1:0] node2479;
	wire [14-1:0] node2481;
	wire [14-1:0] node2482;
	wire [14-1:0] node2483;
	wire [14-1:0] node2485;
	wire [14-1:0] node2488;
	wire [14-1:0] node2490;
	wire [14-1:0] node2495;
	wire [14-1:0] node2496;
	wire [14-1:0] node2497;
	wire [14-1:0] node2498;
	wire [14-1:0] node2499;
	wire [14-1:0] node2501;
	wire [14-1:0] node2504;
	wire [14-1:0] node2505;
	wire [14-1:0] node2508;
	wire [14-1:0] node2511;
	wire [14-1:0] node2512;
	wire [14-1:0] node2513;
	wire [14-1:0] node2516;
	wire [14-1:0] node2520;
	wire [14-1:0] node2521;
	wire [14-1:0] node2522;
	wire [14-1:0] node2523;
	wire [14-1:0] node2526;
	wire [14-1:0] node2529;
	wire [14-1:0] node2530;
	wire [14-1:0] node2532;
	wire [14-1:0] node2535;
	wire [14-1:0] node2536;
	wire [14-1:0] node2539;
	wire [14-1:0] node2542;
	wire [14-1:0] node2543;
	wire [14-1:0] node2544;
	wire [14-1:0] node2547;
	wire [14-1:0] node2550;
	wire [14-1:0] node2551;
	wire [14-1:0] node2555;
	wire [14-1:0] node2556;
	wire [14-1:0] node2557;
	wire [14-1:0] node2558;
	wire [14-1:0] node2559;
	wire [14-1:0] node2562;
	wire [14-1:0] node2565;
	wire [14-1:0] node2566;
	wire [14-1:0] node2569;
	wire [14-1:0] node2572;
	wire [14-1:0] node2574;
	wire [14-1:0] node2575;
	wire [14-1:0] node2578;
	wire [14-1:0] node2582;
	wire [14-1:0] node2583;
	wire [14-1:0] node2584;
	wire [14-1:0] node2585;
	wire [14-1:0] node2586;
	wire [14-1:0] node2587;
	wire [14-1:0] node2588;
	wire [14-1:0] node2589;
	wire [14-1:0] node2598;
	wire [14-1:0] node2599;
	wire [14-1:0] node2600;
	wire [14-1:0] node2601;
	wire [14-1:0] node2602;
	wire [14-1:0] node2603;
	wire [14-1:0] node2606;
	wire [14-1:0] node2609;
	wire [14-1:0] node2610;
	wire [14-1:0] node2613;
	wire [14-1:0] node2616;
	wire [14-1:0] node2617;
	wire [14-1:0] node2618;
	wire [14-1:0] node2621;
	wire [14-1:0] node2624;
	wire [14-1:0] node2625;
	wire [14-1:0] node2628;
	wire [14-1:0] node2631;
	wire [14-1:0] node2632;
	wire [14-1:0] node2633;
	wire [14-1:0] node2634;
	wire [14-1:0] node2637;
	wire [14-1:0] node2640;
	wire [14-1:0] node2641;
	wire [14-1:0] node2644;
	wire [14-1:0] node2648;
	wire [14-1:0] node2649;
	wire [14-1:0] node2650;
	wire [14-1:0] node2651;
	wire [14-1:0] node2652;
	wire [14-1:0] node2655;
	wire [14-1:0] node2658;
	wire [14-1:0] node2659;
	wire [14-1:0] node2662;
	wire [14-1:0] node2667;
	wire [14-1:0] node2668;
	wire [14-1:0] node2669;
	wire [14-1:0] node2670;
	wire [14-1:0] node2671;
	wire [14-1:0] node2673;
	wire [14-1:0] node2674;
	wire [14-1:0] node2675;
	wire [14-1:0] node2676;
	wire [14-1:0] node2677;
	wire [14-1:0] node2680;
	wire [14-1:0] node2683;
	wire [14-1:0] node2684;
	wire [14-1:0] node2688;
	wire [14-1:0] node2689;
	wire [14-1:0] node2691;
	wire [14-1:0] node2694;
	wire [14-1:0] node2695;
	wire [14-1:0] node2698;
	wire [14-1:0] node2701;
	wire [14-1:0] node2702;
	wire [14-1:0] node2704;
	wire [14-1:0] node2705;
	wire [14-1:0] node2709;
	wire [14-1:0] node2710;
	wire [14-1:0] node2711;
	wire [14-1:0] node2714;
	wire [14-1:0] node2718;
	wire [14-1:0] node2719;
	wire [14-1:0] node2720;
	wire [14-1:0] node2721;
	wire [14-1:0] node2722;
	wire [14-1:0] node2723;
	wire [14-1:0] node2727;
	wire [14-1:0] node2728;
	wire [14-1:0] node2731;
	wire [14-1:0] node2734;
	wire [14-1:0] node2735;
	wire [14-1:0] node2737;
	wire [14-1:0] node2740;
	wire [14-1:0] node2741;
	wire [14-1:0] node2744;
	wire [14-1:0] node2747;
	wire [14-1:0] node2748;
	wire [14-1:0] node2750;
	wire [14-1:0] node2752;
	wire [14-1:0] node2755;
	wire [14-1:0] node2756;
	wire [14-1:0] node2757;
	wire [14-1:0] node2762;
	wire [14-1:0] node2763;
	wire [14-1:0] node2764;
	wire [14-1:0] node2765;
	wire [14-1:0] node2767;
	wire [14-1:0] node2770;
	wire [14-1:0] node2771;
	wire [14-1:0] node2774;
	wire [14-1:0] node2777;
	wire [14-1:0] node2778;
	wire [14-1:0] node2779;
	wire [14-1:0] node2783;
	wire [14-1:0] node2785;
	wire [14-1:0] node2788;
	wire [14-1:0] node2789;
	wire [14-1:0] node2790;
	wire [14-1:0] node2792;
	wire [14-1:0] node2797;
	wire [14-1:0] node2798;
	wire [14-1:0] node2799;
	wire [14-1:0] node2800;
	wire [14-1:0] node2802;
	wire [14-1:0] node2804;
	wire [14-1:0] node2807;
	wire [14-1:0] node2808;
	wire [14-1:0] node2809;
	wire [14-1:0] node2810;
	wire [14-1:0] node2813;
	wire [14-1:0] node2816;
	wire [14-1:0] node2817;
	wire [14-1:0] node2820;
	wire [14-1:0] node2823;
	wire [14-1:0] node2824;
	wire [14-1:0] node2827;
	wire [14-1:0] node2828;
	wire [14-1:0] node2831;
	wire [14-1:0] node2834;
	wire [14-1:0] node2835;
	wire [14-1:0] node2836;
	wire [14-1:0] node2837;
	wire [14-1:0] node2838;
	wire [14-1:0] node2843;
	wire [14-1:0] node2844;
	wire [14-1:0] node2847;
	wire [14-1:0] node2849;
	wire [14-1:0] node2854;
	wire [14-1:0] node2855;
	wire [14-1:0] node2856;
	wire [14-1:0] node2857;
	wire [14-1:0] node2859;
	wire [14-1:0] node2860;
	wire [14-1:0] node2863;
	wire [14-1:0] node2866;
	wire [14-1:0] node2867;
	wire [14-1:0] node2868;
	wire [14-1:0] node2874;
	wire [14-1:0] node2875;
	wire [14-1:0] node2877;
	wire [14-1:0] node2879;
	wire [14-1:0] node2881;
	wire [14-1:0] node2886;
	wire [14-1:0] node2887;
	wire [14-1:0] node2888;
	wire [14-1:0] node2889;
	wire [14-1:0] node2890;
	wire [14-1:0] node2891;
	wire [14-1:0] node2892;
	wire [14-1:0] node2893;
	wire [14-1:0] node2894;
	wire [14-1:0] node2895;
	wire [14-1:0] node2897;
	wire [14-1:0] node2900;
	wire [14-1:0] node2901;
	wire [14-1:0] node2902;
	wire [14-1:0] node2905;
	wire [14-1:0] node2908;
	wire [14-1:0] node2909;
	wire [14-1:0] node2913;
	wire [14-1:0] node2914;
	wire [14-1:0] node2915;
	wire [14-1:0] node2916;
	wire [14-1:0] node2919;
	wire [14-1:0] node2922;
	wire [14-1:0] node2923;
	wire [14-1:0] node2926;
	wire [14-1:0] node2929;
	wire [14-1:0] node2930;
	wire [14-1:0] node2933;
	wire [14-1:0] node2934;
	wire [14-1:0] node2938;
	wire [14-1:0] node2939;
	wire [14-1:0] node2940;
	wire [14-1:0] node2943;
	wire [14-1:0] node2944;
	wire [14-1:0] node2945;
	wire [14-1:0] node2949;
	wire [14-1:0] node2951;
	wire [14-1:0] node2954;
	wire [14-1:0] node2955;
	wire [14-1:0] node2956;
	wire [14-1:0] node2957;
	wire [14-1:0] node2960;
	wire [14-1:0] node2963;
	wire [14-1:0] node2964;
	wire [14-1:0] node2967;
	wire [14-1:0] node2970;
	wire [14-1:0] node2971;
	wire [14-1:0] node2972;
	wire [14-1:0] node2976;
	wire [14-1:0] node2979;
	wire [14-1:0] node2980;
	wire [14-1:0] node2981;
	wire [14-1:0] node2982;
	wire [14-1:0] node2983;
	wire [14-1:0] node2984;
	wire [14-1:0] node2987;
	wire [14-1:0] node2990;
	wire [14-1:0] node2991;
	wire [14-1:0] node2994;
	wire [14-1:0] node2997;
	wire [14-1:0] node2998;
	wire [14-1:0] node2999;
	wire [14-1:0] node3004;
	wire [14-1:0] node3005;
	wire [14-1:0] node3006;
	wire [14-1:0] node3007;
	wire [14-1:0] node3010;
	wire [14-1:0] node3013;
	wire [14-1:0] node3015;
	wire [14-1:0] node3018;
	wire [14-1:0] node3020;
	wire [14-1:0] node3021;
	wire [14-1:0] node3024;
	wire [14-1:0] node3027;
	wire [14-1:0] node3028;
	wire [14-1:0] node3029;
	wire [14-1:0] node3031;
	wire [14-1:0] node3032;
	wire [14-1:0] node3036;
	wire [14-1:0] node3037;
	wire [14-1:0] node3042;
	wire [14-1:0] node3043;
	wire [14-1:0] node3044;
	wire [14-1:0] node3045;
	wire [14-1:0] node3046;
	wire [14-1:0] node3047;
	wire [14-1:0] node3049;
	wire [14-1:0] node3052;
	wire [14-1:0] node3053;
	wire [14-1:0] node3057;
	wire [14-1:0] node3058;
	wire [14-1:0] node3061;
	wire [14-1:0] node3064;
	wire [14-1:0] node3065;
	wire [14-1:0] node3066;
	wire [14-1:0] node3067;
	wire [14-1:0] node3070;
	wire [14-1:0] node3073;
	wire [14-1:0] node3074;
	wire [14-1:0] node3078;
	wire [14-1:0] node3079;
	wire [14-1:0] node3080;
	wire [14-1:0] node3083;
	wire [14-1:0] node3086;
	wire [14-1:0] node3089;
	wire [14-1:0] node3090;
	wire [14-1:0] node3092;
	wire [14-1:0] node3093;
	wire [14-1:0] node3094;
	wire [14-1:0] node3098;
	wire [14-1:0] node3099;
	wire [14-1:0] node3105;
	wire [14-1:0] node3106;
	wire [14-1:0] node3107;
	wire [14-1:0] node3108;
	wire [14-1:0] node3110;
	wire [14-1:0] node3111;
	wire [14-1:0] node3114;
	wire [14-1:0] node3117;
	wire [14-1:0] node3118;
	wire [14-1:0] node3119;
	wire [14-1:0] node3122;
	wire [14-1:0] node3126;
	wire [14-1:0] node3127;
	wire [14-1:0] node3128;
	wire [14-1:0] node3129;
	wire [14-1:0] node3132;
	wire [14-1:0] node3135;
	wire [14-1:0] node3136;
	wire [14-1:0] node3139;
	wire [14-1:0] node3142;
	wire [14-1:0] node3143;
	wire [14-1:0] node3144;
	wire [14-1:0] node3147;
	wire [14-1:0] node3151;
	wire [14-1:0] node3152;
	wire [14-1:0] node3153;
	wire [14-1:0] node3154;
	wire [14-1:0] node3155;
	wire [14-1:0] node3158;
	wire [14-1:0] node3161;
	wire [14-1:0] node3162;
	wire [14-1:0] node3165;
	wire [14-1:0] node3168;
	wire [14-1:0] node3170;
	wire [14-1:0] node3171;
	wire [14-1:0] node3174;
	wire [14-1:0] node3178;
	wire [14-1:0] node3179;
	wire [14-1:0] node3180;
	wire [14-1:0] node3181;
	wire [14-1:0] node3182;
	wire [14-1:0] node3183;
	wire [14-1:0] node3184;
	wire [14-1:0] node3186;
	wire [14-1:0] node3188;
	wire [14-1:0] node3191;
	wire [14-1:0] node3192;
	wire [14-1:0] node3193;
	wire [14-1:0] node3196;
	wire [14-1:0] node3199;
	wire [14-1:0] node3200;
	wire [14-1:0] node3203;
	wire [14-1:0] node3206;
	wire [14-1:0] node3207;
	wire [14-1:0] node3208;
	wire [14-1:0] node3209;
	wire [14-1:0] node3212;
	wire [14-1:0] node3215;
	wire [14-1:0] node3217;
	wire [14-1:0] node3220;
	wire [14-1:0] node3221;
	wire [14-1:0] node3222;
	wire [14-1:0] node3226;
	wire [14-1:0] node3229;
	wire [14-1:0] node3230;
	wire [14-1:0] node3231;
	wire [14-1:0] node3232;
	wire [14-1:0] node3236;
	wire [14-1:0] node3237;
	wire [14-1:0] node3238;
	wire [14-1:0] node3241;
	wire [14-1:0] node3244;
	wire [14-1:0] node3247;
	wire [14-1:0] node3248;
	wire [14-1:0] node3249;
	wire [14-1:0] node3251;
	wire [14-1:0] node3254;
	wire [14-1:0] node3258;
	wire [14-1:0] node3259;
	wire [14-1:0] node3260;
	wire [14-1:0] node3261;
	wire [14-1:0] node3262;
	wire [14-1:0] node3265;
	wire [14-1:0] node3267;
	wire [14-1:0] node3270;
	wire [14-1:0] node3271;
	wire [14-1:0] node3272;
	wire [14-1:0] node3275;
	wire [14-1:0] node3278;
	wire [14-1:0] node3279;
	wire [14-1:0] node3283;
	wire [14-1:0] node3285;
	wire [14-1:0] node3286;
	wire [14-1:0] node3288;
	wire [14-1:0] node3293;
	wire [14-1:0] node3294;
	wire [14-1:0] node3296;
	wire [14-1:0] node3297;
	wire [14-1:0] node3299;
	wire [14-1:0] node3303;
	wire [14-1:0] node3304;
	wire [14-1:0] node3305;
	wire [14-1:0] node3306;
	wire [14-1:0] node3309;
	wire [14-1:0] node3312;
	wire [14-1:0] node3313;
	wire [14-1:0] node3316;
	wire [14-1:0] node3319;
	wire [14-1:0] node3320;
	wire [14-1:0] node3321;
	wire [14-1:0] node3324;
	wire [14-1:0] node3329;
	wire [14-1:0] node3330;
	wire [14-1:0] node3331;
	wire [14-1:0] node3332;
	wire [14-1:0] node3333;
	wire [14-1:0] node3334;
	wire [14-1:0] node3335;
	wire [14-1:0] node3336;
	wire [14-1:0] node3337;
	wire [14-1:0] node3338;
	wire [14-1:0] node3342;
	wire [14-1:0] node3343;
	wire [14-1:0] node3347;
	wire [14-1:0] node3348;
	wire [14-1:0] node3349;
	wire [14-1:0] node3352;
	wire [14-1:0] node3355;
	wire [14-1:0] node3358;
	wire [14-1:0] node3359;
	wire [14-1:0] node3360;
	wire [14-1:0] node3361;
	wire [14-1:0] node3364;
	wire [14-1:0] node3367;
	wire [14-1:0] node3368;
	wire [14-1:0] node3371;
	wire [14-1:0] node3374;
	wire [14-1:0] node3375;
	wire [14-1:0] node3376;
	wire [14-1:0] node3381;
	wire [14-1:0] node3382;
	wire [14-1:0] node3383;
	wire [14-1:0] node3384;
	wire [14-1:0] node3385;
	wire [14-1:0] node3388;
	wire [14-1:0] node3391;
	wire [14-1:0] node3392;
	wire [14-1:0] node3395;
	wire [14-1:0] node3398;
	wire [14-1:0] node3399;
	wire [14-1:0] node3401;
	wire [14-1:0] node3404;
	wire [14-1:0] node3406;
	wire [14-1:0] node3409;
	wire [14-1:0] node3410;
	wire [14-1:0] node3411;
	wire [14-1:0] node3414;
	wire [14-1:0] node3417;
	wire [14-1:0] node3418;
	wire [14-1:0] node3421;
	wire [14-1:0] node3424;
	wire [14-1:0] node3425;
	wire [14-1:0] node3426;
	wire [14-1:0] node3427;
	wire [14-1:0] node3428;
	wire [14-1:0] node3430;
	wire [14-1:0] node3433;
	wire [14-1:0] node3434;
	wire [14-1:0] node3438;
	wire [14-1:0] node3439;
	wire [14-1:0] node3440;
	wire [14-1:0] node3443;
	wire [14-1:0] node3446;
	wire [14-1:0] node3448;
	wire [14-1:0] node3451;
	wire [14-1:0] node3452;
	wire [14-1:0] node3454;
	wire [14-1:0] node3455;
	wire [14-1:0] node3458;
	wire [14-1:0] node3463;
	wire [14-1:0] node3465;
	wire [14-1:0] node3466;
	wire [14-1:0] node3467;
	wire [14-1:0] node3468;
	wire [14-1:0] node3469;
	wire [14-1:0] node3472;
	wire [14-1:0] node3474;
	wire [14-1:0] node3477;
	wire [14-1:0] node3478;
	wire [14-1:0] node3479;
	wire [14-1:0] node3482;
	wire [14-1:0] node3485;
	wire [14-1:0] node3486;
	wire [14-1:0] node3490;
	wire [14-1:0] node3491;
	wire [14-1:0] node3492;
	wire [14-1:0] node3494;
	wire [14-1:0] node3498;
	wire [14-1:0] node3500;
	wire [14-1:0] node3503;
	wire [14-1:0] node3504;
	wire [14-1:0] node3505;
	wire [14-1:0] node3506;
	wire [14-1:0] node3507;
	wire [14-1:0] node3510;
	wire [14-1:0] node3513;
	wire [14-1:0] node3516;
	wire [14-1:0] node3517;
	wire [14-1:0] node3519;
	wire [14-1:0] node3524;
	wire [14-1:0] node3525;
	wire [14-1:0] node3526;
	wire [14-1:0] node3527;
	wire [14-1:0] node3529;
	wire [14-1:0] node3531;
	wire [14-1:0] node3532;
	wire [14-1:0] node3537;
	wire [14-1:0] node3538;
	wire [14-1:0] node3539;
	wire [14-1:0] node3540;
	wire [14-1:0] node3541;
	wire [14-1:0] node3544;
	wire [14-1:0] node3545;
	wire [14-1:0] node3548;
	wire [14-1:0] node3551;
	wire [14-1:0] node3552;
	wire [14-1:0] node3554;
	wire [14-1:0] node3557;
	wire [14-1:0] node3559;
	wire [14-1:0] node3562;
	wire [14-1:0] node3563;
	wire [14-1:0] node3564;
	wire [14-1:0] node3567;
	wire [14-1:0] node3568;
	wire [14-1:0] node3572;
	wire [14-1:0] node3573;
	wire [14-1:0] node3574;
	wire [14-1:0] node3577;
	wire [14-1:0] node3581;
	wire [14-1:0] node3582;
	wire [14-1:0] node3583;
	wire [14-1:0] node3584;
	wire [14-1:0] node3585;
	wire [14-1:0] node3588;
	wire [14-1:0] node3591;
	wire [14-1:0] node3592;
	wire [14-1:0] node3595;
	wire [14-1:0] node3598;
	wire [14-1:0] node3600;
	wire [14-1:0] node3601;
	wire [14-1:0] node3607;
	wire [14-1:0] node3608;
	wire [14-1:0] node3609;
	wire [14-1:0] node3610;
	wire [14-1:0] node3611;
	wire [14-1:0] node3613;
	wire [14-1:0] node3614;
	wire [14-1:0] node3618;
	wire [14-1:0] node3619;
	wire [14-1:0] node3621;
	wire [14-1:0] node3625;
	wire [14-1:0] node3626;
	wire [14-1:0] node3627;
	wire [14-1:0] node3629;
	wire [14-1:0] node3634;
	wire [14-1:0] node3636;
	wire [14-1:0] node3637;
	wire [14-1:0] node3638;
	wire [14-1:0] node3639;
	wire [14-1:0] node3646;
	wire [14-1:0] node3648;
	wire [14-1:0] node3649;
	wire [14-1:0] node3650;
	wire [14-1:0] node3651;
	wire [14-1:0] node3652;
	wire [14-1:0] node3653;
	wire [14-1:0] node3654;
	wire [14-1:0] node3655;
	wire [14-1:0] node3658;
	wire [14-1:0] node3661;
	wire [14-1:0] node3662;
	wire [14-1:0] node3665;
	wire [14-1:0] node3668;
	wire [14-1:0] node3669;
	wire [14-1:0] node3670;
	wire [14-1:0] node3673;
	wire [14-1:0] node3676;
	wire [14-1:0] node3677;
	wire [14-1:0] node3680;
	wire [14-1:0] node3683;
	wire [14-1:0] node3684;
	wire [14-1:0] node3685;
	wire [14-1:0] node3686;
	wire [14-1:0] node3689;
	wire [14-1:0] node3692;
	wire [14-1:0] node3693;
	wire [14-1:0] node3696;
	wire [14-1:0] node3700;
	wire [14-1:0] node3701;
	wire [14-1:0] node3702;
	wire [14-1:0] node3703;
	wire [14-1:0] node3704;
	wire [14-1:0] node3707;
	wire [14-1:0] node3710;
	wire [14-1:0] node3711;
	wire [14-1:0] node3714;
	wire [14-1:0] node3719;
	wire [14-1:0] node3721;
	wire [14-1:0] node3722;
	wire [14-1:0] node3723;
	wire [14-1:0] node3724;
	wire [14-1:0] node3725;
	wire [14-1:0] node3728;
	wire [14-1:0] node3731;
	wire [14-1:0] node3732;
	wire [14-1:0] node3736;
	wire [14-1:0] node3737;
	wire [14-1:0] node3738;
	wire [14-1:0] node3744;
	wire [14-1:0] node3746;
	wire [14-1:0] node3748;
	wire [14-1:0] node3750;
	wire [14-1:0] node3752;
	wire [14-1:0] node3754;
	wire [14-1:0] node3755;

	assign outp = (inp[8]) ? node1178 : node1;
		assign node1 = (inp[13]) ? node3 : 14'b00000000000000;
			assign node3 = (inp[10]) ? node817 : node4;
				assign node4 = (inp[0]) ? node554 : node5;
					assign node5 = (inp[6]) ? node351 : node6;
						assign node6 = (inp[4]) ? node218 : node7;
							assign node7 = (inp[7]) ? node117 : node8;
								assign node8 = (inp[12]) ? node60 : node9;
									assign node9 = (inp[2]) ? node31 : node10;
										assign node10 = (inp[5]) ? node18 : node11;
											assign node11 = (inp[1]) ? 14'b00000000000001 : node12;
												assign node12 = (inp[3]) ? 14'b00000000000001 : node13;
													assign node13 = (inp[9]) ? 14'b00000000000001 : 14'b10000000001000;
											assign node18 = (inp[9]) ? node24 : node19;
												assign node19 = (inp[3]) ? 14'b01010110110110 : node20;
													assign node20 = (inp[1]) ? 14'b01010110100110 : 14'b00000000000001;
												assign node24 = (inp[3]) ? node28 : node25;
													assign node25 = (inp[1]) ? 14'b01010110000110 : 14'b01000100000110;
													assign node28 = (inp[11]) ? 14'b01000110000110 : 14'b01010110010110;
										assign node31 = (inp[5]) ? node47 : node32;
											assign node32 = (inp[3]) ? node40 : node33;
												assign node33 = (inp[1]) ? node37 : node34;
													assign node34 = (inp[9]) ? 14'b01100100000110 : 14'b00000000000001;
													assign node37 = (inp[9]) ? 14'b01110110000110 : 14'b01110110100110;
												assign node40 = (inp[1]) ? node44 : node41;
													assign node41 = (inp[9]) ? 14'b01110110010110 : 14'b01110110110110;
													assign node44 = (inp[9]) ? 14'b01100110000110 : 14'b01100110100110;
											assign node47 = (inp[1]) ? node53 : node48;
												assign node48 = (inp[9]) ? node50 : 14'b00000000000001;
													assign node50 = (inp[3]) ? 14'b01010110010010 : 14'b01000100000010;
												assign node53 = (inp[3]) ? node57 : node54;
													assign node54 = (inp[9]) ? 14'b01010110000010 : 14'b01010110100010;
													assign node57 = (inp[9]) ? 14'b01000110000010 : 14'b01000110100010;
									assign node60 = (inp[9]) ? node86 : node61;
										assign node61 = (inp[1]) ? node71 : node62;
											assign node62 = (inp[3]) ? node64 : 14'b00000000000001;
												assign node64 = (inp[5]) ? node68 : node65;
													assign node65 = (inp[2]) ? 14'b01110110110100 : 14'b01010010110100;
													assign node68 = (inp[2]) ? 14'b01010110110000 : 14'b01010110110100;
											assign node71 = (inp[3]) ? node79 : node72;
												assign node72 = (inp[5]) ? node76 : node73;
													assign node73 = (inp[2]) ? 14'b01110110100100 : 14'b01010010100100;
													assign node76 = (inp[2]) ? 14'b01010110100000 : 14'b01010110100100;
												assign node79 = (inp[5]) ? node83 : node80;
													assign node80 = (inp[2]) ? 14'b01100110100100 : 14'b01000010100100;
													assign node83 = (inp[2]) ? 14'b01000110100000 : 14'b01000110100100;
										assign node86 = (inp[2]) ? node102 : node87;
											assign node87 = (inp[5]) ? node95 : node88;
												assign node88 = (inp[1]) ? node92 : node89;
													assign node89 = (inp[3]) ? 14'b01010010010100 : 14'b01000000000100;
													assign node92 = (inp[3]) ? 14'b01000010000100 : 14'b01010010000100;
												assign node95 = (inp[1]) ? node99 : node96;
													assign node96 = (inp[3]) ? 14'b01010110010100 : 14'b01000100000100;
													assign node99 = (inp[3]) ? 14'b01000110000100 : 14'b01010110000100;
											assign node102 = (inp[5]) ? node110 : node103;
												assign node103 = (inp[3]) ? node107 : node104;
													assign node104 = (inp[1]) ? 14'b01110110000100 : 14'b01100100000100;
													assign node107 = (inp[1]) ? 14'b01100110000100 : 14'b01110110010100;
												assign node110 = (inp[3]) ? node114 : node111;
													assign node111 = (inp[1]) ? 14'b01010110000000 : 14'b01000100000000;
													assign node114 = (inp[11]) ? 14'b01010110010000 : 14'b01000110000000;
								assign node117 = (inp[5]) ? node173 : node118;
									assign node118 = (inp[2]) ? node150 : node119;
										assign node119 = (inp[12]) ? node135 : node120;
											assign node120 = (inp[3]) ? node128 : node121;
												assign node121 = (inp[1]) ? node125 : node122;
													assign node122 = (inp[9]) ? 14'b00000000000010 : 14'b00000000000001;
													assign node125 = (inp[9]) ? 14'b00010010000010 : 14'b00010010100010;
												assign node128 = (inp[1]) ? node132 : node129;
													assign node129 = (inp[9]) ? 14'b00010010010010 : 14'b00010010110010;
													assign node132 = (inp[9]) ? 14'b00000010000010 : 14'b00000010100010;
											assign node135 = (inp[1]) ? node143 : node136;
												assign node136 = (inp[3]) ? node140 : node137;
													assign node137 = (inp[9]) ? 14'b00000000000000 : 14'b00000000000001;
													assign node140 = (inp[9]) ? 14'b00010010010000 : 14'b00010010110000;
												assign node143 = (inp[9]) ? node147 : node144;
													assign node144 = (inp[3]) ? 14'b00000010100000 : 14'b00010010100000;
													assign node147 = (inp[3]) ? 14'b00000010000000 : 14'b00010010000000;
										assign node150 = (inp[1]) ? node158 : node151;
											assign node151 = (inp[3]) ? node155 : node152;
												assign node152 = (inp[9]) ? 14'b01100000000100 : 14'b00000000000001;
												assign node155 = (inp[9]) ? 14'b01110010010110 : 14'b01110010110110;
											assign node158 = (inp[9]) ? node166 : node159;
												assign node159 = (inp[3]) ? node163 : node160;
													assign node160 = (inp[12]) ? 14'b01110010100100 : 14'b01110010100110;
													assign node163 = (inp[12]) ? 14'b01100010100100 : 14'b01100010100110;
												assign node166 = (inp[3]) ? node170 : node167;
													assign node167 = (inp[12]) ? 14'b01110010000100 : 14'b01110010000110;
													assign node170 = (inp[12]) ? 14'b01100010000100 : 14'b01100010000110;
									assign node173 = (inp[3]) ? node199 : node174;
										assign node174 = (inp[1]) ? node184 : node175;
											assign node175 = (inp[9]) ? node177 : 14'b00000000000001;
												assign node177 = (inp[2]) ? node181 : node178;
													assign node178 = (inp[12]) ? 14'b00000000000001 : 14'b01000000000110;
													assign node181 = (inp[12]) ? 14'b01000000000000 : 14'b00000000000001;
											assign node184 = (inp[9]) ? node192 : node185;
												assign node185 = (inp[2]) ? node189 : node186;
													assign node186 = (inp[12]) ? 14'b00000000000001 : 14'b01010010100110;
													assign node189 = (inp[12]) ? 14'b01010010100000 : 14'b00000000000001;
												assign node192 = (inp[11]) ? node194 : 14'b00000000000001;
													assign node194 = (inp[2]) ? 14'b00000000000001 : node195;
														assign node195 = (inp[12]) ? 14'b00000000000001 : 14'b01010010000110;
										assign node199 = (inp[2]) ? node209 : node200;
											assign node200 = (inp[12]) ? 14'b00000000000001 : node201;
												assign node201 = (inp[1]) ? node205 : node202;
													assign node202 = (inp[9]) ? 14'b01010010010110 : 14'b01010010110110;
													assign node205 = (inp[9]) ? 14'b01000010000110 : 14'b01000010100110;
											assign node209 = (inp[12]) ? node211 : 14'b00000000000001;
												assign node211 = (inp[1]) ? node215 : node212;
													assign node212 = (inp[9]) ? 14'b01010010010000 : 14'b01010010110000;
													assign node215 = (inp[9]) ? 14'b01000010000000 : 14'b01000010100000;
							assign node218 = (inp[2]) ? node318 : node219;
								assign node219 = (inp[12]) ? node277 : node220;
									assign node220 = (inp[3]) ? node246 : node221;
										assign node221 = (inp[1]) ? node231 : node222;
											assign node222 = (inp[9]) ? node224 : 14'b00000000000001;
												assign node224 = (inp[7]) ? node228 : node225;
													assign node225 = (inp[5]) ? 14'b00000100000110 : 14'b00100100000110;
													assign node228 = (inp[5]) ? 14'b00000000000110 : 14'b00100000000110;
											assign node231 = (inp[7]) ? node239 : node232;
												assign node232 = (inp[5]) ? node236 : node233;
													assign node233 = (inp[9]) ? 14'b00110110000110 : 14'b00110110100110;
													assign node236 = (inp[9]) ? 14'b00010110000110 : 14'b00010110100110;
												assign node239 = (inp[9]) ? node243 : node240;
													assign node240 = (inp[11]) ? 14'b00110010100110 : 14'b00010010100110;
													assign node243 = (inp[5]) ? 14'b00010010000110 : 14'b00110010000110;
										assign node246 = (inp[1]) ? node262 : node247;
											assign node247 = (inp[7]) ? node255 : node248;
												assign node248 = (inp[5]) ? node252 : node249;
													assign node249 = (inp[9]) ? 14'b00110110010110 : 14'b00110110110110;
													assign node252 = (inp[9]) ? 14'b00010110010110 : 14'b00010110110110;
												assign node255 = (inp[9]) ? node259 : node256;
													assign node256 = (inp[5]) ? 14'b00010010110110 : 14'b00110010110110;
													assign node259 = (inp[5]) ? 14'b00010010010110 : 14'b00110010010110;
											assign node262 = (inp[9]) ? node270 : node263;
												assign node263 = (inp[5]) ? node267 : node264;
													assign node264 = (inp[7]) ? 14'b00100010100110 : 14'b00100110100110;
													assign node267 = (inp[7]) ? 14'b00000010100110 : 14'b00000110100110;
												assign node270 = (inp[5]) ? node274 : node271;
													assign node271 = (inp[7]) ? 14'b00100010000110 : 14'b00100110000110;
													assign node274 = (inp[7]) ? 14'b00000010000110 : 14'b00000110000110;
									assign node277 = (inp[5]) ? node303 : node278;
										assign node278 = (inp[1]) ? node290 : node279;
											assign node279 = (inp[3]) ? node285 : node280;
												assign node280 = (inp[9]) ? node282 : 14'b00000000000001;
													assign node282 = (inp[7]) ? 14'b00100000000100 : 14'b00100100000100;
												assign node285 = (inp[7]) ? node287 : 14'b00110110010100;
													assign node287 = (inp[9]) ? 14'b00110010010100 : 14'b00110010110100;
											assign node290 = (inp[9]) ? node298 : node291;
												assign node291 = (inp[3]) ? node295 : node292;
													assign node292 = (inp[7]) ? 14'b00110010100100 : 14'b00110110100100;
													assign node295 = (inp[7]) ? 14'b00100010100100 : 14'b00100110100100;
												assign node298 = (inp[7]) ? 14'b00100010000100 : node299;
													assign node299 = (inp[3]) ? 14'b00100110000100 : 14'b00110110000100;
										assign node303 = (inp[7]) ? node305 : 14'b00000000000001;
											assign node305 = (inp[1]) ? node311 : node306;
												assign node306 = (inp[3]) ? 14'b00010010010100 : node307;
													assign node307 = (inp[9]) ? 14'b00000000000100 : 14'b00000000000001;
												assign node311 = (inp[9]) ? node315 : node312;
													assign node312 = (inp[3]) ? 14'b00000010100100 : 14'b00010010100100;
													assign node315 = (inp[3]) ? 14'b00000010000100 : 14'b00010010000100;
								assign node318 = (inp[7]) ? 14'b00000000000001 : node319;
									assign node319 = (inp[5]) ? node335 : node320;
										assign node320 = (inp[12]) ? node322 : 14'b00000000000001;
											assign node322 = (inp[3]) ? node328 : node323;
												assign node323 = (inp[9]) ? node325 : 14'b00000000000001;
													assign node325 = (inp[1]) ? 14'b00010110000100 : 14'b00000100000100;
												assign node328 = (inp[1]) ? node332 : node329;
													assign node329 = (inp[9]) ? 14'b00010110010100 : 14'b00010110110100;
													assign node332 = (inp[9]) ? 14'b00000110000100 : 14'b00000110100100;
										assign node335 = (inp[12]) ? 14'b00000000000001 : node336;
											assign node336 = (inp[1]) ? node342 : node337;
												assign node337 = (inp[3]) ? 14'b01010010010010 : node338;
													assign node338 = (inp[9]) ? 14'b01000000000010 : 14'b00000000000001;
												assign node342 = (inp[9]) ? node346 : node343;
													assign node343 = (inp[3]) ? 14'b01000010100010 : 14'b01010010100010;
													assign node346 = (inp[3]) ? 14'b01000010000010 : 14'b01010010000010;
						assign node351 = (inp[3]) ? node539 : node352;
							assign node352 = (inp[4]) ? node464 : node353;
								assign node353 = (inp[9]) ? node407 : node354;
									assign node354 = (inp[12]) ? node380 : node355;
										assign node355 = (inp[7]) ? node367 : node356;
											assign node356 = (inp[5]) ? node360 : node357;
												assign node357 = (inp[2]) ? 14'b01110100100110 : 14'b00000000000001;
												assign node360 = (inp[2]) ? node364 : node361;
													assign node361 = (inp[1]) ? 14'b01010100100110 : 14'b01010100110110;
													assign node364 = (inp[1]) ? 14'b01010100100010 : 14'b01010100110010;
											assign node367 = (inp[2]) ? node375 : node368;
												assign node368 = (inp[5]) ? node372 : node369;
													assign node369 = (inp[1]) ? 14'b00010000100010 : 14'b00010000110010;
													assign node372 = (inp[11]) ? 14'b01010000110110 : 14'b01010000100110;
												assign node375 = (inp[5]) ? 14'b00000000000001 : node376;
													assign node376 = (inp[1]) ? 14'b01110000100110 : 14'b01110000110110;
										assign node380 = (inp[1]) ? node394 : node381;
											assign node381 = (inp[7]) ? node389 : node382;
												assign node382 = (inp[2]) ? node386 : node383;
													assign node383 = (inp[5]) ? 14'b01010100110100 : 14'b01010000110100;
													assign node386 = (inp[5]) ? 14'b01010100110000 : 14'b01110100110100;
												assign node389 = (inp[2]) ? node391 : 14'b00010000110000;
													assign node391 = (inp[5]) ? 14'b01010000110000 : 14'b01110000110100;
											assign node394 = (inp[7]) ? node402 : node395;
												assign node395 = (inp[2]) ? node399 : node396;
													assign node396 = (inp[5]) ? 14'b01010100100100 : 14'b01010000100100;
													assign node399 = (inp[5]) ? 14'b01010100100000 : 14'b01110100100100;
												assign node402 = (inp[2]) ? node404 : 14'b00010000100000;
													assign node404 = (inp[5]) ? 14'b01010000100000 : 14'b01110000100100;
									assign node407 = (inp[7]) ? node439 : node408;
										assign node408 = (inp[1]) ? node424 : node409;
											assign node409 = (inp[12]) ? node417 : node410;
												assign node410 = (inp[2]) ? node414 : node411;
													assign node411 = (inp[5]) ? 14'b01010100010110 : 14'b00000000000001;
													assign node414 = (inp[5]) ? 14'b01010100010010 : 14'b01110100010110;
												assign node417 = (inp[2]) ? node421 : node418;
													assign node418 = (inp[5]) ? 14'b01010100010100 : 14'b01010000010100;
													assign node421 = (inp[5]) ? 14'b01010100010000 : 14'b01110100010100;
											assign node424 = (inp[12]) ? node432 : node425;
												assign node425 = (inp[5]) ? node429 : node426;
													assign node426 = (inp[2]) ? 14'b01110100000110 : 14'b00000000000001;
													assign node429 = (inp[2]) ? 14'b01010100000010 : 14'b01010100000110;
												assign node432 = (inp[5]) ? node436 : node433;
													assign node433 = (inp[2]) ? 14'b01110100000100 : 14'b01010000000100;
													assign node436 = (inp[2]) ? 14'b01010100000000 : 14'b01010100000100;
										assign node439 = (inp[5]) ? node455 : node440;
											assign node440 = (inp[2]) ? node448 : node441;
												assign node441 = (inp[12]) ? node445 : node442;
													assign node442 = (inp[1]) ? 14'b00010000000010 : 14'b00010000010010;
													assign node445 = (inp[1]) ? 14'b00010000000000 : 14'b00010000010000;
												assign node448 = (inp[12]) ? node452 : node449;
													assign node449 = (inp[1]) ? 14'b01110000000110 : 14'b01110000010110;
													assign node452 = (inp[1]) ? 14'b01110000000100 : 14'b01110000010100;
											assign node455 = (inp[2]) ? node461 : node456;
												assign node456 = (inp[12]) ? 14'b00000000000001 : node457;
													assign node457 = (inp[1]) ? 14'b01010000000110 : 14'b01010000010110;
												assign node461 = (inp[12]) ? 14'b01010000000000 : 14'b00000000000001;
								assign node464 = (inp[2]) ? node518 : node465;
									assign node465 = (inp[12]) ? node495 : node466;
										assign node466 = (inp[7]) ? node480 : node467;
											assign node467 = (inp[9]) ? node473 : node468;
												assign node468 = (inp[5]) ? 14'b00010100100110 : node469;
													assign node469 = (inp[1]) ? 14'b00110100100110 : 14'b00110100110110;
												assign node473 = (inp[1]) ? node477 : node474;
													assign node474 = (inp[5]) ? 14'b00010100010110 : 14'b00110100010110;
													assign node477 = (inp[5]) ? 14'b00010100000110 : 14'b00110100000110;
											assign node480 = (inp[5]) ? node488 : node481;
												assign node481 = (inp[1]) ? node485 : node482;
													assign node482 = (inp[9]) ? 14'b00110000010110 : 14'b00110000110110;
													assign node485 = (inp[9]) ? 14'b00110000000110 : 14'b00110000100110;
												assign node488 = (inp[1]) ? node492 : node489;
													assign node489 = (inp[9]) ? 14'b00010000010110 : 14'b00010000110110;
													assign node492 = (inp[9]) ? 14'b00010000000110 : 14'b00010000100110;
										assign node495 = (inp[5]) ? node509 : node496;
											assign node496 = (inp[1]) ? node504 : node497;
												assign node497 = (inp[7]) ? node501 : node498;
													assign node498 = (inp[9]) ? 14'b00110100010100 : 14'b00110100110100;
													assign node501 = (inp[9]) ? 14'b00110000010100 : 14'b00110000110100;
												assign node504 = (inp[7]) ? 14'b00110000000100 : node505;
													assign node505 = (inp[9]) ? 14'b00110100000100 : 14'b00110100100100;
											assign node509 = (inp[7]) ? node511 : 14'b00000000000001;
												assign node511 = (inp[9]) ? node515 : node512;
													assign node512 = (inp[1]) ? 14'b00010000100100 : 14'b00010000110100;
													assign node515 = (inp[1]) ? 14'b00010000000100 : 14'b00010000010100;
									assign node518 = (inp[7]) ? 14'b00000000000001 : node519;
										assign node519 = (inp[5]) ? node529 : node520;
											assign node520 = (inp[12]) ? node522 : 14'b00000000000001;
												assign node522 = (inp[1]) ? node526 : node523;
													assign node523 = (inp[9]) ? 14'b00010100010100 : 14'b00010100110100;
													assign node526 = (inp[9]) ? 14'b00010100000100 : 14'b00010100100100;
											assign node529 = (inp[12]) ? 14'b00000000000001 : node530;
												assign node530 = (inp[9]) ? node534 : node531;
													assign node531 = (inp[1]) ? 14'b01010000100010 : 14'b01010000110010;
													assign node534 = (inp[1]) ? 14'b01010000000010 : 14'b01010000010010;
							assign node539 = (inp[9]) ? 14'b00000000000001 : node540;
								assign node540 = (inp[4]) ? node542 : 14'b00000000000001;
									assign node542 = (inp[1]) ? 14'b00000000000001 : node543;
										assign node543 = (inp[2]) ? node545 : 14'b00000000000001;
											assign node545 = (inp[7]) ? 14'b00000000000001 : node546;
												assign node546 = (inp[5]) ? 14'b00000000000001 : node547;
													assign node547 = (inp[12]) ? 14'b00000000000001 : 14'b10000001001010;
					assign node554 = (inp[1]) ? node794 : node555;
						assign node555 = (inp[3]) ? node733 : node556;
							assign node556 = (inp[4]) ? node656 : node557;
								assign node557 = (inp[7]) ? node611 : node558;
									assign node558 = (inp[6]) ? node586 : node559;
										assign node559 = (inp[9]) ? node573 : node560;
											assign node560 = (inp[12]) ? node566 : node561;
												assign node561 = (inp[5]) ? node563 : 14'b01100110110110;
													assign node563 = (inp[2]) ? 14'b01000110110010 : 14'b01000110110110;
												assign node566 = (inp[5]) ? node570 : node567;
													assign node567 = (inp[2]) ? 14'b01100110110100 : 14'b01000010110100;
													assign node570 = (inp[2]) ? 14'b01000110110000 : 14'b01000110110100;
											assign node573 = (inp[2]) ? node581 : node574;
												assign node574 = (inp[5]) ? node578 : node575;
													assign node575 = (inp[12]) ? 14'b01000010010100 : 14'b00000000000001;
													assign node578 = (inp[12]) ? 14'b01000110010100 : 14'b01000110010110;
												assign node581 = (inp[5]) ? 14'b01000110010010 : node582;
													assign node582 = (inp[12]) ? 14'b01100110010100 : 14'b01100110010110;
										assign node586 = (inp[2]) ? node598 : node587;
											assign node587 = (inp[5]) ? node593 : node588;
												assign node588 = (inp[12]) ? node590 : 14'b00000000000001;
													assign node590 = (inp[9]) ? 14'b01000000010100 : 14'b01000000110100;
												assign node593 = (inp[12]) ? 14'b01000100110100 : node594;
													assign node594 = (inp[9]) ? 14'b01000100010110 : 14'b01000100110110;
											assign node598 = (inp[5]) ? node606 : node599;
												assign node599 = (inp[9]) ? node603 : node600;
													assign node600 = (inp[12]) ? 14'b01100100110100 : 14'b01100100110110;
													assign node603 = (inp[12]) ? 14'b01100100010100 : 14'b01100100010110;
												assign node606 = (inp[12]) ? 14'b01000100010000 : node607;
													assign node607 = (inp[9]) ? 14'b01000100010010 : 14'b01000100110010;
									assign node611 = (inp[5]) ? node639 : node612;
										assign node612 = (inp[2]) ? node626 : node613;
											assign node613 = (inp[9]) ? node619 : node614;
												assign node614 = (inp[12]) ? node616 : 14'b00000000110010;
													assign node616 = (inp[6]) ? 14'b00000000110000 : 14'b00000010110000;
												assign node619 = (inp[6]) ? node623 : node620;
													assign node620 = (inp[12]) ? 14'b00000010010000 : 14'b00000010010010;
													assign node623 = (inp[12]) ? 14'b00000000010000 : 14'b00000000010010;
											assign node626 = (inp[9]) ? node632 : node627;
												assign node627 = (inp[12]) ? 14'b01100010110100 : node628;
													assign node628 = (inp[6]) ? 14'b01100000110110 : 14'b01100010110110;
												assign node632 = (inp[6]) ? node636 : node633;
													assign node633 = (inp[12]) ? 14'b01100010010100 : 14'b01100010010110;
													assign node636 = (inp[12]) ? 14'b01100000010100 : 14'b01100000010110;
										assign node639 = (inp[2]) ? node647 : node640;
											assign node640 = (inp[12]) ? 14'b00000000000001 : node641;
												assign node641 = (inp[9]) ? node643 : 14'b01000000110110;
													assign node643 = (inp[6]) ? 14'b01000000010110 : 14'b01000010010110;
											assign node647 = (inp[12]) ? node649 : 14'b00000000000001;
												assign node649 = (inp[9]) ? node653 : node650;
													assign node650 = (inp[6]) ? 14'b01000000110000 : 14'b01000010110000;
													assign node653 = (inp[6]) ? 14'b01000000010000 : 14'b01000010010000;
								assign node656 = (inp[2]) ? node712 : node657;
									assign node657 = (inp[12]) ? node687 : node658;
										assign node658 = (inp[5]) ? node674 : node659;
											assign node659 = (inp[7]) ? node667 : node660;
												assign node660 = (inp[6]) ? node664 : node661;
													assign node661 = (inp[9]) ? 14'b00100110010110 : 14'b00100110110110;
													assign node664 = (inp[9]) ? 14'b00100100010110 : 14'b00100100110110;
												assign node667 = (inp[9]) ? node671 : node668;
													assign node668 = (inp[6]) ? 14'b00100000110110 : 14'b00100010110110;
													assign node671 = (inp[6]) ? 14'b00100000010110 : 14'b00100010010110;
											assign node674 = (inp[7]) ? node680 : node675;
												assign node675 = (inp[6]) ? 14'b00000100110110 : node676;
													assign node676 = (inp[9]) ? 14'b00000110010110 : 14'b00000110110110;
												assign node680 = (inp[6]) ? node684 : node681;
													assign node681 = (inp[9]) ? 14'b00000010010110 : 14'b00000010110110;
													assign node684 = (inp[9]) ? 14'b00000000010110 : 14'b00000000110110;
										assign node687 = (inp[5]) ? node703 : node688;
											assign node688 = (inp[6]) ? node696 : node689;
												assign node689 = (inp[7]) ? node693 : node690;
													assign node690 = (inp[9]) ? 14'b00100110010100 : 14'b00100110110100;
													assign node693 = (inp[9]) ? 14'b00100010010100 : 14'b00100010110100;
												assign node696 = (inp[9]) ? node700 : node697;
													assign node697 = (inp[7]) ? 14'b00100000110100 : 14'b00100100110100;
													assign node700 = (inp[7]) ? 14'b00100000010100 : 14'b00100100010100;
											assign node703 = (inp[7]) ? node705 : 14'b00000000000001;
												assign node705 = (inp[9]) ? node709 : node706;
													assign node706 = (inp[6]) ? 14'b00000000110100 : 14'b00000010110100;
													assign node709 = (inp[11]) ? 14'b00000000010100 : 14'b00000010010100;
									assign node712 = (inp[7]) ? 14'b00000000000001 : node713;
										assign node713 = (inp[5]) ? node723 : node714;
											assign node714 = (inp[12]) ? node716 : 14'b00000000000001;
												assign node716 = (inp[6]) ? node720 : node717;
													assign node717 = (inp[9]) ? 14'b00000110010100 : 14'b00000110110100;
													assign node720 = (inp[9]) ? 14'b00000100010100 : 14'b00000100110100;
											assign node723 = (inp[12]) ? 14'b00000000000001 : node724;
												assign node724 = (inp[9]) ? node728 : node725;
													assign node725 = (inp[6]) ? 14'b01000000110010 : 14'b01000010110010;
													assign node728 = (inp[6]) ? 14'b01000000010010 : 14'b01000010010010;
							assign node733 = (inp[6]) ? node735 : 14'b00000000000001;
								assign node735 = (inp[9]) ? 14'b00000000000001 : node736;
									assign node736 = (inp[4]) ? node768 : node737;
										assign node737 = (inp[7]) ? node753 : node738;
											assign node738 = (inp[2]) ? node746 : node739;
												assign node739 = (inp[5]) ? node743 : node740;
													assign node740 = (inp[12]) ? 14'b01000000100100 : 14'b00000000000001;
													assign node743 = (inp[12]) ? 14'b01000100100100 : 14'b01000100100110;
												assign node746 = (inp[5]) ? node750 : node747;
													assign node747 = (inp[12]) ? 14'b01100100100100 : 14'b01100100100110;
													assign node750 = (inp[12]) ? 14'b01000100100000 : 14'b01000100100010;
											assign node753 = (inp[5]) ? node761 : node754;
												assign node754 = (inp[2]) ? node758 : node755;
													assign node755 = (inp[12]) ? 14'b00000000100000 : 14'b00000000100010;
													assign node758 = (inp[12]) ? 14'b01100000100100 : 14'b01100000100110;
												assign node761 = (inp[2]) ? node765 : node762;
													assign node762 = (inp[12]) ? 14'b00000000000001 : 14'b01000000100110;
													assign node765 = (inp[12]) ? 14'b01000000100000 : 14'b00000000000001;
										assign node768 = (inp[2]) ? node784 : node769;
											assign node769 = (inp[5]) ? node777 : node770;
												assign node770 = (inp[12]) ? node774 : node771;
													assign node771 = (inp[7]) ? 14'b00100000100110 : 14'b00100100100110;
													assign node774 = (inp[7]) ? 14'b00100000100100 : 14'b00100100100100;
												assign node777 = (inp[12]) ? node781 : node778;
													assign node778 = (inp[7]) ? 14'b00000000100110 : 14'b00000100100110;
													assign node781 = (inp[7]) ? 14'b00000000100100 : 14'b00000000000001;
											assign node784 = (inp[7]) ? 14'b00000000000001 : node785;
												assign node785 = (inp[5]) ? node789 : node786;
													assign node786 = (inp[12]) ? 14'b00000100100100 : 14'b00000000000001;
													assign node789 = (inp[12]) ? 14'b00000000000001 : 14'b01000000100010;
						assign node794 = (inp[6]) ? 14'b00000000000001 : node795;
							assign node795 = (inp[5]) ? 14'b00000000000001 : node796;
								assign node796 = (inp[12]) ? 14'b00000000000001 : node797;
									assign node797 = (inp[7]) ? 14'b00000000000001 : node798;
										assign node798 = (inp[3]) ? node806 : node799;
											assign node799 = (inp[2]) ? node801 : 14'b00000000000001;
												assign node801 = (inp[9]) ? 14'b00000000000001 : node802;
													assign node802 = (inp[11]) ? 14'b10000001000010 : 14'b00000000000001;
											assign node806 = (inp[2]) ? 14'b00000000000001 : node807;
												assign node807 = (inp[4]) ? 14'b00000000000001 : node808;
													assign node808 = (inp[9]) ? 14'b10000000000010 : 14'b00000000000001;
				assign node817 = (inp[5]) ? 14'b00000000000001 : node818;
					assign node818 = (inp[2]) ? node1068 : node819;
						assign node819 = (inp[3]) ? node987 : node820;
							assign node820 = (inp[1]) ? node926 : node821;
								assign node821 = (inp[0]) ? node869 : node822;
									assign node822 = (inp[6]) ? node840 : node823;
										assign node823 = (inp[9]) ? node825 : 14'b00000000000001;
											assign node825 = (inp[4]) ? node833 : node826;
												assign node826 = (inp[12]) ? node830 : node827;
													assign node827 = (inp[7]) ? 14'b01100000000010 : 14'b01100100000010;
													assign node830 = (inp[7]) ? 14'b01100000000000 : 14'b01100100000000;
												assign node833 = (inp[12]) ? node837 : node834;
													assign node834 = (inp[11]) ? 14'b00100000000010 : 14'b00100100000010;
													assign node837 = (inp[7]) ? 14'b00100000000000 : 14'b00100100000000;
										assign node840 = (inp[7]) ? node854 : node841;
											assign node841 = (inp[4]) ? node847 : node842;
												assign node842 = (inp[9]) ? 14'b01110100010000 : node843;
													assign node843 = (inp[12]) ? 14'b01110100110000 : 14'b01110100110010;
												assign node847 = (inp[12]) ? node851 : node848;
													assign node848 = (inp[9]) ? 14'b00110100010010 : 14'b00110100110010;
													assign node851 = (inp[9]) ? 14'b00110100010000 : 14'b00110100110000;
											assign node854 = (inp[4]) ? node862 : node855;
												assign node855 = (inp[12]) ? node859 : node856;
													assign node856 = (inp[9]) ? 14'b01110000010010 : 14'b01110000110010;
													assign node859 = (inp[9]) ? 14'b01110000010000 : 14'b01110000110000;
												assign node862 = (inp[12]) ? node866 : node863;
													assign node863 = (inp[11]) ? 14'b00110000110010 : 14'b00110000010010;
													assign node866 = (inp[9]) ? 14'b00110000010000 : 14'b00110000110000;
									assign node869 = (inp[6]) ? node897 : node870;
										assign node870 = (inp[7]) ? node882 : node871;
											assign node871 = (inp[4]) ? node879 : node872;
												assign node872 = (inp[9]) ? node876 : node873;
													assign node873 = (inp[12]) ? 14'b01100110110000 : 14'b01100110110010;
													assign node876 = (inp[12]) ? 14'b01100110010000 : 14'b01100110010010;
												assign node879 = (inp[12]) ? 14'b00100110110000 : 14'b00100110110010;
											assign node882 = (inp[9]) ? node890 : node883;
												assign node883 = (inp[12]) ? node887 : node884;
													assign node884 = (inp[4]) ? 14'b00100010110010 : 14'b01100010110010;
													assign node887 = (inp[4]) ? 14'b00100010110000 : 14'b01100010110000;
												assign node890 = (inp[4]) ? node894 : node891;
													assign node891 = (inp[12]) ? 14'b01100010010000 : 14'b01100010010010;
													assign node894 = (inp[12]) ? 14'b00100010010000 : 14'b00100010010010;
										assign node897 = (inp[4]) ? node911 : node898;
											assign node898 = (inp[12]) ? node904 : node899;
												assign node899 = (inp[7]) ? node901 : 14'b01100100010010;
													assign node901 = (inp[9]) ? 14'b01100000010010 : 14'b01100000110010;
												assign node904 = (inp[7]) ? node908 : node905;
													assign node905 = (inp[9]) ? 14'b01100100010000 : 14'b01100100110000;
													assign node908 = (inp[9]) ? 14'b01100000010000 : 14'b01100000110000;
											assign node911 = (inp[12]) ? node919 : node912;
												assign node912 = (inp[9]) ? node916 : node913;
													assign node913 = (inp[7]) ? 14'b00100000110010 : 14'b00100100110010;
													assign node916 = (inp[7]) ? 14'b00100000010010 : 14'b00100100010010;
												assign node919 = (inp[7]) ? node923 : node920;
													assign node920 = (inp[9]) ? 14'b00100100010000 : 14'b00100100110000;
													assign node923 = (inp[9]) ? 14'b00100000010000 : 14'b00100000110000;
								assign node926 = (inp[0]) ? 14'b00000000000001 : node927;
									assign node927 = (inp[9]) ? node957 : node928;
										assign node928 = (inp[6]) ? node942 : node929;
											assign node929 = (inp[12]) ? node935 : node930;
												assign node930 = (inp[7]) ? node932 : 14'b01110110100010;
													assign node932 = (inp[4]) ? 14'b00110010100010 : 14'b01110010100010;
												assign node935 = (inp[4]) ? node939 : node936;
													assign node936 = (inp[7]) ? 14'b01110010100000 : 14'b01110110100000;
													assign node939 = (inp[7]) ? 14'b00110010100000 : 14'b00110110100000;
											assign node942 = (inp[12]) ? node950 : node943;
												assign node943 = (inp[4]) ? node947 : node944;
													assign node944 = (inp[7]) ? 14'b01110000100010 : 14'b01110100100010;
													assign node947 = (inp[7]) ? 14'b00110000100010 : 14'b00110100100010;
												assign node950 = (inp[7]) ? node954 : node951;
													assign node951 = (inp[4]) ? 14'b00110100100000 : 14'b01110100100000;
													assign node954 = (inp[4]) ? 14'b00110000100000 : 14'b01110000100000;
										assign node957 = (inp[6]) ? node973 : node958;
											assign node958 = (inp[4]) ? node966 : node959;
												assign node959 = (inp[7]) ? node963 : node960;
													assign node960 = (inp[12]) ? 14'b01110110000000 : 14'b01110110000010;
													assign node963 = (inp[12]) ? 14'b01110010000000 : 14'b01110010000010;
												assign node966 = (inp[7]) ? node970 : node967;
													assign node967 = (inp[12]) ? 14'b00110110000000 : 14'b00110110000010;
													assign node970 = (inp[12]) ? 14'b00110010000000 : 14'b00110010000010;
											assign node973 = (inp[4]) ? node979 : node974;
												assign node974 = (inp[7]) ? 14'b01110000000000 : node975;
													assign node975 = (inp[12]) ? 14'b01110100000000 : 14'b01110100000010;
												assign node979 = (inp[12]) ? node983 : node980;
													assign node980 = (inp[7]) ? 14'b00110000000010 : 14'b00110100000010;
													assign node983 = (inp[7]) ? 14'b00110000000000 : 14'b00110100000000;
							assign node987 = (inp[6]) ? node1047 : node988;
								assign node988 = (inp[0]) ? 14'b00000000000001 : node989;
									assign node989 = (inp[1]) ? node1017 : node990;
										assign node990 = (inp[12]) ? node1004 : node991;
											assign node991 = (inp[4]) ? node999 : node992;
												assign node992 = (inp[7]) ? node996 : node993;
													assign node993 = (inp[11]) ? 14'b01110110010010 : 14'b01110110110010;
													assign node996 = (inp[9]) ? 14'b01110010010010 : 14'b01110010110010;
												assign node999 = (inp[7]) ? 14'b00110010110010 : node1000;
													assign node1000 = (inp[9]) ? 14'b00110110010010 : 14'b00110110110010;
											assign node1004 = (inp[7]) ? node1010 : node1005;
												assign node1005 = (inp[9]) ? node1007 : 14'b01110110110000;
													assign node1007 = (inp[4]) ? 14'b00110110010000 : 14'b01110110010000;
												assign node1010 = (inp[9]) ? node1014 : node1011;
													assign node1011 = (inp[4]) ? 14'b00110010110000 : 14'b01110010110000;
													assign node1014 = (inp[11]) ? 14'b01110010010000 : 14'b00110010010000;
										assign node1017 = (inp[9]) ? node1033 : node1018;
											assign node1018 = (inp[12]) ? node1026 : node1019;
												assign node1019 = (inp[4]) ? node1023 : node1020;
													assign node1020 = (inp[7]) ? 14'b01100010100010 : 14'b01100110100010;
													assign node1023 = (inp[7]) ? 14'b00100010100010 : 14'b00100110100010;
												assign node1026 = (inp[4]) ? node1030 : node1027;
													assign node1027 = (inp[7]) ? 14'b01100010100000 : 14'b01100110100000;
													assign node1030 = (inp[7]) ? 14'b00100010100000 : 14'b00100110100000;
											assign node1033 = (inp[4]) ? node1039 : node1034;
												assign node1034 = (inp[12]) ? node1036 : 14'b01100110000010;
													assign node1036 = (inp[11]) ? 14'b01100110000000 : 14'b01100010000000;
												assign node1039 = (inp[7]) ? node1043 : node1040;
													assign node1040 = (inp[12]) ? 14'b00100110000000 : 14'b00100110000010;
													assign node1043 = (inp[12]) ? 14'b00100010000000 : 14'b00100010000010;
								assign node1047 = (inp[1]) ? 14'b00000000000001 : node1048;
									assign node1048 = (inp[0]) ? node1050 : 14'b00000000000001;
										assign node1050 = (inp[9]) ? 14'b00000000000001 : node1051;
											assign node1051 = (inp[4]) ? node1059 : node1052;
												assign node1052 = (inp[12]) ? node1056 : node1053;
													assign node1053 = (inp[7]) ? 14'b01100000100010 : 14'b01100100100010;
													assign node1056 = (inp[7]) ? 14'b01100000100000 : 14'b01100100100000;
												assign node1059 = (inp[12]) ? node1063 : node1060;
													assign node1060 = (inp[7]) ? 14'b00100000100010 : 14'b00100100100010;
													assign node1063 = (inp[7]) ? 14'b00100000100000 : 14'b00100100100000;
						assign node1068 = (inp[7]) ? node1164 : node1069;
							assign node1069 = (inp[4]) ? node1091 : node1070;
								assign node1070 = (inp[9]) ? 14'b00000000000001 : node1071;
									assign node1071 = (inp[12]) ? 14'b00000000000001 : node1072;
										assign node1072 = (inp[1]) ? node1082 : node1073;
											assign node1073 = (inp[3]) ? node1075 : 14'b00000000000001;
												assign node1075 = (inp[6]) ? node1079 : node1076;
													assign node1076 = (inp[0]) ? 14'b10000001000000 : 14'b00000000000001;
													assign node1079 = (inp[0]) ? 14'b00000000000001 : 14'b10000001001000;
											assign node1082 = (inp[3]) ? 14'b00000000000001 : node1083;
												assign node1083 = (inp[0]) ? node1085 : 14'b00000000000001;
													assign node1085 = (inp[6]) ? 14'b00000000000001 : 14'b10000000001010;
								assign node1091 = (inp[0]) ? node1139 : node1092;
									assign node1092 = (inp[6]) ? node1122 : node1093;
										assign node1093 = (inp[3]) ? node1107 : node1094;
											assign node1094 = (inp[1]) ? node1100 : node1095;
												assign node1095 = (inp[9]) ? node1097 : 14'b00000000000001;
													assign node1097 = (inp[12]) ? 14'b00000100000000 : 14'b00000100000010;
												assign node1100 = (inp[12]) ? node1104 : node1101;
													assign node1101 = (inp[9]) ? 14'b00010110000010 : 14'b00010110100010;
													assign node1104 = (inp[9]) ? 14'b00010110000000 : 14'b00010110100000;
											assign node1107 = (inp[1]) ? node1115 : node1108;
												assign node1108 = (inp[12]) ? node1112 : node1109;
													assign node1109 = (inp[9]) ? 14'b00010110010010 : 14'b00010110110010;
													assign node1112 = (inp[9]) ? 14'b00010110010000 : 14'b00010110110000;
												assign node1115 = (inp[9]) ? node1119 : node1116;
													assign node1116 = (inp[12]) ? 14'b00000110100000 : 14'b00000110100010;
													assign node1119 = (inp[12]) ? 14'b00000110000000 : 14'b00000110000010;
										assign node1122 = (inp[3]) ? 14'b00000000000001 : node1123;
											assign node1123 = (inp[12]) ? node1131 : node1124;
												assign node1124 = (inp[1]) ? node1128 : node1125;
													assign node1125 = (inp[9]) ? 14'b00010100010010 : 14'b00010100110010;
													assign node1128 = (inp[9]) ? 14'b00010100000010 : 14'b00010100100010;
												assign node1131 = (inp[9]) ? node1135 : node1132;
													assign node1132 = (inp[1]) ? 14'b00010100100000 : 14'b00010100110000;
													assign node1135 = (inp[1]) ? 14'b00010100000000 : 14'b00010100010000;
									assign node1139 = (inp[1]) ? 14'b00000000000001 : node1140;
										assign node1140 = (inp[3]) ? node1156 : node1141;
											assign node1141 = (inp[12]) ? node1149 : node1142;
												assign node1142 = (inp[6]) ? node1146 : node1143;
													assign node1143 = (inp[9]) ? 14'b00000110010010 : 14'b00000110110010;
													assign node1146 = (inp[9]) ? 14'b00000100010010 : 14'b00000100110010;
												assign node1149 = (inp[9]) ? node1153 : node1150;
													assign node1150 = (inp[6]) ? 14'b00000100110000 : 14'b00000110110000;
													assign node1153 = (inp[6]) ? 14'b00000100010000 : 14'b00000110010000;
											assign node1156 = (inp[9]) ? 14'b00000000000001 : node1157;
												assign node1157 = (inp[6]) ? node1159 : 14'b00000000000001;
													assign node1159 = (inp[12]) ? 14'b00000100100000 : 14'b00000100100010;
							assign node1164 = (inp[11]) ? 14'b00000000000001 : node1165;
								assign node1165 = (inp[4]) ? node1167 : 14'b00000000000001;
									assign node1167 = (inp[12]) ? 14'b00000000000001 : node1168;
										assign node1168 = (inp[9]) ? 14'b00000000000001 : node1169;
											assign node1169 = (inp[6]) ? node1171 : 14'b00000000000001;
												assign node1171 = (inp[0]) ? 14'b00000000000001 : 14'b10000000000000;
		assign node1178 = (inp[0]) ? node2886 : node1179;
			assign node1179 = (inp[3]) ? node2273 : node1180;
				assign node1180 = (inp[12]) ? node1784 : node1181;
					assign node1181 = (inp[2]) ? node1519 : node1182;
						assign node1182 = (inp[13]) ? node1408 : node1183;
							assign node1183 = (inp[11]) ? node1359 : node1184;
								assign node1184 = (inp[4]) ? node1268 : node1185;
									assign node1185 = (inp[10]) ? node1221 : node1186;
										assign node1186 = (inp[5]) ? node1194 : node1187;
											assign node1187 = (inp[7]) ? 14'b00000000000001 : node1188;
												assign node1188 = (inp[6]) ? 14'b00000000000001 : node1189;
													assign node1189 = (inp[9]) ? 14'b00000000000001 : 14'b10000000001000;
											assign node1194 = (inp[7]) ? node1206 : node1195;
												assign node1195 = (inp[6]) ? node1203 : node1196;
													assign node1196 = (inp[1]) ? node1200 : node1197;
														assign node1197 = (inp[9]) ? 14'b00100100000010 : 14'b00000000000001;
														assign node1200 = (inp[9]) ? 14'b00100000000010 : 14'b00110010000010;
													assign node1203 = (inp[1]) ? 14'b00110000010010 : 14'b00110100110010;
												assign node1206 = (inp[1]) ? node1214 : node1207;
													assign node1207 = (inp[6]) ? node1211 : node1208;
														assign node1208 = (inp[9]) ? 14'b00100110010010 : 14'b00100110110010;
														assign node1211 = (inp[9]) ? 14'b00100100010010 : 14'b00100100110010;
													assign node1214 = (inp[9]) ? node1218 : node1215;
														assign node1215 = (inp[6]) ? 14'b00100000110010 : 14'b00100010110010;
														assign node1218 = (inp[6]) ? 14'b00100000010010 : 14'b00100010010010;
										assign node1221 = (inp[1]) ? node1243 : node1222;
											assign node1222 = (inp[7]) ? node1232 : node1223;
												assign node1223 = (inp[6]) ? node1229 : node1224;
													assign node1224 = (inp[9]) ? node1226 : 14'b00000000000001;
														assign node1226 = (inp[5]) ? 14'b01100100000010 : 14'b01101100000010;
													assign node1229 = (inp[9]) ? 14'b01110100010010 : 14'b01110100110010;
												assign node1232 = (inp[6]) ? node1238 : node1233;
													assign node1233 = (inp[5]) ? node1235 : 14'b01101110010010;
														assign node1235 = (inp[9]) ? 14'b01100110010010 : 14'b01100110110010;
													assign node1238 = (inp[5]) ? 14'b01100100010010 : node1239;
														assign node1239 = (inp[9]) ? 14'b01101100010010 : 14'b01101100110010;
											assign node1243 = (inp[5]) ? node1255 : node1244;
												assign node1244 = (inp[9]) ? node1250 : node1245;
													assign node1245 = (inp[6]) ? node1247 : 14'b01101010110010;
														assign node1247 = (inp[7]) ? 14'b01101000110010 : 14'b01111000110010;
													assign node1250 = (inp[6]) ? node1252 : 14'b01101000000010;
														assign node1252 = (inp[7]) ? 14'b01101000010010 : 14'b01111000010010;
												assign node1255 = (inp[6]) ? node1261 : node1256;
													assign node1256 = (inp[7]) ? node1258 : 14'b01110010000010;
														assign node1258 = (inp[9]) ? 14'b01100010010010 : 14'b01100010110010;
													assign node1261 = (inp[9]) ? node1265 : node1262;
														assign node1262 = (inp[7]) ? 14'b01100000110010 : 14'b01110000110010;
														assign node1265 = (inp[7]) ? 14'b01100000010010 : 14'b01110000010010;
									assign node1268 = (inp[10]) ? node1316 : node1269;
										assign node1269 = (inp[6]) ? node1291 : node1270;
											assign node1270 = (inp[7]) ? node1284 : node1271;
												assign node1271 = (inp[1]) ? node1277 : node1272;
													assign node1272 = (inp[9]) ? node1274 : 14'b00000000000001;
														assign node1274 = (inp[5]) ? 14'b01100100000110 : 14'b01101100000110;
													assign node1277 = (inp[9]) ? node1281 : node1278;
														assign node1278 = (inp[5]) ? 14'b01110010000110 : 14'b01111010000110;
														assign node1281 = (inp[5]) ? 14'b01100000000110 : 14'b01101000000110;
												assign node1284 = (inp[9]) ? 14'b01101010010110 : node1285;
													assign node1285 = (inp[5]) ? 14'b01100010110110 : node1286;
														assign node1286 = (inp[1]) ? 14'b01101010110110 : 14'b01101110110110;
											assign node1291 = (inp[1]) ? node1305 : node1292;
												assign node1292 = (inp[5]) ? node1300 : node1293;
													assign node1293 = (inp[7]) ? node1297 : node1294;
														assign node1294 = (inp[9]) ? 14'b01111100010110 : 14'b01111100110110;
														assign node1297 = (inp[9]) ? 14'b01101100010110 : 14'b01101100110110;
													assign node1300 = (inp[7]) ? 14'b01100100110110 : node1301;
														assign node1301 = (inp[9]) ? 14'b01110100010110 : 14'b01110100110110;
												assign node1305 = (inp[9]) ? node1311 : node1306;
													assign node1306 = (inp[5]) ? node1308 : 14'b01101000110110;
														assign node1308 = (inp[7]) ? 14'b01100000110110 : 14'b01110000110110;
													assign node1311 = (inp[7]) ? node1313 : 14'b01111000010110;
														assign node1313 = (inp[5]) ? 14'b01100000010110 : 14'b01101000010110;
										assign node1316 = (inp[6]) ? node1336 : node1317;
											assign node1317 = (inp[7]) ? node1327 : node1318;
												assign node1318 = (inp[9]) ? node1320 : 14'b01110010000000;
													assign node1320 = (inp[5]) ? node1324 : node1321;
														assign node1321 = (inp[1]) ? 14'b01101000000000 : 14'b01101100000000;
														assign node1324 = (inp[1]) ? 14'b01100000000000 : 14'b01100100000000;
												assign node1327 = (inp[9]) ? node1331 : node1328;
													assign node1328 = (inp[1]) ? 14'b01101010110000 : 14'b01101110110000;
													assign node1331 = (inp[5]) ? node1333 : 14'b01101110010000;
														assign node1333 = (inp[1]) ? 14'b01100010010000 : 14'b01100110010000;
											assign node1336 = (inp[9]) ? node1350 : node1337;
												assign node1337 = (inp[7]) ? node1345 : node1338;
													assign node1338 = (inp[5]) ? node1342 : node1339;
														assign node1339 = (inp[1]) ? 14'b01111000110000 : 14'b01111100110000;
														assign node1342 = (inp[1]) ? 14'b01110000110000 : 14'b01110100110000;
													assign node1345 = (inp[5]) ? node1347 : 14'b01101100110000;
														assign node1347 = (inp[1]) ? 14'b01100000110000 : 14'b01100100110000;
												assign node1350 = (inp[1]) ? node1354 : node1351;
													assign node1351 = (inp[5]) ? 14'b01110100010000 : 14'b01111100010000;
													assign node1354 = (inp[7]) ? 14'b01101000010000 : node1355;
														assign node1355 = (inp[5]) ? 14'b01110000010000 : 14'b01111000010000;
								assign node1359 = (inp[10]) ? 14'b00000000000001 : node1360;
									assign node1360 = (inp[4]) ? 14'b00000000000001 : node1361;
										assign node1361 = (inp[1]) ? node1381 : node1362;
											assign node1362 = (inp[5]) ? node1370 : node1363;
												assign node1363 = (inp[6]) ? node1367 : node1364;
													assign node1364 = (inp[9]) ? 14'b01101100000100 : 14'b00000000000001;
													assign node1367 = (inp[9]) ? 14'b01111100010100 : 14'b01101100110100;
												assign node1370 = (inp[9]) ? node1376 : node1371;
													assign node1371 = (inp[6]) ? node1373 : 14'b01100110110100;
														assign node1373 = (inp[7]) ? 14'b01100100110100 : 14'b01110100110100;
													assign node1376 = (inp[7]) ? node1378 : 14'b01100100000100;
														assign node1378 = (inp[6]) ? 14'b01100100010100 : 14'b01100110010100;
											assign node1381 = (inp[5]) ? node1393 : node1382;
												assign node1382 = (inp[7]) ? node1388 : node1383;
													assign node1383 = (inp[6]) ? node1385 : 14'b01111010000100;
														assign node1385 = (inp[9]) ? 14'b01111000010100 : 14'b01111000110100;
													assign node1388 = (inp[6]) ? 14'b01101000010100 : node1389;
														assign node1389 = (inp[9]) ? 14'b01101010010100 : 14'b01101010110100;
												assign node1393 = (inp[6]) ? node1401 : node1394;
													assign node1394 = (inp[7]) ? node1398 : node1395;
														assign node1395 = (inp[9]) ? 14'b01100000000100 : 14'b01110010000100;
														assign node1398 = (inp[9]) ? 14'b01100010010100 : 14'b01100010110100;
													assign node1401 = (inp[7]) ? node1403 : 14'b01110000110100;
														assign node1403 = (inp[9]) ? 14'b01100000010100 : 14'b01100000110100;
							assign node1408 = (inp[6]) ? node1462 : node1409;
								assign node1409 = (inp[1]) ? node1433 : node1410;
									assign node1410 = (inp[9]) ? node1418 : node1411;
										assign node1411 = (inp[7]) ? 14'b00000000000001 : node1412;
											assign node1412 = (inp[4]) ? 14'b00000000000001 : node1413;
												assign node1413 = (inp[5]) ? 14'b00000000000001 : 14'b10000000001000;
										assign node1418 = (inp[4]) ? node1426 : node1419;
											assign node1419 = (inp[5]) ? node1423 : node1420;
												assign node1420 = (inp[7]) ? 14'b00000000000000 : 14'b00000000000001;
												assign node1423 = (inp[7]) ? 14'b01100000000000 : 14'b01100100000000;
											assign node1426 = (inp[5]) ? node1430 : node1427;
												assign node1427 = (inp[7]) ? 14'b00100000000100 : 14'b00100100000100;
												assign node1430 = (inp[7]) ? 14'b00100000000000 : 14'b00100100000000;
									assign node1433 = (inp[4]) ? node1447 : node1434;
										assign node1434 = (inp[5]) ? node1440 : node1435;
											assign node1435 = (inp[7]) ? node1437 : 14'b00000000000001;
												assign node1437 = (inp[9]) ? 14'b00010010000000 : 14'b00010010100000;
											assign node1440 = (inp[9]) ? node1444 : node1441;
												assign node1441 = (inp[7]) ? 14'b01110010100000 : 14'b01110110100000;
												assign node1444 = (inp[7]) ? 14'b01110010000000 : 14'b01110110000000;
										assign node1447 = (inp[7]) ? node1455 : node1448;
											assign node1448 = (inp[9]) ? node1452 : node1449;
												assign node1449 = (inp[5]) ? 14'b00110110100000 : 14'b00110110100100;
												assign node1452 = (inp[5]) ? 14'b00110110000000 : 14'b00110110000100;
											assign node1455 = (inp[5]) ? node1459 : node1456;
												assign node1456 = (inp[9]) ? 14'b00110010000100 : 14'b00110010100100;
												assign node1459 = (inp[9]) ? 14'b00110010000000 : 14'b00110010100000;
								assign node1462 = (inp[4]) ? node1488 : node1463;
									assign node1463 = (inp[5]) ? node1473 : node1464;
										assign node1464 = (inp[7]) ? node1466 : 14'b00000000000001;
											assign node1466 = (inp[1]) ? node1470 : node1467;
												assign node1467 = (inp[9]) ? 14'b00010000010000 : 14'b00010000110000;
												assign node1470 = (inp[9]) ? 14'b00010000000000 : 14'b00010000100000;
										assign node1473 = (inp[1]) ? node1481 : node1474;
											assign node1474 = (inp[9]) ? node1478 : node1475;
												assign node1475 = (inp[7]) ? 14'b01110000110000 : 14'b01110100110000;
												assign node1478 = (inp[7]) ? 14'b01110000010000 : 14'b01110100010000;
											assign node1481 = (inp[7]) ? node1485 : node1482;
												assign node1482 = (inp[9]) ? 14'b01110100000000 : 14'b01110100100000;
												assign node1485 = (inp[9]) ? 14'b01110000000000 : 14'b01110000100000;
									assign node1488 = (inp[9]) ? node1504 : node1489;
										assign node1489 = (inp[7]) ? node1497 : node1490;
											assign node1490 = (inp[1]) ? node1494 : node1491;
												assign node1491 = (inp[5]) ? 14'b00110100110000 : 14'b00110100110100;
												assign node1494 = (inp[5]) ? 14'b00110100100000 : 14'b00110100100100;
											assign node1497 = (inp[1]) ? node1501 : node1498;
												assign node1498 = (inp[5]) ? 14'b00110000110000 : 14'b00110000110100;
												assign node1501 = (inp[5]) ? 14'b00110000100000 : 14'b00110000100100;
										assign node1504 = (inp[5]) ? node1512 : node1505;
											assign node1505 = (inp[1]) ? node1509 : node1506;
												assign node1506 = (inp[7]) ? 14'b00110000010100 : 14'b00110100010100;
												assign node1509 = (inp[7]) ? 14'b00110000000100 : 14'b00110100000100;
											assign node1512 = (inp[1]) ? node1516 : node1513;
												assign node1513 = (inp[7]) ? 14'b00110000010000 : 14'b00110100010000;
												assign node1516 = (inp[7]) ? 14'b00110000000000 : 14'b00110100000000;
						assign node1519 = (inp[4]) ? node1681 : node1520;
							assign node1520 = (inp[5]) ? node1624 : node1521;
								assign node1521 = (inp[13]) ? node1595 : node1522;
									assign node1522 = (inp[11]) ? node1574 : node1523;
										assign node1523 = (inp[10]) ? node1547 : node1524;
											assign node1524 = (inp[6]) ? node1534 : node1525;
												assign node1525 = (inp[7]) ? node1527 : 14'b00000000000001;
													assign node1527 = (inp[1]) ? node1531 : node1528;
														assign node1528 = (inp[9]) ? 14'b00001110010000 : 14'b00001110110000;
														assign node1531 = (inp[9]) ? 14'b00001010010000 : 14'b00001010110000;
												assign node1534 = (inp[1]) ? node1542 : node1535;
													assign node1535 = (inp[7]) ? node1539 : node1536;
														assign node1536 = (inp[9]) ? 14'b00011100010000 : 14'b00011100110000;
														assign node1539 = (inp[9]) ? 14'b00001100010000 : 14'b00001100110000;
													assign node1542 = (inp[7]) ? 14'b00001000010000 : node1543;
														assign node1543 = (inp[9]) ? 14'b00011000010000 : 14'b00011000110000;
											assign node1547 = (inp[1]) ? node1561 : node1548;
												assign node1548 = (inp[9]) ? node1554 : node1549;
													assign node1549 = (inp[7]) ? node1551 : 14'b00111100110010;
														assign node1551 = (inp[6]) ? 14'b00101100110010 : 14'b00101110110010;
													assign node1554 = (inp[7]) ? node1558 : node1555;
														assign node1555 = (inp[6]) ? 14'b00111100010010 : 14'b00101100000010;
														assign node1558 = (inp[6]) ? 14'b00101100010010 : 14'b00101110010010;
												assign node1561 = (inp[7]) ? node1569 : node1562;
													assign node1562 = (inp[6]) ? node1566 : node1563;
														assign node1563 = (inp[9]) ? 14'b00101000000010 : 14'b00111010000010;
														assign node1566 = (inp[9]) ? 14'b00111000010010 : 14'b00111000110010;
													assign node1569 = (inp[6]) ? node1571 : 14'b00101010110010;
														assign node1571 = (inp[9]) ? 14'b00101000010010 : 14'b00101000110010;
										assign node1574 = (inp[10]) ? 14'b00000000000001 : node1575;
											assign node1575 = (inp[7]) ? node1585 : node1576;
												assign node1576 = (inp[6]) ? node1582 : node1577;
													assign node1577 = (inp[9]) ? node1579 : 14'b00000000000001;
														assign node1579 = (inp[1]) ? 14'b00101000000100 : 14'b00101100000100;
													assign node1582 = (inp[9]) ? 14'b00111100010100 : 14'b00111100110100;
												assign node1585 = (inp[9]) ? node1591 : node1586;
													assign node1586 = (inp[6]) ? 14'b00101000110100 : node1587;
														assign node1587 = (inp[1]) ? 14'b00101010110100 : 14'b00101110110100;
													assign node1591 = (inp[6]) ? 14'b00101100010100 : 14'b00101110010100;
									assign node1595 = (inp[1]) ? node1609 : node1596;
										assign node1596 = (inp[6]) ? node1602 : node1597;
											assign node1597 = (inp[9]) ? node1599 : 14'b00000000000001;
												assign node1599 = (inp[7]) ? 14'b01100000000100 : 14'b01100100000100;
											assign node1602 = (inp[9]) ? node1606 : node1603;
												assign node1603 = (inp[7]) ? 14'b01110000110100 : 14'b01110100110100;
												assign node1606 = (inp[7]) ? 14'b01110000010100 : 14'b01110100010100;
										assign node1609 = (inp[6]) ? node1617 : node1610;
											assign node1610 = (inp[7]) ? node1614 : node1611;
												assign node1611 = (inp[9]) ? 14'b01110110000100 : 14'b01110110100100;
												assign node1614 = (inp[9]) ? 14'b01110010000100 : 14'b01110010100100;
											assign node1617 = (inp[7]) ? node1621 : node1618;
												assign node1618 = (inp[9]) ? 14'b01110100000100 : 14'b01110100100100;
												assign node1621 = (inp[9]) ? 14'b01110000000100 : 14'b01110000100100;
								assign node1624 = (inp[13]) ? 14'b00000000000001 : node1625;
									assign node1625 = (inp[10]) ? 14'b00000000000001 : node1626;
										assign node1626 = (inp[11]) ? node1652 : node1627;
											assign node1627 = (inp[6]) ? node1639 : node1628;
												assign node1628 = (inp[7]) ? node1634 : node1629;
													assign node1629 = (inp[9]) ? node1631 : 14'b00000000000001;
														assign node1631 = (inp[1]) ? 14'b00000000000000 : 14'b00000100000000;
													assign node1634 = (inp[9]) ? node1636 : 14'b00000110110000;
														assign node1636 = (inp[1]) ? 14'b00000010010000 : 14'b00000110010000;
												assign node1639 = (inp[7]) ? node1647 : node1640;
													assign node1640 = (inp[1]) ? node1644 : node1641;
														assign node1641 = (inp[9]) ? 14'b00010100010000 : 14'b00010100110000;
														assign node1644 = (inp[9]) ? 14'b00010000010000 : 14'b00010000110000;
													assign node1647 = (inp[9]) ? node1649 : 14'b00000100110000;
														assign node1649 = (inp[1]) ? 14'b00000000010000 : 14'b00000100010000;
											assign node1652 = (inp[6]) ? node1666 : node1653;
												assign node1653 = (inp[7]) ? node1659 : node1654;
													assign node1654 = (inp[9]) ? node1656 : 14'b00000000000001;
														assign node1656 = (inp[1]) ? 14'b00100000000100 : 14'b00100100000100;
													assign node1659 = (inp[9]) ? node1663 : node1660;
														assign node1660 = (inp[1]) ? 14'b00100010110100 : 14'b00100110110100;
														assign node1663 = (inp[1]) ? 14'b00100010010100 : 14'b00100110010100;
												assign node1666 = (inp[1]) ? node1672 : node1667;
													assign node1667 = (inp[9]) ? 14'b00110100010100 : node1668;
														assign node1668 = (inp[7]) ? 14'b00100100110100 : 14'b00110100110100;
													assign node1672 = (inp[9]) ? node1676 : node1673;
														assign node1673 = (inp[7]) ? 14'b00100000110100 : 14'b00110000110100;
														assign node1676 = (inp[7]) ? 14'b00100000010100 : 14'b00110000010100;
							assign node1681 = (inp[11]) ? node1763 : node1682;
								assign node1682 = (inp[13]) ? node1744 : node1683;
									assign node1683 = (inp[10]) ? node1725 : node1684;
										assign node1684 = (inp[5]) ? node1704 : node1685;
											assign node1685 = (inp[1]) ? node1693 : node1686;
												assign node1686 = (inp[9]) ? node1690 : node1687;
													assign node1687 = (inp[7]) ? 14'b00101100110110 : 14'b00111100110110;
													assign node1690 = (inp[7]) ? 14'b00101100010110 : 14'b00111100010110;
												assign node1693 = (inp[7]) ? node1699 : node1694;
													assign node1694 = (inp[6]) ? node1696 : 14'b00111010000110;
														assign node1696 = (inp[9]) ? 14'b00111000010110 : 14'b00111000110110;
													assign node1699 = (inp[6]) ? node1701 : 14'b00101010110110;
														assign node1701 = (inp[9]) ? 14'b00101000010110 : 14'b00101000110110;
											assign node1704 = (inp[7]) ? node1714 : node1705;
												assign node1705 = (inp[9]) ? node1709 : node1706;
													assign node1706 = (inp[1]) ? 14'b00110010000110 : 14'b00000000000001;
													assign node1709 = (inp[6]) ? node1711 : 14'b00100100000110;
														assign node1711 = (inp[1]) ? 14'b00110000010110 : 14'b00110100010110;
												assign node1714 = (inp[6]) ? node1722 : node1715;
													assign node1715 = (inp[9]) ? node1719 : node1716;
														assign node1716 = (inp[1]) ? 14'b00100010110110 : 14'b00100110110110;
														assign node1719 = (inp[1]) ? 14'b00100010010110 : 14'b00100110010110;
													assign node1722 = (inp[9]) ? 14'b00100000010110 : 14'b00100000110110;
										assign node1725 = (inp[5]) ? node1727 : 14'b00000000000001;
											assign node1727 = (inp[6]) ? node1735 : node1728;
												assign node1728 = (inp[1]) ? node1730 : 14'b00000000000001;
													assign node1730 = (inp[7]) ? node1732 : 14'b00110010000000;
														assign node1732 = (inp[9]) ? 14'b00100010010000 : 14'b00100010110000;
												assign node1735 = (inp[7]) ? node1741 : node1736;
													assign node1736 = (inp[1]) ? 14'b00110000110000 : node1737;
														assign node1737 = (inp[9]) ? 14'b00110100010000 : 14'b00110100110000;
													assign node1741 = (inp[9]) ? 14'b00100100010000 : 14'b00100100110000;
									assign node1744 = (inp[5]) ? node1746 : 14'b00000000000001;
										assign node1746 = (inp[7]) ? 14'b00000000000001 : node1747;
											assign node1747 = (inp[1]) ? node1755 : node1748;
												assign node1748 = (inp[6]) ? node1752 : node1749;
													assign node1749 = (inp[9]) ? 14'b00000100000000 : 14'b00000000000001;
													assign node1752 = (inp[10]) ? 14'b00010100010000 : 14'b00010100110000;
												assign node1755 = (inp[6]) ? node1759 : node1756;
													assign node1756 = (inp[9]) ? 14'b00010110000000 : 14'b00010110100000;
													assign node1759 = (inp[9]) ? 14'b00010100000000 : 14'b00010100100000;
								assign node1763 = (inp[13]) ? node1765 : 14'b00000000000001;
									assign node1765 = (inp[7]) ? 14'b00000000000001 : node1766;
										assign node1766 = (inp[5]) ? node1768 : 14'b00000000000001;
											assign node1768 = (inp[6]) ? node1776 : node1769;
												assign node1769 = (inp[1]) ? node1773 : node1770;
													assign node1770 = (inp[9]) ? 14'b00000100000000 : 14'b00000000000001;
													assign node1773 = (inp[9]) ? 14'b00010110000000 : 14'b00010110100000;
												assign node1776 = (inp[1]) ? node1780 : node1777;
													assign node1777 = (inp[9]) ? 14'b00010100010000 : 14'b00010100110000;
													assign node1780 = (inp[9]) ? 14'b00010100000000 : 14'b00010100100000;
					assign node1784 = (inp[4]) ? node2122 : node1785;
						assign node1785 = (inp[5]) ? node1983 : node1786;
							assign node1786 = (inp[13]) ? node1926 : node1787;
								assign node1787 = (inp[10]) ? node1877 : node1788;
									assign node1788 = (inp[11]) ? node1832 : node1789;
										assign node1789 = (inp[7]) ? node1809 : node1790;
											assign node1790 = (inp[6]) ? node1800 : node1791;
												assign node1791 = (inp[1]) ? node1793 : 14'b00000000000001;
													assign node1793 = (inp[9]) ? node1797 : node1794;
														assign node1794 = (inp[2]) ? 14'b00011010000110 : 14'b01011010000110;
														assign node1797 = (inp[2]) ? 14'b00001000000110 : 14'b01001000000110;
												assign node1800 = (inp[9]) ? node1804 : node1801;
													assign node1801 = (inp[1]) ? 14'b00011000110110 : 14'b00011100110110;
													assign node1804 = (inp[1]) ? node1806 : 14'b01011100010110;
														assign node1806 = (inp[2]) ? 14'b00011000010110 : 14'b01011000010110;
											assign node1809 = (inp[2]) ? node1821 : node1810;
												assign node1810 = (inp[9]) ? node1816 : node1811;
													assign node1811 = (inp[6]) ? 14'b01001100110110 : node1812;
														assign node1812 = (inp[1]) ? 14'b01001010110110 : 14'b01001110110110;
													assign node1816 = (inp[6]) ? 14'b01001000010110 : node1817;
														assign node1817 = (inp[1]) ? 14'b01001010010110 : 14'b01001110010110;
												assign node1821 = (inp[1]) ? node1827 : node1822;
													assign node1822 = (inp[9]) ? node1824 : 14'b00001110110110;
														assign node1824 = (inp[6]) ? 14'b00001100010110 : 14'b00001110010110;
													assign node1827 = (inp[9]) ? 14'b00001010010110 : node1828;
														assign node1828 = (inp[6]) ? 14'b00001000110110 : 14'b00001010110110;
										assign node1832 = (inp[1]) ? node1856 : node1833;
											assign node1833 = (inp[6]) ? node1843 : node1834;
												assign node1834 = (inp[7]) ? node1840 : node1835;
													assign node1835 = (inp[9]) ? node1837 : 14'b00000000000001;
														assign node1837 = (inp[2]) ? 14'b00001100000100 : 14'b01001100000100;
													assign node1840 = (inp[9]) ? 14'b00001110010100 : 14'b01001110110100;
												assign node1843 = (inp[2]) ? node1849 : node1844;
													assign node1844 = (inp[7]) ? 14'b01001100010100 : node1845;
														assign node1845 = (inp[9]) ? 14'b01011100010100 : 14'b01011100110100;
													assign node1849 = (inp[7]) ? node1853 : node1850;
														assign node1850 = (inp[9]) ? 14'b00011100010100 : 14'b00011100110100;
														assign node1853 = (inp[9]) ? 14'b00001100010100 : 14'b00001100110100;
											assign node1856 = (inp[7]) ? node1864 : node1857;
												assign node1857 = (inp[6]) ? 14'b01011000010100 : node1858;
													assign node1858 = (inp[9]) ? 14'b00001000000100 : node1859;
														assign node1859 = (inp[2]) ? 14'b00011010000100 : 14'b01011010000100;
												assign node1864 = (inp[2]) ? node1870 : node1865;
													assign node1865 = (inp[9]) ? node1867 : 14'b01001000110100;
														assign node1867 = (inp[6]) ? 14'b01001000010100 : 14'b01001010010100;
													assign node1870 = (inp[6]) ? node1874 : node1871;
														assign node1871 = (inp[9]) ? 14'b00001010010100 : 14'b00001010110100;
														assign node1874 = (inp[9]) ? 14'b00001000010100 : 14'b00001000110100;
									assign node1877 = (inp[11]) ? 14'b00000000000001 : node1878;
										assign node1878 = (inp[7]) ? node1900 : node1879;
											assign node1879 = (inp[6]) ? node1887 : node1880;
												assign node1880 = (inp[9]) ? node1882 : 14'b00000000000001;
													assign node1882 = (inp[1]) ? node1884 : 14'b01001100000010;
														assign node1884 = (inp[2]) ? 14'b00001000000010 : 14'b01001000000010;
												assign node1887 = (inp[1]) ? node1893 : node1888;
													assign node1888 = (inp[9]) ? node1890 : 14'b01011100110010;
														assign node1890 = (inp[2]) ? 14'b00011100010010 : 14'b01011100010010;
													assign node1893 = (inp[2]) ? node1897 : node1894;
														assign node1894 = (inp[9]) ? 14'b01011000010010 : 14'b01011000110010;
														assign node1897 = (inp[9]) ? 14'b00011000010010 : 14'b00011000110010;
											assign node1900 = (inp[6]) ? node1914 : node1901;
												assign node1901 = (inp[2]) ? node1909 : node1902;
													assign node1902 = (inp[9]) ? node1906 : node1903;
														assign node1903 = (inp[1]) ? 14'b01001010110010 : 14'b01001110110010;
														assign node1906 = (inp[1]) ? 14'b01001010010010 : 14'b01001110010010;
													assign node1909 = (inp[1]) ? node1911 : 14'b00001110010010;
														assign node1911 = (inp[9]) ? 14'b00001010010010 : 14'b00001010110010;
												assign node1914 = (inp[2]) ? node1918 : node1915;
													assign node1915 = (inp[9]) ? 14'b01001000010010 : 14'b01001000110010;
													assign node1918 = (inp[9]) ? node1922 : node1919;
														assign node1919 = (inp[1]) ? 14'b00001000110010 : 14'b00001100110010;
														assign node1922 = (inp[1]) ? 14'b00001000010010 : 14'b00001100010010;
								assign node1926 = (inp[1]) ? node1952 : node1927;
									assign node1927 = (inp[6]) ? node1937 : node1928;
										assign node1928 = (inp[9]) ? node1930 : 14'b00000000000001;
											assign node1930 = (inp[7]) ? node1934 : node1931;
												assign node1931 = (inp[2]) ? 14'b01000100000000 : 14'b01000100000100;
												assign node1934 = (inp[2]) ? 14'b01000000000000 : 14'b01000000000100;
										assign node1937 = (inp[7]) ? node1945 : node1938;
											assign node1938 = (inp[9]) ? node1942 : node1939;
												assign node1939 = (inp[2]) ? 14'b01010100110000 : 14'b01010100110100;
												assign node1942 = (inp[2]) ? 14'b01010100010000 : 14'b01010100010100;
											assign node1945 = (inp[9]) ? node1949 : node1946;
												assign node1946 = (inp[2]) ? 14'b01010000110000 : 14'b01010000110100;
												assign node1949 = (inp[2]) ? 14'b01010000010000 : 14'b01010000010100;
									assign node1952 = (inp[9]) ? node1968 : node1953;
										assign node1953 = (inp[7]) ? node1961 : node1954;
											assign node1954 = (inp[2]) ? node1958 : node1955;
												assign node1955 = (inp[6]) ? 14'b01010100100100 : 14'b01010110100100;
												assign node1958 = (inp[6]) ? 14'b01010100100000 : 14'b01010110100000;
											assign node1961 = (inp[6]) ? node1965 : node1962;
												assign node1962 = (inp[2]) ? 14'b01010010100000 : 14'b01010010100100;
												assign node1965 = (inp[2]) ? 14'b01010000100000 : 14'b01010000100100;
										assign node1968 = (inp[7]) ? node1976 : node1969;
											assign node1969 = (inp[2]) ? node1973 : node1970;
												assign node1970 = (inp[6]) ? 14'b01010100000100 : 14'b01010110000100;
												assign node1973 = (inp[6]) ? 14'b01010100000000 : 14'b01010110000000;
											assign node1976 = (inp[6]) ? node1980 : node1977;
												assign node1977 = (inp[2]) ? 14'b01010010000000 : 14'b01010010000100;
												assign node1980 = (inp[2]) ? 14'b01010000000000 : 14'b01010000000100;
							assign node1983 = (inp[13]) ? node2111 : node1984;
								assign node1984 = (inp[10]) ? node2082 : node1985;
									assign node1985 = (inp[6]) ? node2033 : node1986;
										assign node1986 = (inp[7]) ? node2008 : node1987;
											assign node1987 = (inp[1]) ? node1997 : node1988;
												assign node1988 = (inp[9]) ? node1990 : 14'b00000000000001;
													assign node1990 = (inp[11]) ? node1994 : node1991;
														assign node1991 = (inp[2]) ? 14'b00000100000110 : 14'b01000100000110;
														assign node1994 = (inp[2]) ? 14'b00000100000100 : 14'b01000100000100;
												assign node1997 = (inp[9]) ? node2005 : node1998;
													assign node1998 = (inp[2]) ? node2002 : node1999;
														assign node1999 = (inp[11]) ? 14'b01010010000100 : 14'b01010010000110;
														assign node2002 = (inp[11]) ? 14'b00010010000100 : 14'b00010010000110;
													assign node2005 = (inp[2]) ? 14'b00000000000100 : 14'b01000000000100;
											assign node2008 = (inp[1]) ? node2018 : node2009;
												assign node2009 = (inp[9]) ? node2015 : node2010;
													assign node2010 = (inp[2]) ? node2012 : 14'b01000110110110;
														assign node2012 = (inp[11]) ? 14'b00000110110100 : 14'b00000110110110;
													assign node2015 = (inp[11]) ? 14'b00000110010100 : 14'b00000110010110;
												assign node2018 = (inp[11]) ? node2026 : node2019;
													assign node2019 = (inp[9]) ? node2023 : node2020;
														assign node2020 = (inp[2]) ? 14'b00000010110110 : 14'b01000010110110;
														assign node2023 = (inp[2]) ? 14'b00000010010110 : 14'b01000010010110;
													assign node2026 = (inp[9]) ? node2030 : node2027;
														assign node2027 = (inp[2]) ? 14'b00000010110100 : 14'b01000010110100;
														assign node2030 = (inp[2]) ? 14'b00000010010100 : 14'b01000010010100;
										assign node2033 = (inp[9]) ? node2055 : node2034;
											assign node2034 = (inp[1]) ? node2044 : node2035;
												assign node2035 = (inp[11]) ? node2039 : node2036;
													assign node2036 = (inp[7]) ? 14'b01000100110110 : 14'b00010100110110;
													assign node2039 = (inp[2]) ? node2041 : 14'b01010100110100;
														assign node2041 = (inp[7]) ? 14'b00000100110100 : 14'b00010100110100;
												assign node2044 = (inp[11]) ? node2048 : node2045;
													assign node2045 = (inp[2]) ? 14'b00010000110110 : 14'b01010000110110;
													assign node2048 = (inp[7]) ? node2052 : node2049;
														assign node2049 = (inp[2]) ? 14'b00010000110100 : 14'b01010000110100;
														assign node2052 = (inp[2]) ? 14'b00000000110100 : 14'b01000000110100;
											assign node2055 = (inp[2]) ? node2069 : node2056;
												assign node2056 = (inp[7]) ? node2064 : node2057;
													assign node2057 = (inp[11]) ? node2061 : node2058;
														assign node2058 = (inp[1]) ? 14'b01010000010110 : 14'b01010100010110;
														assign node2061 = (inp[1]) ? 14'b01010000010100 : 14'b01010100010100;
													assign node2064 = (inp[1]) ? 14'b01000000010110 : node2065;
														assign node2065 = (inp[11]) ? 14'b01000100010100 : 14'b01000100010110;
												assign node2069 = (inp[1]) ? node2075 : node2070;
													assign node2070 = (inp[7]) ? node2072 : 14'b00010100010100;
														assign node2072 = (inp[11]) ? 14'b00000100010100 : 14'b00000100010110;
													assign node2075 = (inp[7]) ? node2079 : node2076;
														assign node2076 = (inp[11]) ? 14'b00010000010100 : 14'b00010000010110;
														assign node2079 = (inp[11]) ? 14'b00000000010100 : 14'b00000000010110;
									assign node2082 = (inp[2]) ? node2084 : 14'b00000000000001;
										assign node2084 = (inp[11]) ? 14'b00000000000001 : node2085;
											assign node2085 = (inp[6]) ? node2099 : node2086;
												assign node2086 = (inp[7]) ? node2094 : node2087;
													assign node2087 = (inp[1]) ? node2091 : node2088;
														assign node2088 = (inp[9]) ? 14'b00000100000010 : 14'b00000000000001;
														assign node2091 = (inp[9]) ? 14'b00000000000010 : 14'b00010010000010;
													assign node2094 = (inp[1]) ? 14'b00000010010010 : node2095;
														assign node2095 = (inp[9]) ? 14'b00000110010010 : 14'b00000110110010;
												assign node2099 = (inp[7]) ? node2105 : node2100;
													assign node2100 = (inp[1]) ? 14'b00010000010010 : node2101;
														assign node2101 = (inp[9]) ? 14'b00010100010010 : 14'b00010100110010;
													assign node2105 = (inp[9]) ? 14'b00000000010010 : node2106;
														assign node2106 = (inp[1]) ? 14'b00000000110010 : 14'b00000100110010;
								assign node2111 = (inp[7]) ? node2113 : 14'b00000000000001;
									assign node2113 = (inp[9]) ? 14'b00000000000001 : node2114;
										assign node2114 = (inp[1]) ? 14'b00000000000001 : node2115;
											assign node2115 = (inp[2]) ? node2117 : 14'b00000000000001;
												assign node2117 = (inp[6]) ? 14'b00000000000001 : 14'b10001000001000;
						assign node2122 = (inp[2]) ? node2258 : node2123;
							assign node2123 = (inp[5]) ? node2207 : node2124;
								assign node2124 = (inp[13]) ? node2178 : node2125;
									assign node2125 = (inp[11]) ? node2151 : node2126;
										assign node2126 = (inp[10]) ? node2128 : 14'b00000000000001;
											assign node2128 = (inp[7]) ? node2138 : node2129;
												assign node2129 = (inp[6]) ? node2135 : node2130;
													assign node2130 = (inp[9]) ? node2132 : 14'b00000000000001;
														assign node2132 = (inp[1]) ? 14'b00101000000000 : 14'b00101100000000;
													assign node2135 = (inp[9]) ? 14'b00111000010000 : 14'b00111100110000;
												assign node2138 = (inp[9]) ? node2146 : node2139;
													assign node2139 = (inp[6]) ? node2143 : node2140;
														assign node2140 = (inp[1]) ? 14'b00101010110000 : 14'b00101110110000;
														assign node2143 = (inp[1]) ? 14'b00101000110000 : 14'b00101100110000;
													assign node2146 = (inp[1]) ? 14'b00101010010000 : node2147;
														assign node2147 = (inp[6]) ? 14'b00101100010000 : 14'b00101110010000;
										assign node2151 = (inp[10]) ? 14'b00000000000001 : node2152;
											assign node2152 = (inp[7]) ? node2164 : node2153;
												assign node2153 = (inp[6]) ? node2159 : node2154;
													assign node2154 = (inp[9]) ? node2156 : 14'b00000000000001;
														assign node2156 = (inp[1]) ? 14'b01001000000000 : 14'b01001100000000;
													assign node2159 = (inp[1]) ? 14'b01011000010000 : node2160;
														assign node2160 = (inp[9]) ? 14'b01011100010000 : 14'b01011100110000;
												assign node2164 = (inp[6]) ? node2170 : node2165;
													assign node2165 = (inp[9]) ? node2167 : 14'b01001110110000;
														assign node2167 = (inp[1]) ? 14'b01001010010000 : 14'b01001110010000;
													assign node2170 = (inp[9]) ? node2174 : node2171;
														assign node2171 = (inp[1]) ? 14'b01001000110000 : 14'b01001100110000;
														assign node2174 = (inp[1]) ? 14'b01001000010000 : 14'b01001100010000;
									assign node2178 = (inp[6]) ? node2192 : node2179;
										assign node2179 = (inp[1]) ? node2185 : node2180;
											assign node2180 = (inp[9]) ? node2182 : 14'b00000000000001;
												assign node2182 = (inp[7]) ? 14'b00000000000100 : 14'b00000100000100;
											assign node2185 = (inp[7]) ? node2189 : node2186;
												assign node2186 = (inp[9]) ? 14'b00010110000100 : 14'b00010110100100;
												assign node2189 = (inp[9]) ? 14'b00010010000100 : 14'b00010010100100;
										assign node2192 = (inp[7]) ? node2200 : node2193;
											assign node2193 = (inp[1]) ? node2197 : node2194;
												assign node2194 = (inp[9]) ? 14'b00010100010100 : 14'b00010100110100;
												assign node2197 = (inp[9]) ? 14'b00010100000100 : 14'b00010100100100;
											assign node2200 = (inp[9]) ? node2204 : node2201;
												assign node2201 = (inp[1]) ? 14'b00010000100100 : 14'b00010000110100;
												assign node2204 = (inp[1]) ? 14'b00010000000100 : 14'b00010000010100;
								assign node2207 = (inp[10]) ? 14'b00000000000001 : node2208;
									assign node2208 = (inp[13]) ? 14'b00000000000001 : node2209;
										assign node2209 = (inp[7]) ? node2231 : node2210;
											assign node2210 = (inp[6]) ? node2222 : node2211;
												assign node2211 = (inp[1]) ? node2217 : node2212;
													assign node2212 = (inp[9]) ? node2214 : 14'b00000000000001;
														assign node2214 = (inp[11]) ? 14'b01000100000000 : 14'b01000100000010;
													assign node2217 = (inp[9]) ? 14'b01000000000010 : node2218;
														assign node2218 = (inp[11]) ? 14'b01010010000000 : 14'b01010010000010;
												assign node2222 = (inp[11]) ? node2226 : node2223;
													assign node2223 = (inp[9]) ? 14'b01010000010010 : 14'b01010000110010;
													assign node2226 = (inp[9]) ? 14'b01010100010000 : node2227;
														assign node2227 = (inp[1]) ? 14'b01010000110000 : 14'b01010100110000;
											assign node2231 = (inp[1]) ? node2245 : node2232;
												assign node2232 = (inp[11]) ? node2240 : node2233;
													assign node2233 = (inp[9]) ? node2237 : node2234;
														assign node2234 = (inp[6]) ? 14'b01000100110010 : 14'b01000110110010;
														assign node2237 = (inp[6]) ? 14'b01000100010010 : 14'b01000110010010;
													assign node2240 = (inp[6]) ? node2242 : 14'b01000110010000;
														assign node2242 = (inp[9]) ? 14'b01000100010000 : 14'b01000100110000;
												assign node2245 = (inp[6]) ? node2249 : node2246;
													assign node2246 = (inp[11]) ? 14'b01000010110000 : 14'b01000010110010;
													assign node2249 = (inp[9]) ? node2253 : node2250;
														assign node2250 = (inp[11]) ? 14'b01000000110000 : 14'b01000000110010;
														assign node2253 = (inp[11]) ? 14'b01000000010000 : 14'b01000000010010;
							assign node2258 = (inp[9]) ? 14'b00000000000001 : node2259;
								assign node2259 = (inp[10]) ? node2261 : 14'b00000000000001;
									assign node2261 = (inp[5]) ? node2263 : 14'b00000000000001;
										assign node2263 = (inp[7]) ? node2265 : 14'b00000000000001;
											assign node2265 = (inp[13]) ? node2267 : 14'b00000000000001;
												assign node2267 = (inp[1]) ? 14'b00000000000001 : node2268;
													assign node2268 = (inp[6]) ? 14'b00000000000001 : 14'b10001001000010;
				assign node2273 = (inp[6]) ? node2667 : node2274;
					assign node2274 = (inp[7]) ? node2582 : node2275;
						assign node2275 = (inp[13]) ? node2495 : node2276;
							assign node2276 = (inp[11]) ? node2430 : node2277;
								assign node2277 = (inp[12]) ? node2365 : node2278;
									assign node2278 = (inp[2]) ? node2330 : node2279;
										assign node2279 = (inp[5]) ? node2303 : node2280;
											assign node2280 = (inp[4]) ? node2288 : node2281;
												assign node2281 = (inp[10]) ? node2283 : 14'b00000000000001;
													assign node2283 = (inp[9]) ? node2285 : 14'b01111110110010;
														assign node2285 = (inp[1]) ? 14'b01111010010010 : 14'b01111110010010;
												assign node2288 = (inp[10]) ? node2296 : node2289;
													assign node2289 = (inp[1]) ? node2293 : node2290;
														assign node2290 = (inp[9]) ? 14'b01111110010110 : 14'b01111110110110;
														assign node2293 = (inp[9]) ? 14'b01111010010110 : 14'b01111010110110;
													assign node2296 = (inp[1]) ? node2300 : node2297;
														assign node2297 = (inp[9]) ? 14'b01111110010000 : 14'b01111110110000;
														assign node2300 = (inp[9]) ? 14'b01111010010000 : 14'b01111010110000;
											assign node2303 = (inp[9]) ? node2317 : node2304;
												assign node2304 = (inp[1]) ? node2312 : node2305;
													assign node2305 = (inp[10]) ? node2309 : node2306;
														assign node2306 = (inp[4]) ? 14'b01110110110110 : 14'b00110110110010;
														assign node2309 = (inp[4]) ? 14'b01110110110000 : 14'b01110110110010;
													assign node2312 = (inp[4]) ? 14'b01110010110110 : node2313;
														assign node2313 = (inp[10]) ? 14'b01110010110010 : 14'b00110010110010;
												assign node2317 = (inp[1]) ? node2325 : node2318;
													assign node2318 = (inp[4]) ? node2322 : node2319;
														assign node2319 = (inp[10]) ? 14'b01110110010010 : 14'b00110110010010;
														assign node2322 = (inp[10]) ? 14'b01110110010000 : 14'b01110110010110;
													assign node2325 = (inp[10]) ? node2327 : 14'b00110010010010;
														assign node2327 = (inp[4]) ? 14'b01110010010000 : 14'b01110010010010;
										assign node2330 = (inp[10]) ? node2350 : node2331;
											assign node2331 = (inp[4]) ? node2339 : node2332;
												assign node2332 = (inp[9]) ? 14'b00011110010000 : node2333;
													assign node2333 = (inp[5]) ? node2335 : 14'b00011010110000;
														assign node2335 = (inp[1]) ? 14'b00010010110000 : 14'b00010110110000;
												assign node2339 = (inp[5]) ? node2345 : node2340;
													assign node2340 = (inp[9]) ? 14'b00111110010110 : node2341;
														assign node2341 = (inp[1]) ? 14'b00111010110110 : 14'b00111110110110;
													assign node2345 = (inp[9]) ? 14'b00110010010110 : node2346;
														assign node2346 = (inp[1]) ? 14'b00110010110110 : 14'b00110110110110;
											assign node2350 = (inp[5]) ? node2356 : node2351;
												assign node2351 = (inp[4]) ? 14'b00000000000001 : node2352;
													assign node2352 = (inp[9]) ? 14'b00111010010010 : 14'b00111010110010;
												assign node2356 = (inp[4]) ? node2358 : 14'b00000000000001;
													assign node2358 = (inp[1]) ? node2362 : node2359;
														assign node2359 = (inp[9]) ? 14'b00110110010000 : 14'b00110110110000;
														assign node2362 = (inp[9]) ? 14'b00110010010000 : 14'b00110010110000;
									assign node2365 = (inp[4]) ? node2411 : node2366;
										assign node2366 = (inp[10]) ? node2394 : node2367;
											assign node2367 = (inp[1]) ? node2381 : node2368;
												assign node2368 = (inp[2]) ? node2374 : node2369;
													assign node2369 = (inp[9]) ? 14'b01011110010110 : node2370;
														assign node2370 = (inp[5]) ? 14'b01010110110110 : 14'b01011110110110;
													assign node2374 = (inp[9]) ? node2378 : node2375;
														assign node2375 = (inp[5]) ? 14'b00010110110110 : 14'b00011110110110;
														assign node2378 = (inp[5]) ? 14'b00010110010110 : 14'b00011110010110;
												assign node2381 = (inp[2]) ? node2387 : node2382;
													assign node2382 = (inp[9]) ? 14'b01010010010110 : node2383;
														assign node2383 = (inp[5]) ? 14'b01010010110110 : 14'b01011010110110;
													assign node2387 = (inp[5]) ? node2391 : node2388;
														assign node2388 = (inp[9]) ? 14'b00011010010110 : 14'b00011010110110;
														assign node2391 = (inp[9]) ? 14'b00010010010110 : 14'b00010010110110;
											assign node2394 = (inp[5]) ? node2404 : node2395;
												assign node2395 = (inp[9]) ? node2399 : node2396;
													assign node2396 = (inp[2]) ? 14'b00011010110010 : 14'b01011010110010;
													assign node2399 = (inp[2]) ? node2401 : 14'b01011010010010;
														assign node2401 = (inp[1]) ? 14'b00011010010010 : 14'b00011110010010;
												assign node2404 = (inp[2]) ? node2406 : 14'b00000000000001;
													assign node2406 = (inp[1]) ? node2408 : 14'b00010110110010;
														assign node2408 = (inp[9]) ? 14'b00010010010010 : 14'b00010010110010;
										assign node2411 = (inp[2]) ? 14'b00000000000001 : node2412;
											assign node2412 = (inp[10]) ? node2420 : node2413;
												assign node2413 = (inp[5]) ? node2415 : 14'b00000000000001;
													assign node2415 = (inp[9]) ? 14'b01010010010010 : node2416;
														assign node2416 = (inp[1]) ? 14'b01010010110010 : 14'b01010110110010;
												assign node2420 = (inp[5]) ? 14'b00000000000001 : node2421;
													assign node2421 = (inp[1]) ? node2425 : node2422;
														assign node2422 = (inp[9]) ? 14'b00111110010000 : 14'b00111110110000;
														assign node2425 = (inp[9]) ? 14'b00111010010000 : 14'b00111010110000;
								assign node2430 = (inp[10]) ? 14'b00000000000001 : node2431;
									assign node2431 = (inp[4]) ? node2479 : node2432;
										assign node2432 = (inp[5]) ? node2454 : node2433;
											assign node2433 = (inp[12]) ? node2443 : node2434;
												assign node2434 = (inp[9]) ? node2440 : node2435;
													assign node2435 = (inp[2]) ? 14'b00111010110100 : node2436;
														assign node2436 = (inp[1]) ? 14'b01111010110100 : 14'b01111110110100;
													assign node2440 = (inp[2]) ? 14'b00111010010100 : 14'b01111010010100;
												assign node2443 = (inp[1]) ? node2449 : node2444;
													assign node2444 = (inp[9]) ? 14'b00011110010100 : node2445;
														assign node2445 = (inp[2]) ? 14'b00011110110100 : 14'b01011110110100;
													assign node2449 = (inp[9]) ? 14'b01011010010100 : node2450;
														assign node2450 = (inp[2]) ? 14'b00011010110100 : 14'b01011010110100;
											assign node2454 = (inp[9]) ? node2466 : node2455;
												assign node2455 = (inp[2]) ? node2459 : node2456;
													assign node2456 = (inp[1]) ? 14'b01110010110100 : 14'b01110110110100;
													assign node2459 = (inp[12]) ? node2463 : node2460;
														assign node2460 = (inp[1]) ? 14'b00110010110100 : 14'b00110110110100;
														assign node2463 = (inp[1]) ? 14'b00010010110100 : 14'b00010110110100;
												assign node2466 = (inp[1]) ? node2474 : node2467;
													assign node2467 = (inp[2]) ? node2471 : node2468;
														assign node2468 = (inp[12]) ? 14'b01010110010100 : 14'b01110110010100;
														assign node2471 = (inp[12]) ? 14'b00010110010100 : 14'b00110110010100;
													assign node2474 = (inp[12]) ? node2476 : 14'b00110010010100;
														assign node2476 = (inp[2]) ? 14'b00010010010100 : 14'b01010010010100;
										assign node2479 = (inp[12]) ? node2481 : 14'b00000000000001;
											assign node2481 = (inp[2]) ? 14'b00000000000001 : node2482;
												assign node2482 = (inp[5]) ? node2488 : node2483;
													assign node2483 = (inp[9]) ? node2485 : 14'b01011010110000;
														assign node2485 = (inp[1]) ? 14'b01011010010000 : 14'b01011110010000;
													assign node2488 = (inp[1]) ? node2490 : 14'b01010110110000;
														assign node2490 = (inp[9]) ? 14'b01010010010000 : 14'b01010010110000;
							assign node2495 = (inp[5]) ? node2555 : node2496;
								assign node2496 = (inp[1]) ? node2520 : node2497;
									assign node2497 = (inp[4]) ? node2511 : node2498;
										assign node2498 = (inp[12]) ? node2504 : node2499;
											assign node2499 = (inp[2]) ? node2501 : 14'b00000000000001;
												assign node2501 = (inp[9]) ? 14'b01110110010100 : 14'b01110110110100;
											assign node2504 = (inp[2]) ? node2508 : node2505;
												assign node2505 = (inp[9]) ? 14'b01010110010100 : 14'b01010110110100;
												assign node2508 = (inp[9]) ? 14'b01010110010000 : 14'b01010110110000;
										assign node2511 = (inp[2]) ? 14'b00000000000001 : node2512;
											assign node2512 = (inp[12]) ? node2516 : node2513;
												assign node2513 = (inp[9]) ? 14'b00110110010100 : 14'b00110110110100;
												assign node2516 = (inp[9]) ? 14'b00010110010100 : 14'b00010110110100;
									assign node2520 = (inp[12]) ? node2542 : node2521;
										assign node2521 = (inp[9]) ? node2529 : node2522;
											assign node2522 = (inp[4]) ? node2526 : node2523;
												assign node2523 = (inp[2]) ? 14'b01100110100100 : 14'b00000000000001;
												assign node2526 = (inp[2]) ? 14'b00000000000001 : 14'b00100110100100;
											assign node2529 = (inp[10]) ? node2535 : node2530;
												assign node2530 = (inp[4]) ? node2532 : 14'b00000000000001;
													assign node2532 = (inp[2]) ? 14'b00000000000001 : 14'b00100110000100;
												assign node2535 = (inp[4]) ? node2539 : node2536;
													assign node2536 = (inp[2]) ? 14'b01100110000100 : 14'b00000000000001;
													assign node2539 = (inp[2]) ? 14'b00000000000001 : 14'b00100110000100;
										assign node2542 = (inp[2]) ? node2550 : node2543;
											assign node2543 = (inp[9]) ? node2547 : node2544;
												assign node2544 = (inp[4]) ? 14'b00000110100100 : 14'b01000110100100;
												assign node2547 = (inp[4]) ? 14'b00000110000100 : 14'b01000110000100;
											assign node2550 = (inp[4]) ? 14'b00000000000001 : node2551;
												assign node2551 = (inp[9]) ? 14'b01000110000000 : 14'b01000110100000;
								assign node2555 = (inp[12]) ? 14'b00000000000001 : node2556;
									assign node2556 = (inp[2]) ? node2572 : node2557;
										assign node2557 = (inp[1]) ? node2565 : node2558;
											assign node2558 = (inp[9]) ? node2562 : node2559;
												assign node2559 = (inp[4]) ? 14'b00110110110000 : 14'b01110110110000;
												assign node2562 = (inp[4]) ? 14'b00110110010000 : 14'b01110110010000;
											assign node2565 = (inp[9]) ? node2569 : node2566;
												assign node2566 = (inp[4]) ? 14'b00100110100000 : 14'b01100110100000;
												assign node2569 = (inp[4]) ? 14'b00100110000000 : 14'b01100110000000;
										assign node2572 = (inp[4]) ? node2574 : 14'b00000000000001;
											assign node2574 = (inp[1]) ? node2578 : node2575;
												assign node2575 = (inp[9]) ? 14'b00010110010000 : 14'b00010110110000;
												assign node2578 = (inp[9]) ? 14'b00000110000000 : 14'b00000110100000;
						assign node2582 = (inp[13]) ? node2598 : node2583;
							assign node2583 = (inp[12]) ? 14'b00000000000001 : node2584;
								assign node2584 = (inp[5]) ? 14'b00000000000001 : node2585;
									assign node2585 = (inp[10]) ? 14'b00000000000001 : node2586;
										assign node2586 = (inp[2]) ? 14'b00000000000001 : node2587;
											assign node2587 = (inp[9]) ? 14'b00000000000001 : node2588;
												assign node2588 = (inp[1]) ? 14'b00000000000001 : node2589;
													assign node2589 = (inp[4]) ? 14'b10000001000000 : 14'b00000000000001;
							assign node2598 = (inp[5]) ? node2648 : node2599;
								assign node2599 = (inp[4]) ? node2631 : node2600;
									assign node2600 = (inp[1]) ? node2616 : node2601;
										assign node2601 = (inp[9]) ? node2609 : node2602;
											assign node2602 = (inp[2]) ? node2606 : node2603;
												assign node2603 = (inp[12]) ? 14'b01010010110100 : 14'b00010010110000;
												assign node2606 = (inp[12]) ? 14'b01010010110000 : 14'b01110010110100;
											assign node2609 = (inp[2]) ? node2613 : node2610;
												assign node2610 = (inp[12]) ? 14'b01010010010100 : 14'b00010010010000;
												assign node2613 = (inp[12]) ? 14'b01010010010000 : 14'b01110010010100;
										assign node2616 = (inp[9]) ? node2624 : node2617;
											assign node2617 = (inp[12]) ? node2621 : node2618;
												assign node2618 = (inp[2]) ? 14'b01100010100100 : 14'b00000010100000;
												assign node2621 = (inp[2]) ? 14'b01000010100000 : 14'b01000010100100;
											assign node2624 = (inp[12]) ? node2628 : node2625;
												assign node2625 = (inp[2]) ? 14'b01100010000100 : 14'b00000010000000;
												assign node2628 = (inp[2]) ? 14'b01000010000000 : 14'b01000010000100;
									assign node2631 = (inp[2]) ? 14'b00000000000001 : node2632;
										assign node2632 = (inp[1]) ? node2640 : node2633;
											assign node2633 = (inp[12]) ? node2637 : node2634;
												assign node2634 = (inp[9]) ? 14'b00110010010100 : 14'b00110010110100;
												assign node2637 = (inp[9]) ? 14'b00010010010100 : 14'b00010010110100;
											assign node2640 = (inp[12]) ? node2644 : node2641;
												assign node2641 = (inp[9]) ? 14'b00100010000100 : 14'b00100010100100;
												assign node2644 = (inp[9]) ? 14'b00000010000100 : 14'b00000010100100;
								assign node2648 = (inp[12]) ? 14'b00000000000001 : node2649;
									assign node2649 = (inp[2]) ? 14'b00000000000001 : node2650;
										assign node2650 = (inp[1]) ? node2658 : node2651;
											assign node2651 = (inp[9]) ? node2655 : node2652;
												assign node2652 = (inp[4]) ? 14'b00110010110000 : 14'b01110010110000;
												assign node2655 = (inp[4]) ? 14'b00110010010000 : 14'b01110010010000;
											assign node2658 = (inp[9]) ? node2662 : node2659;
												assign node2659 = (inp[4]) ? 14'b00100010100000 : 14'b01100010100000;
												assign node2662 = (inp[4]) ? 14'b00100010000000 : 14'b01100010000000;
					assign node2667 = (inp[9]) ? 14'b00000000000001 : node2668;
						assign node2668 = (inp[13]) ? node2854 : node2669;
							assign node2669 = (inp[11]) ? node2797 : node2670;
								assign node2670 = (inp[7]) ? node2718 : node2671;
									assign node2671 = (inp[1]) ? node2673 : 14'b00000000000001;
										assign node2673 = (inp[4]) ? node2701 : node2674;
											assign node2674 = (inp[5]) ? node2688 : node2675;
												assign node2675 = (inp[12]) ? node2683 : node2676;
													assign node2676 = (inp[10]) ? node2680 : node2677;
														assign node2677 = (inp[2]) ? 14'b00011000100000 : 14'b00000000000001;
														assign node2680 = (inp[2]) ? 14'b00111000100010 : 14'b01111000100010;
													assign node2683 = (inp[10]) ? 14'b00011000100010 : node2684;
														assign node2684 = (inp[2]) ? 14'b00011000100110 : 14'b01011000100110;
												assign node2688 = (inp[10]) ? node2694 : node2689;
													assign node2689 = (inp[2]) ? node2691 : 14'b00110000100010;
														assign node2691 = (inp[12]) ? 14'b00010000100110 : 14'b00010000100000;
													assign node2694 = (inp[12]) ? node2698 : node2695;
														assign node2695 = (inp[2]) ? 14'b00000000000001 : 14'b01110000100010;
														assign node2698 = (inp[2]) ? 14'b00010000100010 : 14'b00000000000001;
											assign node2701 = (inp[12]) ? node2709 : node2702;
												assign node2702 = (inp[5]) ? node2704 : 14'b00000000000001;
													assign node2704 = (inp[10]) ? 14'b00110000100000 : node2705;
														assign node2705 = (inp[2]) ? 14'b00110000100110 : 14'b01110000100110;
												assign node2709 = (inp[2]) ? 14'b00000000000001 : node2710;
													assign node2710 = (inp[10]) ? node2714 : node2711;
														assign node2711 = (inp[5]) ? 14'b01010000100010 : 14'b00000000000001;
														assign node2714 = (inp[5]) ? 14'b00000000000001 : 14'b00111000100000;
									assign node2718 = (inp[2]) ? node2762 : node2719;
										assign node2719 = (inp[12]) ? node2747 : node2720;
											assign node2720 = (inp[1]) ? node2734 : node2721;
												assign node2721 = (inp[4]) ? node2727 : node2722;
													assign node2722 = (inp[10]) ? 14'b01101100100010 : node2723;
														assign node2723 = (inp[5]) ? 14'b00100100100010 : 14'b00000000000001;
													assign node2727 = (inp[10]) ? node2731 : node2728;
														assign node2728 = (inp[5]) ? 14'b01100100100110 : 14'b01101100100110;
														assign node2731 = (inp[5]) ? 14'b01100100100000 : 14'b01101100100000;
												assign node2734 = (inp[5]) ? node2740 : node2735;
													assign node2735 = (inp[10]) ? node2737 : 14'b01101000100110;
														assign node2737 = (inp[4]) ? 14'b01101000100000 : 14'b01101000100010;
													assign node2740 = (inp[10]) ? node2744 : node2741;
														assign node2741 = (inp[4]) ? 14'b01100000100110 : 14'b00100000100010;
														assign node2744 = (inp[4]) ? 14'b01100000100000 : 14'b01100000100010;
											assign node2747 = (inp[10]) ? node2755 : node2748;
												assign node2748 = (inp[5]) ? node2750 : 14'b00000000000001;
													assign node2750 = (inp[4]) ? node2752 : 14'b01000000100110;
														assign node2752 = (inp[1]) ? 14'b01000000100010 : 14'b01000100100010;
												assign node2755 = (inp[5]) ? 14'b00000000000001 : node2756;
													assign node2756 = (inp[4]) ? 14'b00101000100000 : node2757;
														assign node2757 = (inp[1]) ? 14'b01001000100010 : 14'b01001100100010;
										assign node2762 = (inp[4]) ? node2788 : node2763;
											assign node2763 = (inp[5]) ? node2777 : node2764;
												assign node2764 = (inp[1]) ? node2770 : node2765;
													assign node2765 = (inp[12]) ? node2767 : 14'b00001100100000;
														assign node2767 = (inp[10]) ? 14'b00001100100010 : 14'b00001100100110;
													assign node2770 = (inp[10]) ? node2774 : node2771;
														assign node2771 = (inp[12]) ? 14'b00001000100110 : 14'b00001000100000;
														assign node2774 = (inp[12]) ? 14'b00001000100010 : 14'b00101000100010;
												assign node2777 = (inp[12]) ? node2783 : node2778;
													assign node2778 = (inp[10]) ? 14'b00000000000001 : node2779;
														assign node2779 = (inp[1]) ? 14'b00000000100000 : 14'b00000100100000;
													assign node2783 = (inp[10]) ? node2785 : 14'b00000100100110;
														assign node2785 = (inp[1]) ? 14'b00000000100010 : 14'b00000100100010;
											assign node2788 = (inp[12]) ? 14'b00000000000001 : node2789;
												assign node2789 = (inp[10]) ? 14'b00000000000001 : node2790;
													assign node2790 = (inp[5]) ? node2792 : 14'b00101100100110;
														assign node2792 = (inp[1]) ? 14'b00100000100110 : 14'b00100100100110;
								assign node2797 = (inp[10]) ? 14'b00000000000001 : node2798;
									assign node2798 = (inp[4]) ? node2834 : node2799;
										assign node2799 = (inp[1]) ? node2807 : node2800;
											assign node2800 = (inp[7]) ? node2802 : 14'b00000000000001;
												assign node2802 = (inp[2]) ? node2804 : 14'b01101100100100;
													assign node2804 = (inp[12]) ? 14'b00000100100100 : 14'b00100100100100;
											assign node2807 = (inp[2]) ? node2823 : node2808;
												assign node2808 = (inp[12]) ? node2816 : node2809;
													assign node2809 = (inp[5]) ? node2813 : node2810;
														assign node2810 = (inp[7]) ? 14'b01101000100100 : 14'b01111000100100;
														assign node2813 = (inp[7]) ? 14'b01100000100100 : 14'b01110000100100;
													assign node2816 = (inp[7]) ? node2820 : node2817;
														assign node2817 = (inp[5]) ? 14'b01010000100100 : 14'b01011000100100;
														assign node2820 = (inp[5]) ? 14'b01000000100100 : 14'b01001000100100;
												assign node2823 = (inp[5]) ? node2827 : node2824;
													assign node2824 = (inp[12]) ? 14'b00011000100100 : 14'b00111000100100;
													assign node2827 = (inp[12]) ? node2831 : node2828;
														assign node2828 = (inp[7]) ? 14'b00100000100100 : 14'b00110000100100;
														assign node2831 = (inp[7]) ? 14'b00000000100100 : 14'b00010000100100;
										assign node2834 = (inp[2]) ? 14'b00000000000001 : node2835;
											assign node2835 = (inp[12]) ? node2843 : node2836;
												assign node2836 = (inp[1]) ? 14'b00000000000001 : node2837;
													assign node2837 = (inp[5]) ? 14'b00000000000001 : node2838;
														assign node2838 = (inp[7]) ? 14'b00000000000001 : 14'b10000001001000;
												assign node2843 = (inp[7]) ? node2847 : node2844;
													assign node2844 = (inp[5]) ? 14'b01010000100000 : 14'b00000000000001;
													assign node2847 = (inp[5]) ? node2849 : 14'b01001100100000;
														assign node2849 = (inp[1]) ? 14'b01000000100000 : 14'b01000100100000;
							assign node2854 = (inp[7]) ? node2874 : node2855;
								assign node2855 = (inp[1]) ? 14'b00000000000001 : node2856;
									assign node2856 = (inp[12]) ? node2866 : node2857;
										assign node2857 = (inp[2]) ? node2859 : 14'b00000000000001;
											assign node2859 = (inp[5]) ? node2863 : node2860;
												assign node2860 = (inp[4]) ? 14'b10000001001010 : 14'b00000000000001;
												assign node2863 = (inp[4]) ? 14'b00000000000001 : 14'b10000001001000;
										assign node2866 = (inp[2]) ? 14'b00000000000001 : node2867;
											assign node2867 = (inp[4]) ? 14'b00000000000001 : node2868;
												assign node2868 = (inp[5]) ? 14'b10001000000010 : 14'b00000000000001;
								assign node2874 = (inp[12]) ? 14'b00000000000001 : node2875;
									assign node2875 = (inp[4]) ? node2877 : 14'b00000000000001;
										assign node2877 = (inp[1]) ? node2879 : 14'b00000000000001;
											assign node2879 = (inp[2]) ? node2881 : 14'b00000000000001;
												assign node2881 = (inp[5]) ? 14'b00000000000001 : 14'b10000000000000;
			assign node2886 = (inp[7]) ? node3646 : node2887;
				assign node2887 = (inp[1]) ? node3329 : node2888;
					assign node2888 = (inp[3]) ? node3178 : node2889;
						assign node2889 = (inp[13]) ? node3105 : node2890;
							assign node2890 = (inp[11]) ? node3042 : node2891;
								assign node2891 = (inp[12]) ? node2979 : node2892;
									assign node2892 = (inp[9]) ? node2938 : node2893;
										assign node2893 = (inp[4]) ? node2913 : node2894;
											assign node2894 = (inp[10]) ? node2900 : node2895;
												assign node2895 = (inp[5]) ? node2897 : 14'b00000000000001;
													assign node2897 = (inp[2]) ? 14'b00010110100000 : 14'b00110110100010;
												assign node2900 = (inp[2]) ? node2908 : node2901;
													assign node2901 = (inp[6]) ? node2905 : node2902;
														assign node2902 = (inp[5]) ? 14'b01110110100010 : 14'b01111110100010;
														assign node2905 = (inp[5]) ? 14'b01110100100010 : 14'b01111100100010;
													assign node2908 = (inp[5]) ? 14'b00000000000001 : node2909;
														assign node2909 = (inp[6]) ? 14'b00111100100010 : 14'b00111110100010;
											assign node2913 = (inp[10]) ? node2929 : node2914;
												assign node2914 = (inp[2]) ? node2922 : node2915;
													assign node2915 = (inp[6]) ? node2919 : node2916;
														assign node2916 = (inp[5]) ? 14'b01110110100110 : 14'b01111110100110;
														assign node2919 = (inp[5]) ? 14'b01110100100110 : 14'b01111100100110;
													assign node2922 = (inp[5]) ? node2926 : node2923;
														assign node2923 = (inp[6]) ? 14'b00111100100110 : 14'b00111110100110;
														assign node2926 = (inp[6]) ? 14'b00110100100110 : 14'b00110110100110;
												assign node2929 = (inp[6]) ? node2933 : node2930;
													assign node2930 = (inp[2]) ? 14'b00110110100000 : 14'b01110110100000;
													assign node2933 = (inp[2]) ? 14'b00110100100000 : node2934;
														assign node2934 = (inp[5]) ? 14'b01110100100000 : 14'b01111100100000;
										assign node2938 = (inp[2]) ? node2954 : node2939;
											assign node2939 = (inp[10]) ? node2943 : node2940;
												assign node2940 = (inp[5]) ? 14'b01110110000110 : 14'b00000000000001;
												assign node2943 = (inp[6]) ? node2949 : node2944;
													assign node2944 = (inp[4]) ? 14'b01110110000000 : node2945;
														assign node2945 = (inp[5]) ? 14'b01110110000010 : 14'b01111110000010;
													assign node2949 = (inp[4]) ? node2951 : 14'b01111100000010;
														assign node2951 = (inp[5]) ? 14'b01110100000000 : 14'b01111100000000;
											assign node2954 = (inp[10]) ? node2970 : node2955;
												assign node2955 = (inp[4]) ? node2963 : node2956;
													assign node2956 = (inp[6]) ? node2960 : node2957;
														assign node2957 = (inp[5]) ? 14'b00010110000000 : 14'b00011110000000;
														assign node2960 = (inp[5]) ? 14'b00010100000000 : 14'b00011100000000;
													assign node2963 = (inp[6]) ? node2967 : node2964;
														assign node2964 = (inp[5]) ? 14'b00110110000110 : 14'b00111110000110;
														assign node2967 = (inp[5]) ? 14'b00110100000110 : 14'b00111100000110;
												assign node2970 = (inp[5]) ? node2976 : node2971;
													assign node2971 = (inp[4]) ? 14'b00000000000001 : node2972;
														assign node2972 = (inp[6]) ? 14'b00111100000010 : 14'b00111110000010;
													assign node2976 = (inp[4]) ? 14'b00110110000000 : 14'b00000000000001;
									assign node2979 = (inp[4]) ? node3027 : node2980;
										assign node2980 = (inp[5]) ? node3004 : node2981;
											assign node2981 = (inp[10]) ? node2997 : node2982;
												assign node2982 = (inp[9]) ? node2990 : node2983;
													assign node2983 = (inp[2]) ? node2987 : node2984;
														assign node2984 = (inp[6]) ? 14'b01011100100110 : 14'b01011110100110;
														assign node2987 = (inp[6]) ? 14'b00011100100110 : 14'b00011110100110;
													assign node2990 = (inp[6]) ? node2994 : node2991;
														assign node2991 = (inp[2]) ? 14'b00011110000110 : 14'b01011110000110;
														assign node2994 = (inp[2]) ? 14'b00011100000110 : 14'b01011100000110;
												assign node2997 = (inp[9]) ? 14'b01011110000010 : node2998;
													assign node2998 = (inp[2]) ? 14'b00011110100010 : node2999;
														assign node2999 = (inp[6]) ? 14'b01011100100010 : 14'b01011110100010;
											assign node3004 = (inp[10]) ? node3018 : node3005;
												assign node3005 = (inp[6]) ? node3013 : node3006;
													assign node3006 = (inp[9]) ? node3010 : node3007;
														assign node3007 = (inp[2]) ? 14'b00010110100110 : 14'b01010110100110;
														assign node3010 = (inp[2]) ? 14'b00010110000110 : 14'b01010110000110;
													assign node3013 = (inp[9]) ? node3015 : 14'b00010100100110;
														assign node3015 = (inp[2]) ? 14'b00010100000110 : 14'b01010100000110;
												assign node3018 = (inp[2]) ? node3020 : 14'b00000000000001;
													assign node3020 = (inp[9]) ? node3024 : node3021;
														assign node3021 = (inp[6]) ? 14'b00010100100010 : 14'b00010110100010;
														assign node3024 = (inp[6]) ? 14'b00010100000010 : 14'b00010110000010;
										assign node3027 = (inp[2]) ? 14'b00000000000001 : node3028;
											assign node3028 = (inp[5]) ? node3036 : node3029;
												assign node3029 = (inp[10]) ? node3031 : 14'b00000000000001;
													assign node3031 = (inp[9]) ? 14'b00111100000000 : node3032;
														assign node3032 = (inp[6]) ? 14'b00111100100000 : 14'b00111110100000;
												assign node3036 = (inp[10]) ? 14'b00000000000001 : node3037;
													assign node3037 = (inp[6]) ? 14'b01010100100010 : 14'b01010110100010;
								assign node3042 = (inp[10]) ? 14'b00000000000001 : node3043;
									assign node3043 = (inp[4]) ? node3089 : node3044;
										assign node3044 = (inp[12]) ? node3064 : node3045;
											assign node3045 = (inp[2]) ? node3057 : node3046;
												assign node3046 = (inp[6]) ? node3052 : node3047;
													assign node3047 = (inp[9]) ? node3049 : 14'b01110110100100;
														assign node3049 = (inp[5]) ? 14'b01110110000100 : 14'b01111110000100;
													assign node3052 = (inp[5]) ? 14'b01110100000100 : node3053;
														assign node3053 = (inp[9]) ? 14'b01111100000100 : 14'b01111100100100;
												assign node3057 = (inp[9]) ? node3061 : node3058;
													assign node3058 = (inp[6]) ? 14'b00111100100100 : 14'b00111110100100;
													assign node3061 = (inp[6]) ? 14'b00111100000100 : 14'b00111110000100;
											assign node3064 = (inp[2]) ? node3078 : node3065;
												assign node3065 = (inp[9]) ? node3073 : node3066;
													assign node3066 = (inp[5]) ? node3070 : node3067;
														assign node3067 = (inp[6]) ? 14'b01011100100100 : 14'b01011110100100;
														assign node3070 = (inp[6]) ? 14'b01010100100100 : 14'b01010110100100;
													assign node3073 = (inp[5]) ? 14'b01010100000100 : node3074;
														assign node3074 = (inp[6]) ? 14'b01011100000100 : 14'b01011110000100;
												assign node3078 = (inp[6]) ? node3086 : node3079;
													assign node3079 = (inp[9]) ? node3083 : node3080;
														assign node3080 = (inp[5]) ? 14'b00010110100100 : 14'b00011110100100;
														assign node3083 = (inp[5]) ? 14'b00010110000100 : 14'b00011110000100;
													assign node3086 = (inp[9]) ? 14'b00010100000100 : 14'b00010100100100;
										assign node3089 = (inp[2]) ? 14'b00000000000001 : node3090;
											assign node3090 = (inp[12]) ? node3092 : 14'b00000000000001;
												assign node3092 = (inp[9]) ? node3098 : node3093;
													assign node3093 = (inp[5]) ? 14'b01010100100000 : node3094;
														assign node3094 = (inp[6]) ? 14'b01011100100000 : 14'b01011110100000;
													assign node3098 = (inp[6]) ? 14'b01010100000000 : node3099;
														assign node3099 = (inp[5]) ? 14'b01010110000000 : 14'b01011110000000;
							assign node3105 = (inp[5]) ? node3151 : node3106;
								assign node3106 = (inp[12]) ? node3126 : node3107;
									assign node3107 = (inp[4]) ? node3117 : node3108;
										assign node3108 = (inp[2]) ? node3110 : 14'b00000000000001;
											assign node3110 = (inp[6]) ? node3114 : node3111;
												assign node3111 = (inp[9]) ? 14'b01100110010100 : 14'b01100110110100;
												assign node3114 = (inp[9]) ? 14'b01100100010100 : 14'b01100100110100;
										assign node3117 = (inp[2]) ? 14'b00000000000001 : node3118;
											assign node3118 = (inp[9]) ? node3122 : node3119;
												assign node3119 = (inp[6]) ? 14'b00100100110100 : 14'b00100110110100;
												assign node3122 = (inp[6]) ? 14'b00100100010100 : 14'b00100110010100;
									assign node3126 = (inp[2]) ? node3142 : node3127;
										assign node3127 = (inp[6]) ? node3135 : node3128;
											assign node3128 = (inp[4]) ? node3132 : node3129;
												assign node3129 = (inp[9]) ? 14'b01000110010100 : 14'b01000110110100;
												assign node3132 = (inp[9]) ? 14'b00000110010100 : 14'b00000110110100;
											assign node3135 = (inp[9]) ? node3139 : node3136;
												assign node3136 = (inp[4]) ? 14'b00000100110100 : 14'b01000100110100;
												assign node3139 = (inp[4]) ? 14'b00000100010100 : 14'b01000100010100;
										assign node3142 = (inp[4]) ? 14'b00000000000001 : node3143;
											assign node3143 = (inp[6]) ? node3147 : node3144;
												assign node3144 = (inp[9]) ? 14'b01000110010000 : 14'b01000110110000;
												assign node3147 = (inp[9]) ? 14'b01000100010000 : 14'b01000100110000;
								assign node3151 = (inp[12]) ? 14'b00000000000001 : node3152;
									assign node3152 = (inp[2]) ? node3168 : node3153;
										assign node3153 = (inp[9]) ? node3161 : node3154;
											assign node3154 = (inp[6]) ? node3158 : node3155;
												assign node3155 = (inp[4]) ? 14'b00100110110000 : 14'b01100110110000;
												assign node3158 = (inp[4]) ? 14'b00100100110000 : 14'b01100100110000;
											assign node3161 = (inp[6]) ? node3165 : node3162;
												assign node3162 = (inp[4]) ? 14'b00100110010000 : 14'b01100110010000;
												assign node3165 = (inp[4]) ? 14'b00100100010000 : 14'b01100100010000;
										assign node3168 = (inp[4]) ? node3170 : 14'b00000000000001;
											assign node3170 = (inp[9]) ? node3174 : node3171;
												assign node3171 = (inp[6]) ? 14'b00000100110000 : 14'b00000110110000;
												assign node3174 = (inp[6]) ? 14'b00000100010000 : 14'b00000110010000;
						assign node3178 = (inp[9]) ? 14'b00000000000001 : node3179;
							assign node3179 = (inp[13]) ? node3293 : node3180;
								assign node3180 = (inp[11]) ? node3258 : node3181;
									assign node3181 = (inp[4]) ? node3229 : node3182;
										assign node3182 = (inp[5]) ? node3206 : node3183;
											assign node3183 = (inp[12]) ? node3191 : node3184;
												assign node3184 = (inp[10]) ? node3186 : 14'b00000000000001;
													assign node3186 = (inp[2]) ? node3188 : 14'b01101110100010;
														assign node3188 = (inp[6]) ? 14'b00101110000010 : 14'b00101110100010;
												assign node3191 = (inp[2]) ? node3199 : node3192;
													assign node3192 = (inp[6]) ? node3196 : node3193;
														assign node3193 = (inp[10]) ? 14'b01001110100010 : 14'b01001110100110;
														assign node3196 = (inp[10]) ? 14'b01001110000010 : 14'b01001110000110;
													assign node3199 = (inp[6]) ? node3203 : node3200;
														assign node3200 = (inp[10]) ? 14'b00001110100010 : 14'b00001110100110;
														assign node3203 = (inp[10]) ? 14'b00001110000010 : 14'b00001110000110;
											assign node3206 = (inp[10]) ? node3220 : node3207;
												assign node3207 = (inp[12]) ? node3215 : node3208;
													assign node3208 = (inp[2]) ? node3212 : node3209;
														assign node3209 = (inp[6]) ? 14'b00100110000010 : 14'b00100110100010;
														assign node3212 = (inp[6]) ? 14'b00000110000000 : 14'b00000110100000;
													assign node3215 = (inp[2]) ? node3217 : 14'b01000110100110;
														assign node3217 = (inp[6]) ? 14'b00000110000110 : 14'b00000110100110;
												assign node3220 = (inp[2]) ? node3226 : node3221;
													assign node3221 = (inp[12]) ? 14'b00000000000001 : node3222;
														assign node3222 = (inp[6]) ? 14'b01100110000010 : 14'b01100110100010;
													assign node3226 = (inp[12]) ? 14'b00000110000010 : 14'b00000000000001;
										assign node3229 = (inp[12]) ? node3247 : node3230;
											assign node3230 = (inp[10]) ? node3236 : node3231;
												assign node3231 = (inp[2]) ? 14'b00101110000110 : node3232;
													assign node3232 = (inp[5]) ? 14'b01100110000110 : 14'b01101110100110;
												assign node3236 = (inp[2]) ? node3244 : node3237;
													assign node3237 = (inp[5]) ? node3241 : node3238;
														assign node3238 = (inp[6]) ? 14'b01101110000000 : 14'b01101110100000;
														assign node3241 = (inp[6]) ? 14'b01100110000000 : 14'b01100110100000;
													assign node3244 = (inp[5]) ? 14'b00100110100000 : 14'b00000000000001;
											assign node3247 = (inp[2]) ? 14'b00000000000001 : node3248;
												assign node3248 = (inp[5]) ? node3254 : node3249;
													assign node3249 = (inp[10]) ? node3251 : 14'b00000000000001;
														assign node3251 = (inp[6]) ? 14'b00101110000000 : 14'b00101110100000;
													assign node3254 = (inp[10]) ? 14'b00000000000001 : 14'b01000110000010;
									assign node3258 = (inp[10]) ? 14'b00000000000001 : node3259;
										assign node3259 = (inp[4]) ? node3283 : node3260;
											assign node3260 = (inp[5]) ? node3270 : node3261;
												assign node3261 = (inp[2]) ? node3265 : node3262;
													assign node3262 = (inp[12]) ? 14'b01001110100100 : 14'b01101110100100;
													assign node3265 = (inp[12]) ? node3267 : 14'b00101110100100;
														assign node3267 = (inp[6]) ? 14'b00001110000100 : 14'b00001110100100;
												assign node3270 = (inp[12]) ? node3278 : node3271;
													assign node3271 = (inp[6]) ? node3275 : node3272;
														assign node3272 = (inp[2]) ? 14'b00100110100100 : 14'b01100110100100;
														assign node3275 = (inp[2]) ? 14'b00100110000100 : 14'b01100110000100;
													assign node3278 = (inp[2]) ? 14'b00000110100100 : node3279;
														assign node3279 = (inp[6]) ? 14'b01000110000100 : 14'b01000110100100;
											assign node3283 = (inp[12]) ? node3285 : 14'b00000000000001;
												assign node3285 = (inp[2]) ? 14'b00000000000001 : node3286;
													assign node3286 = (inp[5]) ? node3288 : 14'b01001110100000;
														assign node3288 = (inp[6]) ? 14'b01000110000000 : 14'b01000110100000;
								assign node3293 = (inp[6]) ? node3303 : node3294;
									assign node3294 = (inp[2]) ? node3296 : 14'b00000000000001;
										assign node3296 = (inp[12]) ? 14'b00000000000001 : node3297;
											assign node3297 = (inp[5]) ? node3299 : 14'b00000000000001;
												assign node3299 = (inp[11]) ? 14'b00000000000001 : 14'b10000001000000;
									assign node3303 = (inp[12]) ? node3319 : node3304;
										assign node3304 = (inp[5]) ? node3312 : node3305;
											assign node3305 = (inp[4]) ? node3309 : node3306;
												assign node3306 = (inp[2]) ? 14'b01100100100100 : 14'b00000000000001;
												assign node3309 = (inp[2]) ? 14'b00000000000001 : 14'b00100100100100;
											assign node3312 = (inp[2]) ? node3316 : node3313;
												assign node3313 = (inp[4]) ? 14'b00100100100000 : 14'b01100100100000;
												assign node3316 = (inp[4]) ? 14'b00000100100000 : 14'b00000000000001;
										assign node3319 = (inp[5]) ? 14'b00000000000001 : node3320;
											assign node3320 = (inp[4]) ? node3324 : node3321;
												assign node3321 = (inp[2]) ? 14'b01000100100000 : 14'b01000100100100;
												assign node3324 = (inp[2]) ? 14'b00000000000001 : 14'b00000100100100;
					assign node3329 = (inp[13]) ? node3607 : node3330;
						assign node3330 = (inp[6]) ? node3524 : node3331;
							assign node3331 = (inp[9]) ? node3463 : node3332;
								assign node3332 = (inp[11]) ? node3424 : node3333;
									assign node3333 = (inp[3]) ? node3381 : node3334;
										assign node3334 = (inp[12]) ? node3358 : node3335;
											assign node3335 = (inp[5]) ? node3347 : node3336;
												assign node3336 = (inp[10]) ? node3342 : node3337;
													assign node3337 = (inp[4]) ? 14'b01111010100110 : node3338;
														assign node3338 = (inp[2]) ? 14'b00011010100000 : 14'b00000000000001;
													assign node3342 = (inp[4]) ? 14'b01111010100000 : node3343;
														assign node3343 = (inp[2]) ? 14'b00111010100010 : 14'b01111010100010;
												assign node3347 = (inp[10]) ? node3355 : node3348;
													assign node3348 = (inp[4]) ? node3352 : node3349;
														assign node3349 = (inp[2]) ? 14'b00010010100000 : 14'b00110010100010;
														assign node3352 = (inp[2]) ? 14'b00110010100110 : 14'b01110010100110;
													assign node3355 = (inp[2]) ? 14'b00110010100000 : 14'b01110010100000;
											assign node3358 = (inp[4]) ? node3374 : node3359;
												assign node3359 = (inp[5]) ? node3367 : node3360;
													assign node3360 = (inp[10]) ? node3364 : node3361;
														assign node3361 = (inp[2]) ? 14'b00011010100110 : 14'b01011010100110;
														assign node3364 = (inp[2]) ? 14'b00011010100010 : 14'b01011010100010;
													assign node3367 = (inp[10]) ? node3371 : node3368;
														assign node3368 = (inp[2]) ? 14'b00010010100110 : 14'b01010010100110;
														assign node3371 = (inp[2]) ? 14'b00010010100010 : 14'b00000000000001;
												assign node3374 = (inp[2]) ? 14'b00000000000001 : node3375;
													assign node3375 = (inp[5]) ? 14'b01010010100010 : node3376;
														assign node3376 = (inp[10]) ? 14'b00111010100000 : 14'b00000000000001;
										assign node3381 = (inp[5]) ? node3409 : node3382;
											assign node3382 = (inp[4]) ? node3398 : node3383;
												assign node3383 = (inp[10]) ? node3391 : node3384;
													assign node3384 = (inp[12]) ? node3388 : node3385;
														assign node3385 = (inp[2]) ? 14'b00001010100000 : 14'b00000000000001;
														assign node3388 = (inp[2]) ? 14'b00001010100110 : 14'b01001010100110;
													assign node3391 = (inp[2]) ? node3395 : node3392;
														assign node3392 = (inp[12]) ? 14'b01001010100010 : 14'b01101010100010;
														assign node3395 = (inp[12]) ? 14'b00001010100010 : 14'b00101010100010;
												assign node3398 = (inp[12]) ? node3404 : node3399;
													assign node3399 = (inp[10]) ? node3401 : 14'b00101010100110;
														assign node3401 = (inp[2]) ? 14'b00000000000001 : 14'b01101010100000;
													assign node3404 = (inp[10]) ? node3406 : 14'b00000000000001;
														assign node3406 = (inp[2]) ? 14'b00000000000001 : 14'b00101010100000;
											assign node3409 = (inp[12]) ? node3417 : node3410;
												assign node3410 = (inp[2]) ? node3414 : node3411;
													assign node3411 = (inp[4]) ? 14'b01100010100110 : 14'b01100010100010;
													assign node3414 = (inp[4]) ? 14'b00100010100110 : 14'b00000010100000;
												assign node3417 = (inp[10]) ? node3421 : node3418;
													assign node3418 = (inp[4]) ? 14'b01000010100010 : 14'b01000010100110;
													assign node3421 = (inp[2]) ? 14'b00000010100010 : 14'b00000000000001;
									assign node3424 = (inp[10]) ? 14'b00000000000001 : node3425;
										assign node3425 = (inp[4]) ? node3451 : node3426;
											assign node3426 = (inp[12]) ? node3438 : node3427;
												assign node3427 = (inp[5]) ? node3433 : node3428;
													assign node3428 = (inp[2]) ? node3430 : 14'b01101010100100;
														assign node3430 = (inp[3]) ? 14'b00101010100100 : 14'b00111010100100;
													assign node3433 = (inp[3]) ? 14'b00100010100100 : node3434;
														assign node3434 = (inp[2]) ? 14'b00110010100100 : 14'b01110010100100;
												assign node3438 = (inp[5]) ? node3446 : node3439;
													assign node3439 = (inp[3]) ? node3443 : node3440;
														assign node3440 = (inp[2]) ? 14'b00011010100100 : 14'b01011010100100;
														assign node3443 = (inp[2]) ? 14'b00001010100100 : 14'b01001010100100;
													assign node3446 = (inp[2]) ? node3448 : 14'b01000010100100;
														assign node3448 = (inp[3]) ? 14'b00000010100100 : 14'b00010010100100;
											assign node3451 = (inp[2]) ? 14'b00000000000001 : node3452;
												assign node3452 = (inp[12]) ? node3454 : 14'b00000000000001;
													assign node3454 = (inp[3]) ? node3458 : node3455;
														assign node3455 = (inp[5]) ? 14'b01010010100000 : 14'b01011010100000;
														assign node3458 = (inp[5]) ? 14'b01000010100000 : 14'b01001010100000;
								assign node3463 = (inp[3]) ? node3465 : 14'b00000000000001;
									assign node3465 = (inp[10]) ? node3503 : node3466;
										assign node3466 = (inp[4]) ? node3490 : node3467;
											assign node3467 = (inp[5]) ? node3477 : node3468;
												assign node3468 = (inp[2]) ? node3472 : node3469;
													assign node3469 = (inp[11]) ? 14'b01001010000100 : 14'b01001010000110;
													assign node3472 = (inp[11]) ? node3474 : 14'b00001010000000;
														assign node3474 = (inp[12]) ? 14'b00001010000100 : 14'b00101010000100;
												assign node3477 = (inp[11]) ? node3485 : node3478;
													assign node3478 = (inp[12]) ? node3482 : node3479;
														assign node3479 = (inp[2]) ? 14'b00000010000000 : 14'b00100010000010;
														assign node3482 = (inp[2]) ? 14'b00000010000110 : 14'b01000010000110;
													assign node3485 = (inp[2]) ? 14'b00000010000100 : node3486;
														assign node3486 = (inp[12]) ? 14'b01000010000100 : 14'b01100010000100;
											assign node3490 = (inp[11]) ? node3498 : node3491;
												assign node3491 = (inp[12]) ? 14'b00000000000001 : node3492;
													assign node3492 = (inp[2]) ? node3494 : 14'b01101010000110;
														assign node3494 = (inp[5]) ? 14'b00100010000110 : 14'b00101010000110;
												assign node3498 = (inp[12]) ? node3500 : 14'b00000000000001;
													assign node3500 = (inp[5]) ? 14'b01000010000000 : 14'b01001010000000;
										assign node3503 = (inp[11]) ? 14'b00000000000001 : node3504;
											assign node3504 = (inp[4]) ? node3516 : node3505;
												assign node3505 = (inp[5]) ? node3513 : node3506;
													assign node3506 = (inp[12]) ? node3510 : node3507;
														assign node3507 = (inp[2]) ? 14'b00101010000010 : 14'b01101010000010;
														assign node3510 = (inp[2]) ? 14'b00001010000010 : 14'b01001010000010;
													assign node3513 = (inp[12]) ? 14'b00000000000001 : 14'b01100010000010;
												assign node3516 = (inp[12]) ? 14'b00000000000001 : node3517;
													assign node3517 = (inp[5]) ? node3519 : 14'b00000000000001;
														assign node3519 = (inp[2]) ? 14'b00100010000000 : 14'b01100010000000;
							assign node3524 = (inp[3]) ? 14'b00000000000001 : node3525;
								assign node3525 = (inp[9]) ? node3537 : node3526;
									assign node3526 = (inp[5]) ? 14'b00000000000001 : node3527;
										assign node3527 = (inp[2]) ? node3529 : 14'b00000000000001;
											assign node3529 = (inp[11]) ? node3531 : 14'b00000000000001;
												assign node3531 = (inp[10]) ? 14'b00000000000001 : node3532;
													assign node3532 = (inp[4]) ? 14'b10000000000000 : 14'b00000000000001;
									assign node3537 = (inp[11]) ? node3581 : node3538;
										assign node3538 = (inp[12]) ? node3562 : node3539;
											assign node3539 = (inp[2]) ? node3551 : node3540;
												assign node3540 = (inp[5]) ? node3544 : node3541;
													assign node3541 = (inp[10]) ? 14'b01111000000000 : 14'b01111000000110;
													assign node3544 = (inp[4]) ? node3548 : node3545;
														assign node3545 = (inp[10]) ? 14'b01110000000010 : 14'b00110000000010;
														assign node3548 = (inp[10]) ? 14'b01110000000000 : 14'b01110000000110;
												assign node3551 = (inp[10]) ? node3557 : node3552;
													assign node3552 = (inp[4]) ? node3554 : 14'b00010000000000;
														assign node3554 = (inp[5]) ? 14'b00110000000110 : 14'b00111000000110;
													assign node3557 = (inp[4]) ? node3559 : 14'b00111000000010;
														assign node3559 = (inp[5]) ? 14'b00110000000000 : 14'b00000000000001;
											assign node3562 = (inp[4]) ? node3572 : node3563;
												assign node3563 = (inp[2]) ? node3567 : node3564;
													assign node3564 = (inp[10]) ? 14'b01011000000010 : 14'b01010000000110;
													assign node3567 = (inp[5]) ? 14'b00010000000010 : node3568;
														assign node3568 = (inp[10]) ? 14'b00011000000010 : 14'b00011000000110;
												assign node3572 = (inp[2]) ? 14'b00000000000001 : node3573;
													assign node3573 = (inp[10]) ? node3577 : node3574;
														assign node3574 = (inp[5]) ? 14'b01010000000010 : 14'b00000000000001;
														assign node3577 = (inp[5]) ? 14'b00000000000001 : 14'b00111000000000;
										assign node3581 = (inp[10]) ? 14'b00000000000001 : node3582;
											assign node3582 = (inp[4]) ? node3598 : node3583;
												assign node3583 = (inp[2]) ? node3591 : node3584;
													assign node3584 = (inp[5]) ? node3588 : node3585;
														assign node3585 = (inp[12]) ? 14'b01011000000100 : 14'b01111000000100;
														assign node3588 = (inp[12]) ? 14'b01010000000100 : 14'b01110000000100;
													assign node3591 = (inp[5]) ? node3595 : node3592;
														assign node3592 = (inp[12]) ? 14'b00011000000100 : 14'b00111000000100;
														assign node3595 = (inp[12]) ? 14'b00010000000100 : 14'b00110000000100;
												assign node3598 = (inp[12]) ? node3600 : 14'b00000000000001;
													assign node3600 = (inp[2]) ? 14'b00000000000001 : node3601;
														assign node3601 = (inp[5]) ? 14'b01010000000000 : 14'b01011000000000;
						assign node3607 = (inp[6]) ? 14'b00000000000001 : node3608;
							assign node3608 = (inp[12]) ? node3634 : node3609;
								assign node3609 = (inp[5]) ? node3625 : node3610;
									assign node3610 = (inp[9]) ? node3618 : node3611;
										assign node3611 = (inp[4]) ? node3613 : 14'b00000000000001;
											assign node3613 = (inp[3]) ? 14'b00000000000001 : node3614;
												assign node3614 = (inp[2]) ? 14'b10000001000010 : 14'b00000000000001;
										assign node3618 = (inp[4]) ? 14'b00000000000001 : node3619;
											assign node3619 = (inp[3]) ? node3621 : 14'b00000000000001;
												assign node3621 = (inp[2]) ? 14'b00000000000001 : 14'b10000000000010;
									assign node3625 = (inp[3]) ? 14'b00000000000001 : node3626;
										assign node3626 = (inp[9]) ? 14'b00000000000001 : node3627;
											assign node3627 = (inp[2]) ? node3629 : 14'b00000000000001;
												assign node3629 = (inp[4]) ? 14'b00000000000001 : 14'b10000000001010;
								assign node3634 = (inp[5]) ? node3636 : 14'b00000000000001;
									assign node3636 = (inp[2]) ? 14'b00000000000001 : node3637;
										assign node3637 = (inp[3]) ? 14'b00000000000001 : node3638;
											assign node3638 = (inp[9]) ? 14'b00000000000001 : node3639;
												assign node3639 = (inp[4]) ? 14'b00000000000001 : 14'b10001001001000;
				assign node3646 = (inp[13]) ? node3648 : 14'b00000000000001;
					assign node3648 = (inp[1]) ? node3744 : node3649;
						assign node3649 = (inp[3]) ? node3719 : node3650;
							assign node3650 = (inp[5]) ? node3700 : node3651;
								assign node3651 = (inp[4]) ? node3683 : node3652;
									assign node3652 = (inp[6]) ? node3668 : node3653;
										assign node3653 = (inp[9]) ? node3661 : node3654;
											assign node3654 = (inp[12]) ? node3658 : node3655;
												assign node3655 = (inp[2]) ? 14'b01100010110100 : 14'b00000010110000;
												assign node3658 = (inp[2]) ? 14'b01000010110000 : 14'b01000010110100;
											assign node3661 = (inp[12]) ? node3665 : node3662;
												assign node3662 = (inp[2]) ? 14'b01100010010100 : 14'b00000010010000;
												assign node3665 = (inp[2]) ? 14'b01000010010000 : 14'b01000010010100;
										assign node3668 = (inp[9]) ? node3676 : node3669;
											assign node3669 = (inp[12]) ? node3673 : node3670;
												assign node3670 = (inp[2]) ? 14'b01100000110100 : 14'b00000000110000;
												assign node3673 = (inp[2]) ? 14'b01000000110000 : 14'b01000000110100;
											assign node3676 = (inp[12]) ? node3680 : node3677;
												assign node3677 = (inp[2]) ? 14'b01100000010100 : 14'b00000000010000;
												assign node3680 = (inp[2]) ? 14'b01000000010000 : 14'b01000000010100;
									assign node3683 = (inp[2]) ? 14'b00000000000001 : node3684;
										assign node3684 = (inp[12]) ? node3692 : node3685;
											assign node3685 = (inp[9]) ? node3689 : node3686;
												assign node3686 = (inp[6]) ? 14'b00100000110100 : 14'b00100010110100;
												assign node3689 = (inp[6]) ? 14'b00100000010100 : 14'b00100010010100;
											assign node3692 = (inp[6]) ? node3696 : node3693;
												assign node3693 = (inp[9]) ? 14'b00000010010100 : 14'b00000010110100;
												assign node3696 = (inp[9]) ? 14'b00000000010100 : 14'b00000000110100;
								assign node3700 = (inp[2]) ? 14'b00000000000001 : node3701;
									assign node3701 = (inp[12]) ? 14'b00000000000001 : node3702;
										assign node3702 = (inp[4]) ? node3710 : node3703;
											assign node3703 = (inp[6]) ? node3707 : node3704;
												assign node3704 = (inp[9]) ? 14'b01100010010000 : 14'b01100010110000;
												assign node3707 = (inp[9]) ? 14'b01100000010000 : 14'b01100000110000;
											assign node3710 = (inp[6]) ? node3714 : node3711;
												assign node3711 = (inp[9]) ? 14'b00100010010000 : 14'b00100010110000;
												assign node3714 = (inp[9]) ? 14'b00100000010000 : 14'b00100000110000;
							assign node3719 = (inp[6]) ? node3721 : 14'b00000000000001;
								assign node3721 = (inp[9]) ? 14'b00000000000001 : node3722;
									assign node3722 = (inp[5]) ? node3736 : node3723;
										assign node3723 = (inp[4]) ? node3731 : node3724;
											assign node3724 = (inp[2]) ? node3728 : node3725;
												assign node3725 = (inp[12]) ? 14'b01000000100100 : 14'b00000000100000;
												assign node3728 = (inp[12]) ? 14'b01000000100000 : 14'b01100000100100;
											assign node3731 = (inp[2]) ? 14'b00000000000001 : node3732;
												assign node3732 = (inp[12]) ? 14'b00000000100100 : 14'b00100000100100;
										assign node3736 = (inp[12]) ? 14'b00000000000001 : node3737;
											assign node3737 = (inp[2]) ? 14'b00000000000001 : node3738;
												assign node3738 = (inp[4]) ? 14'b00100000100000 : 14'b01100000100000;
						assign node3744 = (inp[12]) ? node3746 : 14'b00000000000001;
							assign node3746 = (inp[2]) ? node3748 : 14'b00000000000001;
								assign node3748 = (inp[3]) ? node3750 : 14'b00000000000001;
									assign node3750 = (inp[9]) ? node3752 : 14'b00000000000001;
										assign node3752 = (inp[5]) ? node3754 : 14'b00000000000001;
											assign node3754 = (inp[4]) ? 14'b10001001001010 : node3755;
												assign node3755 = (inp[6]) ? 14'b10001001000000 : 14'b10001000000000;

endmodule