module dtc_split5_bm76 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node41;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node50;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node92;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node111;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node141;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node241;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node247;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node264;
	wire [3-1:0] node268;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node283;
	wire [3-1:0] node287;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node304;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node322;
	wire [3-1:0] node325;
	wire [3-1:0] node327;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node333;
	wire [3-1:0] node336;
	wire [3-1:0] node338;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node347;
	wire [3-1:0] node349;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node356;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node367;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node385;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node406;
	wire [3-1:0] node408;
	wire [3-1:0] node410;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node425;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node433;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node446;
	wire [3-1:0] node450;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node469;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node493;
	wire [3-1:0] node497;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node502;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node518;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node527;
	wire [3-1:0] node532;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node537;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node547;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node554;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node575;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node592;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node611;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node618;
	wire [3-1:0] node620;
	wire [3-1:0] node622;
	wire [3-1:0] node625;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node638;

	assign outp = (inp[9]) ? node438 : node1;
		assign node1 = (inp[6]) ? node187 : node2;
			assign node2 = (inp[10]) ? node72 : node3;
				assign node3 = (inp[7]) ? node17 : node4;
					assign node4 = (inp[8]) ? node6 : 3'b111;
						assign node6 = (inp[3]) ? node8 : 3'b111;
							assign node8 = (inp[11]) ? node10 : 3'b111;
								assign node10 = (inp[4]) ? 3'b011 : node11;
									assign node11 = (inp[0]) ? node13 : 3'b111;
										assign node13 = (inp[5]) ? 3'b011 : 3'b111;
					assign node17 = (inp[11]) ? node45 : node18;
						assign node18 = (inp[3]) ? node30 : node19;
							assign node19 = (inp[4]) ? node21 : 3'b111;
								assign node21 = (inp[8]) ? node23 : 3'b111;
									assign node23 = (inp[5]) ? 3'b011 : node24;
										assign node24 = (inp[1]) ? node26 : 3'b111;
											assign node26 = (inp[0]) ? 3'b011 : 3'b111;
							assign node30 = (inp[8]) ? 3'b011 : node31;
								assign node31 = (inp[4]) ? node33 : 3'b111;
									assign node33 = (inp[0]) ? node39 : node34;
										assign node34 = (inp[1]) ? node36 : 3'b111;
											assign node36 = (inp[2]) ? 3'b111 : 3'b011;
										assign node39 = (inp[1]) ? node41 : 3'b011;
											assign node41 = (inp[2]) ? 3'b011 : 3'b111;
						assign node45 = (inp[8]) ? node63 : node46;
							assign node46 = (inp[4]) ? node54 : node47;
								assign node47 = (inp[3]) ? 3'b011 : node48;
									assign node48 = (inp[5]) ? node50 : 3'b111;
										assign node50 = (inp[0]) ? 3'b011 : 3'b111;
								assign node54 = (inp[3]) ? node56 : 3'b011;
									assign node56 = (inp[5]) ? node58 : 3'b011;
										assign node58 = (inp[2]) ? 3'b101 : node59;
											assign node59 = (inp[0]) ? 3'b101 : 3'b011;
							assign node63 = (inp[3]) ? 3'b101 : node64;
								assign node64 = (inp[4]) ? node66 : 3'b011;
									assign node66 = (inp[0]) ? 3'b101 : node67;
										assign node67 = (inp[5]) ? 3'b101 : 3'b011;
				assign node72 = (inp[7]) ? node118 : node73;
					assign node73 = (inp[11]) ? node101 : node74;
						assign node74 = (inp[8]) ? node92 : node75;
							assign node75 = (inp[3]) ? node85 : node76;
								assign node76 = (inp[1]) ? node78 : 3'b111;
									assign node78 = (inp[0]) ? node80 : 3'b111;
										assign node80 = (inp[5]) ? node82 : 3'b111;
											assign node82 = (inp[4]) ? 3'b011 : 3'b111;
								assign node85 = (inp[2]) ? 3'b011 : node86;
									assign node86 = (inp[5]) ? 3'b011 : node87;
										assign node87 = (inp[0]) ? 3'b011 : 3'b111;
							assign node92 = (inp[3]) ? node94 : 3'b011;
								assign node94 = (inp[4]) ? 3'b101 : node95;
									assign node95 = (inp[0]) ? node97 : 3'b011;
										assign node97 = (inp[5]) ? 3'b101 : 3'b011;
						assign node101 = (inp[3]) ? node111 : node102;
							assign node102 = (inp[8]) ? 3'b101 : node103;
								assign node103 = (inp[0]) ? node105 : 3'b011;
									assign node105 = (inp[5]) ? node107 : 3'b011;
										assign node107 = (inp[4]) ? 3'b101 : 3'b011;
							assign node111 = (inp[8]) ? node113 : 3'b101;
								assign node113 = (inp[1]) ? 3'b001 : node114;
									assign node114 = (inp[4]) ? 3'b001 : 3'b101;
					assign node118 = (inp[11]) ? node150 : node119;
						assign node119 = (inp[8]) ? node137 : node120;
							assign node120 = (inp[3]) ? node130 : node121;
								assign node121 = (inp[4]) ? 3'b101 : node122;
									assign node122 = (inp[5]) ? node124 : 3'b011;
										assign node124 = (inp[0]) ? 3'b101 : node125;
											assign node125 = (inp[1]) ? 3'b111 : 3'b011;
								assign node130 = (inp[4]) ? node132 : 3'b101;
									assign node132 = (inp[5]) ? 3'b001 : node133;
										assign node133 = (inp[0]) ? 3'b001 : 3'b101;
							assign node137 = (inp[3]) ? 3'b001 : node138;
								assign node138 = (inp[4]) ? node144 : node139;
									assign node139 = (inp[0]) ? node141 : 3'b101;
										assign node141 = (inp[5]) ? 3'b001 : 3'b101;
									assign node144 = (inp[5]) ? 3'b001 : node145;
										assign node145 = (inp[2]) ? 3'b001 : 3'b101;
						assign node150 = (inp[8]) ? node168 : node151;
							assign node151 = (inp[3]) ? node157 : node152;
								assign node152 = (inp[5]) ? 3'b001 : node153;
									assign node153 = (inp[0]) ? 3'b001 : 3'b101;
								assign node157 = (inp[5]) ? node163 : node158;
									assign node158 = (inp[0]) ? node160 : 3'b001;
										assign node160 = (inp[4]) ? 3'b110 : 3'b001;
									assign node163 = (inp[4]) ? 3'b110 : node164;
										assign node164 = (inp[0]) ? 3'b110 : 3'b001;
							assign node168 = (inp[3]) ? node178 : node169;
								assign node169 = (inp[4]) ? node171 : 3'b001;
									assign node171 = (inp[2]) ? 3'b110 : node172;
										assign node172 = (inp[5]) ? 3'b110 : node173;
											assign node173 = (inp[1]) ? 3'b110 : 3'b001;
								assign node178 = (inp[2]) ? 3'b110 : node179;
									assign node179 = (inp[4]) ? node181 : 3'b110;
										assign node181 = (inp[5]) ? node183 : 3'b110;
											assign node183 = (inp[1]) ? 3'b010 : 3'b110;
			assign node187 = (inp[10]) ? node341 : node188;
				assign node188 = (inp[7]) ? node258 : node189;
					assign node189 = (inp[11]) ? node231 : node190;
						assign node190 = (inp[2]) ? node212 : node191;
							assign node191 = (inp[8]) ? node199 : node192;
								assign node192 = (inp[3]) ? node194 : 3'b011;
									assign node194 = (inp[0]) ? 3'b101 : node195;
										assign node195 = (inp[4]) ? 3'b101 : 3'b011;
								assign node199 = (inp[3]) ? node205 : node200;
									assign node200 = (inp[4]) ? 3'b101 : node201;
										assign node201 = (inp[5]) ? 3'b101 : 3'b011;
									assign node205 = (inp[4]) ? 3'b001 : node206;
										assign node206 = (inp[5]) ? node208 : 3'b101;
											assign node208 = (inp[0]) ? 3'b001 : 3'b101;
							assign node212 = (inp[1]) ? node218 : node213;
								assign node213 = (inp[8]) ? node215 : 3'b101;
									assign node215 = (inp[3]) ? 3'b001 : 3'b101;
								assign node218 = (inp[3]) ? node226 : node219;
									assign node219 = (inp[8]) ? 3'b101 : node220;
										assign node220 = (inp[0]) ? node222 : 3'b011;
											assign node222 = (inp[5]) ? 3'b101 : 3'b011;
									assign node226 = (inp[4]) ? node228 : 3'b101;
										assign node228 = (inp[8]) ? 3'b001 : 3'b101;
						assign node231 = (inp[3]) ? node241 : node232;
							assign node232 = (inp[8]) ? 3'b001 : node233;
								assign node233 = (inp[5]) ? node235 : 3'b101;
									assign node235 = (inp[0]) ? node237 : 3'b101;
										assign node237 = (inp[4]) ? 3'b001 : 3'b101;
							assign node241 = (inp[8]) ? node243 : 3'b001;
								assign node243 = (inp[5]) ? node251 : node244;
									assign node244 = (inp[4]) ? 3'b110 : node245;
										assign node245 = (inp[2]) ? node247 : 3'b001;
											assign node247 = (inp[1]) ? 3'b001 : 3'b110;
									assign node251 = (inp[0]) ? 3'b110 : node252;
										assign node252 = (inp[2]) ? 3'b110 : node253;
											assign node253 = (inp[1]) ? 3'b110 : 3'b001;
					assign node258 = (inp[11]) ? node294 : node259;
						assign node259 = (inp[3]) ? node275 : node260;
							assign node260 = (inp[4]) ? node268 : node261;
								assign node261 = (inp[8]) ? 3'b001 : node262;
									assign node262 = (inp[5]) ? node264 : 3'b101;
										assign node264 = (inp[2]) ? 3'b101 : 3'b001;
								assign node268 = (inp[8]) ? node270 : 3'b001;
									assign node270 = (inp[0]) ? 3'b110 : node271;
										assign node271 = (inp[5]) ? 3'b110 : 3'b001;
							assign node275 = (inp[8]) ? node287 : node276;
								assign node276 = (inp[4]) ? node278 : 3'b001;
									assign node278 = (inp[1]) ? 3'b110 : node279;
										assign node279 = (inp[5]) ? node283 : node280;
											assign node280 = (inp[0]) ? 3'b111 : 3'b001;
											assign node283 = (inp[0]) ? 3'b110 : 3'b111;
								assign node287 = (inp[0]) ? node289 : 3'b110;
									assign node289 = (inp[5]) ? node291 : 3'b110;
										assign node291 = (inp[2]) ? 3'b110 : 3'b010;
						assign node294 = (inp[0]) ? node318 : node295;
							assign node295 = (inp[8]) ? node309 : node296;
								assign node296 = (inp[3]) ? node304 : node297;
									assign node297 = (inp[4]) ? 3'b110 : node298;
										assign node298 = (inp[5]) ? node300 : 3'b001;
											assign node300 = (inp[1]) ? 3'b110 : 3'b001;
									assign node304 = (inp[4]) ? node306 : 3'b110;
										assign node306 = (inp[5]) ? 3'b010 : 3'b110;
								assign node309 = (inp[3]) ? 3'b010 : node310;
									assign node310 = (inp[1]) ? node314 : node311;
										assign node311 = (inp[2]) ? 3'b110 : 3'b010;
										assign node314 = (inp[2]) ? 3'b010 : 3'b110;
							assign node318 = (inp[4]) ? node330 : node319;
								assign node319 = (inp[2]) ? node325 : node320;
									assign node320 = (inp[8]) ? node322 : 3'b110;
										assign node322 = (inp[3]) ? 3'b100 : 3'b110;
									assign node325 = (inp[1]) ? node327 : 3'b110;
										assign node327 = (inp[8]) ? 3'b010 : 3'b110;
								assign node330 = (inp[3]) ? node336 : node331;
									assign node331 = (inp[8]) ? node333 : 3'b110;
										assign node333 = (inp[1]) ? 3'b010 : 3'b110;
									assign node336 = (inp[8]) ? node338 : 3'b010;
										assign node338 = (inp[5]) ? 3'b100 : 3'b010;
				assign node341 = (inp[7]) ? node381 : node342;
					assign node342 = (inp[8]) ? node360 : node343;
						assign node343 = (inp[11]) ? node353 : node344;
							assign node344 = (inp[3]) ? 3'b110 : node345;
								assign node345 = (inp[4]) ? node347 : 3'b001;
									assign node347 = (inp[5]) ? node349 : 3'b001;
										assign node349 = (inp[0]) ? 3'b110 : 3'b001;
							assign node353 = (inp[3]) ? 3'b010 : node354;
								assign node354 = (inp[4]) ? node356 : 3'b110;
									assign node356 = (inp[2]) ? 3'b010 : 3'b110;
						assign node360 = (inp[11]) ? node372 : node361;
							assign node361 = (inp[3]) ? node363 : 3'b110;
								assign node363 = (inp[4]) ? 3'b010 : node364;
									assign node364 = (inp[5]) ? 3'b010 : node365;
										assign node365 = (inp[2]) ? node367 : 3'b110;
											assign node367 = (inp[0]) ? 3'b010 : 3'b110;
							assign node372 = (inp[3]) ? node374 : 3'b010;
								assign node374 = (inp[0]) ? 3'b100 : node375;
									assign node375 = (inp[4]) ? 3'b100 : node376;
										assign node376 = (inp[5]) ? 3'b100 : 3'b010;
					assign node381 = (inp[11]) ? node413 : node382;
						assign node382 = (inp[8]) ? node392 : node383;
							assign node383 = (inp[3]) ? node385 : 3'b010;
								assign node385 = (inp[4]) ? node387 : 3'b010;
									assign node387 = (inp[2]) ? 3'b100 : node388;
										assign node388 = (inp[5]) ? 3'b100 : 3'b010;
							assign node392 = (inp[3]) ? node406 : node393;
								assign node393 = (inp[4]) ? node399 : node394;
									assign node394 = (inp[1]) ? 3'b010 : node395;
										assign node395 = (inp[5]) ? 3'b100 : 3'b010;
									assign node399 = (inp[5]) ? 3'b100 : node400;
										assign node400 = (inp[1]) ? 3'b100 : node401;
											assign node401 = (inp[2]) ? 3'b100 : 3'b010;
								assign node406 = (inp[4]) ? node408 : 3'b100;
									assign node408 = (inp[0]) ? node410 : 3'b100;
										assign node410 = (inp[5]) ? 3'b000 : 3'b100;
						assign node413 = (inp[3]) ? node429 : node414;
							assign node414 = (inp[8]) ? node422 : node415;
								assign node415 = (inp[4]) ? 3'b100 : node416;
									assign node416 = (inp[5]) ? 3'b100 : node417;
										assign node417 = (inp[0]) ? 3'b100 : 3'b010;
								assign node422 = (inp[4]) ? 3'b000 : node423;
									assign node423 = (inp[0]) ? node425 : 3'b100;
										assign node425 = (inp[2]) ? 3'b000 : 3'b100;
							assign node429 = (inp[8]) ? 3'b000 : node430;
								assign node430 = (inp[1]) ? 3'b000 : node431;
									assign node431 = (inp[5]) ? node433 : 3'b100;
										assign node433 = (inp[4]) ? 3'b000 : 3'b100;
		assign node438 = (inp[6]) ? node604 : node439;
			assign node439 = (inp[10]) ? node541 : node440;
				assign node440 = (inp[7]) ? node472 : node441;
					assign node441 = (inp[11]) ? node459 : node442;
						assign node442 = (inp[8]) ? node450 : node443;
							assign node443 = (inp[3]) ? 3'b001 : node444;
								assign node444 = (inp[4]) ? node446 : 3'b101;
									assign node446 = (inp[5]) ? 3'b001 : 3'b101;
							assign node450 = (inp[3]) ? node452 : 3'b001;
								assign node452 = (inp[0]) ? 3'b110 : node453;
									assign node453 = (inp[4]) ? 3'b110 : node454;
										assign node454 = (inp[5]) ? 3'b110 : 3'b001;
						assign node459 = (inp[3]) ? node469 : node460;
							assign node460 = (inp[8]) ? 3'b110 : node461;
								assign node461 = (inp[4]) ? node463 : 3'b001;
									assign node463 = (inp[5]) ? 3'b110 : node464;
										assign node464 = (inp[0]) ? 3'b110 : 3'b001;
							assign node469 = (inp[8]) ? 3'b010 : 3'b110;
					assign node472 = (inp[11]) ? node510 : node473;
						assign node473 = (inp[8]) ? node489 : node474;
							assign node474 = (inp[3]) ? node482 : node475;
								assign node475 = (inp[4]) ? 3'b110 : node476;
									assign node476 = (inp[0]) ? 3'b110 : node477;
										assign node477 = (inp[5]) ? 3'b110 : 3'b001;
								assign node482 = (inp[2]) ? 3'b110 : node483;
									assign node483 = (inp[4]) ? 3'b010 : node484;
										assign node484 = (inp[1]) ? 3'b010 : 3'b110;
							assign node489 = (inp[4]) ? node497 : node490;
								assign node490 = (inp[3]) ? 3'b010 : node491;
									assign node491 = (inp[0]) ? node493 : 3'b110;
										assign node493 = (inp[5]) ? 3'b010 : 3'b110;
								assign node497 = (inp[3]) ? node499 : 3'b010;
									assign node499 = (inp[5]) ? node505 : node500;
										assign node500 = (inp[0]) ? node502 : 3'b010;
											assign node502 = (inp[2]) ? 3'b100 : 3'b010;
										assign node505 = (inp[2]) ? 3'b100 : node506;
											assign node506 = (inp[0]) ? 3'b100 : 3'b010;
						assign node510 = (inp[8]) ? node522 : node511;
							assign node511 = (inp[3]) ? node515 : node512;
								assign node512 = (inp[4]) ? 3'b010 : 3'b110;
								assign node515 = (inp[4]) ? 3'b100 : node516;
									assign node516 = (inp[0]) ? node518 : 3'b010;
										assign node518 = (inp[5]) ? 3'b100 : 3'b010;
							assign node522 = (inp[4]) ? node532 : node523;
								assign node523 = (inp[3]) ? 3'b100 : node524;
									assign node524 = (inp[1]) ? 3'b010 : node525;
										assign node525 = (inp[2]) ? node527 : 3'b100;
											assign node527 = (inp[5]) ? 3'b000 : 3'b010;
								assign node532 = (inp[3]) ? node534 : 3'b100;
									assign node534 = (inp[0]) ? 3'b000 : node535;
										assign node535 = (inp[1]) ? node537 : 3'b100;
											assign node537 = (inp[2]) ? 3'b000 : 3'b100;
				assign node541 = (inp[7]) ? node585 : node542;
					assign node542 = (inp[11]) ? node558 : node543;
						assign node543 = (inp[8]) ? node551 : node544;
							assign node544 = (inp[3]) ? 3'b010 : node545;
								assign node545 = (inp[1]) ? node547 : 3'b110;
									assign node547 = (inp[4]) ? 3'b010 : 3'b110;
							assign node551 = (inp[3]) ? 3'b100 : node552;
								assign node552 = (inp[2]) ? node554 : 3'b010;
									assign node554 = (inp[1]) ? 3'b010 : 3'b100;
						assign node558 = (inp[8]) ? node572 : node559;
							assign node559 = (inp[3]) ? 3'b100 : node560;
								assign node560 = (inp[4]) ? node566 : node561;
									assign node561 = (inp[5]) ? node563 : 3'b000;
										assign node563 = (inp[0]) ? 3'b100 : 3'b000;
									assign node566 = (inp[2]) ? 3'b100 : node567;
										assign node567 = (inp[5]) ? 3'b100 : 3'b000;
							assign node572 = (inp[3]) ? node578 : node573;
								assign node573 = (inp[2]) ? node575 : 3'b100;
									assign node575 = (inp[1]) ? 3'b100 : 3'b000;
								assign node578 = (inp[5]) ? 3'b000 : node579;
									assign node579 = (inp[0]) ? 3'b000 : node580;
										assign node580 = (inp[4]) ? 3'b000 : 3'b100;
					assign node585 = (inp[11]) ? 3'b000 : node586;
						assign node586 = (inp[8]) ? node596 : node587;
							assign node587 = (inp[3]) ? node589 : 3'b100;
								assign node589 = (inp[4]) ? 3'b000 : node590;
									assign node590 = (inp[0]) ? node592 : 3'b100;
										assign node592 = (inp[5]) ? 3'b000 : 3'b100;
							assign node596 = (inp[0]) ? 3'b000 : node597;
								assign node597 = (inp[5]) ? 3'b000 : node598;
									assign node598 = (inp[4]) ? 3'b000 : 3'b100;
			assign node604 = (inp[10]) ? 3'b000 : node605;
				assign node605 = (inp[7]) ? 3'b000 : node606;
					assign node606 = (inp[11]) ? node634 : node607;
						assign node607 = (inp[8]) ? node615 : node608;
							assign node608 = (inp[3]) ? 3'b100 : node609;
								assign node609 = (inp[1]) ? node611 : 3'b010;
									assign node611 = (inp[4]) ? 3'b100 : 3'b010;
							assign node615 = (inp[3]) ? node625 : node616;
								assign node616 = (inp[2]) ? node618 : 3'b100;
									assign node618 = (inp[1]) ? node620 : 3'b000;
										assign node620 = (inp[4]) ? node622 : 3'b100;
											assign node622 = (inp[5]) ? 3'b000 : 3'b100;
								assign node625 = (inp[1]) ? node627 : 3'b000;
									assign node627 = (inp[0]) ? 3'b000 : node628;
										assign node628 = (inp[4]) ? 3'b000 : node629;
											assign node629 = (inp[5]) ? 3'b000 : 3'b100;
						assign node634 = (inp[3]) ? 3'b000 : node635;
							assign node635 = (inp[8]) ? 3'b000 : node636;
								assign node636 = (inp[2]) ? node638 : 3'b100;
									assign node638 = (inp[4]) ? 3'b000 : 3'b100;

endmodule