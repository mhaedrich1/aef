module dtc_split75_bm5 (
	input  wire [10-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node6;
	wire [1-1:0] node7;
	wire [1-1:0] node8;
	wire [1-1:0] node9;
	wire [1-1:0] node14;
	wire [1-1:0] node15;
	wire [1-1:0] node19;
	wire [1-1:0] node20;
	wire [1-1:0] node21;
	wire [1-1:0] node22;
	wire [1-1:0] node25;
	wire [1-1:0] node29;
	wire [1-1:0] node30;
	wire [1-1:0] node33;
	wire [1-1:0] node36;
	wire [1-1:0] node37;
	wire [1-1:0] node38;
	wire [1-1:0] node41;
	wire [1-1:0] node43;
	wire [1-1:0] node46;
	wire [1-1:0] node47;
	wire [1-1:0] node48;
	wire [1-1:0] node52;
	wire [1-1:0] node53;
	wire [1-1:0] node56;
	wire [1-1:0] node59;
	wire [1-1:0] node60;
	wire [1-1:0] node61;
	wire [1-1:0] node62;
	wire [1-1:0] node63;
	wire [1-1:0] node65;
	wire [1-1:0] node69;
	wire [1-1:0] node70;
	wire [1-1:0] node73;
	wire [1-1:0] node76;
	wire [1-1:0] node77;
	wire [1-1:0] node78;
	wire [1-1:0] node83;
	wire [1-1:0] node84;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node90;
	wire [1-1:0] node91;
	wire [1-1:0] node94;
	wire [1-1:0] node97;
	wire [1-1:0] node98;
	wire [1-1:0] node99;
	wire [1-1:0] node103;
	wire [1-1:0] node104;
	wire [1-1:0] node107;
	wire [1-1:0] node110;
	wire [1-1:0] node111;
	wire [1-1:0] node112;
	wire [1-1:0] node114;
	wire [1-1:0] node118;
	wire [1-1:0] node119;
	wire [1-1:0] node121;
	wire [1-1:0] node122;
	wire [1-1:0] node126;
	wire [1-1:0] node127;
	wire [1-1:0] node128;
	wire [1-1:0] node130;
	wire [1-1:0] node133;
	wire [1-1:0] node134;
	wire [1-1:0] node138;
	wire [1-1:0] node140;
	wire [1-1:0] node142;
	wire [1-1:0] node145;
	wire [1-1:0] node146;
	wire [1-1:0] node147;
	wire [1-1:0] node148;
	wire [1-1:0] node149;
	wire [1-1:0] node150;
	wire [1-1:0] node151;
	wire [1-1:0] node153;
	wire [1-1:0] node156;
	wire [1-1:0] node160;
	wire [1-1:0] node161;
	wire [1-1:0] node163;
	wire [1-1:0] node167;
	wire [1-1:0] node168;
	wire [1-1:0] node169;
	wire [1-1:0] node170;
	wire [1-1:0] node173;
	wire [1-1:0] node174;
	wire [1-1:0] node179;
	wire [1-1:0] node180;
	wire [1-1:0] node181;
	wire [1-1:0] node184;
	wire [1-1:0] node185;
	wire [1-1:0] node190;
	wire [1-1:0] node191;
	wire [1-1:0] node192;
	wire [1-1:0] node193;
	wire [1-1:0] node194;
	wire [1-1:0] node198;
	wire [1-1:0] node200;
	wire [1-1:0] node201;
	wire [1-1:0] node204;
	wire [1-1:0] node207;
	wire [1-1:0] node208;
	wire [1-1:0] node209;
	wire [1-1:0] node212;
	wire [1-1:0] node214;
	wire [1-1:0] node217;
	wire [1-1:0] node218;
	wire [1-1:0] node219;
	wire [1-1:0] node222;
	wire [1-1:0] node225;
	wire [1-1:0] node226;
	wire [1-1:0] node229;
	wire [1-1:0] node232;
	wire [1-1:0] node233;
	wire [1-1:0] node234;
	wire [1-1:0] node235;
	wire [1-1:0] node239;
	wire [1-1:0] node240;
	wire [1-1:0] node241;
	wire [1-1:0] node244;
	wire [1-1:0] node247;
	wire [1-1:0] node248;
	wire [1-1:0] node251;
	wire [1-1:0] node254;
	wire [1-1:0] node255;
	wire [1-1:0] node256;
	wire [1-1:0] node259;
	wire [1-1:0] node260;
	wire [1-1:0] node264;
	wire [1-1:0] node266;
	wire [1-1:0] node267;
	wire [1-1:0] node270;
	wire [1-1:0] node273;
	wire [1-1:0] node274;
	wire [1-1:0] node275;
	wire [1-1:0] node276;
	wire [1-1:0] node277;
	wire [1-1:0] node279;
	wire [1-1:0] node282;
	wire [1-1:0] node284;
	wire [1-1:0] node287;
	wire [1-1:0] node288;
	wire [1-1:0] node290;
	wire [1-1:0] node293;
	wire [1-1:0] node295;
	wire [1-1:0] node298;
	wire [1-1:0] node299;
	wire [1-1:0] node301;
	wire [1-1:0] node302;
	wire [1-1:0] node303;
	wire [1-1:0] node307;
	wire [1-1:0] node309;
	wire [1-1:0] node312;
	wire [1-1:0] node313;
	wire [1-1:0] node314;
	wire [1-1:0] node316;
	wire [1-1:0] node319;
	wire [1-1:0] node320;
	wire [1-1:0] node323;
	wire [1-1:0] node326;
	wire [1-1:0] node327;
	wire [1-1:0] node330;
	wire [1-1:0] node333;
	wire [1-1:0] node335;
	wire [1-1:0] node337;
	wire [1-1:0] node338;
	wire [1-1:0] node342;
	wire [1-1:0] node343;
	wire [1-1:0] node344;
	wire [1-1:0] node345;
	wire [1-1:0] node346;
	wire [1-1:0] node348;
	wire [1-1:0] node351;
	wire [1-1:0] node352;
	wire [1-1:0] node353;
	wire [1-1:0] node355;
	wire [1-1:0] node359;
	wire [1-1:0] node360;
	wire [1-1:0] node363;
	wire [1-1:0] node366;
	wire [1-1:0] node367;
	wire [1-1:0] node368;
	wire [1-1:0] node370;
	wire [1-1:0] node371;
	wire [1-1:0] node372;
	wire [1-1:0] node377;
	wire [1-1:0] node378;
	wire [1-1:0] node379;
	wire [1-1:0] node380;
	wire [1-1:0] node385;
	wire [1-1:0] node386;
	wire [1-1:0] node390;
	wire [1-1:0] node391;
	wire [1-1:0] node393;
	wire [1-1:0] node396;
	wire [1-1:0] node397;
	wire [1-1:0] node400;
	wire [1-1:0] node403;
	wire [1-1:0] node404;
	wire [1-1:0] node405;
	wire [1-1:0] node407;
	wire [1-1:0] node410;
	wire [1-1:0] node413;
	wire [1-1:0] node414;
	wire [1-1:0] node415;
	wire [1-1:0] node416;
	wire [1-1:0] node420;
	wire [1-1:0] node421;
	wire [1-1:0] node423;
	wire [1-1:0] node424;
	wire [1-1:0] node427;
	wire [1-1:0] node430;
	wire [1-1:0] node431;
	wire [1-1:0] node434;
	wire [1-1:0] node437;
	wire [1-1:0] node438;
	wire [1-1:0] node439;
	wire [1-1:0] node443;
	wire [1-1:0] node444;
	wire [1-1:0] node446;
	wire [1-1:0] node449;
	wire [1-1:0] node451;
	wire [1-1:0] node454;
	wire [1-1:0] node455;
	wire [1-1:0] node456;
	wire [1-1:0] node458;
	wire [1-1:0] node459;
	wire [1-1:0] node463;
	wire [1-1:0] node464;
	wire [1-1:0] node467;
	wire [1-1:0] node469;
	wire [1-1:0] node472;
	wire [1-1:0] node473;
	wire [1-1:0] node474;
	wire [1-1:0] node475;
	wire [1-1:0] node477;
	wire [1-1:0] node481;
	wire [1-1:0] node482;
	wire [1-1:0] node485;
	wire [1-1:0] node487;
	wire [1-1:0] node490;
	wire [1-1:0] node491;
	wire [1-1:0] node492;
	wire [1-1:0] node493;
	wire [1-1:0] node494;
	wire [1-1:0] node496;
	wire [1-1:0] node499;
	wire [1-1:0] node502;
	wire [1-1:0] node504;
	wire [1-1:0] node506;
	wire [1-1:0] node509;
	wire [1-1:0] node511;
	wire [1-1:0] node513;
	wire [1-1:0] node514;
	wire [1-1:0] node517;
	wire [1-1:0] node520;
	wire [1-1:0] node521;
	wire [1-1:0] node523;

	assign outp = (inp[8]) ? node342 : node1;
		assign node1 = (inp[6]) ? node145 : node2;
			assign node2 = (inp[4]) ? node110 : node3;
				assign node3 = (inp[2]) ? node59 : node4;
					assign node4 = (inp[9]) ? node36 : node5;
						assign node5 = (inp[3]) ? node19 : node6;
							assign node6 = (inp[7]) ? node14 : node7;
								assign node7 = (inp[5]) ? 1'b0 : node8;
									assign node8 = (inp[0]) ? 1'b1 : node9;
										assign node9 = (inp[1]) ? 1'b0 : 1'b1;
								assign node14 = (inp[0]) ? 1'b0 : node15;
									assign node15 = (inp[1]) ? 1'b1 : 1'b0;
							assign node19 = (inp[7]) ? node29 : node20;
								assign node20 = (inp[1]) ? 1'b0 : node21;
									assign node21 = (inp[5]) ? node25 : node22;
										assign node22 = (inp[0]) ? 1'b0 : 1'b1;
										assign node25 = (inp[0]) ? 1'b1 : 1'b0;
								assign node29 = (inp[0]) ? node33 : node30;
									assign node30 = (inp[1]) ? 1'b1 : 1'b0;
									assign node33 = (inp[1]) ? 1'b0 : 1'b1;
						assign node36 = (inp[5]) ? node46 : node37;
							assign node37 = (inp[0]) ? node41 : node38;
								assign node38 = (inp[1]) ? 1'b1 : 1'b0;
								assign node41 = (inp[3]) ? node43 : 1'b0;
									assign node43 = (inp[1]) ? 1'b0 : 1'b1;
							assign node46 = (inp[3]) ? node52 : node47;
								assign node47 = (inp[0]) ? 1'b1 : node48;
									assign node48 = (inp[1]) ? 1'b0 : 1'b1;
								assign node52 = (inp[0]) ? node56 : node53;
									assign node53 = (inp[1]) ? 1'b0 : 1'b1;
									assign node56 = (inp[1]) ? 1'b1 : 1'b0;
					assign node59 = (inp[5]) ? node83 : node60;
						assign node60 = (inp[1]) ? node76 : node61;
							assign node61 = (inp[9]) ? node69 : node62;
								assign node62 = (inp[0]) ? 1'b1 : node63;
									assign node63 = (inp[7]) ? node65 : 1'b1;
										assign node65 = (inp[3]) ? 1'b1 : 1'b0;
								assign node69 = (inp[3]) ? node73 : node70;
									assign node70 = (inp[0]) ? 1'b1 : 1'b0;
									assign node73 = (inp[0]) ? 1'b0 : 1'b1;
							assign node76 = (inp[9]) ? 1'b1 : node77;
								assign node77 = (inp[7]) ? 1'b1 : node78;
									assign node78 = (inp[0]) ? 1'b0 : 1'b1;
						assign node83 = (inp[9]) ? node97 : node84;
							assign node84 = (inp[3]) ? node90 : node85;
								assign node85 = (inp[0]) ? 1'b1 : node86;
									assign node86 = (inp[1]) ? 1'b1 : 1'b0;
								assign node90 = (inp[0]) ? node94 : node91;
									assign node91 = (inp[1]) ? 1'b0 : 1'b1;
									assign node94 = (inp[1]) ? 1'b1 : 1'b0;
							assign node97 = (inp[3]) ? node103 : node98;
								assign node98 = (inp[0]) ? 1'b0 : node99;
									assign node99 = (inp[7]) ? 1'b0 : 1'b1;
								assign node103 = (inp[1]) ? node107 : node104;
									assign node104 = (inp[0]) ? 1'b1 : 1'b0;
									assign node107 = (inp[0]) ? 1'b0 : 1'b1;
				assign node110 = (inp[3]) ? node118 : node111;
					assign node111 = (inp[5]) ? 1'b1 : node112;
						assign node112 = (inp[9]) ? node114 : 1'b1;
							assign node114 = (inp[7]) ? 1'b0 : 1'b1;
					assign node118 = (inp[2]) ? node126 : node119;
						assign node119 = (inp[9]) ? node121 : 1'b1;
							assign node121 = (inp[5]) ? 1'b1 : node122;
								assign node122 = (inp[7]) ? 1'b0 : 1'b1;
						assign node126 = (inp[1]) ? node138 : node127;
							assign node127 = (inp[0]) ? node133 : node128;
								assign node128 = (inp[9]) ? node130 : 1'b0;
									assign node130 = (inp[7]) ? 1'b1 : 1'b0;
								assign node133 = (inp[5]) ? 1'b1 : node134;
									assign node134 = (inp[9]) ? 1'b0 : 1'b1;
							assign node138 = (inp[9]) ? node140 : 1'b0;
								assign node140 = (inp[7]) ? node142 : 1'b0;
									assign node142 = (inp[5]) ? 1'b0 : 1'b1;
			assign node145 = (inp[5]) ? node273 : node146;
				assign node146 = (inp[2]) ? node190 : node147;
					assign node147 = (inp[9]) ? node167 : node148;
						assign node148 = (inp[7]) ? node160 : node149;
							assign node149 = (inp[4]) ? 1'b1 : node150;
								assign node150 = (inp[1]) ? node156 : node151;
									assign node151 = (inp[0]) ? node153 : 1'b1;
										assign node153 = (inp[3]) ? 1'b0 : 1'b1;
									assign node156 = (inp[0]) ? 1'b1 : 1'b0;
							assign node160 = (inp[4]) ? 1'b0 : node161;
								assign node161 = (inp[3]) ? node163 : 1'b1;
									assign node163 = (inp[0]) ? 1'b0 : 1'b1;
						assign node167 = (inp[7]) ? node179 : node168;
							assign node168 = (inp[4]) ? 1'b0 : node169;
								assign node169 = (inp[0]) ? node173 : node170;
									assign node170 = (inp[1]) ? 1'b1 : 1'b0;
									assign node173 = (inp[1]) ? 1'b0 : node174;
										assign node174 = (inp[3]) ? 1'b1 : 1'b0;
							assign node179 = (inp[4]) ? 1'b1 : node180;
								assign node180 = (inp[3]) ? node184 : node181;
									assign node181 = (inp[0]) ? 1'b1 : 1'b0;
									assign node184 = (inp[1]) ? 1'b0 : node185;
										assign node185 = (inp[0]) ? 1'b0 : 1'b1;
					assign node190 = (inp[0]) ? node232 : node191;
						assign node191 = (inp[1]) ? node207 : node192;
							assign node192 = (inp[3]) ? node198 : node193;
								assign node193 = (inp[7]) ? 1'b1 : node194;
									assign node194 = (inp[9]) ? 1'b0 : 1'b1;
								assign node198 = (inp[4]) ? node200 : 1'b0;
									assign node200 = (inp[7]) ? node204 : node201;
										assign node201 = (inp[9]) ? 1'b1 : 1'b0;
										assign node204 = (inp[9]) ? 1'b0 : 1'b1;
							assign node207 = (inp[4]) ? node217 : node208;
								assign node208 = (inp[3]) ? node212 : node209;
									assign node209 = (inp[7]) ? 1'b0 : 1'b1;
									assign node212 = (inp[9]) ? node214 : 1'b1;
										assign node214 = (inp[7]) ? 1'b1 : 1'b0;
								assign node217 = (inp[7]) ? node225 : node218;
									assign node218 = (inp[3]) ? node222 : node219;
										assign node219 = (inp[9]) ? 1'b0 : 1'b1;
										assign node222 = (inp[9]) ? 1'b1 : 1'b0;
									assign node225 = (inp[3]) ? node229 : node226;
										assign node226 = (inp[9]) ? 1'b1 : 1'b0;
										assign node229 = (inp[9]) ? 1'b0 : 1'b1;
						assign node232 = (inp[3]) ? node254 : node233;
							assign node233 = (inp[9]) ? node239 : node234;
								assign node234 = (inp[7]) ? 1'b0 : node235;
									assign node235 = (inp[4]) ? 1'b1 : 1'b0;
								assign node239 = (inp[1]) ? node247 : node240;
									assign node240 = (inp[4]) ? node244 : node241;
										assign node241 = (inp[7]) ? 1'b0 : 1'b1;
										assign node244 = (inp[7]) ? 1'b1 : 1'b0;
									assign node247 = (inp[4]) ? node251 : node248;
										assign node248 = (inp[7]) ? 1'b0 : 1'b1;
										assign node251 = (inp[7]) ? 1'b1 : 1'b0;
							assign node254 = (inp[1]) ? node264 : node255;
								assign node255 = (inp[7]) ? node259 : node256;
									assign node256 = (inp[9]) ? 1'b0 : 1'b1;
									assign node259 = (inp[9]) ? 1'b1 : node260;
										assign node260 = (inp[4]) ? 1'b0 : 1'b1;
								assign node264 = (inp[4]) ? node266 : 1'b0;
									assign node266 = (inp[7]) ? node270 : node267;
										assign node267 = (inp[9]) ? 1'b1 : 1'b0;
										assign node270 = (inp[9]) ? 1'b0 : 1'b1;
				assign node273 = (inp[4]) ? node333 : node274;
					assign node274 = (inp[3]) ? node298 : node275;
						assign node275 = (inp[7]) ? node287 : node276;
							assign node276 = (inp[1]) ? node282 : node277;
								assign node277 = (inp[2]) ? node279 : 1'b1;
									assign node279 = (inp[0]) ? 1'b0 : 1'b1;
								assign node282 = (inp[0]) ? node284 : 1'b0;
									assign node284 = (inp[2]) ? 1'b0 : 1'b1;
							assign node287 = (inp[1]) ? node293 : node288;
								assign node288 = (inp[2]) ? node290 : 1'b0;
									assign node290 = (inp[0]) ? 1'b1 : 1'b0;
								assign node293 = (inp[0]) ? node295 : 1'b1;
									assign node295 = (inp[2]) ? 1'b1 : 1'b0;
						assign node298 = (inp[0]) ? node312 : node299;
							assign node299 = (inp[2]) ? node301 : 1'b0;
								assign node301 = (inp[9]) ? node307 : node302;
									assign node302 = (inp[7]) ? 1'b0 : node303;
										assign node303 = (inp[1]) ? 1'b1 : 1'b0;
									assign node307 = (inp[7]) ? node309 : 1'b0;
										assign node309 = (inp[1]) ? 1'b0 : 1'b1;
							assign node312 = (inp[1]) ? node326 : node313;
								assign node313 = (inp[9]) ? node319 : node314;
									assign node314 = (inp[2]) ? node316 : 1'b0;
										assign node316 = (inp[7]) ? 1'b0 : 1'b1;
									assign node319 = (inp[7]) ? node323 : node320;
										assign node320 = (inp[2]) ? 1'b1 : 1'b0;
										assign node323 = (inp[2]) ? 1'b0 : 1'b1;
								assign node326 = (inp[7]) ? node330 : node327;
									assign node327 = (inp[2]) ? 1'b0 : 1'b1;
									assign node330 = (inp[2]) ? 1'b1 : 1'b0;
					assign node333 = (inp[3]) ? node335 : 1'b0;
						assign node335 = (inp[2]) ? node337 : 1'b0;
							assign node337 = (inp[1]) ? 1'b1 : node338;
								assign node338 = (inp[0]) ? 1'b0 : 1'b1;
		assign node342 = (inp[4]) ? node454 : node343;
			assign node343 = (inp[1]) ? node403 : node344;
				assign node344 = (inp[6]) ? node366 : node345;
					assign node345 = (inp[3]) ? node351 : node346;
						assign node346 = (inp[2]) ? node348 : 1'b1;
							assign node348 = (inp[0]) ? 1'b0 : 1'b1;
						assign node351 = (inp[7]) ? node359 : node352;
							assign node352 = (inp[5]) ? 1'b0 : node353;
								assign node353 = (inp[0]) ? node355 : 1'b1;
									assign node355 = (inp[2]) ? 1'b1 : 1'b0;
							assign node359 = (inp[2]) ? node363 : node360;
								assign node360 = (inp[0]) ? 1'b0 : 1'b1;
								assign node363 = (inp[0]) ? 1'b1 : 1'b0;
					assign node366 = (inp[7]) ? node390 : node367;
						assign node367 = (inp[0]) ? node377 : node368;
							assign node368 = (inp[3]) ? node370 : 1'b1;
								assign node370 = (inp[2]) ? 1'b0 : node371;
									assign node371 = (inp[5]) ? 1'b1 : node372;
										assign node372 = (inp[9]) ? 1'b1 : 1'b0;
							assign node377 = (inp[3]) ? node385 : node378;
								assign node378 = (inp[5]) ? 1'b0 : node379;
									assign node379 = (inp[9]) ? 1'b0 : node380;
										assign node380 = (inp[2]) ? 1'b1 : 1'b0;
								assign node385 = (inp[2]) ? 1'b1 : node386;
									assign node386 = (inp[5]) ? 1'b0 : 1'b1;
						assign node390 = (inp[3]) ? node396 : node391;
							assign node391 = (inp[0]) ? node393 : 1'b0;
								assign node393 = (inp[2]) ? 1'b1 : 1'b0;
							assign node396 = (inp[0]) ? node400 : node397;
								assign node397 = (inp[2]) ? 1'b1 : 1'b0;
								assign node400 = (inp[2]) ? 1'b0 : 1'b1;
				assign node403 = (inp[6]) ? node413 : node404;
					assign node404 = (inp[0]) ? node410 : node405;
						assign node405 = (inp[3]) ? node407 : 1'b0;
							assign node407 = (inp[2]) ? 1'b1 : 1'b0;
						assign node410 = (inp[2]) ? 1'b0 : 1'b1;
					assign node413 = (inp[7]) ? node437 : node414;
						assign node414 = (inp[3]) ? node420 : node415;
							assign node415 = (inp[5]) ? 1'b0 : node416;
								assign node416 = (inp[9]) ? 1'b0 : 1'b1;
							assign node420 = (inp[9]) ? node430 : node421;
								assign node421 = (inp[0]) ? node423 : 1'b0;
									assign node423 = (inp[2]) ? node427 : node424;
										assign node424 = (inp[5]) ? 1'b1 : 1'b0;
										assign node427 = (inp[5]) ? 1'b0 : 1'b1;
								assign node430 = (inp[0]) ? node434 : node431;
									assign node431 = (inp[2]) ? 1'b1 : 1'b0;
									assign node434 = (inp[2]) ? 1'b0 : 1'b1;
						assign node437 = (inp[3]) ? node443 : node438;
							assign node438 = (inp[2]) ? 1'b1 : node439;
								assign node439 = (inp[0]) ? 1'b0 : 1'b1;
							assign node443 = (inp[5]) ? node449 : node444;
								assign node444 = (inp[2]) ? node446 : 1'b0;
									assign node446 = (inp[0]) ? 1'b1 : 1'b0;
								assign node449 = (inp[0]) ? node451 : 1'b1;
									assign node451 = (inp[2]) ? 1'b1 : 1'b0;
			assign node454 = (inp[3]) ? node472 : node455;
				assign node455 = (inp[6]) ? node463 : node456;
					assign node456 = (inp[7]) ? node458 : 1'b0;
						assign node458 = (inp[5]) ? 1'b0 : node459;
							assign node459 = (inp[9]) ? 1'b0 : 1'b1;
					assign node463 = (inp[9]) ? node467 : node464;
						assign node464 = (inp[7]) ? 1'b0 : 1'b1;
						assign node467 = (inp[7]) ? node469 : 1'b0;
							assign node469 = (inp[5]) ? 1'b1 : 1'b0;
				assign node472 = (inp[2]) ? node490 : node473;
					assign node473 = (inp[6]) ? node481 : node474;
						assign node474 = (inp[5]) ? 1'b0 : node475;
							assign node475 = (inp[7]) ? node477 : 1'b0;
								assign node477 = (inp[9]) ? 1'b0 : 1'b1;
						assign node481 = (inp[9]) ? node485 : node482;
							assign node482 = (inp[7]) ? 1'b0 : 1'b1;
							assign node485 = (inp[7]) ? node487 : 1'b0;
								assign node487 = (inp[5]) ? 1'b1 : 1'b0;
					assign node490 = (inp[1]) ? node520 : node491;
						assign node491 = (inp[0]) ? node509 : node492;
							assign node492 = (inp[9]) ? node502 : node493;
								assign node493 = (inp[6]) ? node499 : node494;
									assign node494 = (inp[7]) ? node496 : 1'b1;
										assign node496 = (inp[5]) ? 1'b1 : 1'b0;
									assign node499 = (inp[7]) ? 1'b1 : 1'b0;
								assign node502 = (inp[6]) ? node504 : 1'b1;
									assign node504 = (inp[7]) ? node506 : 1'b1;
										assign node506 = (inp[5]) ? 1'b0 : 1'b1;
							assign node509 = (inp[6]) ? node511 : 1'b0;
								assign node511 = (inp[5]) ? node513 : 1'b0;
									assign node513 = (inp[7]) ? node517 : node514;
										assign node514 = (inp[9]) ? 1'b0 : 1'b1;
										assign node517 = (inp[9]) ? 1'b1 : 1'b0;
						assign node520 = (inp[9]) ? 1'b1 : node521;
							assign node521 = (inp[6]) ? node523 : 1'b1;
								assign node523 = (inp[7]) ? 1'b1 : 1'b0;

endmodule