module dtc_split66_bm79 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node125;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node177;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node229;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node266;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node290;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node312;
	wire [3-1:0] node316;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node339;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node344;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node363;
	wire [3-1:0] node365;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node375;
	wire [3-1:0] node377;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node396;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node409;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node419;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node430;
	wire [3-1:0] node432;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node444;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node451;
	wire [3-1:0] node453;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node459;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node466;
	wire [3-1:0] node468;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node480;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node487;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node528;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node535;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node541;
	wire [3-1:0] node543;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node554;
	wire [3-1:0] node558;
	wire [3-1:0] node560;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node566;
	wire [3-1:0] node568;
	wire [3-1:0] node571;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node583;
	wire [3-1:0] node586;
	wire [3-1:0] node588;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node594;
	wire [3-1:0] node597;
	wire [3-1:0] node599;
	wire [3-1:0] node601;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node609;
	wire [3-1:0] node612;
	wire [3-1:0] node613;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node626;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node639;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node650;
	wire [3-1:0] node652;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node658;
	wire [3-1:0] node660;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node669;
	wire [3-1:0] node671;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node683;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node694;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node711;
	wire [3-1:0] node713;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node723;
	wire [3-1:0] node725;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node735;
	wire [3-1:0] node737;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node744;
	wire [3-1:0] node746;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node758;
	wire [3-1:0] node760;
	wire [3-1:0] node761;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node773;
	wire [3-1:0] node775;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node787;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node794;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node802;
	wire [3-1:0] node805;
	wire [3-1:0] node807;
	wire [3-1:0] node810;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node825;
	wire [3-1:0] node827;
	wire [3-1:0] node829;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node839;
	wire [3-1:0] node843;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node855;
	wire [3-1:0] node858;
	wire [3-1:0] node861;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node869;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node897;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node913;
	wire [3-1:0] node915;
	wire [3-1:0] node916;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node930;
	wire [3-1:0] node934;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node938;
	wire [3-1:0] node939;
	wire [3-1:0] node944;
	wire [3-1:0] node945;
	wire [3-1:0] node947;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node961;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node966;
	wire [3-1:0] node970;
	wire [3-1:0] node971;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node976;
	wire [3-1:0] node980;
	wire [3-1:0] node982;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node988;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node995;
	wire [3-1:0] node999;
	wire [3-1:0] node1000;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1011;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1015;
	wire [3-1:0] node1016;
	wire [3-1:0] node1020;
	wire [3-1:0] node1026;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1031;
	wire [3-1:0] node1034;
	wire [3-1:0] node1035;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1043;
	wire [3-1:0] node1045;
	wire [3-1:0] node1048;
	wire [3-1:0] node1049;
	wire [3-1:0] node1050;
	wire [3-1:0] node1051;
	wire [3-1:0] node1053;
	wire [3-1:0] node1057;
	wire [3-1:0] node1060;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1064;
	wire [3-1:0] node1068;
	wire [3-1:0] node1069;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1077;
	wire [3-1:0] node1078;
	wire [3-1:0] node1080;
	wire [3-1:0] node1084;
	wire [3-1:0] node1086;
	wire [3-1:0] node1089;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1095;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1109;
	wire [3-1:0] node1110;

	assign outp = (inp[6]) ? node322 : node1;
		assign node1 = (inp[9]) ? node295 : node2;
			assign node2 = (inp[0]) ? node220 : node3;
				assign node3 = (inp[7]) ? node91 : node4;
					assign node4 = (inp[10]) ? node64 : node5;
						assign node5 = (inp[1]) ? node43 : node6;
							assign node6 = (inp[11]) ? node22 : node7;
								assign node7 = (inp[2]) ? node15 : node8;
									assign node8 = (inp[3]) ? 3'b110 : node9;
										assign node9 = (inp[4]) ? 3'b110 : node10;
											assign node10 = (inp[5]) ? 3'b110 : 3'b010;
									assign node15 = (inp[3]) ? 3'b010 : node16;
										assign node16 = (inp[8]) ? 3'b110 : node17;
											assign node17 = (inp[4]) ? 3'b010 : 3'b110;
								assign node22 = (inp[8]) ? node36 : node23;
									assign node23 = (inp[2]) ? node29 : node24;
										assign node24 = (inp[5]) ? node26 : 3'b100;
											assign node26 = (inp[3]) ? 3'b100 : 3'b110;
										assign node29 = (inp[3]) ? 3'b000 : node30;
											assign node30 = (inp[4]) ? node32 : 3'b100;
												assign node32 = (inp[5]) ? 3'b000 : 3'b100;
									assign node36 = (inp[4]) ? 3'b010 : node37;
										assign node37 = (inp[2]) ? 3'b010 : node38;
											assign node38 = (inp[3]) ? 3'b010 : 3'b110;
							assign node43 = (inp[11]) ? node55 : node44;
								assign node44 = (inp[8]) ? node50 : node45;
									assign node45 = (inp[2]) ? node47 : 3'b100;
										assign node47 = (inp[3]) ? 3'b000 : 3'b100;
									assign node50 = (inp[3]) ? node52 : 3'b010;
										assign node52 = (inp[2]) ? 3'b100 : 3'b010;
								assign node55 = (inp[8]) ? node57 : 3'b000;
									assign node57 = (inp[2]) ? node59 : 3'b100;
										assign node59 = (inp[5]) ? 3'b000 : node60;
											assign node60 = (inp[3]) ? 3'b000 : 3'b100;
						assign node64 = (inp[1]) ? 3'b000 : node65;
							assign node65 = (inp[8]) ? node67 : 3'b000;
								assign node67 = (inp[11]) ? node83 : node68;
									assign node68 = (inp[3]) ? node76 : node69;
										assign node69 = (inp[2]) ? 3'b100 : node70;
											assign node70 = (inp[4]) ? node72 : 3'b000;
												assign node72 = (inp[5]) ? 3'b100 : 3'b000;
										assign node76 = (inp[5]) ? node78 : 3'b100;
											assign node78 = (inp[2]) ? node80 : 3'b100;
												assign node80 = (inp[4]) ? 3'b000 : 3'b100;
									assign node83 = (inp[3]) ? 3'b000 : node84;
										assign node84 = (inp[5]) ? node86 : 3'b100;
											assign node86 = (inp[4]) ? 3'b000 : 3'b100;
					assign node91 = (inp[10]) ? node153 : node92;
						assign node92 = (inp[8]) ? node130 : node93;
							assign node93 = (inp[1]) ? node117 : node94;
								assign node94 = (inp[11]) ? node106 : node95;
									assign node95 = (inp[2]) ? node101 : node96;
										assign node96 = (inp[4]) ? 3'b001 : node97;
											assign node97 = (inp[3]) ? 3'b001 : 3'b101;
										assign node101 = (inp[4]) ? node103 : 3'b001;
											assign node103 = (inp[5]) ? 3'b001 : 3'b110;
									assign node106 = (inp[2]) ? node112 : node107;
										assign node107 = (inp[3]) ? 3'b110 : node108;
											assign node108 = (inp[4]) ? 3'b110 : 3'b001;
										assign node112 = (inp[4]) ? node114 : 3'b110;
											assign node114 = (inp[3]) ? 3'b010 : 3'b110;
								assign node117 = (inp[11]) ? node125 : node118;
									assign node118 = (inp[2]) ? node120 : 3'b110;
										assign node120 = (inp[5]) ? 3'b010 : node121;
											assign node121 = (inp[4]) ? 3'b010 : 3'b110;
									assign node125 = (inp[2]) ? node127 : 3'b010;
										assign node127 = (inp[3]) ? 3'b100 : 3'b010;
							assign node130 = (inp[1]) ? node138 : node131;
								assign node131 = (inp[11]) ? node133 : 3'b101;
									assign node133 = (inp[3]) ? 3'b001 : node134;
										assign node134 = (inp[2]) ? 3'b001 : 3'b101;
								assign node138 = (inp[11]) ? node148 : node139;
									assign node139 = (inp[3]) ? node145 : node140;
										assign node140 = (inp[5]) ? 3'b001 : node141;
											assign node141 = (inp[2]) ? 3'b001 : 3'b101;
										assign node145 = (inp[2]) ? 3'b110 : 3'b001;
									assign node148 = (inp[2]) ? node150 : 3'b110;
										assign node150 = (inp[3]) ? 3'b010 : 3'b110;
						assign node153 = (inp[1]) ? node187 : node154;
							assign node154 = (inp[11]) ? node170 : node155;
								assign node155 = (inp[8]) ? node165 : node156;
									assign node156 = (inp[3]) ? 3'b010 : node157;
										assign node157 = (inp[2]) ? 3'b010 : node158;
											assign node158 = (inp[4]) ? node160 : 3'b110;
												assign node160 = (inp[5]) ? 3'b010 : 3'b110;
									assign node165 = (inp[3]) ? 3'b110 : node166;
										assign node166 = (inp[2]) ? 3'b110 : 3'b001;
								assign node170 = (inp[8]) ? node182 : node171;
									assign node171 = (inp[2]) ? node175 : node172;
										assign node172 = (inp[3]) ? 3'b100 : 3'b010;
										assign node175 = (inp[4]) ? node177 : 3'b100;
											assign node177 = (inp[5]) ? node179 : 3'b100;
												assign node179 = (inp[3]) ? 3'b000 : 3'b100;
									assign node182 = (inp[2]) ? 3'b010 : node183;
										assign node183 = (inp[3]) ? 3'b010 : 3'b110;
							assign node187 = (inp[8]) ? node195 : node188;
								assign node188 = (inp[11]) ? 3'b000 : node189;
									assign node189 = (inp[3]) ? node191 : 3'b100;
										assign node191 = (inp[2]) ? 3'b000 : 3'b100;
								assign node195 = (inp[11]) ? node207 : node196;
									assign node196 = (inp[3]) ? node202 : node197;
										assign node197 = (inp[2]) ? 3'b010 : node198;
											assign node198 = (inp[4]) ? 3'b010 : 3'b110;
										assign node202 = (inp[2]) ? node204 : 3'b010;
											assign node204 = (inp[4]) ? 3'b100 : 3'b010;
									assign node207 = (inp[4]) ? node213 : node208;
										assign node208 = (inp[2]) ? node210 : 3'b010;
											assign node210 = (inp[3]) ? 3'b000 : 3'b100;
										assign node213 = (inp[5]) ? node215 : 3'b100;
											assign node215 = (inp[2]) ? node217 : 3'b100;
												assign node217 = (inp[3]) ? 3'b000 : 3'b100;
				assign node220 = (inp[10]) ? node284 : node221;
					assign node221 = (inp[7]) ? node235 : node222;
						assign node222 = (inp[11]) ? 3'b000 : node223;
							assign node223 = (inp[8]) ? node225 : 3'b000;
								assign node225 = (inp[1]) ? 3'b000 : node226;
									assign node226 = (inp[2]) ? 3'b000 : node227;
										assign node227 = (inp[3]) ? node229 : 3'b100;
											assign node229 = (inp[4]) ? 3'b000 : 3'b100;
						assign node235 = (inp[8]) ? node257 : node236;
							assign node236 = (inp[1]) ? node250 : node237;
								assign node237 = (inp[11]) ? node247 : node238;
									assign node238 = (inp[5]) ? 3'b100 : node239;
										assign node239 = (inp[2]) ? node241 : 3'b010;
											assign node241 = (inp[4]) ? 3'b100 : node242;
												assign node242 = (inp[3]) ? 3'b100 : 3'b010;
									assign node247 = (inp[2]) ? 3'b000 : 3'b100;
								assign node250 = (inp[3]) ? 3'b000 : node251;
									assign node251 = (inp[2]) ? 3'b000 : node252;
										assign node252 = (inp[11]) ? 3'b000 : 3'b100;
							assign node257 = (inp[1]) ? node273 : node258;
								assign node258 = (inp[11]) ? node266 : node259;
									assign node259 = (inp[2]) ? node261 : 3'b110;
										assign node261 = (inp[3]) ? 3'b010 : node262;
											assign node262 = (inp[4]) ? 3'b010 : 3'b110;
									assign node266 = (inp[2]) ? node268 : 3'b010;
										assign node268 = (inp[4]) ? 3'b100 : node269;
											assign node269 = (inp[3]) ? 3'b100 : 3'b010;
								assign node273 = (inp[11]) ? node279 : node274;
									assign node274 = (inp[2]) ? 3'b100 : node275;
										assign node275 = (inp[3]) ? 3'b100 : 3'b010;
									assign node279 = (inp[2]) ? 3'b000 : node280;
										assign node280 = (inp[3]) ? 3'b000 : 3'b100;
					assign node284 = (inp[1]) ? 3'b000 : node285;
						assign node285 = (inp[7]) ? node287 : 3'b000;
							assign node287 = (inp[2]) ? 3'b000 : node288;
								assign node288 = (inp[8]) ? node290 : 3'b000;
									assign node290 = (inp[11]) ? 3'b000 : 3'b100;
			assign node295 = (inp[0]) ? 3'b000 : node296;
				assign node296 = (inp[1]) ? 3'b000 : node297;
					assign node297 = (inp[7]) ? node299 : 3'b000;
						assign node299 = (inp[10]) ? 3'b000 : node300;
							assign node300 = (inp[8]) ? node308 : node301;
								assign node301 = (inp[3]) ? 3'b000 : node302;
									assign node302 = (inp[11]) ? 3'b000 : node303;
										assign node303 = (inp[2]) ? 3'b000 : 3'b100;
								assign node308 = (inp[2]) ? node316 : node309;
									assign node309 = (inp[11]) ? 3'b100 : node310;
										assign node310 = (inp[3]) ? node312 : 3'b010;
											assign node312 = (inp[4]) ? 3'b100 : 3'b010;
									assign node316 = (inp[11]) ? 3'b000 : 3'b100;
		assign node322 = (inp[9]) ? node778 : node323;
			assign node323 = (inp[0]) ? node513 : node324;
				assign node324 = (inp[7]) ? node456 : node325;
					assign node325 = (inp[10]) ? node381 : node326;
						assign node326 = (inp[1]) ? node348 : node327;
							assign node327 = (inp[8]) ? node339 : node328;
								assign node328 = (inp[11]) ? node334 : node329;
									assign node329 = (inp[3]) ? 3'b011 : node330;
										assign node330 = (inp[2]) ? 3'b011 : 3'b111;
									assign node334 = (inp[2]) ? 3'b101 : node335;
										assign node335 = (inp[3]) ? 3'b101 : 3'b011;
								assign node339 = (inp[11]) ? node341 : 3'b111;
									assign node341 = (inp[2]) ? 3'b011 : node342;
										assign node342 = (inp[3]) ? node344 : 3'b111;
											assign node344 = (inp[5]) ? 3'b011 : 3'b111;
							assign node348 = (inp[11]) ? node368 : node349;
								assign node349 = (inp[8]) ? node357 : node350;
									assign node350 = (inp[3]) ? 3'b101 : node351;
										assign node351 = (inp[4]) ? 3'b101 : node352;
											assign node352 = (inp[5]) ? 3'b101 : 3'b011;
									assign node357 = (inp[2]) ? node363 : node358;
										assign node358 = (inp[4]) ? 3'b011 : node359;
											assign node359 = (inp[3]) ? 3'b011 : 3'b111;
										assign node363 = (inp[3]) ? node365 : 3'b011;
											assign node365 = (inp[4]) ? 3'b101 : 3'b011;
								assign node368 = (inp[8]) ? 3'b101 : node369;
									assign node369 = (inp[2]) ? node375 : node370;
										assign node370 = (inp[4]) ? 3'b001 : node371;
											assign node371 = (inp[3]) ? 3'b001 : 3'b101;
										assign node375 = (inp[3]) ? node377 : 3'b001;
											assign node377 = (inp[4]) ? 3'b110 : 3'b001;
						assign node381 = (inp[1]) ? node413 : node382;
							assign node382 = (inp[11]) ? node400 : node383;
								assign node383 = (inp[8]) ? node393 : node384;
									assign node384 = (inp[2]) ? 3'b001 : node385;
										assign node385 = (inp[3]) ? node387 : 3'b101;
											assign node387 = (inp[4]) ? 3'b001 : node388;
												assign node388 = (inp[5]) ? 3'b001 : 3'b101;
									assign node393 = (inp[2]) ? 3'b101 : node394;
										assign node394 = (inp[3]) ? node396 : 3'b011;
											assign node396 = (inp[4]) ? 3'b101 : 3'b011;
								assign node400 = (inp[8]) ? node406 : node401;
									assign node401 = (inp[2]) ? 3'b110 : node402;
										assign node402 = (inp[4]) ? 3'b110 : 3'b001;
									assign node406 = (inp[2]) ? 3'b001 : node407;
										assign node407 = (inp[4]) ? node409 : 3'b101;
											assign node409 = (inp[3]) ? 3'b001 : 3'b101;
							assign node413 = (inp[8]) ? node435 : node414;
								assign node414 = (inp[11]) ? node424 : node415;
									assign node415 = (inp[4]) ? node419 : node416;
										assign node416 = (inp[2]) ? 3'b110 : 3'b001;
										assign node419 = (inp[2]) ? node421 : 3'b110;
											assign node421 = (inp[3]) ? 3'b010 : 3'b110;
									assign node424 = (inp[4]) ? node430 : node425;
										assign node425 = (inp[2]) ? 3'b010 : node426;
											assign node426 = (inp[3]) ? 3'b010 : 3'b110;
										assign node430 = (inp[2]) ? node432 : 3'b010;
											assign node432 = (inp[3]) ? 3'b100 : 3'b010;
								assign node435 = (inp[11]) ? node447 : node436;
									assign node436 = (inp[4]) ? node438 : 3'b001;
										assign node438 = (inp[3]) ? node444 : node439;
											assign node439 = (inp[2]) ? 3'b001 : node440;
												assign node440 = (inp[5]) ? 3'b001 : 3'b101;
											assign node444 = (inp[2]) ? 3'b110 : 3'b001;
									assign node447 = (inp[3]) ? node451 : node448;
										assign node448 = (inp[2]) ? 3'b110 : 3'b001;
										assign node451 = (inp[4]) ? node453 : 3'b110;
											assign node453 = (inp[2]) ? 3'b010 : 3'b110;
					assign node456 = (inp[10]) ? node472 : node457;
						assign node457 = (inp[11]) ? node459 : 3'b111;
							assign node459 = (inp[1]) ? node461 : 3'b111;
								assign node461 = (inp[8]) ? 3'b111 : node462;
									assign node462 = (inp[2]) ? node466 : node463;
										assign node463 = (inp[3]) ? 3'b011 : 3'b111;
										assign node466 = (inp[3]) ? node468 : 3'b011;
											assign node468 = (inp[5]) ? 3'b101 : 3'b011;
						assign node472 = (inp[1]) ? node490 : node473;
							assign node473 = (inp[8]) ? node483 : node474;
								assign node474 = (inp[11]) ? node478 : node475;
									assign node475 = (inp[2]) ? 3'b011 : 3'b111;
									assign node478 = (inp[2]) ? node480 : 3'b011;
										assign node480 = (inp[5]) ? 3'b101 : 3'b011;
								assign node483 = (inp[11]) ? node485 : 3'b111;
									assign node485 = (inp[2]) ? node487 : 3'b111;
										assign node487 = (inp[3]) ? 3'b011 : 3'b111;
							assign node490 = (inp[8]) ? node502 : node491;
								assign node491 = (inp[11]) ? node497 : node492;
									assign node492 = (inp[3]) ? 3'b101 : node493;
										assign node493 = (inp[2]) ? 3'b101 : 3'b011;
									assign node497 = (inp[3]) ? 3'b001 : node498;
										assign node498 = (inp[2]) ? 3'b001 : 3'b101;
								assign node502 = (inp[11]) ? node508 : node503;
									assign node503 = (inp[5]) ? 3'b011 : node504;
										assign node504 = (inp[2]) ? 3'b011 : 3'b111;
									assign node508 = (inp[2]) ? 3'b101 : node509;
										assign node509 = (inp[3]) ? 3'b101 : 3'b011;
				assign node513 = (inp[7]) ? node633 : node514;
					assign node514 = (inp[10]) ? node578 : node515;
						assign node515 = (inp[8]) ? node547 : node516;
							assign node516 = (inp[11]) ? node532 : node517;
								assign node517 = (inp[1]) ? node525 : node518;
									assign node518 = (inp[2]) ? node520 : 3'b001;
										assign node520 = (inp[4]) ? 3'b110 : node521;
											assign node521 = (inp[3]) ? 3'b110 : 3'b001;
									assign node525 = (inp[2]) ? 3'b010 : node526;
										assign node526 = (inp[3]) ? node528 : 3'b110;
											assign node528 = (inp[4]) ? 3'b010 : 3'b110;
								assign node532 = (inp[1]) ? node538 : node533;
									assign node533 = (inp[3]) ? node535 : 3'b110;
										assign node535 = (inp[2]) ? 3'b010 : 3'b110;
									assign node538 = (inp[2]) ? 3'b100 : node539;
										assign node539 = (inp[3]) ? node541 : 3'b010;
											assign node541 = (inp[4]) ? node543 : 3'b010;
												assign node543 = (inp[5]) ? 3'b100 : 3'b010;
							assign node547 = (inp[1]) ? node563 : node548;
								assign node548 = (inp[11]) ? node558 : node549;
									assign node549 = (inp[2]) ? node551 : 3'b101;
										assign node551 = (inp[3]) ? 3'b001 : node552;
											assign node552 = (inp[4]) ? node554 : 3'b101;
												assign node554 = (inp[5]) ? 3'b001 : 3'b101;
									assign node558 = (inp[2]) ? node560 : 3'b001;
										assign node560 = (inp[3]) ? 3'b110 : 3'b001;
								assign node563 = (inp[2]) ? node571 : node564;
									assign node564 = (inp[11]) ? node566 : 3'b001;
										assign node566 = (inp[3]) ? node568 : 3'b110;
											assign node568 = (inp[5]) ? 3'b010 : 3'b110;
									assign node571 = (inp[11]) ? node573 : 3'b110;
										assign node573 = (inp[4]) ? 3'b010 : node574;
											assign node574 = (inp[5]) ? 3'b010 : 3'b110;
						assign node578 = (inp[1]) ? node604 : node579;
							assign node579 = (inp[8]) ? node591 : node580;
								assign node580 = (inp[11]) ? node586 : node581;
									assign node581 = (inp[3]) ? node583 : 3'b010;
										assign node583 = (inp[2]) ? 3'b100 : 3'b010;
									assign node586 = (inp[3]) ? node588 : 3'b100;
										assign node588 = (inp[2]) ? 3'b000 : 3'b100;
								assign node591 = (inp[11]) ? node597 : node592;
									assign node592 = (inp[3]) ? node594 : 3'b110;
										assign node594 = (inp[2]) ? 3'b010 : 3'b110;
									assign node597 = (inp[3]) ? node599 : 3'b010;
										assign node599 = (inp[2]) ? node601 : 3'b010;
											assign node601 = (inp[5]) ? 3'b100 : 3'b010;
							assign node604 = (inp[8]) ? node618 : node605;
								assign node605 = (inp[11]) ? 3'b000 : node606;
									assign node606 = (inp[4]) ? node612 : node607;
										assign node607 = (inp[2]) ? node609 : 3'b100;
											assign node609 = (inp[5]) ? 3'b000 : 3'b100;
										assign node612 = (inp[3]) ? 3'b000 : node613;
											assign node613 = (inp[2]) ? 3'b000 : 3'b100;
								assign node618 = (inp[11]) ? node626 : node619;
									assign node619 = (inp[2]) ? node621 : 3'b010;
										assign node621 = (inp[5]) ? 3'b100 : node622;
											assign node622 = (inp[3]) ? 3'b100 : 3'b010;
									assign node626 = (inp[2]) ? node628 : 3'b100;
										assign node628 = (inp[3]) ? 3'b000 : node629;
											assign node629 = (inp[5]) ? 3'b000 : 3'b100;
					assign node633 = (inp[10]) ? node701 : node634;
						assign node634 = (inp[1]) ? node674 : node635;
							assign node635 = (inp[8]) ? node655 : node636;
								assign node636 = (inp[11]) ? node642 : node637;
									assign node637 = (inp[2]) ? node639 : 3'b011;
										assign node639 = (inp[3]) ? 3'b101 : 3'b011;
									assign node642 = (inp[5]) ? node650 : node643;
										assign node643 = (inp[4]) ? 3'b001 : node644;
											assign node644 = (inp[2]) ? 3'b101 : node645;
												assign node645 = (inp[3]) ? 3'b101 : 3'b011;
										assign node650 = (inp[3]) ? node652 : 3'b101;
											assign node652 = (inp[2]) ? 3'b001 : 3'b101;
								assign node655 = (inp[11]) ? node663 : node656;
									assign node656 = (inp[2]) ? node658 : 3'b111;
										assign node658 = (inp[3]) ? node660 : 3'b111;
											assign node660 = (inp[4]) ? 3'b011 : 3'b111;
									assign node663 = (inp[3]) ? node669 : node664;
										assign node664 = (inp[2]) ? 3'b011 : node665;
											assign node665 = (inp[4]) ? 3'b011 : 3'b111;
										assign node669 = (inp[4]) ? node671 : 3'b011;
											assign node671 = (inp[2]) ? 3'b101 : 3'b011;
							assign node674 = (inp[8]) ? node686 : node675;
								assign node675 = (inp[11]) ? node683 : node676;
									assign node676 = (inp[2]) ? node678 : 3'b101;
										assign node678 = (inp[4]) ? 3'b001 : node679;
											assign node679 = (inp[3]) ? 3'b001 : 3'b101;
									assign node683 = (inp[2]) ? 3'b110 : 3'b001;
								assign node686 = (inp[11]) ? node694 : node687;
									assign node687 = (inp[2]) ? node689 : 3'b011;
										assign node689 = (inp[4]) ? 3'b101 : node690;
											assign node690 = (inp[3]) ? 3'b101 : 3'b011;
									assign node694 = (inp[2]) ? node696 : 3'b101;
										assign node696 = (inp[3]) ? 3'b001 : node697;
											assign node697 = (inp[4]) ? 3'b001 : 3'b101;
						assign node701 = (inp[1]) ? node749 : node702;
							assign node702 = (inp[11]) ? node728 : node703;
								assign node703 = (inp[8]) ? node717 : node704;
									assign node704 = (inp[4]) ? 3'b001 : node705;
										assign node705 = (inp[5]) ? node711 : node706;
											assign node706 = (inp[2]) ? 3'b001 : node707;
												assign node707 = (inp[3]) ? 3'b001 : 3'b101;
											assign node711 = (inp[2]) ? node713 : 3'b001;
												assign node713 = (inp[3]) ? 3'b110 : 3'b001;
									assign node717 = (inp[2]) ? node723 : node718;
										assign node718 = (inp[3]) ? 3'b101 : node719;
											assign node719 = (inp[4]) ? 3'b101 : 3'b011;
										assign node723 = (inp[3]) ? node725 : 3'b101;
											assign node725 = (inp[4]) ? 3'b001 : 3'b101;
								assign node728 = (inp[8]) ? node740 : node729;
									assign node729 = (inp[4]) ? node735 : node730;
										assign node730 = (inp[2]) ? 3'b110 : node731;
											assign node731 = (inp[3]) ? 3'b110 : 3'b001;
										assign node735 = (inp[2]) ? node737 : 3'b110;
											assign node737 = (inp[3]) ? 3'b010 : 3'b110;
									assign node740 = (inp[2]) ? node744 : node741;
										assign node741 = (inp[3]) ? 3'b001 : 3'b101;
										assign node744 = (inp[3]) ? node746 : 3'b011;
											assign node746 = (inp[4]) ? 3'b110 : 3'b001;
							assign node749 = (inp[8]) ? node765 : node750;
								assign node750 = (inp[11]) ? node758 : node751;
									assign node751 = (inp[2]) ? node753 : 3'b110;
										assign node753 = (inp[4]) ? 3'b010 : node754;
											assign node754 = (inp[3]) ? 3'b010 : 3'b110;
									assign node758 = (inp[2]) ? node760 : 3'b010;
										assign node760 = (inp[4]) ? 3'b100 : node761;
											assign node761 = (inp[3]) ? 3'b100 : 3'b010;
								assign node765 = (inp[11]) ? node773 : node766;
									assign node766 = (inp[2]) ? node768 : 3'b001;
										assign node768 = (inp[3]) ? 3'b110 : node769;
											assign node769 = (inp[5]) ? 3'b110 : 3'b001;
									assign node773 = (inp[2]) ? node775 : 3'b110;
										assign node775 = (inp[3]) ? 3'b010 : 3'b110;
			assign node778 = (inp[0]) ? node1008 : node779;
				assign node779 = (inp[7]) ? node889 : node780;
					assign node780 = (inp[10]) ? node850 : node781;
						assign node781 = (inp[1]) ? node817 : node782;
							assign node782 = (inp[8]) ? node798 : node783;
								assign node783 = (inp[11]) ? node791 : node784;
									assign node784 = (inp[2]) ? 3'b010 : node785;
										assign node785 = (inp[4]) ? node787 : 3'b110;
											assign node787 = (inp[3]) ? 3'b010 : 3'b110;
									assign node791 = (inp[2]) ? 3'b100 : node792;
										assign node792 = (inp[3]) ? node794 : 3'b010;
											assign node794 = (inp[5]) ? 3'b100 : 3'b010;
								assign node798 = (inp[2]) ? node810 : node799;
									assign node799 = (inp[11]) ? node805 : node800;
										assign node800 = (inp[3]) ? node802 : 3'b001;
											assign node802 = (inp[5]) ? 3'b110 : 3'b001;
										assign node805 = (inp[5]) ? node807 : 3'b110;
											assign node807 = (inp[4]) ? 3'b010 : 3'b110;
									assign node810 = (inp[11]) ? node812 : 3'b110;
										assign node812 = (inp[4]) ? 3'b010 : node813;
											assign node813 = (inp[3]) ? 3'b010 : 3'b110;
							assign node817 = (inp[8]) ? node837 : node818;
								assign node818 = (inp[11]) ? node832 : node819;
									assign node819 = (inp[2]) ? node825 : node820;
										assign node820 = (inp[3]) ? 3'b100 : node821;
											assign node821 = (inp[5]) ? 3'b100 : 3'b010;
										assign node825 = (inp[4]) ? node827 : 3'b100;
											assign node827 = (inp[3]) ? node829 : 3'b100;
												assign node829 = (inp[5]) ? 3'b000 : 3'b100;
									assign node832 = (inp[2]) ? 3'b000 : node833;
										assign node833 = (inp[3]) ? 3'b000 : 3'b100;
								assign node837 = (inp[11]) ? node843 : node838;
									assign node838 = (inp[2]) ? 3'b010 : node839;
										assign node839 = (inp[3]) ? 3'b010 : 3'b110;
									assign node843 = (inp[5]) ? node845 : 3'b100;
										assign node845 = (inp[3]) ? 3'b100 : node846;
											assign node846 = (inp[2]) ? 3'b100 : 3'b010;
						assign node850 = (inp[1]) ? node876 : node851;
							assign node851 = (inp[2]) ? node861 : node852;
								assign node852 = (inp[11]) ? node858 : node853;
									assign node853 = (inp[8]) ? node855 : 3'b100;
										assign node855 = (inp[3]) ? 3'b100 : 3'b010;
									assign node858 = (inp[8]) ? 3'b100 : 3'b000;
								assign node861 = (inp[8]) ? node863 : 3'b000;
									assign node863 = (inp[11]) ? node869 : node864;
										assign node864 = (inp[3]) ? 3'b100 : node865;
											assign node865 = (inp[5]) ? 3'b100 : 3'b010;
										assign node869 = (inp[4]) ? 3'b000 : node870;
											assign node870 = (inp[5]) ? 3'b000 : node871;
												assign node871 = (inp[3]) ? 3'b000 : 3'b100;
							assign node876 = (inp[2]) ? 3'b000 : node877;
								assign node877 = (inp[8]) ? node879 : 3'b000;
									assign node879 = (inp[11]) ? 3'b000 : node880;
										assign node880 = (inp[3]) ? node882 : 3'b100;
											assign node882 = (inp[4]) ? 3'b000 : node883;
												assign node883 = (inp[5]) ? 3'b000 : 3'b100;
					assign node889 = (inp[10]) ? node951 : node890;
						assign node890 = (inp[1]) ? node920 : node891;
							assign node891 = (inp[8]) ? node905 : node892;
								assign node892 = (inp[5]) ? node900 : node893;
									assign node893 = (inp[2]) ? node897 : node894;
										assign node894 = (inp[11]) ? 3'b001 : 3'b101;
										assign node897 = (inp[3]) ? 3'b110 : 3'b001;
									assign node900 = (inp[2]) ? 3'b001 : node901;
										assign node901 = (inp[11]) ? 3'b001 : 3'b101;
								assign node905 = (inp[11]) ? node913 : node906;
									assign node906 = (inp[2]) ? node908 : 3'b011;
										assign node908 = (inp[3]) ? 3'b101 : node909;
											assign node909 = (inp[4]) ? 3'b101 : 3'b011;
									assign node913 = (inp[2]) ? node915 : 3'b101;
										assign node915 = (inp[3]) ? 3'b001 : node916;
											assign node916 = (inp[4]) ? 3'b001 : 3'b101;
							assign node920 = (inp[11]) ? node934 : node921;
								assign node921 = (inp[8]) ? node927 : node922;
									assign node922 = (inp[2]) ? 3'b110 : node923;
										assign node923 = (inp[3]) ? 3'b110 : 3'b001;
									assign node927 = (inp[2]) ? 3'b001 : node928;
										assign node928 = (inp[3]) ? node930 : 3'b101;
											assign node930 = (inp[4]) ? 3'b001 : 3'b101;
								assign node934 = (inp[8]) ? node944 : node935;
									assign node935 = (inp[2]) ? 3'b010 : node936;
										assign node936 = (inp[3]) ? node938 : 3'b110;
											assign node938 = (inp[4]) ? 3'b010 : node939;
												assign node939 = (inp[5]) ? 3'b010 : 3'b110;
									assign node944 = (inp[2]) ? 3'b110 : node945;
										assign node945 = (inp[4]) ? node947 : 3'b001;
											assign node947 = (inp[3]) ? 3'b110 : 3'b001;
						assign node951 = (inp[1]) ? node985 : node952;
							assign node952 = (inp[8]) ? node970 : node953;
								assign node953 = (inp[11]) ? node961 : node954;
									assign node954 = (inp[2]) ? node956 : 3'b110;
										assign node956 = (inp[4]) ? 3'b010 : node957;
											assign node957 = (inp[3]) ? 3'b010 : 3'b110;
									assign node961 = (inp[2]) ? node963 : 3'b010;
										assign node963 = (inp[3]) ? 3'b100 : node964;
											assign node964 = (inp[5]) ? node966 : 3'b010;
												assign node966 = (inp[4]) ? 3'b100 : 3'b010;
								assign node970 = (inp[11]) ? node980 : node971;
									assign node971 = (inp[2]) ? node973 : 3'b001;
										assign node973 = (inp[3]) ? 3'b110 : node974;
											assign node974 = (inp[5]) ? node976 : 3'b001;
												assign node976 = (inp[4]) ? 3'b110 : 3'b001;
									assign node980 = (inp[3]) ? node982 : 3'b110;
										assign node982 = (inp[2]) ? 3'b010 : 3'b110;
							assign node985 = (inp[8]) ? node999 : node986;
								assign node986 = (inp[11]) ? node992 : node987;
									assign node987 = (inp[2]) ? 3'b100 : node988;
										assign node988 = (inp[3]) ? 3'b100 : 3'b010;
									assign node992 = (inp[2]) ? 3'b000 : node993;
										assign node993 = (inp[3]) ? node995 : 3'b100;
											assign node995 = (inp[4]) ? 3'b000 : 3'b100;
								assign node999 = (inp[11]) ? node1003 : node1000;
									assign node1000 = (inp[2]) ? 3'b010 : 3'b110;
									assign node1003 = (inp[2]) ? 3'b100 : node1004;
										assign node1004 = (inp[4]) ? 3'b100 : 3'b010;
				assign node1008 = (inp[7]) ? node1026 : node1009;
					assign node1009 = (inp[11]) ? 3'b000 : node1010;
						assign node1010 = (inp[1]) ? 3'b000 : node1011;
							assign node1011 = (inp[8]) ? node1013 : 3'b000;
								assign node1013 = (inp[10]) ? 3'b000 : node1014;
									assign node1014 = (inp[3]) ? node1020 : node1015;
										assign node1015 = (inp[4]) ? 3'b100 : node1016;
											assign node1016 = (inp[5]) ? 3'b100 : 3'b010;
										assign node1020 = (inp[2]) ? 3'b000 : 3'b100;
					assign node1026 = (inp[10]) ? node1098 : node1027;
						assign node1027 = (inp[1]) ? node1073 : node1028;
							assign node1028 = (inp[11]) ? node1048 : node1029;
								assign node1029 = (inp[8]) ? node1039 : node1030;
									assign node1030 = (inp[5]) ? node1034 : node1031;
										assign node1031 = (inp[3]) ? 3'b100 : 3'b010;
										assign node1034 = (inp[3]) ? 3'b010 : node1035;
											assign node1035 = (inp[2]) ? 3'b010 : 3'b110;
									assign node1039 = (inp[3]) ? node1043 : node1040;
										assign node1040 = (inp[2]) ? 3'b110 : 3'b001;
										assign node1043 = (inp[2]) ? node1045 : 3'b110;
											assign node1045 = (inp[4]) ? 3'b010 : 3'b110;
								assign node1048 = (inp[8]) ? node1060 : node1049;
									assign node1049 = (inp[2]) ? node1057 : node1050;
										assign node1050 = (inp[3]) ? 3'b100 : node1051;
											assign node1051 = (inp[4]) ? node1053 : 3'b010;
												assign node1053 = (inp[5]) ? 3'b100 : 3'b010;
										assign node1057 = (inp[3]) ? 3'b000 : 3'b100;
									assign node1060 = (inp[2]) ? node1068 : node1061;
										assign node1061 = (inp[3]) ? 3'b010 : node1062;
											assign node1062 = (inp[5]) ? node1064 : 3'b110;
												assign node1064 = (inp[4]) ? 3'b010 : 3'b110;
										assign node1068 = (inp[4]) ? 3'b100 : node1069;
											assign node1069 = (inp[3]) ? 3'b000 : 3'b010;
							assign node1073 = (inp[11]) ? node1089 : node1074;
								assign node1074 = (inp[8]) ? node1084 : node1075;
									assign node1075 = (inp[2]) ? node1077 : 3'b100;
										assign node1077 = (inp[3]) ? 3'b000 : node1078;
											assign node1078 = (inp[4]) ? node1080 : 3'b100;
												assign node1080 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1084 = (inp[2]) ? node1086 : 3'b010;
										assign node1086 = (inp[3]) ? 3'b100 : 3'b010;
								assign node1089 = (inp[8]) ? node1091 : 3'b000;
									assign node1091 = (inp[3]) ? node1095 : node1092;
										assign node1092 = (inp[2]) ? 3'b100 : 3'b000;
										assign node1095 = (inp[2]) ? 3'b000 : 3'b100;
						assign node1098 = (inp[1]) ? 3'b000 : node1099;
							assign node1099 = (inp[8]) ? node1101 : 3'b000;
								assign node1101 = (inp[11]) ? node1109 : node1102;
									assign node1102 = (inp[2]) ? 3'b100 : node1103;
										assign node1103 = (inp[3]) ? 3'b100 : node1104;
											assign node1104 = (inp[4]) ? 3'b010 : 3'b011;
									assign node1109 = (inp[3]) ? 3'b000 : node1110;
										assign node1110 = (inp[2]) ? 3'b000 : 3'b100;

endmodule