module dtc_split33_bm32 (
	input  wire [15-1:0] inp,
	output wire [9-1:0] outp
);

	wire [9-1:0] node1;
	wire [9-1:0] node2;
	wire [9-1:0] node5;
	wire [9-1:0] node6;
	wire [9-1:0] node7;
	wire [9-1:0] node9;
	wire [9-1:0] node10;
	wire [9-1:0] node12;
	wire [9-1:0] node14;
	wire [9-1:0] node18;
	wire [9-1:0] node21;
	wire [9-1:0] node22;
	wire [9-1:0] node24;
	wire [9-1:0] node26;
	wire [9-1:0] node29;
	wire [9-1:0] node30;
	wire [9-1:0] node32;
	wire [9-1:0] node34;
	wire [9-1:0] node35;
	wire [9-1:0] node39;
	wire [9-1:0] node41;
	wire [9-1:0] node42;
	wire [9-1:0] node45;
	wire [9-1:0] node48;
	wire [9-1:0] node49;
	wire [9-1:0] node50;
	wire [9-1:0] node51;
	wire [9-1:0] node52;
	wire [9-1:0] node53;
	wire [9-1:0] node54;
	wire [9-1:0] node55;
	wire [9-1:0] node60;
	wire [9-1:0] node61;
	wire [9-1:0] node62;
	wire [9-1:0] node63;
	wire [9-1:0] node68;
	wire [9-1:0] node71;
	wire [9-1:0] node72;
	wire [9-1:0] node73;
	wire [9-1:0] node74;
	wire [9-1:0] node79;
	wire [9-1:0] node80;
	wire [9-1:0] node81;
	wire [9-1:0] node82;
	wire [9-1:0] node87;
	wire [9-1:0] node90;
	wire [9-1:0] node91;
	wire [9-1:0] node92;
	wire [9-1:0] node93;
	wire [9-1:0] node94;
	wire [9-1:0] node99;
	wire [9-1:0] node100;
	wire [9-1:0] node101;
	wire [9-1:0] node102;
	wire [9-1:0] node107;
	wire [9-1:0] node110;
	wire [9-1:0] node111;
	wire [9-1:0] node112;
	wire [9-1:0] node113;
	wire [9-1:0] node114;
	wire [9-1:0] node116;
	wire [9-1:0] node118;
	wire [9-1:0] node121;
	wire [9-1:0] node123;
	wire [9-1:0] node126;
	wire [9-1:0] node127;
	wire [9-1:0] node129;
	wire [9-1:0] node131;
	wire [9-1:0] node134;
	wire [9-1:0] node136;
	wire [9-1:0] node139;
	wire [9-1:0] node141;
	wire [9-1:0] node144;
	wire [9-1:0] node145;
	wire [9-1:0] node146;
	wire [9-1:0] node147;
	wire [9-1:0] node148;
	wire [9-1:0] node152;
	wire [9-1:0] node153;
	wire [9-1:0] node155;
	wire [9-1:0] node159;
	wire [9-1:0] node160;
	wire [9-1:0] node162;
	wire [9-1:0] node163;
	wire [9-1:0] node167;
	wire [9-1:0] node169;
	wire [9-1:0] node172;
	wire [9-1:0] node174;
	wire [9-1:0] node177;
	wire [9-1:0] node178;
	wire [9-1:0] node179;
	wire [9-1:0] node180;
	wire [9-1:0] node181;
	wire [9-1:0] node182;
	wire [9-1:0] node187;
	wire [9-1:0] node188;
	wire [9-1:0] node189;
	wire [9-1:0] node190;
	wire [9-1:0] node195;
	wire [9-1:0] node198;
	wire [9-1:0] node199;
	wire [9-1:0] node200;
	wire [9-1:0] node201;
	wire [9-1:0] node206;
	wire [9-1:0] node207;
	wire [9-1:0] node208;
	wire [9-1:0] node209;
	wire [9-1:0] node214;
	wire [9-1:0] node217;
	wire [9-1:0] node218;
	wire [9-1:0] node219;
	wire [9-1:0] node220;
	wire [9-1:0] node221;
	wire [9-1:0] node226;
	wire [9-1:0] node227;
	wire [9-1:0] node228;
	wire [9-1:0] node229;
	wire [9-1:0] node234;
	wire [9-1:0] node237;
	wire [9-1:0] node238;
	wire [9-1:0] node239;
	wire [9-1:0] node240;
	wire [9-1:0] node241;
	wire [9-1:0] node242;
	wire [9-1:0] node244;
	wire [9-1:0] node246;
	wire [9-1:0] node249;
	wire [9-1:0] node251;
	wire [9-1:0] node254;
	wire [9-1:0] node255;
	wire [9-1:0] node257;
	wire [9-1:0] node259;
	wire [9-1:0] node262;
	wire [9-1:0] node264;
	wire [9-1:0] node267;
	wire [9-1:0] node269;
	wire [9-1:0] node272;
	wire [9-1:0] node273;
	wire [9-1:0] node274;
	wire [9-1:0] node275;
	wire [9-1:0] node276;
	wire [9-1:0] node280;
	wire [9-1:0] node284;
	wire [9-1:0] node285;
	wire [9-1:0] node286;
	wire [9-1:0] node287;
	wire [9-1:0] node292;
	wire [9-1:0] node293;
	wire [9-1:0] node297;
	wire [9-1:0] node298;
	wire [9-1:0] node299;
	wire [9-1:0] node300;
	wire [9-1:0] node301;
	wire [9-1:0] node302;
	wire [9-1:0] node306;
	wire [9-1:0] node307;
	wire [9-1:0] node311;
	wire [9-1:0] node312;
	wire [9-1:0] node313;
	wire [9-1:0] node317;
	wire [9-1:0] node319;
	wire [9-1:0] node322;
	wire [9-1:0] node324;
	wire [9-1:0] node327;
	wire [9-1:0] node328;
	wire [9-1:0] node329;
	wire [9-1:0] node330;
	wire [9-1:0] node332;
	wire [9-1:0] node334;
	wire [9-1:0] node337;
	wire [9-1:0] node340;
	wire [9-1:0] node341;
	wire [9-1:0] node342;
	wire [9-1:0] node346;
	wire [9-1:0] node347;
	wire [9-1:0] node351;
	wire [9-1:0] node353;
	wire [9-1:0] node356;
	wire [9-1:0] node357;
	wire [9-1:0] node358;
	wire [9-1:0] node359;
	wire [9-1:0] node361;
	wire [9-1:0] node364;
	wire [9-1:0] node365;
	wire [9-1:0] node368;
	wire [9-1:0] node369;
	wire [9-1:0] node372;
	wire [9-1:0] node373;
	wire [9-1:0] node376;
	wire [9-1:0] node379;
	wire [9-1:0] node380;
	wire [9-1:0] node382;
	wire [9-1:0] node385;
	wire [9-1:0] node386;
	wire [9-1:0] node389;
	wire [9-1:0] node390;
	wire [9-1:0] node393;
	wire [9-1:0] node394;
	wire [9-1:0] node397;
	wire [9-1:0] node400;
	wire [9-1:0] node401;
	wire [9-1:0] node402;
	wire [9-1:0] node403;
	wire [9-1:0] node406;
	wire [9-1:0] node408;
	wire [9-1:0] node411;
	wire [9-1:0] node412;
	wire [9-1:0] node415;
	wire [9-1:0] node417;
	wire [9-1:0] node418;
	wire [9-1:0] node421;
	wire [9-1:0] node424;
	wire [9-1:0] node425;
	wire [9-1:0] node426;
	wire [9-1:0] node429;
	wire [9-1:0] node432;
	wire [9-1:0] node433;
	wire [9-1:0] node436;
	wire [9-1:0] node437;
	wire [9-1:0] node438;
	wire [9-1:0] node441;
	wire [9-1:0] node442;
	wire [9-1:0] node445;
	wire [9-1:0] node448;
	wire [9-1:0] node449;
	wire [9-1:0] node452;
	wire [9-1:0] node453;
	wire [9-1:0] node456;

	assign outp = (inp[12]) ? node48 : node1;
		assign node1 = (inp[13]) ? node5 : node2;
			assign node2 = (inp[11]) ? 9'b101010101 : 9'b101010000;
			assign node5 = (inp[14]) ? node21 : node6;
				assign node6 = (inp[0]) ? node18 : node7;
					assign node7 = (inp[3]) ? node9 : 9'b101010001;
						assign node9 = (inp[4]) ? 9'b100010001 : node10;
							assign node10 = (inp[9]) ? node12 : 9'b100010001;
								assign node12 = (inp[8]) ? node14 : 9'b100010001;
									assign node14 = (inp[6]) ? 9'b001010001 : 9'b101010001;
					assign node18 = (inp[3]) ? 9'b000010101 : 9'b101010101;
				assign node21 = (inp[3]) ? node29 : node22;
					assign node22 = (inp[8]) ? node24 : 9'b111010101;
						assign node24 = (inp[9]) ? node26 : 9'b101010101;
							assign node26 = (inp[4]) ? 9'b111010101 : 9'b101010101;
					assign node29 = (inp[0]) ? node39 : node30;
						assign node30 = (inp[8]) ? node32 : 9'b111010111;
							assign node32 = (inp[9]) ? node34 : 9'b101010111;
								assign node34 = (inp[4]) ? 9'b111010111 : node35;
									assign node35 = (inp[6]) ? 9'b011010101 : 9'b111010101;
						assign node39 = (inp[8]) ? node41 : 9'b011010111;
							assign node41 = (inp[4]) ? node45 : node42;
								assign node42 = (inp[9]) ? 9'b000010111 : 9'b001010111;
								assign node45 = (inp[9]) ? 9'b001010101 : 9'b001010111;
		assign node48 = (inp[8]) ? node356 : node49;
			assign node49 = (inp[6]) ? node177 : node50;
				assign node50 = (inp[13]) ? node90 : node51;
					assign node51 = (inp[11]) ? node71 : node52;
						assign node52 = (inp[7]) ? node60 : node53;
							assign node53 = (inp[1]) ? 9'b111011000 : node54;
								assign node54 = (inp[9]) ? 9'b111011000 : node55;
									assign node55 = (inp[2]) ? 9'b111111000 : 9'b111110000;
							assign node60 = (inp[4]) ? node68 : node61;
								assign node61 = (inp[9]) ? 9'b111111000 : node62;
									assign node62 = (inp[2]) ? 9'b111111000 : node63;
										assign node63 = (inp[1]) ? 9'b111111000 : 9'b111110000;
								assign node68 = (inp[9]) ? 9'b111010000 : 9'b111110000;
						assign node71 = (inp[7]) ? node79 : node72;
							assign node72 = (inp[9]) ? 9'b111011100 : node73;
								assign node73 = (inp[1]) ? 9'b111011100 : node74;
									assign node74 = (inp[2]) ? 9'b111111100 : 9'b111110100;
							assign node79 = (inp[4]) ? node87 : node80;
								assign node80 = (inp[9]) ? 9'b111111100 : node81;
									assign node81 = (inp[1]) ? 9'b111111100 : node82;
										assign node82 = (inp[2]) ? 9'b111111100 : 9'b111110100;
								assign node87 = (inp[9]) ? 9'b111010100 : 9'b111110100;
					assign node90 = (inp[3]) ? node110 : node91;
						assign node91 = (inp[7]) ? node99 : node92;
							assign node92 = (inp[1]) ? 9'b111011100 : node93;
								assign node93 = (inp[9]) ? 9'b111011100 : node94;
									assign node94 = (inp[2]) ? 9'b111111100 : 9'b111110100;
							assign node99 = (inp[4]) ? node107 : node100;
								assign node100 = (inp[9]) ? 9'b111111100 : node101;
									assign node101 = (inp[2]) ? 9'b111111100 : node102;
										assign node102 = (inp[1]) ? 9'b111111100 : 9'b111110100;
								assign node107 = (inp[9]) ? 9'b111010100 : 9'b111110100;
						assign node110 = (inp[14]) ? node144 : node111;
							assign node111 = (inp[9]) ? node139 : node112;
								assign node112 = (inp[10]) ? node126 : node113;
									assign node113 = (inp[1]) ? node121 : node114;
										assign node114 = (inp[2]) ? node116 : 9'b110110100;
											assign node116 = (inp[7]) ? node118 : 9'b110111100;
												assign node118 = (inp[4]) ? 9'b110110100 : 9'b110111100;
										assign node121 = (inp[7]) ? node123 : 9'b110011100;
											assign node123 = (inp[4]) ? 9'b110110100 : 9'b110111100;
									assign node126 = (inp[1]) ? node134 : node127;
										assign node127 = (inp[2]) ? node129 : 9'b110110110;
											assign node129 = (inp[7]) ? node131 : 9'b110111110;
												assign node131 = (inp[4]) ? 9'b110110110 : 9'b110111110;
										assign node134 = (inp[7]) ? node136 : 9'b110011110;
											assign node136 = (inp[4]) ? 9'b110110110 : 9'b110111110;
								assign node139 = (inp[7]) ? node141 : 9'b110011110;
									assign node141 = (inp[4]) ? 9'b110010110 : 9'b110111110;
							assign node144 = (inp[9]) ? node172 : node145;
								assign node145 = (inp[10]) ? node159 : node146;
									assign node146 = (inp[7]) ? node152 : node147;
										assign node147 = (inp[1]) ? 9'b111011100 : node148;
											assign node148 = (inp[2]) ? 9'b111111100 : 9'b111110100;
										assign node152 = (inp[4]) ? 9'b111110100 : node153;
											assign node153 = (inp[11]) ? node155 : 9'b111111100;
												assign node155 = (inp[1]) ? 9'b111111100 : 9'b111110100;
									assign node159 = (inp[1]) ? node167 : node160;
										assign node160 = (inp[2]) ? node162 : 9'b111110110;
											assign node162 = (inp[5]) ? 9'b111111110 : node163;
												assign node163 = (inp[4]) ? 9'b111110110 : 9'b111111110;
										assign node167 = (inp[7]) ? node169 : 9'b111011110;
											assign node169 = (inp[4]) ? 9'b111110110 : 9'b111111110;
								assign node172 = (inp[7]) ? node174 : 9'b111011110;
									assign node174 = (inp[4]) ? 9'b111010110 : 9'b111111110;
				assign node177 = (inp[13]) ? node217 : node178;
					assign node178 = (inp[11]) ? node198 : node179;
						assign node179 = (inp[7]) ? node187 : node180;
							assign node180 = (inp[9]) ? 9'b111011000 : node181;
								assign node181 = (inp[1]) ? 9'b111011000 : node182;
									assign node182 = (inp[2]) ? 9'b111111000 : 9'b111110000;
							assign node187 = (inp[4]) ? node195 : node188;
								assign node188 = (inp[2]) ? 9'b111111000 : node189;
									assign node189 = (inp[9]) ? 9'b111111000 : node190;
										assign node190 = (inp[1]) ? 9'b111111000 : 9'b111110000;
								assign node195 = (inp[9]) ? 9'b111010000 : 9'b111110000;
						assign node198 = (inp[7]) ? node206 : node199;
							assign node199 = (inp[9]) ? 9'b111011101 : node200;
								assign node200 = (inp[1]) ? 9'b111011101 : node201;
									assign node201 = (inp[2]) ? 9'b111111101 : 9'b111110101;
							assign node206 = (inp[4]) ? node214 : node207;
								assign node207 = (inp[9]) ? 9'b111111101 : node208;
									assign node208 = (inp[1]) ? 9'b111111101 : node209;
										assign node209 = (inp[2]) ? 9'b111111101 : 9'b111110101;
								assign node214 = (inp[9]) ? 9'b111010101 : 9'b111110101;
					assign node217 = (inp[3]) ? node237 : node218;
						assign node218 = (inp[7]) ? node226 : node219;
							assign node219 = (inp[1]) ? 9'b111011101 : node220;
								assign node220 = (inp[9]) ? 9'b111011101 : node221;
									assign node221 = (inp[2]) ? 9'b111111101 : 9'b111110101;
							assign node226 = (inp[4]) ? node234 : node227;
								assign node227 = (inp[1]) ? 9'b111111101 : node228;
									assign node228 = (inp[9]) ? 9'b111111101 : node229;
										assign node229 = (inp[2]) ? 9'b111111101 : 9'b111110101;
								assign node234 = (inp[9]) ? 9'b111010101 : 9'b111110101;
						assign node237 = (inp[5]) ? node297 : node238;
							assign node238 = (inp[14]) ? node272 : node239;
								assign node239 = (inp[9]) ? node267 : node240;
									assign node240 = (inp[10]) ? node254 : node241;
										assign node241 = (inp[1]) ? node249 : node242;
											assign node242 = (inp[2]) ? node244 : 9'b110100101;
												assign node244 = (inp[7]) ? node246 : 9'b110101101;
													assign node246 = (inp[4]) ? 9'b110100101 : 9'b110101101;
											assign node249 = (inp[7]) ? node251 : 9'b110001101;
												assign node251 = (inp[4]) ? 9'b110100101 : 9'b110101101;
										assign node254 = (inp[1]) ? node262 : node255;
											assign node255 = (inp[2]) ? node257 : 9'b110100111;
												assign node257 = (inp[4]) ? node259 : 9'b110101111;
													assign node259 = (inp[7]) ? 9'b110100111 : 9'b110101111;
											assign node262 = (inp[7]) ? node264 : 9'b110001111;
												assign node264 = (inp[4]) ? 9'b110100111 : 9'b110101111;
									assign node267 = (inp[7]) ? node269 : 9'b110001111;
										assign node269 = (inp[4]) ? 9'b110000111 : 9'b110101111;
								assign node272 = (inp[7]) ? node284 : node273;
									assign node273 = (inp[9]) ? 9'b111001111 : node274;
										assign node274 = (inp[1]) ? node280 : node275;
											assign node275 = (inp[2]) ? 9'b111101101 : node276;
												assign node276 = (inp[10]) ? 9'b111100111 : 9'b111100101;
											assign node280 = (inp[10]) ? 9'b111001111 : 9'b111001101;
									assign node284 = (inp[4]) ? node292 : node285;
										assign node285 = (inp[10]) ? 9'b111101111 : node286;
											assign node286 = (inp[9]) ? 9'b111101111 : node287;
												assign node287 = (inp[2]) ? 9'b111101101 : 9'b111100101;
										assign node292 = (inp[9]) ? 9'b111000111 : node293;
											assign node293 = (inp[10]) ? 9'b111100111 : 9'b111100101;
							assign node297 = (inp[14]) ? node327 : node298;
								assign node298 = (inp[9]) ? node322 : node299;
									assign node299 = (inp[10]) ? node311 : node300;
										assign node300 = (inp[7]) ? node306 : node301;
											assign node301 = (inp[1]) ? 9'b110011101 : node302;
												assign node302 = (inp[4]) ? 9'b110111101 : 9'b110110101;
											assign node306 = (inp[4]) ? 9'b110110101 : node307;
												assign node307 = (inp[1]) ? 9'b110111101 : 9'b110110101;
										assign node311 = (inp[1]) ? node317 : node312;
											assign node312 = (inp[7]) ? 9'b110110111 : node313;
												assign node313 = (inp[2]) ? 9'b110111111 : 9'b110110111;
											assign node317 = (inp[7]) ? node319 : 9'b110011111;
												assign node319 = (inp[4]) ? 9'b110110111 : 9'b110111111;
									assign node322 = (inp[7]) ? node324 : 9'b110011111;
										assign node324 = (inp[4]) ? 9'b110010111 : 9'b110111111;
								assign node327 = (inp[9]) ? node351 : node328;
									assign node328 = (inp[10]) ? node340 : node329;
										assign node329 = (inp[1]) ? node337 : node330;
											assign node330 = (inp[2]) ? node332 : 9'b111110101;
												assign node332 = (inp[7]) ? node334 : 9'b111111101;
													assign node334 = (inp[4]) ? 9'b111110101 : 9'b111111101;
											assign node337 = (inp[7]) ? 9'b111111101 : 9'b111011101;
										assign node340 = (inp[7]) ? node346 : node341;
											assign node341 = (inp[1]) ? 9'b111011111 : node342;
												assign node342 = (inp[2]) ? 9'b111111111 : 9'b111110111;
											assign node346 = (inp[4]) ? 9'b111110111 : node347;
												assign node347 = (inp[2]) ? 9'b111111111 : 9'b111110111;
									assign node351 = (inp[7]) ? node353 : 9'b111011111;
										assign node353 = (inp[4]) ? 9'b111010111 : 9'b111111111;
			assign node356 = (inp[9]) ? node400 : node357;
				assign node357 = (inp[4]) ? node379 : node358;
					assign node358 = (inp[13]) ? node364 : node359;
						assign node359 = (inp[11]) ? node361 : 9'b101111000;
							assign node361 = (inp[6]) ? 9'b101111101 : 9'b101111100;
						assign node364 = (inp[3]) ? node368 : node365;
							assign node365 = (inp[6]) ? 9'b101111101 : 9'b101111100;
							assign node368 = (inp[6]) ? node372 : node369;
								assign node369 = (inp[14]) ? 9'b101111110 : 9'b100111110;
								assign node372 = (inp[5]) ? node376 : node373;
									assign node373 = (inp[14]) ? 9'b101101111 : 9'b100101111;
									assign node376 = (inp[14]) ? 9'b101111111 : 9'b100111111;
					assign node379 = (inp[13]) ? node385 : node380;
						assign node380 = (inp[11]) ? node382 : 9'b101010000;
							assign node382 = (inp[6]) ? 9'b101010101 : 9'b101010100;
						assign node385 = (inp[3]) ? node389 : node386;
							assign node386 = (inp[6]) ? 9'b101010101 : 9'b101010100;
							assign node389 = (inp[6]) ? node393 : node390;
								assign node390 = (inp[14]) ? 9'b101010110 : 9'b100010110;
								assign node393 = (inp[5]) ? node397 : node394;
									assign node394 = (inp[14]) ? 9'b101000111 : 9'b100000111;
									assign node397 = (inp[14]) ? 9'b101010111 : 9'b100010111;
				assign node400 = (inp[6]) ? node424 : node401;
					assign node401 = (inp[4]) ? node411 : node402;
						assign node402 = (inp[13]) ? node406 : node403;
							assign node403 = (inp[11]) ? 9'b101010100 : 9'b101010000;
							assign node406 = (inp[3]) ? node408 : 9'b101010100;
								assign node408 = (inp[0]) ? 9'b100010110 : 9'b111010100;
						assign node411 = (inp[13]) ? node415 : node412;
							assign node412 = (inp[11]) ? 9'b111010100 : 9'b111010000;
							assign node415 = (inp[3]) ? node417 : 9'b111010100;
								assign node417 = (inp[0]) ? node421 : node418;
									assign node418 = (inp[14]) ? 9'b111010110 : 9'b110010110;
									assign node421 = (inp[14]) ? 9'b101010100 : 9'b100010100;
					assign node424 = (inp[13]) ? node432 : node425;
						assign node425 = (inp[11]) ? node429 : node426;
							assign node426 = (inp[4]) ? 9'b111010000 : 9'b101010000;
							assign node429 = (inp[4]) ? 9'b111010101 : 9'b101010101;
						assign node432 = (inp[3]) ? node436 : node433;
							assign node433 = (inp[4]) ? 9'b111010101 : 9'b101010101;
							assign node436 = (inp[0]) ? node448 : node437;
								assign node437 = (inp[4]) ? node441 : node438;
									assign node438 = (inp[5]) ? 9'b011010101 : 9'b011000101;
									assign node441 = (inp[14]) ? node445 : node442;
										assign node442 = (inp[5]) ? 9'b110010111 : 9'b110000111;
										assign node445 = (inp[5]) ? 9'b111010111 : 9'b111000111;
								assign node448 = (inp[4]) ? node452 : node449;
									assign node449 = (inp[5]) ? 9'b100010111 : 9'b100000111;
									assign node452 = (inp[5]) ? node456 : node453;
										assign node453 = (inp[14]) ? 9'b101000101 : 9'b100000101;
										assign node456 = (inp[14]) ? 9'b101010101 : 9'b100010101;

endmodule