module dtc_split75_bm77 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node25;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node236;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node253;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node258;
	wire [3-1:0] node260;
	wire [3-1:0] node262;
	wire [3-1:0] node264;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node292;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node299;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node337;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node352;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node364;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node387;
	wire [3-1:0] node389;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node404;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node426;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node446;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node455;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node469;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node482;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node498;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node511;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node549;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node557;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node564;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node580;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node586;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node593;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node602;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node609;
	wire [3-1:0] node612;
	wire [3-1:0] node613;
	wire [3-1:0] node614;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node629;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node637;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node648;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node654;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node661;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node668;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node681;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node695;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node700;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node707;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node714;
	wire [3-1:0] node717;
	wire [3-1:0] node719;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node727;
	wire [3-1:0] node730;
	wire [3-1:0] node732;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node743;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node751;
	wire [3-1:0] node754;
	wire [3-1:0] node756;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node762;
	wire [3-1:0] node764;
	wire [3-1:0] node767;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node773;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node779;
	wire [3-1:0] node781;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node787;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node794;
	wire [3-1:0] node796;
	wire [3-1:0] node799;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node805;
	wire [3-1:0] node808;
	wire [3-1:0] node810;
	wire [3-1:0] node812;
	wire [3-1:0] node814;

	assign outp = (inp[3]) ? node104 : node1;
		assign node1 = (inp[0]) ? node3 : 3'b000;
			assign node3 = (inp[4]) ? node5 : 3'b000;
				assign node5 = (inp[6]) ? 3'b000 : node6;
					assign node6 = (inp[7]) ? node88 : node7;
						assign node7 = (inp[1]) ? node41 : node8;
							assign node8 = (inp[9]) ? node30 : node9;
								assign node9 = (inp[10]) ? node19 : node10;
									assign node10 = (inp[5]) ? node16 : node11;
										assign node11 = (inp[11]) ? node13 : 3'b100;
											assign node13 = (inp[8]) ? 3'b100 : 3'b000;
										assign node16 = (inp[8]) ? 3'b000 : 3'b100;
									assign node19 = (inp[8]) ? node25 : node20;
										assign node20 = (inp[5]) ? 3'b010 : node21;
											assign node21 = (inp[2]) ? 3'b000 : 3'b100;
										assign node25 = (inp[11]) ? node27 : 3'b100;
											assign node27 = (inp[5]) ? 3'b100 : 3'b000;
								assign node30 = (inp[2]) ? node32 : 3'b000;
									assign node32 = (inp[8]) ? 3'b000 : node33;
										assign node33 = (inp[10]) ? node37 : node34;
											assign node34 = (inp[11]) ? 3'b000 : 3'b100;
											assign node37 = (inp[5]) ? 3'b010 : 3'b000;
							assign node41 = (inp[5]) ? node65 : node42;
								assign node42 = (inp[9]) ? node52 : node43;
									assign node43 = (inp[8]) ? 3'b100 : node44;
										assign node44 = (inp[11]) ? node48 : node45;
											assign node45 = (inp[10]) ? 3'b000 : 3'b100;
											assign node48 = (inp[10]) ? 3'b100 : 3'b000;
									assign node52 = (inp[2]) ? node58 : node53;
										assign node53 = (inp[11]) ? 3'b100 : node54;
											assign node54 = (inp[10]) ? 3'b000 : 3'b000;
										assign node58 = (inp[11]) ? node62 : node59;
											assign node59 = (inp[8]) ? 3'b000 : 3'b000;
											assign node62 = (inp[8]) ? 3'b010 : 3'b010;
								assign node65 = (inp[9]) ? node73 : node66;
									assign node66 = (inp[8]) ? node70 : node67;
										assign node67 = (inp[10]) ? 3'b010 : 3'b100;
										assign node70 = (inp[10]) ? 3'b100 : 3'b000;
									assign node73 = (inp[2]) ? node81 : node74;
										assign node74 = (inp[8]) ? node78 : node75;
											assign node75 = (inp[10]) ? 3'b110 : 3'b010;
											assign node78 = (inp[10]) ? 3'b010 : 3'b100;
										assign node81 = (inp[10]) ? node85 : node82;
											assign node82 = (inp[8]) ? 3'b010 : 3'b110;
											assign node85 = (inp[8]) ? 3'b110 : 3'b001;
						assign node88 = (inp[2]) ? node90 : 3'b000;
							assign node90 = (inp[1]) ? node92 : 3'b000;
								assign node92 = (inp[8]) ? 3'b000 : node93;
									assign node93 = (inp[9]) ? node95 : 3'b000;
										assign node95 = (inp[10]) ? node99 : node96;
											assign node96 = (inp[5]) ? 3'b100 : 3'b000;
											assign node99 = (inp[5]) ? 3'b010 : 3'b000;
		assign node104 = (inp[0]) ? node268 : node105;
			assign node105 = (inp[6]) ? node253 : node106;
				assign node106 = (inp[4]) ? node142 : node107;
					assign node107 = (inp[7]) ? 3'b000 : node108;
						assign node108 = (inp[9]) ? node110 : 3'b000;
							assign node110 = (inp[1]) ? node120 : node111;
								assign node111 = (inp[2]) ? node113 : 3'b000;
									assign node113 = (inp[11]) ? node115 : 3'b000;
										assign node115 = (inp[10]) ? node117 : 3'b000;
											assign node117 = (inp[8]) ? 3'b000 : 3'b100;
								assign node120 = (inp[5]) ? node128 : node121;
									assign node121 = (inp[10]) ? node123 : 3'b000;
										assign node123 = (inp[8]) ? 3'b000 : node124;
											assign node124 = (inp[2]) ? 3'b100 : 3'b000;
									assign node128 = (inp[10]) ? node136 : node129;
										assign node129 = (inp[8]) ? node133 : node130;
											assign node130 = (inp[2]) ? 3'b000 : 3'b100;
											assign node133 = (inp[11]) ? 3'b100 : 3'b000;
										assign node136 = (inp[8]) ? node138 : 3'b010;
											assign node138 = (inp[2]) ? 3'b000 : 3'b000;
					assign node142 = (inp[7]) ? node220 : node143;
						assign node143 = (inp[1]) ? node171 : node144;
							assign node144 = (inp[9]) ? node146 : 3'b000;
								assign node146 = (inp[2]) ? node156 : node147;
									assign node147 = (inp[5]) ? node149 : 3'b000;
										assign node149 = (inp[10]) ? node153 : node150;
											assign node150 = (inp[8]) ? 3'b000 : 3'b100;
											assign node153 = (inp[8]) ? 3'b100 : 3'b010;
									assign node156 = (inp[10]) ? node164 : node157;
										assign node157 = (inp[8]) ? node161 : node158;
											assign node158 = (inp[5]) ? 3'b010 : 3'b000;
											assign node161 = (inp[5]) ? 3'b100 : 3'b110;
										assign node164 = (inp[8]) ? node168 : node165;
											assign node165 = (inp[5]) ? 3'b110 : 3'b010;
											assign node168 = (inp[5]) ? 3'b010 : 3'b000;
							assign node171 = (inp[9]) ? node193 : node172;
								assign node172 = (inp[10]) ? node180 : node173;
									assign node173 = (inp[5]) ? node175 : 3'b100;
										assign node175 = (inp[8]) ? 3'b100 : node176;
											assign node176 = (inp[2]) ? 3'b110 : 3'b100;
									assign node180 = (inp[5]) ? node186 : node181;
										assign node181 = (inp[8]) ? 3'b100 : node182;
											assign node182 = (inp[2]) ? 3'b110 : 3'b100;
										assign node186 = (inp[8]) ? node190 : node187;
											assign node187 = (inp[2]) ? 3'b100 : 3'b110;
											assign node190 = (inp[2]) ? 3'b110 : 3'b100;
								assign node193 = (inp[2]) ? node205 : node194;
									assign node194 = (inp[10]) ? node200 : node195;
										assign node195 = (inp[8]) ? node197 : 3'b110;
											assign node197 = (inp[5]) ? 3'b010 : 3'b000;
										assign node200 = (inp[11]) ? node202 : 3'b110;
											assign node202 = (inp[8]) ? 3'b110 : 3'b100;
									assign node205 = (inp[5]) ? node213 : node206;
										assign node206 = (inp[10]) ? node210 : node207;
											assign node207 = (inp[8]) ? 3'b010 : 3'b110;
											assign node210 = (inp[8]) ? 3'b110 : 3'b001;
										assign node213 = (inp[10]) ? node217 : node214;
											assign node214 = (inp[8]) ? 3'b000 : 3'b001;
											assign node217 = (inp[11]) ? 3'b001 : 3'b001;
						assign node220 = (inp[9]) ? node222 : 3'b000;
							assign node222 = (inp[1]) ? node232 : node223;
								assign node223 = (inp[2]) ? node225 : 3'b000;
									assign node225 = (inp[10]) ? node227 : 3'b000;
										assign node227 = (inp[8]) ? 3'b000 : node228;
											assign node228 = (inp[5]) ? 3'b100 : 3'b000;
								assign node232 = (inp[10]) ? node240 : node233;
									assign node233 = (inp[5]) ? 3'b100 : node234;
										assign node234 = (inp[11]) ? node236 : 3'b000;
											assign node236 = (inp[8]) ? 3'b000 : 3'b100;
									assign node240 = (inp[2]) ? node248 : node241;
										assign node241 = (inp[8]) ? node245 : node242;
											assign node242 = (inp[5]) ? 3'b010 : 3'b100;
											assign node245 = (inp[5]) ? 3'b100 : 3'b000;
										assign node248 = (inp[8]) ? 3'b010 : node249;
											assign node249 = (inp[11]) ? 3'b010 : 3'b100;
				assign node253 = (inp[10]) ? node255 : 3'b000;
					assign node255 = (inp[8]) ? 3'b000 : node256;
						assign node256 = (inp[4]) ? node258 : 3'b000;
							assign node258 = (inp[5]) ? node260 : 3'b000;
								assign node260 = (inp[1]) ? node262 : 3'b000;
									assign node262 = (inp[2]) ? node264 : 3'b000;
										assign node264 = (inp[7]) ? 3'b000 : 3'b100;
			assign node268 = (inp[6]) ? node664 : node269;
				assign node269 = (inp[7]) ? node477 : node270;
					assign node270 = (inp[4]) ? node378 : node271;
						assign node271 = (inp[11]) ? node331 : node272;
							assign node272 = (inp[1]) ? node302 : node273;
								assign node273 = (inp[9]) ? node287 : node274;
									assign node274 = (inp[2]) ? node282 : node275;
										assign node275 = (inp[10]) ? node279 : node276;
											assign node276 = (inp[5]) ? 3'b000 : 3'b000;
											assign node279 = (inp[8]) ? 3'b001 : 3'b100;
										assign node282 = (inp[5]) ? 3'b010 : node283;
											assign node283 = (inp[10]) ? 3'b001 : 3'b000;
									assign node287 = (inp[10]) ? node295 : node288;
										assign node288 = (inp[5]) ? node292 : node289;
											assign node289 = (inp[2]) ? 3'b000 : 3'b000;
											assign node292 = (inp[2]) ? 3'b010 : 3'b000;
										assign node295 = (inp[8]) ? node299 : node296;
											assign node296 = (inp[2]) ? 3'b100 : 3'b110;
											assign node299 = (inp[5]) ? 3'b010 : 3'b000;
								assign node302 = (inp[2]) ? node316 : node303;
									assign node303 = (inp[5]) ? node309 : node304;
										assign node304 = (inp[8]) ? node306 : 3'b110;
											assign node306 = (inp[10]) ? 3'b000 : 3'b010;
										assign node309 = (inp[9]) ? node313 : node310;
											assign node310 = (inp[8]) ? 3'b000 : 3'b000;
											assign node313 = (inp[8]) ? 3'b101 : 3'b011;
									assign node316 = (inp[9]) ? node324 : node317;
										assign node317 = (inp[10]) ? node321 : node318;
											assign node318 = (inp[5]) ? 3'b101 : 3'b000;
											assign node321 = (inp[8]) ? 3'b010 : 3'b100;
										assign node324 = (inp[5]) ? node328 : node325;
											assign node325 = (inp[10]) ? 3'b001 : 3'b001;
											assign node328 = (inp[8]) ? 3'b001 : 3'b011;
							assign node331 = (inp[8]) ? node355 : node332;
								assign node332 = (inp[9]) ? node340 : node333;
									assign node333 = (inp[5]) ? node337 : node334;
										assign node334 = (inp[10]) ? 3'b001 : 3'b101;
										assign node337 = (inp[10]) ? 3'b101 : 3'b001;
									assign node340 = (inp[1]) ? node348 : node341;
										assign node341 = (inp[2]) ? node345 : node342;
											assign node342 = (inp[10]) ? 3'b110 : 3'b100;
											assign node345 = (inp[5]) ? 3'b001 : 3'b001;
										assign node348 = (inp[5]) ? node352 : node349;
											assign node349 = (inp[2]) ? 3'b001 : 3'b001;
											assign node352 = (inp[2]) ? 3'b011 : 3'b001;
								assign node355 = (inp[10]) ? node367 : node356;
									assign node356 = (inp[9]) ? node360 : node357;
										assign node357 = (inp[5]) ? 3'b110 : 3'b010;
										assign node360 = (inp[1]) ? node364 : node361;
											assign node361 = (inp[5]) ? 3'b010 : 3'b100;
											assign node364 = (inp[2]) ? 3'b101 : 3'b001;
									assign node367 = (inp[9]) ? node371 : node368;
										assign node368 = (inp[5]) ? 3'b001 : 3'b101;
										assign node371 = (inp[1]) ? node375 : node372;
											assign node372 = (inp[2]) ? 3'b000 : 3'b110;
											assign node375 = (inp[5]) ? 3'b101 : 3'b001;
						assign node378 = (inp[2]) ? node434 : node379;
							assign node379 = (inp[1]) ? node407 : node380;
								assign node380 = (inp[9]) ? node392 : node381;
									assign node381 = (inp[10]) ? node387 : node382;
										assign node382 = (inp[11]) ? 3'b101 : node383;
											assign node383 = (inp[8]) ? 3'b101 : 3'b101;
										assign node387 = (inp[8]) ? node389 : 3'b111;
											assign node389 = (inp[11]) ? 3'b101 : 3'b111;
									assign node392 = (inp[5]) ? node400 : node393;
										assign node393 = (inp[8]) ? node397 : node394;
											assign node394 = (inp[10]) ? 3'b101 : 3'b001;
											assign node397 = (inp[10]) ? 3'b001 : 3'b110;
										assign node400 = (inp[8]) ? node404 : node401;
											assign node401 = (inp[10]) ? 3'b011 : 3'b011;
											assign node404 = (inp[11]) ? 3'b101 : 3'b001;
								assign node407 = (inp[9]) ? node421 : node408;
									assign node408 = (inp[5]) ? node414 : node409;
										assign node409 = (inp[11]) ? 3'b011 : node410;
											assign node410 = (inp[8]) ? 3'b001 : 3'b011;
										assign node414 = (inp[11]) ? node418 : node415;
											assign node415 = (inp[8]) ? 3'b001 : 3'b001;
											assign node418 = (inp[10]) ? 3'b001 : 3'b001;
									assign node421 = (inp[11]) ? node429 : node422;
										assign node422 = (inp[8]) ? node426 : node423;
											assign node423 = (inp[5]) ? 3'b111 : 3'b011;
											assign node426 = (inp[10]) ? 3'b011 : 3'b001;
										assign node429 = (inp[5]) ? 3'b111 : node430;
											assign node430 = (inp[8]) ? 3'b011 : 3'b111;
							assign node434 = (inp[9]) ? node458 : node435;
								assign node435 = (inp[8]) ? node449 : node436;
									assign node436 = (inp[10]) ? node442 : node437;
										assign node437 = (inp[11]) ? 3'b111 : node438;
											assign node438 = (inp[5]) ? 3'b101 : 3'b111;
										assign node442 = (inp[1]) ? node446 : node443;
											assign node443 = (inp[5]) ? 3'b101 : 3'b101;
											assign node446 = (inp[11]) ? 3'b111 : 3'b101;
									assign node449 = (inp[10]) ? node455 : node450;
										assign node450 = (inp[11]) ? 3'b101 : node451;
											assign node451 = (inp[1]) ? 3'b101 : 3'b101;
										assign node455 = (inp[11]) ? 3'b111 : 3'b101;
								assign node458 = (inp[1]) ? node472 : node459;
									assign node459 = (inp[8]) ? node465 : node460;
										assign node460 = (inp[5]) ? 3'b111 : node461;
											assign node461 = (inp[11]) ? 3'b011 : 3'b001;
										assign node465 = (inp[5]) ? node469 : node466;
											assign node466 = (inp[10]) ? 3'b101 : 3'b001;
											assign node469 = (inp[11]) ? 3'b011 : 3'b001;
									assign node472 = (inp[5]) ? 3'b111 : node473;
										assign node473 = (inp[11]) ? 3'b111 : 3'b011;
					assign node477 = (inp[4]) ? node567 : node478;
						assign node478 = (inp[9]) ? node514 : node479;
							assign node479 = (inp[10]) ? node485 : node480;
								assign node480 = (inp[11]) ? node482 : 3'b110;
									assign node482 = (inp[8]) ? 3'b110 : 3'b010;
								assign node485 = (inp[1]) ? node501 : node486;
									assign node486 = (inp[2]) ? node494 : node487;
										assign node487 = (inp[8]) ? node491 : node488;
											assign node488 = (inp[11]) ? 3'b110 : 3'b010;
											assign node491 = (inp[11]) ? 3'b010 : 3'b110;
										assign node494 = (inp[8]) ? node498 : node495;
											assign node495 = (inp[11]) ? 3'b110 : 3'b010;
											assign node498 = (inp[11]) ? 3'b010 : 3'b110;
									assign node501 = (inp[5]) ? node507 : node502;
										assign node502 = (inp[2]) ? 3'b010 : node503;
											assign node503 = (inp[11]) ? 3'b010 : 3'b010;
										assign node507 = (inp[11]) ? node511 : node508;
											assign node508 = (inp[8]) ? 3'b110 : 3'b010;
											assign node511 = (inp[8]) ? 3'b010 : 3'b110;
							assign node514 = (inp[1]) ? node538 : node515;
								assign node515 = (inp[2]) ? node523 : node516;
									assign node516 = (inp[5]) ? node518 : 3'b000;
										assign node518 = (inp[11]) ? 3'b000 : node519;
											assign node519 = (inp[10]) ? 3'b100 : 3'b000;
									assign node523 = (inp[8]) ? node531 : node524;
										assign node524 = (inp[5]) ? node528 : node525;
											assign node525 = (inp[11]) ? 3'b000 : 3'b100;
											assign node528 = (inp[11]) ? 3'b010 : 3'b010;
										assign node531 = (inp[10]) ? node535 : node532;
											assign node532 = (inp[5]) ? 3'b100 : 3'b110;
											assign node535 = (inp[11]) ? 3'b000 : 3'b100;
								assign node538 = (inp[5]) ? node552 : node539;
									assign node539 = (inp[2]) ? node545 : node540;
										assign node540 = (inp[11]) ? 3'b100 : node541;
											assign node541 = (inp[8]) ? 3'b100 : 3'b000;
										assign node545 = (inp[8]) ? node549 : node546;
											assign node546 = (inp[11]) ? 3'b110 : 3'b010;
											assign node549 = (inp[10]) ? 3'b010 : 3'b100;
									assign node552 = (inp[2]) ? node560 : node553;
										assign node553 = (inp[11]) ? node557 : node554;
											assign node554 = (inp[8]) ? 3'b010 : 3'b010;
											assign node557 = (inp[10]) ? 3'b000 : 3'b100;
										assign node560 = (inp[10]) ? node564 : node561;
											assign node561 = (inp[11]) ? 3'b000 : 3'b110;
											assign node564 = (inp[8]) ? 3'b001 : 3'b101;
						assign node567 = (inp[5]) ? node623 : node568;
							assign node568 = (inp[1]) ? node596 : node569;
								assign node569 = (inp[2]) ? node583 : node570;
									assign node570 = (inp[10]) ? node576 : node571;
										assign node571 = (inp[9]) ? 3'b010 : node572;
											assign node572 = (inp[8]) ? 3'b010 : 3'b010;
										assign node576 = (inp[9]) ? node580 : node577;
											assign node577 = (inp[8]) ? 3'b010 : 3'b001;
											assign node580 = (inp[8]) ? 3'b000 : 3'b110;
									assign node583 = (inp[8]) ? node589 : node584;
										assign node584 = (inp[10]) ? node586 : 3'b110;
											assign node586 = (inp[11]) ? 3'b001 : 3'b000;
										assign node589 = (inp[10]) ? node593 : node590;
											assign node590 = (inp[11]) ? 3'b010 : 3'b000;
											assign node593 = (inp[11]) ? 3'b110 : 3'b010;
								assign node596 = (inp[9]) ? node612 : node597;
									assign node597 = (inp[11]) ? node605 : node598;
										assign node598 = (inp[8]) ? node602 : node599;
											assign node599 = (inp[10]) ? 3'b100 : 3'b010;
											assign node602 = (inp[10]) ? 3'b010 : 3'b000;
										assign node605 = (inp[8]) ? node609 : node606;
											assign node606 = (inp[10]) ? 3'b001 : 3'b110;
											assign node609 = (inp[10]) ? 3'b110 : 3'b010;
									assign node612 = (inp[10]) ? node618 : node613;
										assign node613 = (inp[11]) ? 3'b001 : node614;
											assign node614 = (inp[8]) ? 3'b000 : 3'b001;
										assign node618 = (inp[11]) ? 3'b101 : node619;
											assign node619 = (inp[2]) ? 3'b001 : 3'b001;
							assign node623 = (inp[8]) ? node645 : node624;
								assign node624 = (inp[9]) ? node632 : node625;
									assign node625 = (inp[11]) ? node629 : node626;
										assign node626 = (inp[10]) ? 3'b101 : 3'b001;
										assign node629 = (inp[10]) ? 3'b011 : 3'b101;
									assign node632 = (inp[1]) ? node640 : node633;
										assign node633 = (inp[11]) ? node637 : node634;
											assign node634 = (inp[2]) ? 3'b001 : 3'b110;
											assign node637 = (inp[2]) ? 3'b011 : 3'b001;
										assign node640 = (inp[2]) ? 3'b111 : node641;
											assign node641 = (inp[11]) ? 3'b011 : 3'b001;
								assign node645 = (inp[10]) ? node653 : node646;
									assign node646 = (inp[9]) ? node648 : 3'b010;
										assign node648 = (inp[1]) ? node650 : 3'b010;
											assign node650 = (inp[11]) ? 3'b101 : 3'b001;
									assign node653 = (inp[9]) ? node657 : node654;
										assign node654 = (inp[11]) ? 3'b101 : 3'b001;
										assign node657 = (inp[2]) ? node661 : node658;
											assign node658 = (inp[1]) ? 3'b011 : 3'b110;
											assign node661 = (inp[1]) ? 3'b011 : 3'b001;
				assign node664 = (inp[4]) ? node692 : node665;
					assign node665 = (inp[7]) ? 3'b000 : node666;
						assign node666 = (inp[1]) ? node668 : 3'b000;
							assign node668 = (inp[9]) ? node670 : 3'b000;
								assign node670 = (inp[10]) ? node678 : node671;
									assign node671 = (inp[2]) ? node673 : 3'b000;
										assign node673 = (inp[8]) ? 3'b000 : node674;
											assign node674 = (inp[5]) ? 3'b010 : 3'b000;
									assign node678 = (inp[2]) ? node684 : node679;
										assign node679 = (inp[5]) ? node681 : 3'b000;
											assign node681 = (inp[8]) ? 3'b000 : 3'b100;
										assign node684 = (inp[5]) ? node688 : node685;
											assign node685 = (inp[8]) ? 3'b000 : 3'b100;
											assign node688 = (inp[8]) ? 3'b100 : 3'b010;
					assign node692 = (inp[7]) ? node776 : node693;
						assign node693 = (inp[10]) ? node735 : node694;
							assign node694 = (inp[9]) ? node710 : node695;
								assign node695 = (inp[11]) ? node703 : node696;
									assign node696 = (inp[8]) ? node700 : node697;
										assign node697 = (inp[5]) ? 3'b010 : 3'b100;
										assign node700 = (inp[5]) ? 3'b100 : 3'b110;
									assign node703 = (inp[8]) ? node707 : node704;
										assign node704 = (inp[5]) ? 3'b110 : 3'b100;
										assign node707 = (inp[5]) ? 3'b100 : 3'b000;
								assign node710 = (inp[1]) ? node722 : node711;
									assign node711 = (inp[11]) ? node717 : node712;
										assign node712 = (inp[5]) ? node714 : 3'b000;
											assign node714 = (inp[2]) ? 3'b100 : 3'b000;
										assign node717 = (inp[2]) ? node719 : 3'b100;
											assign node719 = (inp[5]) ? 3'b000 : 3'b000;
									assign node722 = (inp[11]) ? node730 : node723;
										assign node723 = (inp[5]) ? node727 : node724;
											assign node724 = (inp[2]) ? 3'b100 : 3'b000;
											assign node727 = (inp[2]) ? 3'b000 : 3'b110;
										assign node730 = (inp[8]) ? node732 : 3'b010;
											assign node732 = (inp[2]) ? 3'b010 : 3'b010;
							assign node735 = (inp[8]) ? node759 : node736;
								assign node736 = (inp[5]) ? node746 : node737;
									assign node737 = (inp[9]) ? node739 : 3'b010;
										assign node739 = (inp[2]) ? node743 : node740;
											assign node740 = (inp[1]) ? 3'b010 : 3'b100;
											assign node743 = (inp[1]) ? 3'b001 : 3'b000;
									assign node746 = (inp[1]) ? node754 : node747;
										assign node747 = (inp[9]) ? node751 : node748;
											assign node748 = (inp[11]) ? 3'b001 : 3'b110;
											assign node751 = (inp[2]) ? 3'b110 : 3'b010;
										assign node754 = (inp[2]) ? node756 : 3'b001;
											assign node756 = (inp[11]) ? 3'b011 : 3'b100;
								assign node759 = (inp[5]) ? node767 : node760;
									assign node760 = (inp[11]) ? node762 : 3'b000;
										assign node762 = (inp[9]) ? node764 : 3'b100;
											assign node764 = (inp[2]) ? 3'b100 : 3'b010;
									assign node767 = (inp[9]) ? node769 : 3'b010;
										assign node769 = (inp[2]) ? node773 : node770;
											assign node770 = (inp[1]) ? 3'b110 : 3'b100;
											assign node773 = (inp[1]) ? 3'b001 : 3'b010;
						assign node776 = (inp[10]) ? node790 : node777;
							assign node777 = (inp[9]) ? node779 : 3'b000;
								assign node779 = (inp[5]) ? node781 : 3'b000;
									assign node781 = (inp[1]) ? node783 : 3'b000;
										assign node783 = (inp[2]) ? node787 : node784;
											assign node784 = (inp[8]) ? 3'b000 : 3'b100;
											assign node787 = (inp[8]) ? 3'b100 : 3'b010;
							assign node790 = (inp[8]) ? node808 : node791;
								assign node791 = (inp[5]) ? node799 : node792;
									assign node792 = (inp[1]) ? node794 : 3'b000;
										assign node794 = (inp[9]) ? node796 : 3'b000;
											assign node796 = (inp[11]) ? 3'b010 : 3'b000;
									assign node799 = (inp[9]) ? node801 : 3'b100;
										assign node801 = (inp[2]) ? node805 : node802;
											assign node802 = (inp[1]) ? 3'b010 : 3'b000;
											assign node805 = (inp[1]) ? 3'b110 : 3'b100;
								assign node808 = (inp[9]) ? node810 : 3'b000;
									assign node810 = (inp[1]) ? node812 : 3'b000;
										assign node812 = (inp[11]) ? node814 : 3'b000;
											assign node814 = (inp[5]) ? 3'b000 : 3'b000;

endmodule