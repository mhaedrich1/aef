module dtc_split875_bm28 (
	input  wire [7-1:0] inp,
	output wire [10-1:0] outp
);

	wire [10-1:0] node1;
	wire [10-1:0] node2;
	wire [10-1:0] node3;
	wire [10-1:0] node4;
	wire [10-1:0] node5;
	wire [10-1:0] node6;
	wire [10-1:0] node9;
	wire [10-1:0] node12;
	wire [10-1:0] node13;
	wire [10-1:0] node17;
	wire [10-1:0] node18;
	wire [10-1:0] node19;
	wire [10-1:0] node22;
	wire [10-1:0] node25;
	wire [10-1:0] node26;
	wire [10-1:0] node29;
	wire [10-1:0] node32;
	wire [10-1:0] node33;
	wire [10-1:0] node34;
	wire [10-1:0] node35;
	wire [10-1:0] node38;
	wire [10-1:0] node41;
	wire [10-1:0] node42;
	wire [10-1:0] node45;
	wire [10-1:0] node48;
	wire [10-1:0] node49;
	wire [10-1:0] node50;
	wire [10-1:0] node54;
	wire [10-1:0] node55;
	wire [10-1:0] node58;
	wire [10-1:0] node61;
	wire [10-1:0] node62;
	wire [10-1:0] node63;
	wire [10-1:0] node64;
	wire [10-1:0] node65;
	wire [10-1:0] node68;
	wire [10-1:0] node71;
	wire [10-1:0] node72;
	wire [10-1:0] node76;
	wire [10-1:0] node77;
	wire [10-1:0] node78;
	wire [10-1:0] node81;
	wire [10-1:0] node84;
	wire [10-1:0] node85;
	wire [10-1:0] node89;
	wire [10-1:0] node90;
	wire [10-1:0] node91;
	wire [10-1:0] node92;
	wire [10-1:0] node96;
	wire [10-1:0] node97;
	wire [10-1:0] node100;
	wire [10-1:0] node103;
	wire [10-1:0] node104;
	wire [10-1:0] node105;
	wire [10-1:0] node108;
	wire [10-1:0] node111;
	wire [10-1:0] node112;
	wire [10-1:0] node115;
	wire [10-1:0] node118;
	wire [10-1:0] node119;
	wire [10-1:0] node120;
	wire [10-1:0] node121;
	wire [10-1:0] node122;
	wire [10-1:0] node123;
	wire [10-1:0] node126;
	wire [10-1:0] node129;
	wire [10-1:0] node130;
	wire [10-1:0] node133;
	wire [10-1:0] node136;
	wire [10-1:0] node137;
	wire [10-1:0] node138;
	wire [10-1:0] node141;
	wire [10-1:0] node144;
	wire [10-1:0] node146;
	wire [10-1:0] node149;
	wire [10-1:0] node150;
	wire [10-1:0] node151;
	wire [10-1:0] node152;
	wire [10-1:0] node156;
	wire [10-1:0] node158;
	wire [10-1:0] node161;
	wire [10-1:0] node162;
	wire [10-1:0] node163;
	wire [10-1:0] node166;
	wire [10-1:0] node169;
	wire [10-1:0] node171;
	wire [10-1:0] node174;
	wire [10-1:0] node175;
	wire [10-1:0] node176;
	wire [10-1:0] node177;
	wire [10-1:0] node178;
	wire [10-1:0] node181;
	wire [10-1:0] node184;
	wire [10-1:0] node186;
	wire [10-1:0] node189;
	wire [10-1:0] node190;
	wire [10-1:0] node191;
	wire [10-1:0] node194;
	wire [10-1:0] node197;
	wire [10-1:0] node200;
	wire [10-1:0] node201;
	wire [10-1:0] node202;
	wire [10-1:0] node204;
	wire [10-1:0] node207;
	wire [10-1:0] node208;
	wire [10-1:0] node211;
	wire [10-1:0] node214;
	wire [10-1:0] node215;
	wire [10-1:0] node218;
	wire [10-1:0] node220;

	assign outp = (inp[4]) ? node118 : node1;
		assign node1 = (inp[2]) ? node61 : node2;
			assign node2 = (inp[5]) ? node32 : node3;
				assign node3 = (inp[3]) ? node17 : node4;
					assign node4 = (inp[6]) ? node12 : node5;
						assign node5 = (inp[1]) ? node9 : node6;
							assign node6 = (inp[0]) ? 10'b0101011001 : 10'b0001111101;
							assign node9 = (inp[0]) ? 10'b0011110001 : 10'b0001010101;
						assign node12 = (inp[1]) ? 10'b0111010000 : node13;
							assign node13 = (inp[0]) ? 10'b0011011000 : 10'b0111111000;
					assign node17 = (inp[1]) ? node25 : node18;
						assign node18 = (inp[6]) ? node22 : node19;
							assign node19 = (inp[0]) ? 10'b0101000001 : 10'b0001100101;
							assign node22 = (inp[0]) ? 10'b0011000000 : 10'b0111100000;
						assign node25 = (inp[6]) ? node29 : node26;
							assign node26 = (inp[0]) ? 10'b0011101000 : 10'b0001001100;
							assign node29 = (inp[0]) ? 10'b0001001001 : 10'b0101101001;
				assign node32 = (inp[3]) ? node48 : node33;
					assign node33 = (inp[6]) ? node41 : node34;
						assign node34 = (inp[1]) ? node38 : node35;
							assign node35 = (inp[0]) ? 10'b0100011000 : 10'b0000111100;
							assign node38 = (inp[0]) ? 10'b0010110000 : 10'b0000010100;
						assign node41 = (inp[1]) ? node45 : node42;
							assign node42 = (inp[0]) ? 10'b0000111001 : 10'b0110011001;
							assign node45 = (inp[0]) ? 10'b0000010001 : 10'b0100110001;
					assign node48 = (inp[1]) ? node54 : node49;
						assign node49 = (inp[6]) ? 10'b0000100001 : node50;
							assign node50 = (inp[0]) ? 10'b0100000000 : 10'b0000100100;
						assign node54 = (inp[6]) ? node58 : node55;
							assign node55 = (inp[0]) ? 10'b0010001001 : 10'b0110101001;
							assign node58 = (inp[0]) ? 10'b0000001000 : 10'b0100101000;
			assign node61 = (inp[3]) ? node89 : node62;
				assign node62 = (inp[5]) ? node76 : node63;
					assign node63 = (inp[6]) ? node71 : node64;
						assign node64 = (inp[1]) ? node68 : node65;
							assign node65 = (inp[0]) ? 10'b1100001001 : 10'b1000101101;
							assign node68 = (inp[0]) ? 10'b1010100001 : 10'b1000000101;
						assign node71 = (inp[1]) ? 10'b1110000000 : node72;
							assign node72 = (inp[0]) ? 10'b1010001000 : 10'b1110101000;
					assign node76 = (inp[1]) ? node84 : node77;
						assign node77 = (inp[6]) ? node81 : node78;
							assign node78 = (inp[0]) ? 10'b1101000000 : 10'b1001100100;
							assign node81 = (inp[0]) ? 10'b1001100001 : 10'b1111000001;
						assign node84 = (inp[6]) ? 10'b1101101000 : node85;
							assign node85 = (inp[0]) ? 10'b1011001001 : 10'b1111101001;
				assign node89 = (inp[5]) ? node103 : node90;
					assign node90 = (inp[6]) ? node96 : node91;
						assign node91 = (inp[0]) ? 10'b1011110000 : node92;
							assign node92 = (inp[1]) ? 10'b1001010100 : 10'b1001111100;
						assign node96 = (inp[1]) ? node100 : node97;
							assign node97 = (inp[0]) ? 10'b1001111001 : 10'b1111011001;
							assign node100 = (inp[0]) ? 10'b1001010001 : 10'b1101110001;
					assign node103 = (inp[6]) ? node111 : node104;
						assign node104 = (inp[1]) ? node108 : node105;
							assign node105 = (inp[0]) ? 10'b1010111001 : 10'b1000011101;
							assign node108 = (inp[0]) ? 10'b1010010001 : 10'b1110110001;
						assign node111 = (inp[0]) ? node115 : node112;
							assign node112 = (inp[1]) ? 10'b1100110000 : 10'b1110011000;
							assign node115 = (inp[1]) ? 10'b1000010000 : 10'b1000111000;
		assign node118 = (inp[2]) ? node174 : node119;
			assign node119 = (inp[3]) ? node149 : node120;
				assign node120 = (inp[5]) ? node136 : node121;
					assign node121 = (inp[6]) ? node129 : node122;
						assign node122 = (inp[1]) ? node126 : node123;
							assign node123 = (inp[0]) ? 10'b1100011011 : 10'b1000111111;
							assign node126 = (inp[0]) ? 10'b1010110011 : 10'b1000010111;
						assign node129 = (inp[0]) ? node133 : node130;
							assign node130 = (inp[1]) ? 10'b1110010010 : 10'b1110111010;
							assign node133 = (inp[1]) ? 10'b1000110010 : 10'b1010011010;
					assign node136 = (inp[1]) ? node144 : node137;
						assign node137 = (inp[6]) ? node141 : node138;
							assign node138 = (inp[0]) ? 10'b1101010010 : 10'b1001110110;
							assign node141 = (inp[0]) ? 10'b1001110011 : 10'b1111010011;
						assign node144 = (inp[0]) ? node146 : 10'b1101111010;
							assign node146 = (inp[6]) ? 10'b1001011010 : 10'b1011011011;
				assign node149 = (inp[5]) ? node161 : node150;
					assign node150 = (inp[0]) ? node156 : node151;
						assign node151 = (inp[6]) ? 10'b1100101011 : node152;
							assign node152 = (inp[1]) ? 10'b1000001110 : 10'b1000100111;
						assign node156 = (inp[1]) ? node158 : 10'b1010000010;
							assign node158 = (inp[6]) ? 10'b1000001011 : 10'b1010101010;
					assign node161 = (inp[6]) ? node169 : node162;
						assign node162 = (inp[1]) ? node166 : node163;
							assign node163 = (inp[0]) ? 10'b1011101011 : 10'b1001001111;
							assign node166 = (inp[0]) ? 10'b1011000011 : 10'b1111100011;
						assign node169 = (inp[0]) ? node171 : 10'b1111001010;
							assign node171 = (inp[1]) ? 10'b1001000010 : 10'b1001101010;
			assign node174 = (inp[5]) ? node200 : node175;
				assign node175 = (inp[3]) ? node189 : node176;
					assign node176 = (inp[1]) ? node184 : node177;
						assign node177 = (inp[6]) ? node181 : node178;
							assign node178 = (inp[0]) ? 10'b0101010011 : 10'b0001110111;
							assign node181 = (inp[0]) ? 10'b0011010010 : 10'b0111110010;
						assign node184 = (inp[6]) ? node186 : 10'b0001011110;
							assign node186 = (inp[0]) ? 10'b0001011011 : 10'b0101111011;
					assign node189 = (inp[6]) ? node197 : node190;
						assign node190 = (inp[1]) ? node194 : node191;
							assign node191 = (inp[0]) ? 10'b0101001010 : 10'b0001101110;
							assign node194 = (inp[0]) ? 10'b0011100010 : 10'b0001000110;
						assign node197 = (inp[0]) ? 10'b0001101011 : 10'b0111001011;
				assign node200 = (inp[3]) ? node214 : node201;
					assign node201 = (inp[1]) ? node207 : node202;
						assign node202 = (inp[6]) ? node204 : 10'b0100010010;
							assign node204 = (inp[0]) ? 10'b0000110011 : 10'b0110010011;
						assign node207 = (inp[0]) ? node211 : node208;
							assign node208 = (inp[6]) ? 10'b0100111010 : 10'b0110111011;
							assign node211 = (inp[6]) ? 10'b0000011010 : 10'b0010011011;
					assign node214 = (inp[6]) ? node218 : node215;
						assign node215 = (inp[0]) ? 10'b0010000011 : 10'b0110100011;
						assign node218 = (inp[1]) ? node220 : 10'b0110001010;
							assign node220 = (inp[0]) ? 10'b0000000010 : 10'b0100100010;

endmodule