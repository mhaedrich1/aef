module dtc_split66_bm73 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node260;
	wire [3-1:0] node263;
	wire [3-1:0] node265;
	wire [3-1:0] node268;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node281;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node302;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node316;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node341;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node348;
	wire [3-1:0] node350;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node430;
	wire [3-1:0] node432;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node442;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node448;
	wire [3-1:0] node451;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node474;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node493;
	wire [3-1:0] node495;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node517;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node524;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node542;
	wire [3-1:0] node545;
	wire [3-1:0] node547;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node555;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node562;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node569;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node576;
	wire [3-1:0] node579;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node587;
	wire [3-1:0] node590;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node604;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node628;
	wire [3-1:0] node630;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node649;
	wire [3-1:0] node652;
	wire [3-1:0] node653;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node661;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node668;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node681;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node692;
	wire [3-1:0] node695;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node704;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node718;
	wire [3-1:0] node721;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node734;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node780;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node788;
	wire [3-1:0] node790;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node812;
	wire [3-1:0] node815;
	wire [3-1:0] node817;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node833;
	wire [3-1:0] node834;
	wire [3-1:0] node837;
	wire [3-1:0] node840;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node843;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node851;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node858;
	wire [3-1:0] node860;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node870;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node878;
	wire [3-1:0] node881;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node888;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node901;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node908;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node915;
	wire [3-1:0] node919;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node926;
	wire [3-1:0] node929;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node932;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node941;
	wire [3-1:0] node942;
	wire [3-1:0] node944;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node951;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node965;
	wire [3-1:0] node966;
	wire [3-1:0] node970;
	wire [3-1:0] node971;
	wire [3-1:0] node972;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node984;
	wire [3-1:0] node986;
	wire [3-1:0] node989;
	wire [3-1:0] node990;
	wire [3-1:0] node992;
	wire [3-1:0] node995;
	wire [3-1:0] node998;
	wire [3-1:0] node1000;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1009;
	wire [3-1:0] node1011;
	wire [3-1:0] node1012;
	wire [3-1:0] node1014;
	wire [3-1:0] node1015;
	wire [3-1:0] node1016;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1027;
	wire [3-1:0] node1030;
	wire [3-1:0] node1033;
	wire [3-1:0] node1034;
	wire [3-1:0] node1035;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1043;
	wire [3-1:0] node1046;
	wire [3-1:0] node1047;
	wire [3-1:0] node1048;
	wire [3-1:0] node1050;
	wire [3-1:0] node1054;
	wire [3-1:0] node1055;
	wire [3-1:0] node1057;
	wire [3-1:0] node1060;
	wire [3-1:0] node1062;
	wire [3-1:0] node1065;
	wire [3-1:0] node1066;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1070;
	wire [3-1:0] node1073;
	wire [3-1:0] node1075;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1081;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1089;
	wire [3-1:0] node1090;
	wire [3-1:0] node1092;
	wire [3-1:0] node1096;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1100;
	wire [3-1:0] node1102;
	wire [3-1:0] node1105;
	wire [3-1:0] node1107;
	wire [3-1:0] node1110;
	wire [3-1:0] node1111;
	wire [3-1:0] node1113;
	wire [3-1:0] node1117;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1121;
	wire [3-1:0] node1124;
	wire [3-1:0] node1126;
	wire [3-1:0] node1129;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1135;
	wire [3-1:0] node1137;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1142;
	wire [3-1:0] node1144;
	wire [3-1:0] node1146;

	assign outp = (inp[9]) ? node286 : node1;
		assign node1 = (inp[3]) ? node213 : node2;
			assign node2 = (inp[6]) ? node126 : node3;
				assign node3 = (inp[7]) ? node65 : node4;
					assign node4 = (inp[10]) ? node36 : node5;
						assign node5 = (inp[4]) ? node21 : node6;
							assign node6 = (inp[11]) ? node14 : node7;
								assign node7 = (inp[8]) ? node11 : node8;
									assign node8 = (inp[5]) ? 3'b001 : 3'b101;
									assign node11 = (inp[5]) ? 3'b110 : 3'b001;
								assign node14 = (inp[5]) ? node18 : node15;
									assign node15 = (inp[8]) ? 3'b101 : 3'b011;
									assign node18 = (inp[8]) ? 3'b001 : 3'b101;
							assign node21 = (inp[8]) ? node29 : node22;
								assign node22 = (inp[5]) ? node26 : node23;
									assign node23 = (inp[11]) ? 3'b001 : 3'b110;
									assign node26 = (inp[11]) ? 3'b110 : 3'b010;
								assign node29 = (inp[11]) ? node33 : node30;
									assign node30 = (inp[5]) ? 3'b100 : 3'b010;
									assign node33 = (inp[5]) ? 3'b010 : 3'b110;
						assign node36 = (inp[4]) ? node50 : node37;
							assign node37 = (inp[5]) ? node43 : node38;
								assign node38 = (inp[11]) ? 3'b111 : node39;
									assign node39 = (inp[8]) ? 3'b011 : 3'b111;
								assign node43 = (inp[11]) ? node47 : node44;
									assign node44 = (inp[8]) ? 3'b101 : 3'b011;
									assign node47 = (inp[8]) ? 3'b011 : 3'b111;
							assign node50 = (inp[11]) ? node58 : node51;
								assign node51 = (inp[8]) ? node55 : node52;
									assign node52 = (inp[5]) ? 3'b001 : 3'b101;
									assign node55 = (inp[5]) ? 3'b110 : 3'b001;
								assign node58 = (inp[8]) ? node62 : node59;
									assign node59 = (inp[5]) ? 3'b101 : 3'b011;
									assign node62 = (inp[5]) ? 3'b001 : 3'b101;
					assign node65 = (inp[4]) ? node97 : node66;
						assign node66 = (inp[10]) ? node82 : node67;
							assign node67 = (inp[11]) ? node75 : node68;
								assign node68 = (inp[8]) ? node72 : node69;
									assign node69 = (inp[5]) ? 3'b010 : 3'b110;
									assign node72 = (inp[5]) ? 3'b100 : 3'b010;
								assign node75 = (inp[8]) ? node79 : node76;
									assign node76 = (inp[5]) ? 3'b110 : 3'b001;
									assign node79 = (inp[5]) ? 3'b010 : 3'b110;
							assign node82 = (inp[5]) ? node90 : node83;
								assign node83 = (inp[8]) ? node87 : node84;
									assign node84 = (inp[11]) ? 3'b011 : 3'b101;
									assign node87 = (inp[11]) ? 3'b101 : 3'b001;
								assign node90 = (inp[11]) ? node94 : node91;
									assign node91 = (inp[8]) ? 3'b110 : 3'b001;
									assign node94 = (inp[8]) ? 3'b001 : 3'b101;
						assign node97 = (inp[10]) ? node111 : node98;
							assign node98 = (inp[8]) ? node106 : node99;
								assign node99 = (inp[5]) ? node103 : node100;
									assign node100 = (inp[11]) ? 3'b010 : 3'b100;
									assign node103 = (inp[11]) ? 3'b100 : 3'b000;
								assign node106 = (inp[5]) ? 3'b000 : node107;
									assign node107 = (inp[11]) ? 3'b100 : 3'b000;
							assign node111 = (inp[8]) ? node119 : node112;
								assign node112 = (inp[11]) ? node116 : node113;
									assign node113 = (inp[5]) ? 3'b010 : 3'b110;
									assign node116 = (inp[5]) ? 3'b110 : 3'b001;
								assign node119 = (inp[11]) ? node123 : node120;
									assign node120 = (inp[5]) ? 3'b100 : 3'b010;
									assign node123 = (inp[5]) ? 3'b010 : 3'b110;
				assign node126 = (inp[7]) ? node182 : node127;
					assign node127 = (inp[10]) ? node149 : node128;
						assign node128 = (inp[4]) ? 3'b000 : node129;
							assign node129 = (inp[8]) ? node143 : node130;
								assign node130 = (inp[2]) ? node136 : node131;
									assign node131 = (inp[5]) ? node133 : 3'b100;
										assign node133 = (inp[11]) ? 3'b100 : 3'b000;
									assign node136 = (inp[11]) ? node140 : node137;
										assign node137 = (inp[5]) ? 3'b000 : 3'b100;
										assign node140 = (inp[5]) ? 3'b100 : 3'b010;
								assign node143 = (inp[5]) ? 3'b000 : node144;
									assign node144 = (inp[11]) ? 3'b100 : 3'b000;
						assign node149 = (inp[4]) ? node165 : node150;
							assign node150 = (inp[8]) ? node158 : node151;
								assign node151 = (inp[5]) ? node155 : node152;
									assign node152 = (inp[11]) ? 3'b001 : 3'b110;
									assign node155 = (inp[11]) ? 3'b110 : 3'b010;
								assign node158 = (inp[5]) ? node162 : node159;
									assign node159 = (inp[11]) ? 3'b110 : 3'b010;
									assign node162 = (inp[11]) ? 3'b010 : 3'b100;
							assign node165 = (inp[11]) ? node171 : node166;
								assign node166 = (inp[8]) ? 3'b000 : node167;
									assign node167 = (inp[5]) ? 3'b000 : 3'b100;
								assign node171 = (inp[8]) ? node175 : node172;
									assign node172 = (inp[5]) ? 3'b100 : 3'b010;
									assign node175 = (inp[5]) ? node177 : 3'b100;
										assign node177 = (inp[2]) ? 3'b000 : node178;
											assign node178 = (inp[1]) ? 3'b000 : 3'b000;
					assign node182 = (inp[10]) ? node184 : 3'b000;
						assign node184 = (inp[4]) ? node202 : node185;
							assign node185 = (inp[11]) ? node191 : node186;
								assign node186 = (inp[8]) ? 3'b000 : node187;
									assign node187 = (inp[5]) ? 3'b000 : 3'b100;
								assign node191 = (inp[8]) ? node199 : node192;
									assign node192 = (inp[5]) ? node194 : 3'b010;
										assign node194 = (inp[0]) ? 3'b100 : node195;
											assign node195 = (inp[1]) ? 3'b100 : 3'b010;
									assign node199 = (inp[5]) ? 3'b000 : 3'b100;
							assign node202 = (inp[1]) ? 3'b000 : node203;
								assign node203 = (inp[8]) ? 3'b000 : node204;
									assign node204 = (inp[2]) ? 3'b000 : node205;
										assign node205 = (inp[0]) ? 3'b000 : node206;
											assign node206 = (inp[5]) ? 3'b000 : 3'b100;
			assign node213 = (inp[6]) ? 3'b000 : node214;
				assign node214 = (inp[4]) ? node268 : node215;
					assign node215 = (inp[10]) ? node239 : node216;
						assign node216 = (inp[7]) ? 3'b000 : node217;
							assign node217 = (inp[5]) ? node233 : node218;
								assign node218 = (inp[2]) ? node226 : node219;
									assign node219 = (inp[11]) ? node223 : node220;
										assign node220 = (inp[8]) ? 3'b000 : 3'b100;
										assign node223 = (inp[8]) ? 3'b100 : 3'b010;
									assign node226 = (inp[1]) ? 3'b100 : node227;
										assign node227 = (inp[11]) ? 3'b100 : node228;
											assign node228 = (inp[8]) ? 3'b000 : 3'b100;
								assign node233 = (inp[11]) ? node235 : 3'b000;
									assign node235 = (inp[8]) ? 3'b000 : 3'b100;
						assign node239 = (inp[7]) ? node255 : node240;
							assign node240 = (inp[8]) ? node248 : node241;
								assign node241 = (inp[5]) ? node245 : node242;
									assign node242 = (inp[11]) ? 3'b001 : 3'b110;
									assign node245 = (inp[11]) ? 3'b110 : 3'b010;
								assign node248 = (inp[5]) ? node252 : node249;
									assign node249 = (inp[11]) ? 3'b110 : 3'b010;
									assign node252 = (inp[11]) ? 3'b010 : 3'b100;
							assign node255 = (inp[5]) ? node263 : node256;
								assign node256 = (inp[8]) ? node260 : node257;
									assign node257 = (inp[11]) ? 3'b010 : 3'b100;
									assign node260 = (inp[11]) ? 3'b100 : 3'b000;
								assign node263 = (inp[11]) ? node265 : 3'b000;
									assign node265 = (inp[8]) ? 3'b000 : 3'b100;
					assign node268 = (inp[10]) ? node270 : 3'b000;
						assign node270 = (inp[7]) ? 3'b000 : node271;
							assign node271 = (inp[8]) ? node279 : node272;
								assign node272 = (inp[11]) ? node276 : node273;
									assign node273 = (inp[5]) ? 3'b000 : 3'b100;
									assign node276 = (inp[5]) ? 3'b100 : 3'b010;
								assign node279 = (inp[11]) ? node281 : 3'b000;
									assign node281 = (inp[5]) ? 3'b000 : 3'b100;
		assign node286 = (inp[3]) ? node672 : node287;
			assign node287 = (inp[6]) ? node379 : node288;
				assign node288 = (inp[10]) ? node348 : node289;
					assign node289 = (inp[4]) ? node305 : node290;
						assign node290 = (inp[7]) ? node292 : 3'b111;
							assign node292 = (inp[5]) ? node298 : node293;
								assign node293 = (inp[11]) ? 3'b111 : node294;
									assign node294 = (inp[8]) ? 3'b011 : 3'b111;
								assign node298 = (inp[8]) ? node302 : node299;
									assign node299 = (inp[11]) ? 3'b111 : 3'b011;
									assign node302 = (inp[11]) ? 3'b011 : 3'b101;
						assign node305 = (inp[7]) ? node319 : node306;
							assign node306 = (inp[11]) ? node314 : node307;
								assign node307 = (inp[5]) ? node311 : node308;
									assign node308 = (inp[8]) ? 3'b011 : 3'b111;
									assign node311 = (inp[8]) ? 3'b101 : 3'b011;
								assign node314 = (inp[8]) ? node316 : 3'b111;
									assign node316 = (inp[5]) ? 3'b011 : 3'b111;
							assign node319 = (inp[5]) ? node333 : node320;
								assign node320 = (inp[11]) ? node324 : node321;
									assign node321 = (inp[8]) ? 3'b001 : 3'b101;
									assign node324 = (inp[8]) ? node328 : node325;
										assign node325 = (inp[0]) ? 3'b011 : 3'b111;
										assign node328 = (inp[1]) ? 3'b101 : node329;
											assign node329 = (inp[0]) ? 3'b101 : 3'b011;
								assign node333 = (inp[11]) ? node341 : node334;
									assign node334 = (inp[8]) ? node336 : 3'b001;
										assign node336 = (inp[2]) ? 3'b110 : node337;
											assign node337 = (inp[0]) ? 3'b110 : 3'b000;
									assign node341 = (inp[8]) ? node343 : 3'b101;
										assign node343 = (inp[1]) ? 3'b001 : node344;
											assign node344 = (inp[0]) ? 3'b001 : 3'b101;
					assign node348 = (inp[7]) ? node350 : 3'b111;
						assign node350 = (inp[4]) ? node352 : 3'b111;
							assign node352 = (inp[8]) ? node362 : node353;
								assign node353 = (inp[11]) ? 3'b111 : node354;
									assign node354 = (inp[5]) ? node356 : 3'b111;
										assign node356 = (inp[0]) ? 3'b011 : node357;
											assign node357 = (inp[1]) ? 3'b011 : 3'b111;
								assign node362 = (inp[5]) ? node370 : node363;
									assign node363 = (inp[11]) ? 3'b111 : node364;
										assign node364 = (inp[1]) ? 3'b011 : node365;
											assign node365 = (inp[0]) ? 3'b011 : 3'b111;
									assign node370 = (inp[11]) ? node376 : node371;
										assign node371 = (inp[0]) ? 3'b101 : node372;
											assign node372 = (inp[1]) ? 3'b101 : 3'b011;
										assign node376 = (inp[0]) ? 3'b011 : 3'b111;
				assign node379 = (inp[10]) ? node527 : node380;
					assign node380 = (inp[7]) ? node454 : node381;
						assign node381 = (inp[4]) ? node421 : node382;
							assign node382 = (inp[11]) ? node398 : node383;
								assign node383 = (inp[5]) ? node391 : node384;
									assign node384 = (inp[8]) ? node386 : 3'b101;
										assign node386 = (inp[0]) ? 3'b001 : node387;
											assign node387 = (inp[2]) ? 3'b001 : 3'b101;
									assign node391 = (inp[8]) ? 3'b110 : node392;
										assign node392 = (inp[0]) ? 3'b001 : node393;
											assign node393 = (inp[2]) ? 3'b001 : 3'b001;
								assign node398 = (inp[5]) ? node410 : node399;
									assign node399 = (inp[8]) ? node405 : node400;
										assign node400 = (inp[1]) ? 3'b011 : node401;
											assign node401 = (inp[0]) ? 3'b011 : 3'b111;
										assign node405 = (inp[0]) ? 3'b101 : node406;
											assign node406 = (inp[1]) ? 3'b101 : 3'b011;
									assign node410 = (inp[8]) ? node416 : node411;
										assign node411 = (inp[0]) ? 3'b101 : node412;
											assign node412 = (inp[1]) ? 3'b101 : 3'b011;
										assign node416 = (inp[0]) ? 3'b001 : node417;
											assign node417 = (inp[2]) ? 3'b001 : 3'b101;
							assign node421 = (inp[11]) ? node435 : node422;
								assign node422 = (inp[8]) ? node430 : node423;
									assign node423 = (inp[5]) ? 3'b010 : node424;
										assign node424 = (inp[2]) ? 3'b110 : node425;
											assign node425 = (inp[1]) ? 3'b110 : 3'b001;
									assign node430 = (inp[5]) ? node432 : 3'b010;
										assign node432 = (inp[1]) ? 3'b100 : 3'b010;
								assign node435 = (inp[5]) ? node445 : node436;
									assign node436 = (inp[2]) ? node438 : 3'b001;
										assign node438 = (inp[8]) ? node442 : node439;
											assign node439 = (inp[1]) ? 3'b001 : 3'b101;
											assign node442 = (inp[1]) ? 3'b110 : 3'b000;
									assign node445 = (inp[0]) ? node451 : node446;
										assign node446 = (inp[2]) ? node448 : 3'b001;
											assign node448 = (inp[1]) ? 3'b010 : 3'b000;
										assign node451 = (inp[8]) ? 3'b010 : 3'b110;
						assign node454 = (inp[4]) ? node498 : node455;
							assign node455 = (inp[11]) ? node477 : node456;
								assign node456 = (inp[8]) ? node468 : node457;
									assign node457 = (inp[5]) ? node463 : node458;
										assign node458 = (inp[0]) ? 3'b110 : node459;
											assign node459 = (inp[1]) ? 3'b110 : 3'b001;
										assign node463 = (inp[0]) ? 3'b010 : node464;
											assign node464 = (inp[1]) ? 3'b010 : 3'b110;
									assign node468 = (inp[5]) ? node474 : node469;
										assign node469 = (inp[1]) ? 3'b010 : node470;
											assign node470 = (inp[0]) ? 3'b010 : 3'b110;
										assign node474 = (inp[0]) ? 3'b100 : 3'b010;
								assign node477 = (inp[5]) ? node487 : node478;
									assign node478 = (inp[0]) ? node484 : node479;
										assign node479 = (inp[8]) ? 3'b001 : node480;
											assign node480 = (inp[1]) ? 3'b001 : 3'b101;
										assign node484 = (inp[8]) ? 3'b110 : 3'b001;
									assign node487 = (inp[1]) ? node493 : node488;
										assign node488 = (inp[8]) ? 3'b110 : node489;
											assign node489 = (inp[0]) ? 3'b110 : 3'b001;
										assign node493 = (inp[0]) ? node495 : 3'b110;
											assign node495 = (inp[8]) ? 3'b010 : 3'b110;
							assign node498 = (inp[11]) ? node512 : node499;
								assign node499 = (inp[0]) ? node507 : node500;
									assign node500 = (inp[2]) ? node502 : 3'b100;
										assign node502 = (inp[1]) ? 3'b000 : node503;
											assign node503 = (inp[5]) ? 3'b100 : 3'b000;
									assign node507 = (inp[8]) ? 3'b000 : node508;
										assign node508 = (inp[5]) ? 3'b000 : 3'b100;
								assign node512 = (inp[8]) ? node520 : node513;
									assign node513 = (inp[0]) ? node517 : node514;
										assign node514 = (inp[5]) ? 3'b010 : 3'b110;
										assign node517 = (inp[5]) ? 3'b100 : 3'b010;
									assign node520 = (inp[0]) ? node524 : node521;
										assign node521 = (inp[5]) ? 3'b100 : 3'b010;
										assign node524 = (inp[5]) ? 3'b000 : 3'b100;
					assign node527 = (inp[4]) ? node595 : node528;
						assign node528 = (inp[7]) ? node550 : node529;
							assign node529 = (inp[5]) ? node537 : node530;
								assign node530 = (inp[8]) ? node532 : 3'b111;
									assign node532 = (inp[11]) ? 3'b111 : node533;
										assign node533 = (inp[0]) ? 3'b011 : 3'b111;
								assign node537 = (inp[11]) ? node545 : node538;
									assign node538 = (inp[0]) ? node542 : node539;
										assign node539 = (inp[8]) ? 3'b011 : 3'b111;
										assign node542 = (inp[8]) ? 3'b101 : 3'b011;
									assign node545 = (inp[8]) ? node547 : 3'b111;
										assign node547 = (inp[0]) ? 3'b011 : 3'b111;
							assign node550 = (inp[11]) ? node572 : node551;
								assign node551 = (inp[5]) ? node565 : node552;
									assign node552 = (inp[1]) ? node558 : node553;
										assign node553 = (inp[2]) ? node555 : 3'b101;
											assign node555 = (inp[0]) ? 3'b001 : 3'b101;
										assign node558 = (inp[8]) ? node562 : node559;
											assign node559 = (inp[0]) ? 3'b101 : 3'b011;
											assign node562 = (inp[0]) ? 3'b001 : 3'b101;
									assign node565 = (inp[8]) ? node569 : node566;
										assign node566 = (inp[0]) ? 3'b001 : 3'b101;
										assign node569 = (inp[0]) ? 3'b110 : 3'b001;
								assign node572 = (inp[8]) ? node584 : node573;
									assign node573 = (inp[5]) ? node579 : node574;
										assign node574 = (inp[0]) ? node576 : 3'b111;
											assign node576 = (inp[1]) ? 3'b011 : 3'b011;
										assign node579 = (inp[2]) ? node581 : 3'b011;
											assign node581 = (inp[0]) ? 3'b001 : 3'b011;
									assign node584 = (inp[5]) ? node590 : node585;
										assign node585 = (inp[1]) ? node587 : 3'b011;
											assign node587 = (inp[0]) ? 3'b101 : 3'b011;
										assign node590 = (inp[0]) ? node592 : 3'b101;
											assign node592 = (inp[1]) ? 3'b001 : 3'b101;
						assign node595 = (inp[7]) ? node633 : node596;
							assign node596 = (inp[11]) ? node614 : node597;
								assign node597 = (inp[8]) ? node607 : node598;
									assign node598 = (inp[5]) ? node604 : node599;
										assign node599 = (inp[0]) ? 3'b101 : node600;
											assign node600 = (inp[1]) ? 3'b101 : 3'b011;
										assign node604 = (inp[0]) ? 3'b001 : 3'b101;
									assign node607 = (inp[5]) ? node611 : node608;
										assign node608 = (inp[0]) ? 3'b001 : 3'b101;
										assign node611 = (inp[0]) ? 3'b110 : 3'b001;
								assign node614 = (inp[0]) ? node622 : node615;
									assign node615 = (inp[8]) ? node619 : node616;
										assign node616 = (inp[5]) ? 3'b011 : 3'b111;
										assign node619 = (inp[5]) ? 3'b101 : 3'b011;
									assign node622 = (inp[5]) ? node628 : node623;
										assign node623 = (inp[8]) ? 3'b101 : node624;
											assign node624 = (inp[2]) ? 3'b011 : 3'b111;
										assign node628 = (inp[1]) ? node630 : 3'b101;
											assign node630 = (inp[8]) ? 3'b001 : 3'b101;
							assign node633 = (inp[11]) ? node657 : node634;
								assign node634 = (inp[1]) ? node646 : node635;
									assign node635 = (inp[8]) ? node641 : node636;
										assign node636 = (inp[5]) ? 3'b110 : node637;
											assign node637 = (inp[0]) ? 3'b110 : 3'b001;
										assign node641 = (inp[5]) ? 3'b010 : node642;
											assign node642 = (inp[0]) ? 3'b010 : 3'b110;
									assign node646 = (inp[8]) ? node652 : node647;
										assign node647 = (inp[5]) ? node649 : 3'b001;
											assign node649 = (inp[0]) ? 3'b010 : 3'b110;
										assign node652 = (inp[5]) ? 3'b100 : node653;
											assign node653 = (inp[2]) ? 3'b110 : 3'b010;
								assign node657 = (inp[8]) ? node665 : node658;
									assign node658 = (inp[2]) ? 3'b001 : node659;
										assign node659 = (inp[0]) ? node661 : 3'b001;
											assign node661 = (inp[1]) ? 3'b110 : 3'b101;
									assign node665 = (inp[5]) ? 3'b110 : node666;
										assign node666 = (inp[1]) ? node668 : 3'b001;
											assign node668 = (inp[0]) ? 3'b110 : 3'b001;
			assign node672 = (inp[6]) ? node954 : node673;
				assign node673 = (inp[10]) ? node793 : node674;
					assign node674 = (inp[4]) ? node728 : node675;
						assign node675 = (inp[7]) ? node695 : node676;
							assign node676 = (inp[8]) ? node688 : node677;
								assign node677 = (inp[11]) ? node681 : node678;
									assign node678 = (inp[5]) ? 3'b001 : 3'b101;
									assign node681 = (inp[5]) ? node683 : 3'b011;
										assign node683 = (inp[2]) ? 3'b101 : node684;
											assign node684 = (inp[0]) ? 3'b101 : 3'b001;
								assign node688 = (inp[11]) ? node692 : node689;
									assign node689 = (inp[5]) ? 3'b110 : 3'b001;
									assign node692 = (inp[5]) ? 3'b001 : 3'b101;
							assign node695 = (inp[11]) ? node711 : node696;
								assign node696 = (inp[8]) ? node704 : node697;
									assign node697 = (inp[5]) ? node699 : 3'b110;
										assign node699 = (inp[2]) ? 3'b010 : node700;
											assign node700 = (inp[1]) ? 3'b010 : 3'b110;
									assign node704 = (inp[5]) ? node706 : 3'b010;
										assign node706 = (inp[1]) ? 3'b100 : node707;
											assign node707 = (inp[0]) ? 3'b100 : 3'b010;
								assign node711 = (inp[8]) ? node721 : node712;
									assign node712 = (inp[5]) ? node718 : node713;
										assign node713 = (inp[0]) ? 3'b001 : node714;
											assign node714 = (inp[1]) ? 3'b001 : 3'b101;
										assign node718 = (inp[2]) ? 3'b110 : 3'b001;
									assign node721 = (inp[5]) ? node723 : 3'b110;
										assign node723 = (inp[0]) ? 3'b010 : node724;
											assign node724 = (inp[1]) ? 3'b010 : 3'b110;
						assign node728 = (inp[7]) ? node758 : node729;
							assign node729 = (inp[11]) ? node737 : node730;
								assign node730 = (inp[8]) ? node734 : node731;
									assign node731 = (inp[5]) ? 3'b010 : 3'b110;
									assign node734 = (inp[5]) ? 3'b100 : 3'b010;
								assign node737 = (inp[5]) ? node747 : node738;
									assign node738 = (inp[8]) ? node744 : node739;
										assign node739 = (inp[0]) ? 3'b001 : node740;
											assign node740 = (inp[1]) ? 3'b001 : 3'b001;
										assign node744 = (inp[0]) ? 3'b110 : 3'b001;
									assign node747 = (inp[8]) ? node753 : node748;
										assign node748 = (inp[1]) ? 3'b110 : node749;
											assign node749 = (inp[2]) ? 3'b110 : 3'b001;
										assign node753 = (inp[0]) ? 3'b010 : node754;
											assign node754 = (inp[1]) ? 3'b010 : 3'b110;
							assign node758 = (inp[11]) ? node774 : node759;
								assign node759 = (inp[8]) ? node767 : node760;
									assign node760 = (inp[5]) ? node762 : 3'b100;
										assign node762 = (inp[0]) ? 3'b000 : node763;
											assign node763 = (inp[1]) ? 3'b000 : 3'b100;
									assign node767 = (inp[1]) ? 3'b000 : node768;
										assign node768 = (inp[5]) ? 3'b000 : node769;
											assign node769 = (inp[2]) ? 3'b000 : 3'b100;
								assign node774 = (inp[8]) ? node788 : node775;
									assign node775 = (inp[1]) ? node783 : node776;
										assign node776 = (inp[2]) ? node780 : node777;
											assign node777 = (inp[0]) ? 3'b010 : 3'b010;
											assign node780 = (inp[0]) ? 3'b100 : 3'b010;
										assign node783 = (inp[2]) ? 3'b100 : node784;
											assign node784 = (inp[0]) ? 3'b100 : 3'b010;
									assign node788 = (inp[5]) ? node790 : 3'b100;
										assign node790 = (inp[0]) ? 3'b000 : 3'b100;
					assign node793 = (inp[4]) ? node863 : node794;
						assign node794 = (inp[7]) ? node820 : node795;
							assign node795 = (inp[5]) ? node805 : node796;
								assign node796 = (inp[8]) ? node798 : 3'b111;
									assign node798 = (inp[11]) ? 3'b111 : node799;
										assign node799 = (inp[1]) ? 3'b011 : node800;
											assign node800 = (inp[0]) ? 3'b011 : 3'b111;
								assign node805 = (inp[11]) ? node815 : node806;
									assign node806 = (inp[8]) ? node812 : node807;
										assign node807 = (inp[0]) ? 3'b011 : node808;
											assign node808 = (inp[1]) ? 3'b011 : 3'b111;
										assign node812 = (inp[0]) ? 3'b101 : 3'b011;
									assign node815 = (inp[0]) ? node817 : 3'b111;
										assign node817 = (inp[8]) ? 3'b011 : 3'b111;
							assign node820 = (inp[11]) ? node840 : node821;
								assign node821 = (inp[5]) ? node833 : node822;
									assign node822 = (inp[8]) ? node828 : node823;
										assign node823 = (inp[0]) ? 3'b101 : node824;
											assign node824 = (inp[2]) ? 3'b001 : 3'b011;
										assign node828 = (inp[0]) ? 3'b001 : node829;
											assign node829 = (inp[2]) ? 3'b001 : 3'b101;
									assign node833 = (inp[8]) ? node837 : node834;
										assign node834 = (inp[0]) ? 3'b001 : 3'b101;
										assign node837 = (inp[0]) ? 3'b110 : 3'b001;
								assign node840 = (inp[5]) ? node854 : node841;
									assign node841 = (inp[1]) ? node847 : node842;
										assign node842 = (inp[0]) ? 3'b011 : node843;
											assign node843 = (inp[8]) ? 3'b011 : 3'b111;
										assign node847 = (inp[0]) ? node851 : node848;
											assign node848 = (inp[8]) ? 3'b011 : 3'b111;
											assign node851 = (inp[8]) ? 3'b101 : 3'b011;
									assign node854 = (inp[0]) ? node858 : node855;
										assign node855 = (inp[8]) ? 3'b101 : 3'b011;
										assign node858 = (inp[8]) ? node860 : 3'b101;
											assign node860 = (inp[2]) ? 3'b001 : 3'b001;
						assign node863 = (inp[7]) ? node911 : node864;
							assign node864 = (inp[0]) ? node884 : node865;
								assign node865 = (inp[5]) ? node873 : node866;
									assign node866 = (inp[11]) ? node870 : node867;
										assign node867 = (inp[2]) ? 3'b101 : 3'b011;
										assign node870 = (inp[8]) ? 3'b011 : 3'b111;
									assign node873 = (inp[11]) ? node881 : node874;
										assign node874 = (inp[8]) ? node878 : node875;
											assign node875 = (inp[2]) ? 3'b001 : 3'b101;
											assign node878 = (inp[2]) ? 3'b000 : 3'b001;
										assign node881 = (inp[8]) ? 3'b101 : 3'b011;
								assign node884 = (inp[2]) ? node896 : node885;
									assign node885 = (inp[5]) ? node891 : node886;
										assign node886 = (inp[8]) ? node888 : 3'b101;
											assign node888 = (inp[11]) ? 3'b101 : 3'b001;
										assign node891 = (inp[8]) ? 3'b001 : node892;
											assign node892 = (inp[11]) ? 3'b101 : 3'b001;
									assign node896 = (inp[5]) ? node904 : node897;
										assign node897 = (inp[11]) ? node901 : node898;
											assign node898 = (inp[8]) ? 3'b001 : 3'b101;
											assign node901 = (inp[8]) ? 3'b101 : 3'b011;
										assign node904 = (inp[8]) ? node908 : node905;
											assign node905 = (inp[11]) ? 3'b101 : 3'b001;
											assign node908 = (inp[11]) ? 3'b001 : 3'b110;
							assign node911 = (inp[11]) ? node929 : node912;
								assign node912 = (inp[0]) ? node922 : node913;
									assign node913 = (inp[5]) ? node919 : node914;
										assign node914 = (inp[8]) ? 3'b110 : node915;
											assign node915 = (inp[1]) ? 3'b000 : 3'b001;
										assign node919 = (inp[8]) ? 3'b010 : 3'b110;
									assign node922 = (inp[5]) ? node926 : node923;
										assign node923 = (inp[8]) ? 3'b010 : 3'b110;
										assign node926 = (inp[8]) ? 3'b100 : 3'b010;
								assign node929 = (inp[0]) ? node941 : node930;
									assign node930 = (inp[2]) ? node936 : node931;
										assign node931 = (inp[8]) ? 3'b001 : node932;
											assign node932 = (inp[5]) ? 3'b001 : 3'b101;
										assign node936 = (inp[8]) ? 3'b110 : node937;
											assign node937 = (inp[5]) ? 3'b001 : 3'b101;
									assign node941 = (inp[8]) ? node947 : node942;
										assign node942 = (inp[5]) ? node944 : 3'b001;
											assign node944 = (inp[1]) ? 3'b110 : 3'b001;
										assign node947 = (inp[1]) ? node951 : node948;
											assign node948 = (inp[5]) ? 3'b110 : 3'b001;
											assign node951 = (inp[5]) ? 3'b010 : 3'b110;
				assign node954 = (inp[10]) ? node1022 : node955;
					assign node955 = (inp[7]) ? node1009 : node956;
						assign node956 = (inp[4]) ? node998 : node957;
							assign node957 = (inp[11]) ? node977 : node958;
								assign node958 = (inp[5]) ? node970 : node959;
									assign node959 = (inp[8]) ? node965 : node960;
										assign node960 = (inp[0]) ? 3'b100 : node961;
											assign node961 = (inp[1]) ? 3'b100 : 3'b010;
										assign node965 = (inp[1]) ? 3'b000 : node966;
											assign node966 = (inp[0]) ? 3'b000 : 3'b100;
									assign node970 = (inp[0]) ? 3'b000 : node971;
										assign node971 = (inp[1]) ? 3'b000 : node972;
											assign node972 = (inp[8]) ? 3'b000 : 3'b100;
								assign node977 = (inp[8]) ? node989 : node978;
									assign node978 = (inp[5]) ? node984 : node979;
										assign node979 = (inp[0]) ? 3'b010 : node980;
											assign node980 = (inp[1]) ? 3'b010 : 3'b110;
										assign node984 = (inp[1]) ? node986 : 3'b010;
											assign node986 = (inp[0]) ? 3'b100 : 3'b000;
									assign node989 = (inp[0]) ? node995 : node990;
										assign node990 = (inp[2]) ? node992 : 3'b010;
											assign node992 = (inp[5]) ? 3'b100 : 3'b000;
										assign node995 = (inp[5]) ? 3'b000 : 3'b100;
							assign node998 = (inp[11]) ? node1000 : 3'b000;
								assign node1000 = (inp[1]) ? node1002 : 3'b000;
									assign node1002 = (inp[0]) ? 3'b000 : node1003;
										assign node1003 = (inp[5]) ? 3'b000 : node1004;
											assign node1004 = (inp[8]) ? 3'b000 : 3'b100;
						assign node1009 = (inp[11]) ? node1011 : 3'b000;
							assign node1011 = (inp[5]) ? 3'b000 : node1012;
								assign node1012 = (inp[2]) ? node1014 : 3'b000;
									assign node1014 = (inp[4]) ? 3'b000 : node1015;
										assign node1015 = (inp[8]) ? 3'b000 : node1016;
											assign node1016 = (inp[1]) ? 3'b000 : 3'b100;
					assign node1022 = (inp[4]) ? node1096 : node1023;
						assign node1023 = (inp[7]) ? node1065 : node1024;
							assign node1024 = (inp[8]) ? node1046 : node1025;
								assign node1025 = (inp[11]) ? node1033 : node1026;
									assign node1026 = (inp[5]) ? node1030 : node1027;
										assign node1027 = (inp[0]) ? 3'b110 : 3'b001;
										assign node1030 = (inp[0]) ? 3'b010 : 3'b110;
									assign node1033 = (inp[1]) ? node1039 : node1034;
										assign node1034 = (inp[5]) ? 3'b001 : node1035;
											assign node1035 = (inp[0]) ? 3'b001 : 3'b101;
										assign node1039 = (inp[5]) ? node1043 : node1040;
											assign node1040 = (inp[0]) ? 3'b001 : 3'b101;
											assign node1043 = (inp[0]) ? 3'b110 : 3'b001;
								assign node1046 = (inp[11]) ? node1054 : node1047;
									assign node1047 = (inp[5]) ? 3'b010 : node1048;
										assign node1048 = (inp[0]) ? node1050 : 3'b110;
											assign node1050 = (inp[1]) ? 3'b010 : 3'b010;
									assign node1054 = (inp[5]) ? node1060 : node1055;
										assign node1055 = (inp[0]) ? node1057 : 3'b001;
											assign node1057 = (inp[1]) ? 3'b110 : 3'b001;
										assign node1060 = (inp[0]) ? node1062 : 3'b110;
											assign node1062 = (inp[1]) ? 3'b010 : 3'b110;
							assign node1065 = (inp[11]) ? node1085 : node1066;
								assign node1066 = (inp[5]) ? node1078 : node1067;
									assign node1067 = (inp[8]) ? node1073 : node1068;
										assign node1068 = (inp[0]) ? node1070 : 3'b010;
											assign node1070 = (inp[1]) ? 3'b100 : 3'b010;
										assign node1073 = (inp[0]) ? node1075 : 3'b100;
											assign node1075 = (inp[1]) ? 3'b000 : 3'b100;
									assign node1078 = (inp[8]) ? 3'b000 : node1079;
										assign node1079 = (inp[1]) ? node1081 : 3'b100;
											assign node1081 = (inp[0]) ? 3'b000 : 3'b100;
								assign node1085 = (inp[8]) ? node1089 : node1086;
									assign node1086 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1089 = (inp[5]) ? 3'b100 : node1090;
										assign node1090 = (inp[2]) ? node1092 : 3'b010;
											assign node1092 = (inp[1]) ? 3'b100 : 3'b010;
						assign node1096 = (inp[7]) ? node1140 : node1097;
							assign node1097 = (inp[11]) ? node1117 : node1098;
								assign node1098 = (inp[5]) ? node1110 : node1099;
									assign node1099 = (inp[8]) ? node1105 : node1100;
										assign node1100 = (inp[1]) ? node1102 : 3'b010;
											assign node1102 = (inp[0]) ? 3'b100 : 3'b010;
										assign node1105 = (inp[0]) ? node1107 : 3'b100;
											assign node1107 = (inp[2]) ? 3'b000 : 3'b000;
									assign node1110 = (inp[8]) ? 3'b000 : node1111;
										assign node1111 = (inp[0]) ? node1113 : 3'b100;
											assign node1113 = (inp[2]) ? 3'b000 : 3'b000;
								assign node1117 = (inp[5]) ? node1129 : node1118;
									assign node1118 = (inp[8]) ? node1124 : node1119;
										assign node1119 = (inp[2]) ? node1121 : 3'b110;
											assign node1121 = (inp[0]) ? 3'b010 : 3'b110;
										assign node1124 = (inp[1]) ? node1126 : 3'b010;
											assign node1126 = (inp[0]) ? 3'b100 : 3'b010;
									assign node1129 = (inp[8]) ? node1135 : node1130;
										assign node1130 = (inp[2]) ? 3'b010 : node1131;
											assign node1131 = (inp[1]) ? 3'b000 : 3'b010;
										assign node1135 = (inp[2]) ? node1137 : 3'b100;
											assign node1137 = (inp[1]) ? 3'b000 : 3'b100;
							assign node1140 = (inp[8]) ? 3'b000 : node1141;
								assign node1141 = (inp[5]) ? 3'b000 : node1142;
									assign node1142 = (inp[11]) ? node1144 : 3'b000;
										assign node1144 = (inp[0]) ? node1146 : 3'b100;
											assign node1146 = (inp[1]) ? 3'b000 : 3'b100;

endmodule