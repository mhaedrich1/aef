module dtc_split25_bm61 (
	input  wire [12-1:0] inp,
	output wire [11-1:0] outp
);

	wire [11-1:0] node1;
	wire [11-1:0] node2;
	wire [11-1:0] node3;
	wire [11-1:0] node4;
	wire [11-1:0] node5;
	wire [11-1:0] node6;
	wire [11-1:0] node7;
	wire [11-1:0] node8;
	wire [11-1:0] node10;
	wire [11-1:0] node13;
	wire [11-1:0] node14;
	wire [11-1:0] node18;
	wire [11-1:0] node19;
	wire [11-1:0] node20;
	wire [11-1:0] node21;
	wire [11-1:0] node22;
	wire [11-1:0] node28;
	wire [11-1:0] node29;
	wire [11-1:0] node30;
	wire [11-1:0] node31;
	wire [11-1:0] node36;
	wire [11-1:0] node39;
	wire [11-1:0] node40;
	wire [11-1:0] node41;
	wire [11-1:0] node42;
	wire [11-1:0] node43;
	wire [11-1:0] node47;
	wire [11-1:0] node50;
	wire [11-1:0] node51;
	wire [11-1:0] node55;
	wire [11-1:0] node56;
	wire [11-1:0] node57;
	wire [11-1:0] node59;
	wire [11-1:0] node62;
	wire [11-1:0] node65;
	wire [11-1:0] node67;
	wire [11-1:0] node70;
	wire [11-1:0] node71;
	wire [11-1:0] node72;
	wire [11-1:0] node73;
	wire [11-1:0] node74;
	wire [11-1:0] node79;
	wire [11-1:0] node80;
	wire [11-1:0] node82;
	wire [11-1:0] node83;
	wire [11-1:0] node87;
	wire [11-1:0] node88;
	wire [11-1:0] node91;
	wire [11-1:0] node92;
	wire [11-1:0] node93;
	wire [11-1:0] node98;
	wire [11-1:0] node99;
	wire [11-1:0] node101;
	wire [11-1:0] node102;
	wire [11-1:0] node105;
	wire [11-1:0] node106;
	wire [11-1:0] node109;
	wire [11-1:0] node112;
	wire [11-1:0] node113;
	wire [11-1:0] node114;
	wire [11-1:0] node117;
	wire [11-1:0] node118;
	wire [11-1:0] node121;
	wire [11-1:0] node123;
	wire [11-1:0] node126;
	wire [11-1:0] node127;
	wire [11-1:0] node128;
	wire [11-1:0] node133;
	wire [11-1:0] node134;
	wire [11-1:0] node135;
	wire [11-1:0] node136;
	wire [11-1:0] node137;
	wire [11-1:0] node139;
	wire [11-1:0] node142;
	wire [11-1:0] node143;
	wire [11-1:0] node146;
	wire [11-1:0] node149;
	wire [11-1:0] node150;
	wire [11-1:0] node153;
	wire [11-1:0] node154;
	wire [11-1:0] node157;
	wire [11-1:0] node160;
	wire [11-1:0] node161;
	wire [11-1:0] node162;
	wire [11-1:0] node163;
	wire [11-1:0] node164;
	wire [11-1:0] node168;
	wire [11-1:0] node171;
	wire [11-1:0] node172;
	wire [11-1:0] node174;
	wire [11-1:0] node177;
	wire [11-1:0] node178;
	wire [11-1:0] node181;
	wire [11-1:0] node184;
	wire [11-1:0] node185;
	wire [11-1:0] node186;
	wire [11-1:0] node188;
	wire [11-1:0] node192;
	wire [11-1:0] node193;
	wire [11-1:0] node194;
	wire [11-1:0] node198;
	wire [11-1:0] node199;
	wire [11-1:0] node202;
	wire [11-1:0] node203;
	wire [11-1:0] node207;
	wire [11-1:0] node208;
	wire [11-1:0] node209;
	wire [11-1:0] node210;
	wire [11-1:0] node213;
	wire [11-1:0] node216;
	wire [11-1:0] node217;
	wire [11-1:0] node218;
	wire [11-1:0] node221;
	wire [11-1:0] node224;
	wire [11-1:0] node225;
	wire [11-1:0] node226;
	wire [11-1:0] node230;
	wire [11-1:0] node233;
	wire [11-1:0] node234;
	wire [11-1:0] node235;
	wire [11-1:0] node236;
	wire [11-1:0] node237;
	wire [11-1:0] node239;
	wire [11-1:0] node243;
	wire [11-1:0] node245;
	wire [11-1:0] node248;
	wire [11-1:0] node249;
	wire [11-1:0] node251;
	wire [11-1:0] node254;
	wire [11-1:0] node255;
	wire [11-1:0] node258;
	wire [11-1:0] node261;
	wire [11-1:0] node262;
	wire [11-1:0] node263;
	wire [11-1:0] node266;
	wire [11-1:0] node268;
	wire [11-1:0] node269;
	wire [11-1:0] node273;
	wire [11-1:0] node274;
	wire [11-1:0] node276;
	wire [11-1:0] node280;
	wire [11-1:0] node281;
	wire [11-1:0] node282;
	wire [11-1:0] node283;
	wire [11-1:0] node284;
	wire [11-1:0] node285;
	wire [11-1:0] node286;
	wire [11-1:0] node289;
	wire [11-1:0] node292;
	wire [11-1:0] node294;
	wire [11-1:0] node297;
	wire [11-1:0] node298;
	wire [11-1:0] node300;
	wire [11-1:0] node301;
	wire [11-1:0] node305;
	wire [11-1:0] node306;
	wire [11-1:0] node308;
	wire [11-1:0] node309;
	wire [11-1:0] node312;
	wire [11-1:0] node315;
	wire [11-1:0] node317;
	wire [11-1:0] node320;
	wire [11-1:0] node321;
	wire [11-1:0] node322;
	wire [11-1:0] node323;
	wire [11-1:0] node326;
	wire [11-1:0] node329;
	wire [11-1:0] node331;
	wire [11-1:0] node332;
	wire [11-1:0] node336;
	wire [11-1:0] node338;
	wire [11-1:0] node341;
	wire [11-1:0] node342;
	wire [11-1:0] node343;
	wire [11-1:0] node345;
	wire [11-1:0] node347;
	wire [11-1:0] node348;
	wire [11-1:0] node350;
	wire [11-1:0] node353;
	wire [11-1:0] node355;
	wire [11-1:0] node358;
	wire [11-1:0] node360;
	wire [11-1:0] node362;
	wire [11-1:0] node365;
	wire [11-1:0] node366;
	wire [11-1:0] node367;
	wire [11-1:0] node369;
	wire [11-1:0] node370;
	wire [11-1:0] node373;
	wire [11-1:0] node376;
	wire [11-1:0] node378;
	wire [11-1:0] node381;
	wire [11-1:0] node382;
	wire [11-1:0] node384;
	wire [11-1:0] node387;
	wire [11-1:0] node388;
	wire [11-1:0] node390;
	wire [11-1:0] node392;
	wire [11-1:0] node395;
	wire [11-1:0] node397;
	wire [11-1:0] node400;
	wire [11-1:0] node401;
	wire [11-1:0] node402;
	wire [11-1:0] node403;
	wire [11-1:0] node404;
	wire [11-1:0] node405;
	wire [11-1:0] node407;
	wire [11-1:0] node410;
	wire [11-1:0] node412;
	wire [11-1:0] node415;
	wire [11-1:0] node416;
	wire [11-1:0] node419;
	wire [11-1:0] node422;
	wire [11-1:0] node423;
	wire [11-1:0] node425;
	wire [11-1:0] node428;
	wire [11-1:0] node429;
	wire [11-1:0] node432;
	wire [11-1:0] node435;
	wire [11-1:0] node436;
	wire [11-1:0] node437;
	wire [11-1:0] node438;
	wire [11-1:0] node439;
	wire [11-1:0] node443;
	wire [11-1:0] node444;
	wire [11-1:0] node447;
	wire [11-1:0] node450;
	wire [11-1:0] node451;
	wire [11-1:0] node453;
	wire [11-1:0] node456;
	wire [11-1:0] node459;
	wire [11-1:0] node460;
	wire [11-1:0] node462;
	wire [11-1:0] node464;
	wire [11-1:0] node467;
	wire [11-1:0] node470;
	wire [11-1:0] node471;
	wire [11-1:0] node472;
	wire [11-1:0] node473;
	wire [11-1:0] node475;
	wire [11-1:0] node479;
	wire [11-1:0] node480;
	wire [11-1:0] node481;
	wire [11-1:0] node483;
	wire [11-1:0] node486;
	wire [11-1:0] node489;
	wire [11-1:0] node492;
	wire [11-1:0] node493;
	wire [11-1:0] node494;
	wire [11-1:0] node495;
	wire [11-1:0] node498;
	wire [11-1:0] node501;
	wire [11-1:0] node502;
	wire [11-1:0] node503;
	wire [11-1:0] node507;
	wire [11-1:0] node509;
	wire [11-1:0] node512;
	wire [11-1:0] node513;
	wire [11-1:0] node514;
	wire [11-1:0] node516;
	wire [11-1:0] node519;
	wire [11-1:0] node520;
	wire [11-1:0] node524;
	wire [11-1:0] node525;
	wire [11-1:0] node528;
	wire [11-1:0] node530;
	wire [11-1:0] node533;
	wire [11-1:0] node534;
	wire [11-1:0] node535;
	wire [11-1:0] node536;
	wire [11-1:0] node537;
	wire [11-1:0] node538;
	wire [11-1:0] node539;
	wire [11-1:0] node541;
	wire [11-1:0] node544;
	wire [11-1:0] node545;
	wire [11-1:0] node549;
	wire [11-1:0] node550;
	wire [11-1:0] node551;
	wire [11-1:0] node552;
	wire [11-1:0] node557;
	wire [11-1:0] node558;
	wire [11-1:0] node559;
	wire [11-1:0] node562;
	wire [11-1:0] node564;
	wire [11-1:0] node567;
	wire [11-1:0] node568;
	wire [11-1:0] node572;
	wire [11-1:0] node573;
	wire [11-1:0] node574;
	wire [11-1:0] node575;
	wire [11-1:0] node578;
	wire [11-1:0] node582;
	wire [11-1:0] node583;
	wire [11-1:0] node584;
	wire [11-1:0] node587;
	wire [11-1:0] node590;
	wire [11-1:0] node591;
	wire [11-1:0] node592;
	wire [11-1:0] node596;
	wire [11-1:0] node598;
	wire [11-1:0] node601;
	wire [11-1:0] node602;
	wire [11-1:0] node603;
	wire [11-1:0] node604;
	wire [11-1:0] node605;
	wire [11-1:0] node606;
	wire [11-1:0] node609;
	wire [11-1:0] node610;
	wire [11-1:0] node615;
	wire [11-1:0] node616;
	wire [11-1:0] node617;
	wire [11-1:0] node621;
	wire [11-1:0] node624;
	wire [11-1:0] node625;
	wire [11-1:0] node627;
	wire [11-1:0] node629;
	wire [11-1:0] node632;
	wire [11-1:0] node633;
	wire [11-1:0] node635;
	wire [11-1:0] node639;
	wire [11-1:0] node640;
	wire [11-1:0] node642;
	wire [11-1:0] node643;
	wire [11-1:0] node644;
	wire [11-1:0] node647;
	wire [11-1:0] node650;
	wire [11-1:0] node653;
	wire [11-1:0] node655;
	wire [11-1:0] node658;
	wire [11-1:0] node659;
	wire [11-1:0] node660;
	wire [11-1:0] node661;
	wire [11-1:0] node662;
	wire [11-1:0] node663;
	wire [11-1:0] node666;
	wire [11-1:0] node667;
	wire [11-1:0] node670;
	wire [11-1:0] node673;
	wire [11-1:0] node674;
	wire [11-1:0] node675;
	wire [11-1:0] node678;
	wire [11-1:0] node682;
	wire [11-1:0] node683;
	wire [11-1:0] node684;
	wire [11-1:0] node685;
	wire [11-1:0] node690;
	wire [11-1:0] node692;
	wire [11-1:0] node695;
	wire [11-1:0] node696;
	wire [11-1:0] node697;
	wire [11-1:0] node698;
	wire [11-1:0] node700;
	wire [11-1:0] node704;
	wire [11-1:0] node707;
	wire [11-1:0] node708;
	wire [11-1:0] node709;
	wire [11-1:0] node712;
	wire [11-1:0] node715;
	wire [11-1:0] node717;
	wire [11-1:0] node719;
	wire [11-1:0] node722;
	wire [11-1:0] node723;
	wire [11-1:0] node724;
	wire [11-1:0] node725;
	wire [11-1:0] node727;
	wire [11-1:0] node729;
	wire [11-1:0] node732;
	wire [11-1:0] node733;
	wire [11-1:0] node736;
	wire [11-1:0] node739;
	wire [11-1:0] node740;
	wire [11-1:0] node741;
	wire [11-1:0] node744;
	wire [11-1:0] node745;
	wire [11-1:0] node749;
	wire [11-1:0] node751;
	wire [11-1:0] node753;
	wire [11-1:0] node756;
	wire [11-1:0] node757;
	wire [11-1:0] node758;
	wire [11-1:0] node760;
	wire [11-1:0] node763;
	wire [11-1:0] node764;
	wire [11-1:0] node768;
	wire [11-1:0] node769;
	wire [11-1:0] node770;
	wire [11-1:0] node771;
	wire [11-1:0] node775;
	wire [11-1:0] node776;
	wire [11-1:0] node780;
	wire [11-1:0] node781;
	wire [11-1:0] node782;
	wire [11-1:0] node785;
	wire [11-1:0] node788;
	wire [11-1:0] node791;
	wire [11-1:0] node792;
	wire [11-1:0] node793;
	wire [11-1:0] node794;
	wire [11-1:0] node795;
	wire [11-1:0] node796;
	wire [11-1:0] node797;
	wire [11-1:0] node801;
	wire [11-1:0] node802;
	wire [11-1:0] node804;
	wire [11-1:0] node807;
	wire [11-1:0] node810;
	wire [11-1:0] node811;
	wire [11-1:0] node812;
	wire [11-1:0] node813;
	wire [11-1:0] node816;
	wire [11-1:0] node819;
	wire [11-1:0] node822;
	wire [11-1:0] node825;
	wire [11-1:0] node826;
	wire [11-1:0] node827;
	wire [11-1:0] node828;
	wire [11-1:0] node831;
	wire [11-1:0] node832;
	wire [11-1:0] node836;
	wire [11-1:0] node837;
	wire [11-1:0] node841;
	wire [11-1:0] node842;
	wire [11-1:0] node843;
	wire [11-1:0] node847;
	wire [11-1:0] node848;
	wire [11-1:0] node852;
	wire [11-1:0] node853;
	wire [11-1:0] node854;
	wire [11-1:0] node855;
	wire [11-1:0] node858;
	wire [11-1:0] node861;
	wire [11-1:0] node862;
	wire [11-1:0] node863;
	wire [11-1:0] node865;
	wire [11-1:0] node868;
	wire [11-1:0] node870;
	wire [11-1:0] node873;
	wire [11-1:0] node874;
	wire [11-1:0] node875;
	wire [11-1:0] node879;
	wire [11-1:0] node880;
	wire [11-1:0] node884;
	wire [11-1:0] node885;
	wire [11-1:0] node886;
	wire [11-1:0] node888;
	wire [11-1:0] node889;
	wire [11-1:0] node891;
	wire [11-1:0] node894;
	wire [11-1:0] node897;
	wire [11-1:0] node900;
	wire [11-1:0] node901;
	wire [11-1:0] node902;
	wire [11-1:0] node903;
	wire [11-1:0] node904;
	wire [11-1:0] node910;
	wire [11-1:0] node913;
	wire [11-1:0] node914;
	wire [11-1:0] node915;
	wire [11-1:0] node916;
	wire [11-1:0] node917;
	wire [11-1:0] node920;
	wire [11-1:0] node923;
	wire [11-1:0] node924;
	wire [11-1:0] node925;
	wire [11-1:0] node928;
	wire [11-1:0] node929;
	wire [11-1:0] node933;
	wire [11-1:0] node934;
	wire [11-1:0] node938;
	wire [11-1:0] node939;
	wire [11-1:0] node940;
	wire [11-1:0] node941;
	wire [11-1:0] node943;
	wire [11-1:0] node947;
	wire [11-1:0] node950;
	wire [11-1:0] node951;
	wire [11-1:0] node953;
	wire [11-1:0] node956;
	wire [11-1:0] node957;
	wire [11-1:0] node958;
	wire [11-1:0] node961;
	wire [11-1:0] node964;
	wire [11-1:0] node965;
	wire [11-1:0] node969;
	wire [11-1:0] node970;
	wire [11-1:0] node971;
	wire [11-1:0] node972;
	wire [11-1:0] node974;
	wire [11-1:0] node977;
	wire [11-1:0] node978;
	wire [11-1:0] node980;
	wire [11-1:0] node983;
	wire [11-1:0] node984;
	wire [11-1:0] node988;
	wire [11-1:0] node989;
	wire [11-1:0] node992;
	wire [11-1:0] node993;
	wire [11-1:0] node996;
	wire [11-1:0] node999;
	wire [11-1:0] node1000;
	wire [11-1:0] node1001;
	wire [11-1:0] node1003;
	wire [11-1:0] node1005;
	wire [11-1:0] node1008;
	wire [11-1:0] node1009;
	wire [11-1:0] node1012;
	wire [11-1:0] node1014;
	wire [11-1:0] node1017;
	wire [11-1:0] node1018;
	wire [11-1:0] node1019;
	wire [11-1:0] node1023;
	wire [11-1:0] node1024;
	wire [11-1:0] node1027;
	wire [11-1:0] node1028;
	wire [11-1:0] node1032;
	wire [11-1:0] node1033;
	wire [11-1:0] node1034;
	wire [11-1:0] node1035;
	wire [11-1:0] node1036;
	wire [11-1:0] node1037;
	wire [11-1:0] node1038;
	wire [11-1:0] node1040;
	wire [11-1:0] node1042;
	wire [11-1:0] node1045;
	wire [11-1:0] node1046;
	wire [11-1:0] node1047;
	wire [11-1:0] node1048;
	wire [11-1:0] node1052;
	wire [11-1:0] node1054;
	wire [11-1:0] node1057;
	wire [11-1:0] node1059;
	wire [11-1:0] node1060;
	wire [11-1:0] node1064;
	wire [11-1:0] node1065;
	wire [11-1:0] node1066;
	wire [11-1:0] node1068;
	wire [11-1:0] node1071;
	wire [11-1:0] node1073;
	wire [11-1:0] node1076;
	wire [11-1:0] node1077;
	wire [11-1:0] node1080;
	wire [11-1:0] node1081;
	wire [11-1:0] node1082;
	wire [11-1:0] node1083;
	wire [11-1:0] node1087;
	wire [11-1:0] node1090;
	wire [11-1:0] node1093;
	wire [11-1:0] node1094;
	wire [11-1:0] node1095;
	wire [11-1:0] node1096;
	wire [11-1:0] node1097;
	wire [11-1:0] node1101;
	wire [11-1:0] node1102;
	wire [11-1:0] node1106;
	wire [11-1:0] node1108;
	wire [11-1:0] node1111;
	wire [11-1:0] node1112;
	wire [11-1:0] node1113;
	wire [11-1:0] node1114;
	wire [11-1:0] node1116;
	wire [11-1:0] node1117;
	wire [11-1:0] node1122;
	wire [11-1:0] node1124;
	wire [11-1:0] node1125;
	wire [11-1:0] node1128;
	wire [11-1:0] node1131;
	wire [11-1:0] node1132;
	wire [11-1:0] node1133;
	wire [11-1:0] node1136;
	wire [11-1:0] node1139;
	wire [11-1:0] node1140;
	wire [11-1:0] node1142;
	wire [11-1:0] node1145;
	wire [11-1:0] node1148;
	wire [11-1:0] node1149;
	wire [11-1:0] node1150;
	wire [11-1:0] node1151;
	wire [11-1:0] node1152;
	wire [11-1:0] node1153;
	wire [11-1:0] node1157;
	wire [11-1:0] node1159;
	wire [11-1:0] node1162;
	wire [11-1:0] node1163;
	wire [11-1:0] node1166;
	wire [11-1:0] node1167;
	wire [11-1:0] node1170;
	wire [11-1:0] node1173;
	wire [11-1:0] node1174;
	wire [11-1:0] node1175;
	wire [11-1:0] node1176;
	wire [11-1:0] node1179;
	wire [11-1:0] node1181;
	wire [11-1:0] node1183;
	wire [11-1:0] node1186;
	wire [11-1:0] node1189;
	wire [11-1:0] node1190;
	wire [11-1:0] node1193;
	wire [11-1:0] node1196;
	wire [11-1:0] node1197;
	wire [11-1:0] node1198;
	wire [11-1:0] node1199;
	wire [11-1:0] node1200;
	wire [11-1:0] node1204;
	wire [11-1:0] node1205;
	wire [11-1:0] node1209;
	wire [11-1:0] node1210;
	wire [11-1:0] node1211;
	wire [11-1:0] node1214;
	wire [11-1:0] node1217;
	wire [11-1:0] node1220;
	wire [11-1:0] node1221;
	wire [11-1:0] node1222;
	wire [11-1:0] node1224;
	wire [11-1:0] node1227;
	wire [11-1:0] node1228;
	wire [11-1:0] node1229;
	wire [11-1:0] node1232;
	wire [11-1:0] node1235;
	wire [11-1:0] node1236;
	wire [11-1:0] node1239;
	wire [11-1:0] node1240;
	wire [11-1:0] node1244;
	wire [11-1:0] node1245;
	wire [11-1:0] node1246;
	wire [11-1:0] node1247;
	wire [11-1:0] node1250;
	wire [11-1:0] node1253;
	wire [11-1:0] node1256;
	wire [11-1:0] node1258;
	wire [11-1:0] node1259;
	wire [11-1:0] node1261;
	wire [11-1:0] node1265;
	wire [11-1:0] node1266;
	wire [11-1:0] node1267;
	wire [11-1:0] node1268;
	wire [11-1:0] node1269;
	wire [11-1:0] node1270;
	wire [11-1:0] node1271;
	wire [11-1:0] node1275;
	wire [11-1:0] node1277;
	wire [11-1:0] node1279;
	wire [11-1:0] node1282;
	wire [11-1:0] node1284;
	wire [11-1:0] node1285;
	wire [11-1:0] node1286;
	wire [11-1:0] node1287;
	wire [11-1:0] node1291;
	wire [11-1:0] node1295;
	wire [11-1:0] node1296;
	wire [11-1:0] node1297;
	wire [11-1:0] node1298;
	wire [11-1:0] node1302;
	wire [11-1:0] node1304;
	wire [11-1:0] node1305;
	wire [11-1:0] node1309;
	wire [11-1:0] node1310;
	wire [11-1:0] node1312;
	wire [11-1:0] node1313;
	wire [11-1:0] node1317;
	wire [11-1:0] node1319;
	wire [11-1:0] node1322;
	wire [11-1:0] node1323;
	wire [11-1:0] node1324;
	wire [11-1:0] node1325;
	wire [11-1:0] node1327;
	wire [11-1:0] node1328;
	wire [11-1:0] node1332;
	wire [11-1:0] node1333;
	wire [11-1:0] node1336;
	wire [11-1:0] node1339;
	wire [11-1:0] node1341;
	wire [11-1:0] node1344;
	wire [11-1:0] node1345;
	wire [11-1:0] node1346;
	wire [11-1:0] node1348;
	wire [11-1:0] node1349;
	wire [11-1:0] node1352;
	wire [11-1:0] node1355;
	wire [11-1:0] node1358;
	wire [11-1:0] node1359;
	wire [11-1:0] node1362;
	wire [11-1:0] node1365;
	wire [11-1:0] node1366;
	wire [11-1:0] node1367;
	wire [11-1:0] node1368;
	wire [11-1:0] node1369;
	wire [11-1:0] node1370;
	wire [11-1:0] node1374;
	wire [11-1:0] node1375;
	wire [11-1:0] node1378;
	wire [11-1:0] node1380;
	wire [11-1:0] node1383;
	wire [11-1:0] node1384;
	wire [11-1:0] node1387;
	wire [11-1:0] node1389;
	wire [11-1:0] node1390;
	wire [11-1:0] node1394;
	wire [11-1:0] node1395;
	wire [11-1:0] node1396;
	wire [11-1:0] node1399;
	wire [11-1:0] node1400;
	wire [11-1:0] node1401;
	wire [11-1:0] node1405;
	wire [11-1:0] node1407;
	wire [11-1:0] node1408;
	wire [11-1:0] node1412;
	wire [11-1:0] node1413;
	wire [11-1:0] node1414;
	wire [11-1:0] node1416;
	wire [11-1:0] node1419;
	wire [11-1:0] node1422;
	wire [11-1:0] node1423;
	wire [11-1:0] node1424;
	wire [11-1:0] node1428;
	wire [11-1:0] node1430;
	wire [11-1:0] node1433;
	wire [11-1:0] node1434;
	wire [11-1:0] node1435;
	wire [11-1:0] node1436;
	wire [11-1:0] node1439;
	wire [11-1:0] node1441;
	wire [11-1:0] node1442;
	wire [11-1:0] node1446;
	wire [11-1:0] node1447;
	wire [11-1:0] node1448;
	wire [11-1:0] node1452;
	wire [11-1:0] node1453;
	wire [11-1:0] node1454;
	wire [11-1:0] node1458;
	wire [11-1:0] node1460;
	wire [11-1:0] node1463;
	wire [11-1:0] node1464;
	wire [11-1:0] node1465;
	wire [11-1:0] node1466;
	wire [11-1:0] node1468;
	wire [11-1:0] node1472;
	wire [11-1:0] node1474;
	wire [11-1:0] node1477;
	wire [11-1:0] node1478;
	wire [11-1:0] node1479;
	wire [11-1:0] node1481;
	wire [11-1:0] node1484;
	wire [11-1:0] node1488;
	wire [11-1:0] node1489;
	wire [11-1:0] node1490;
	wire [11-1:0] node1491;
	wire [11-1:0] node1492;
	wire [11-1:0] node1493;
	wire [11-1:0] node1494;
	wire [11-1:0] node1497;
	wire [11-1:0] node1499;
	wire [11-1:0] node1500;
	wire [11-1:0] node1504;
	wire [11-1:0] node1506;
	wire [11-1:0] node1509;
	wire [11-1:0] node1510;
	wire [11-1:0] node1511;
	wire [11-1:0] node1512;
	wire [11-1:0] node1514;
	wire [11-1:0] node1517;
	wire [11-1:0] node1518;
	wire [11-1:0] node1522;
	wire [11-1:0] node1523;
	wire [11-1:0] node1526;
	wire [11-1:0] node1529;
	wire [11-1:0] node1530;
	wire [11-1:0] node1531;
	wire [11-1:0] node1534;
	wire [11-1:0] node1537;
	wire [11-1:0] node1538;
	wire [11-1:0] node1539;
	wire [11-1:0] node1542;
	wire [11-1:0] node1545;
	wire [11-1:0] node1546;
	wire [11-1:0] node1549;
	wire [11-1:0] node1552;
	wire [11-1:0] node1553;
	wire [11-1:0] node1554;
	wire [11-1:0] node1555;
	wire [11-1:0] node1556;
	wire [11-1:0] node1561;
	wire [11-1:0] node1562;
	wire [11-1:0] node1563;
	wire [11-1:0] node1566;
	wire [11-1:0] node1568;
	wire [11-1:0] node1569;
	wire [11-1:0] node1573;
	wire [11-1:0] node1574;
	wire [11-1:0] node1577;
	wire [11-1:0] node1578;
	wire [11-1:0] node1579;
	wire [11-1:0] node1584;
	wire [11-1:0] node1585;
	wire [11-1:0] node1586;
	wire [11-1:0] node1587;
	wire [11-1:0] node1590;
	wire [11-1:0] node1593;
	wire [11-1:0] node1596;
	wire [11-1:0] node1597;
	wire [11-1:0] node1600;
	wire [11-1:0] node1601;
	wire [11-1:0] node1602;
	wire [11-1:0] node1606;
	wire [11-1:0] node1608;
	wire [11-1:0] node1609;
	wire [11-1:0] node1613;
	wire [11-1:0] node1614;
	wire [11-1:0] node1615;
	wire [11-1:0] node1616;
	wire [11-1:0] node1617;
	wire [11-1:0] node1618;
	wire [11-1:0] node1619;
	wire [11-1:0] node1621;
	wire [11-1:0] node1625;
	wire [11-1:0] node1628;
	wire [11-1:0] node1629;
	wire [11-1:0] node1631;
	wire [11-1:0] node1633;
	wire [11-1:0] node1636;
	wire [11-1:0] node1639;
	wire [11-1:0] node1640;
	wire [11-1:0] node1641;
	wire [11-1:0] node1643;
	wire [11-1:0] node1645;
	wire [11-1:0] node1648;
	wire [11-1:0] node1649;
	wire [11-1:0] node1652;
	wire [11-1:0] node1654;
	wire [11-1:0] node1657;
	wire [11-1:0] node1658;
	wire [11-1:0] node1660;
	wire [11-1:0] node1663;
	wire [11-1:0] node1666;
	wire [11-1:0] node1667;
	wire [11-1:0] node1668;
	wire [11-1:0] node1669;
	wire [11-1:0] node1670;
	wire [11-1:0] node1673;
	wire [11-1:0] node1676;
	wire [11-1:0] node1678;
	wire [11-1:0] node1681;
	wire [11-1:0] node1682;
	wire [11-1:0] node1685;
	wire [11-1:0] node1687;
	wire [11-1:0] node1688;
	wire [11-1:0] node1692;
	wire [11-1:0] node1693;
	wire [11-1:0] node1694;
	wire [11-1:0] node1697;
	wire [11-1:0] node1700;
	wire [11-1:0] node1701;
	wire [11-1:0] node1702;
	wire [11-1:0] node1703;
	wire [11-1:0] node1709;
	wire [11-1:0] node1710;
	wire [11-1:0] node1711;
	wire [11-1:0] node1712;
	wire [11-1:0] node1713;
	wire [11-1:0] node1717;
	wire [11-1:0] node1718;
	wire [11-1:0] node1721;
	wire [11-1:0] node1724;
	wire [11-1:0] node1725;
	wire [11-1:0] node1726;
	wire [11-1:0] node1727;
	wire [11-1:0] node1732;
	wire [11-1:0] node1733;
	wire [11-1:0] node1737;
	wire [11-1:0] node1738;
	wire [11-1:0] node1739;
	wire [11-1:0] node1740;
	wire [11-1:0] node1744;
	wire [11-1:0] node1747;
	wire [11-1:0] node1748;
	wire [11-1:0] node1749;
	wire [11-1:0] node1753;
	wire [11-1:0] node1754;
	wire [11-1:0] node1757;
	wire [11-1:0] node1758;
	wire [11-1:0] node1762;
	wire [11-1:0] node1763;
	wire [11-1:0] node1764;
	wire [11-1:0] node1765;
	wire [11-1:0] node1766;
	wire [11-1:0] node1767;
	wire [11-1:0] node1769;
	wire [11-1:0] node1770;
	wire [11-1:0] node1774;
	wire [11-1:0] node1776;
	wire [11-1:0] node1779;
	wire [11-1:0] node1780;
	wire [11-1:0] node1781;
	wire [11-1:0] node1782;
	wire [11-1:0] node1786;
	wire [11-1:0] node1790;
	wire [11-1:0] node1791;
	wire [11-1:0] node1792;
	wire [11-1:0] node1793;
	wire [11-1:0] node1796;
	wire [11-1:0] node1800;
	wire [11-1:0] node1801;
	wire [11-1:0] node1802;
	wire [11-1:0] node1803;
	wire [11-1:0] node1808;
	wire [11-1:0] node1809;
	wire [11-1:0] node1810;
	wire [11-1:0] node1811;
	wire [11-1:0] node1816;
	wire [11-1:0] node1819;
	wire [11-1:0] node1820;
	wire [11-1:0] node1821;
	wire [11-1:0] node1822;
	wire [11-1:0] node1825;
	wire [11-1:0] node1826;
	wire [11-1:0] node1827;
	wire [11-1:0] node1832;
	wire [11-1:0] node1833;
	wire [11-1:0] node1834;
	wire [11-1:0] node1837;
	wire [11-1:0] node1840;
	wire [11-1:0] node1841;
	wire [11-1:0] node1844;
	wire [11-1:0] node1846;
	wire [11-1:0] node1848;
	wire [11-1:0] node1851;
	wire [11-1:0] node1852;
	wire [11-1:0] node1853;
	wire [11-1:0] node1855;
	wire [11-1:0] node1857;
	wire [11-1:0] node1860;
	wire [11-1:0] node1861;
	wire [11-1:0] node1863;
	wire [11-1:0] node1865;
	wire [11-1:0] node1868;
	wire [11-1:0] node1871;
	wire [11-1:0] node1873;
	wire [11-1:0] node1875;
	wire [11-1:0] node1877;
	wire [11-1:0] node1880;
	wire [11-1:0] node1881;
	wire [11-1:0] node1882;
	wire [11-1:0] node1883;
	wire [11-1:0] node1884;
	wire [11-1:0] node1886;
	wire [11-1:0] node1888;
	wire [11-1:0] node1891;
	wire [11-1:0] node1892;
	wire [11-1:0] node1893;
	wire [11-1:0] node1897;
	wire [11-1:0] node1900;
	wire [11-1:0] node1901;
	wire [11-1:0] node1902;
	wire [11-1:0] node1905;
	wire [11-1:0] node1908;
	wire [11-1:0] node1910;
	wire [11-1:0] node1913;
	wire [11-1:0] node1914;
	wire [11-1:0] node1915;
	wire [11-1:0] node1916;
	wire [11-1:0] node1917;
	wire [11-1:0] node1921;
	wire [11-1:0] node1925;
	wire [11-1:0] node1926;
	wire [11-1:0] node1927;
	wire [11-1:0] node1931;
	wire [11-1:0] node1932;
	wire [11-1:0] node1934;
	wire [11-1:0] node1938;
	wire [11-1:0] node1939;
	wire [11-1:0] node1940;
	wire [11-1:0] node1941;
	wire [11-1:0] node1942;
	wire [11-1:0] node1945;
	wire [11-1:0] node1947;
	wire [11-1:0] node1950;
	wire [11-1:0] node1951;
	wire [11-1:0] node1952;
	wire [11-1:0] node1956;
	wire [11-1:0] node1959;
	wire [11-1:0] node1960;
	wire [11-1:0] node1961;
	wire [11-1:0] node1962;
	wire [11-1:0] node1967;
	wire [11-1:0] node1968;
	wire [11-1:0] node1971;
	wire [11-1:0] node1974;
	wire [11-1:0] node1975;
	wire [11-1:0] node1976;
	wire [11-1:0] node1977;
	wire [11-1:0] node1981;
	wire [11-1:0] node1982;
	wire [11-1:0] node1984;
	wire [11-1:0] node1988;
	wire [11-1:0] node1989;
	wire [11-1:0] node1992;

	assign outp = (inp[1]) ? node1032 : node1;
		assign node1 = (inp[7]) ? node533 : node2;
			assign node2 = (inp[2]) ? node280 : node3;
				assign node3 = (inp[0]) ? node133 : node4;
					assign node4 = (inp[11]) ? node70 : node5;
						assign node5 = (inp[5]) ? node39 : node6;
							assign node6 = (inp[6]) ? node18 : node7;
								assign node7 = (inp[10]) ? node13 : node8;
									assign node8 = (inp[4]) ? node10 : 11'b11001101011;
										assign node10 = (inp[8]) ? 11'b11001001111 : 11'b01001001111;
									assign node13 = (inp[4]) ? 11'b11100001011 : node14;
										assign node14 = (inp[8]) ? 11'b01100101111 : 11'b11000111111;
								assign node18 = (inp[8]) ? node28 : node19;
									assign node19 = (inp[10]) ? 11'b11001010110 : node20;
										assign node20 = (inp[3]) ? 11'b11011100010 : node21;
											assign node21 = (inp[4]) ? 11'b01000100110 : node22;
												assign node22 = (inp[9]) ? 11'b01000100000 : 11'b01001100010;
									assign node28 = (inp[3]) ? node36 : node29;
										assign node29 = (inp[10]) ? 11'b11000101010 : node30;
											assign node30 = (inp[4]) ? 11'b01111101100 : node31;
												assign node31 = (inp[9]) ? 11'b01010001000 : 11'b01000101010;
										assign node36 = (inp[4]) ? 11'b11010111010 : 11'b01111011110;
							assign node39 = (inp[6]) ? node55 : node40;
								assign node40 = (inp[4]) ? node50 : node41;
									assign node41 = (inp[10]) ? node47 : node42;
										assign node42 = (inp[3]) ? 11'b11001111010 : node43;
											assign node43 = (inp[9]) ? 11'b01010111010 : 11'b01000011011;
										assign node47 = (inp[3]) ? 11'b01101101100 : 11'b11100111010;
									assign node50 = (inp[10]) ? 11'b01010011010 : node51;
										assign node51 = (inp[3]) ? 11'b11111011110 : 11'b01011011110;
								assign node55 = (inp[8]) ? node65 : node56;
									assign node56 = (inp[10]) ? node62 : node57;
										assign node57 = (inp[3]) ? node59 : 11'b01010111111;
											assign node59 = (inp[9]) ? 11'b11001111111 : 11'b11100111101;
										assign node62 = (inp[9]) ? 11'b11111101111 : 11'b11001101101;
									assign node65 = (inp[4]) ? node67 : 11'b11110111001;
										assign node67 = (inp[3]) ? 11'b01110001001 : 11'b11000001111;
						assign node70 = (inp[10]) ? node98 : node71;
							assign node71 = (inp[3]) ? node79 : node72;
								assign node72 = (inp[9]) ? 11'b01111111001 : node73;
									assign node73 = (inp[4]) ? 11'b01011001111 : node74;
										assign node74 = (inp[6]) ? 11'b01010011011 : 11'b01000001001;
								assign node79 = (inp[5]) ? node87 : node80;
									assign node80 = (inp[9]) ? node82 : 11'b11010101101;
										assign node82 = (inp[6]) ? 11'b11011011001 : node83;
											assign node83 = (inp[8]) ? 11'b11010011011 : 11'b11011011011;
									assign node87 = (inp[4]) ? node91 : node88;
										assign node88 = (inp[9]) ? 11'b11010011111 : 11'b11100001001;
										assign node91 = (inp[8]) ? 11'b11100111101 : node92;
											assign node92 = (inp[9]) ? 11'b11101101000 : node93;
												assign node93 = (inp[6]) ? 11'b11111111100 : 11'b11101011100;
							assign node98 = (inp[3]) ? node112 : node99;
								assign node99 = (inp[6]) ? node101 : 11'b11010011010;
									assign node101 = (inp[8]) ? node105 : node102;
										assign node102 = (inp[5]) ? 11'b11110011001 : 11'b11100011011;
										assign node105 = (inp[5]) ? node109 : node106;
											assign node106 = (inp[9]) ? 11'b11111111001 : 11'b11110101000;
											assign node109 = (inp[4]) ? 11'b11110101101 : 11'b11001111001;
								assign node112 = (inp[4]) ? node126 : node113;
									assign node113 = (inp[5]) ? node117 : node114;
										assign node114 = (inp[8]) ? 11'b01100011100 : 11'b01000111111;
										assign node117 = (inp[8]) ? node121 : node118;
											assign node118 = (inp[9]) ? 11'b01000101100 : 11'b01001001111;
											assign node121 = (inp[9]) ? node123 : 11'b01011101101;
												assign node123 = (inp[6]) ? 11'b01111101111 : 11'b01111101110;
									assign node126 = (inp[6]) ? 11'b01110101000 : node127;
										assign node127 = (inp[8]) ? 11'b01110101000 : node128;
											assign node128 = (inp[9]) ? 11'b01110001000 : 11'b01100001000;
					assign node133 = (inp[3]) ? node207 : node134;
						assign node134 = (inp[4]) ? node160 : node135;
							assign node135 = (inp[11]) ? node149 : node136;
								assign node136 = (inp[5]) ? node142 : node137;
									assign node137 = (inp[8]) ? node139 : 11'b01011100000;
										assign node139 = (inp[6]) ? 11'b01111001100 : 11'b01101101101;
									assign node142 = (inp[10]) ? node146 : node143;
										assign node143 = (inp[9]) ? 11'b01110101100 : 11'b01110101001;
										assign node146 = (inp[8]) ? 11'b01001111010 : 11'b01100111000;
								assign node149 = (inp[5]) ? node153 : node150;
									assign node150 = (inp[8]) ? 11'b01000111111 : 11'b01101111101;
									assign node153 = (inp[6]) ? node157 : node154;
										assign node154 = (inp[9]) ? 11'b01111111110 : 11'b01110011100;
										assign node157 = (inp[8]) ? 11'b01101111111 : 11'b01000011101;
							assign node160 = (inp[11]) ? node184 : node161;
								assign node161 = (inp[10]) ? node171 : node162;
									assign node162 = (inp[9]) ? node168 : node163;
										assign node163 = (inp[8]) ? 11'b01010101010 : node164;
											assign node164 = (inp[6]) ? 11'b01010100000 : 11'b01111001000;
										assign node168 = (inp[8]) ? 11'b01001111100 : 11'b01110010110;
									assign node171 = (inp[9]) ? node177 : node172;
										assign node172 = (inp[6]) ? node174 : 11'b01000011101;
											assign node174 = (inp[5]) ? 11'b01001111111 : 11'b01111111110;
										assign node177 = (inp[8]) ? node181 : node178;
											assign node178 = (inp[5]) ? 11'b01111011001 : 11'b01111010010;
											assign node181 = (inp[5]) ? 11'b01010011011 : 11'b01010111000;
								assign node184 = (inp[9]) ? node192 : node185;
									assign node185 = (inp[10]) ? 11'b01110001101 : node186;
										assign node186 = (inp[8]) ? node188 : 11'b01111111010;
											assign node188 = (inp[6]) ? 11'b01010111011 : 11'b01001111010;
									assign node192 = (inp[10]) ? node198 : node193;
										assign node193 = (inp[8]) ? 11'b01011001101 : node194;
											assign node194 = (inp[6]) ? 11'b01001001111 : 11'b01011001101;
										assign node198 = (inp[8]) ? node202 : node199;
											assign node199 = (inp[6]) ? 11'b01100001001 : 11'b01110001001;
											assign node202 = (inp[5]) ? 11'b01000001011 : node203;
												assign node203 = (inp[6]) ? 11'b01001101001 : 11'b01011001001;
						assign node207 = (inp[10]) ? node233 : node208;
							assign node208 = (inp[6]) ? node216 : node209;
								assign node209 = (inp[9]) ? node213 : node210;
									assign node210 = (inp[11]) ? 11'b01011101011 : 11'b01001101001;
									assign node213 = (inp[11]) ? 11'b01101111011 : 11'b01101001001;
								assign node216 = (inp[9]) ? node224 : node217;
									assign node217 = (inp[4]) ? node221 : node218;
										assign node218 = (inp[11]) ? 11'b01100001011 : 11'b01100101011;
										assign node221 = (inp[8]) ? 11'b01110011011 : 11'b01111111011;
									assign node224 = (inp[4]) ? node230 : node225;
										assign node225 = (inp[8]) ? 11'b01101011010 : node226;
											assign node226 = (inp[5]) ? 11'b01101111001 : 11'b01100111011;
										assign node230 = (inp[8]) ? 11'b01110101000 : 11'b01101000010;
							assign node233 = (inp[9]) ? node261 : node234;
								assign node234 = (inp[5]) ? node248 : node235;
									assign node235 = (inp[6]) ? node243 : node236;
										assign node236 = (inp[4]) ? 11'b01010001001 : node237;
											assign node237 = (inp[8]) ? node239 : 11'b01100101001;
												assign node239 = (inp[11]) ? 11'b01110101011 : 11'b01010101001;
										assign node243 = (inp[8]) ? node245 : 11'b01000100010;
											assign node245 = (inp[4]) ? 11'b01111101010 : 11'b01110101000;
									assign node248 = (inp[6]) ? node254 : node249;
										assign node249 = (inp[8]) ? node251 : 11'b01010001010;
											assign node251 = (inp[11]) ? 11'b01001001010 : 11'b01101001010;
										assign node254 = (inp[4]) ? node258 : node255;
											assign node255 = (inp[8]) ? 11'b01011101011 : 11'b01000001011;
											assign node258 = (inp[8]) ? 11'b01100001001 : 11'b01110101011;
								assign node261 = (inp[4]) ? node273 : node262;
									assign node262 = (inp[8]) ? node266 : node263;
										assign node263 = (inp[5]) ? 11'b01010101000 : 11'b01000101001;
										assign node266 = (inp[6]) ? node268 : 11'b01001101010;
											assign node268 = (inp[5]) ? 11'b01011001011 : node269;
												assign node269 = (inp[11]) ? 11'b01010001010 : 11'b01001001000;
									assign node273 = (inp[11]) ? 11'b01000001000 : node274;
										assign node274 = (inp[8]) ? node276 : 11'b01000001001;
											assign node276 = (inp[5]) ? 11'b01000001001 : 11'b01000001011;
				assign node280 = (inp[0]) ? node400 : node281;
					assign node281 = (inp[8]) ? node341 : node282;
						assign node282 = (inp[4]) ? node320 : node283;
							assign node283 = (inp[9]) ? node297 : node284;
								assign node284 = (inp[5]) ? node292 : node285;
									assign node285 = (inp[3]) ? node289 : node286;
										assign node286 = (inp[6]) ? 11'b01101001011 : 11'b01101001010;
										assign node289 = (inp[11]) ? 11'b11100011010 : 11'b01110001110;
									assign node292 = (inp[6]) ? node294 : 11'b01101010000;
										assign node294 = (inp[3]) ? 11'b11010100001 : 11'b01110110001;
								assign node297 = (inp[3]) ? node305 : node298;
									assign node298 = (inp[10]) ? node300 : 11'b01010010011;
										assign node300 = (inp[5]) ? 11'b11010100101 : node301;
											assign node301 = (inp[6]) ? 11'b11000011110 : 11'b11110110111;
									assign node305 = (inp[10]) ? node315 : node306;
										assign node306 = (inp[5]) ? node308 : 11'b11101100111;
											assign node308 = (inp[11]) ? node312 : node309;
												assign node309 = (inp[6]) ? 11'b11100011110 : 11'b11110010101;
												assign node312 = (inp[6]) ? 11'b11110110101 : 11'b11101010110;
										assign node315 = (inp[11]) ? node317 : 11'b01110111110;
											assign node317 = (inp[6]) ? 11'b01111000111 : 11'b01110000110;
							assign node320 = (inp[5]) ? node336 : node321;
								assign node321 = (inp[10]) ? node329 : node322;
									assign node322 = (inp[9]) ? node326 : node323;
										assign node323 = (inp[3]) ? 11'b11100101100 : 11'b01100101100;
										assign node326 = (inp[11]) ? 11'b11110111000 : 11'b11000111000;
									assign node329 = (inp[6]) ? node331 : 11'b11001110101;
										assign node331 = (inp[3]) ? 11'b01000111010 : node332;
											assign node332 = (inp[9]) ? 11'b11011111000 : 11'b11011111110;
								assign node336 = (inp[10]) ? node338 : 11'b11100100010;
									assign node338 = (inp[11]) ? 11'b01010000001 : 11'b01000100000;
						assign node341 = (inp[5]) ? node365 : node342;
							assign node342 = (inp[3]) ? node358 : node343;
								assign node343 = (inp[10]) ? node345 : 11'b01000000100;
									assign node345 = (inp[4]) ? node347 : 11'b11011000011;
										assign node347 = (inp[11]) ? node353 : node348;
											assign node348 = (inp[9]) ? node350 : 11'b11000110111;
												assign node350 = (inp[6]) ? 11'b11110000011 : 11'b11111100011;
											assign node353 = (inp[6]) ? node355 : 11'b11000110011;
												assign node355 = (inp[9]) ? 11'b11010110000 : 11'b11010110100;
								assign node358 = (inp[10]) ? node360 : 11'b11010110001;
									assign node360 = (inp[4]) ? node362 : 11'b01011010100;
										assign node362 = (inp[9]) ? 11'b01010010011 : 11'b01000010001;
							assign node365 = (inp[11]) ? node381 : node366;
								assign node366 = (inp[6]) ? node376 : node367;
									assign node367 = (inp[3]) ? node369 : 11'b11011110000;
										assign node369 = (inp[10]) ? node373 : node370;
											assign node370 = (inp[4]) ? 11'b11000000001 : 11'b11101010101;
											assign node373 = (inp[9]) ? 11'b01000000111 : 11'b01010110101;
									assign node376 = (inp[4]) ? node378 : 11'b01100010010;
										assign node378 = (inp[3]) ? 11'b01111110000 : 11'b01011110110;
								assign node381 = (inp[3]) ? node387 : node382;
									assign node382 = (inp[9]) ? node384 : 11'b11111110000;
										assign node384 = (inp[10]) ? 11'b11000100100 : 11'b01001000100;
									assign node387 = (inp[10]) ? node395 : node388;
										assign node388 = (inp[9]) ? node390 : 11'b11010010110;
											assign node390 = (inp[4]) ? node392 : 11'b11011010110;
												assign node392 = (inp[6]) ? 11'b11010000010 : 11'b11011000000;
										assign node395 = (inp[4]) ? node397 : 11'b01011000100;
											assign node397 = (inp[6]) ? 11'b01011000000 : 11'b01011000010;
					assign node400 = (inp[3]) ? node470 : node401;
						assign node401 = (inp[11]) ? node435 : node402;
							assign node402 = (inp[6]) ? node422 : node403;
								assign node403 = (inp[4]) ? node415 : node404;
									assign node404 = (inp[5]) ? node410 : node405;
										assign node405 = (inp[8]) ? node407 : 11'b01001100101;
											assign node407 = (inp[9]) ? 11'b01110000100 : 11'b01101000100;
										assign node410 = (inp[8]) ? node412 : 11'b01111000101;
											assign node412 = (inp[9]) ? 11'b01101000111 : 11'b01000100111;
									assign node415 = (inp[9]) ? node419 : node416;
										assign node416 = (inp[8]) ? 11'b01000000001 : 11'b01001100011;
										assign node419 = (inp[10]) ? 11'b01011110001 : 11'b01101010111;
								assign node422 = (inp[9]) ? node428 : node423;
									assign node423 = (inp[10]) ? node425 : 11'b01110000001;
										assign node425 = (inp[4]) ? 11'b01101110110 : 11'b01111100111;
									assign node428 = (inp[5]) ? node432 : node429;
										assign node429 = (inp[10]) ? 11'b01001111000 : 11'b01011101110;
										assign node432 = (inp[8]) ? 11'b01011010010 : 11'b01110011010;
							assign node435 = (inp[10]) ? node459 : node436;
								assign node436 = (inp[9]) ? node450 : node437;
									assign node437 = (inp[5]) ? node443 : node438;
										assign node438 = (inp[6]) ? 11'b01100110010 : node439;
											assign node439 = (inp[4]) ? 11'b01010110011 : 11'b01110110011;
										assign node443 = (inp[8]) ? node447 : node444;
											assign node444 = (inp[4]) ? 11'b01101110000 : 11'b01011010010;
											assign node447 = (inp[6]) ? 11'b01101110000 : 11'b01110110000;
									assign node450 = (inp[4]) ? node456 : node451;
										assign node451 = (inp[8]) ? node453 : 11'b01100110111;
											assign node453 = (inp[6]) ? 11'b01010010111 : 11'b01010110110;
										assign node456 = (inp[5]) ? 11'b01001000100 : 11'b01000100101;
								assign node459 = (inp[9]) ? node467 : node460;
									assign node460 = (inp[4]) ? node462 : 11'b01111010101;
										assign node462 = (inp[8]) ? node464 : 11'b01110000111;
											assign node464 = (inp[6]) ? 11'b01001000110 : 11'b01010000111;
									assign node467 = (inp[5]) ? 11'b01010000010 : 11'b01001100011;
						assign node470 = (inp[10]) ? node492 : node471;
							assign node471 = (inp[5]) ? node479 : node472;
								assign node472 = (inp[6]) ? 11'b01011111000 : node473;
									assign node473 = (inp[9]) ? node475 : 11'b01011110011;
										assign node475 = (inp[11]) ? 11'b01111110001 : 11'b01011110001;
								assign node479 = (inp[11]) ? node489 : node480;
									assign node480 = (inp[8]) ? node486 : node481;
										assign node481 = (inp[6]) ? node483 : 11'b01100110000;
											assign node483 = (inp[9]) ? 11'b01110011000 : 11'b01101011000;
										assign node486 = (inp[4]) ? 11'b01101010001 : 11'b01111100001;
									assign node489 = (inp[6]) ? 11'b01000010010 : 11'b01000010000;
							assign node492 = (inp[9]) ? node512 : node493;
								assign node493 = (inp[6]) ? node501 : node494;
									assign node494 = (inp[11]) ? node498 : node495;
										assign node495 = (inp[8]) ? 11'b01111100001 : 11'b01111100000;
										assign node498 = (inp[5]) ? 11'b01001000010 : 11'b01111000011;
									assign node501 = (inp[8]) ? node507 : node502;
										assign node502 = (inp[11]) ? 11'b01010000001 : node503;
											assign node503 = (inp[5]) ? 11'b01001001000 : 11'b01000001011;
										assign node507 = (inp[11]) ? node509 : 11'b01111000011;
											assign node509 = (inp[5]) ? 11'b01100100000 : 11'b01001100000;
								assign node512 = (inp[11]) ? node524 : node513;
									assign node513 = (inp[5]) ? node519 : node514;
										assign node514 = (inp[8]) ? node516 : 11'b01000100011;
											assign node516 = (inp[6]) ? 11'b01000000011 : 11'b01000000010;
										assign node519 = (inp[8]) ? 11'b01000100000 : node520;
											assign node520 = (inp[4]) ? 11'b01001000010 : 11'b01011001010;
									assign node524 = (inp[5]) ? node528 : node525;
										assign node525 = (inp[4]) ? 11'b01001101000 : 11'b01011000001;
										assign node528 = (inp[6]) ? node530 : 11'b01000000000;
											assign node530 = (inp[4]) ? 11'b01000000000 : 11'b01001000001;
			assign node533 = (inp[6]) ? node791 : node534;
				assign node534 = (inp[2]) ? node658 : node535;
					assign node535 = (inp[8]) ? node601 : node536;
						assign node536 = (inp[5]) ? node572 : node537;
							assign node537 = (inp[4]) ? node549 : node538;
								assign node538 = (inp[0]) ? node544 : node539;
									assign node539 = (inp[9]) ? node541 : 11'b01011000011;
										assign node541 = (inp[11]) ? 11'b11111100111 : 11'b11011100111;
									assign node544 = (inp[11]) ? 11'b01001000011 : node545;
										assign node545 = (inp[3]) ? 11'b01001100011 : 11'b01001110011;
								assign node549 = (inp[11]) ? node557 : node550;
									assign node550 = (inp[10]) ? 11'b11110000001 : node551;
										assign node551 = (inp[3]) ? 11'b01100000011 : node552;
											assign node552 = (inp[0]) ? 11'b01101010101 : 11'b01111000111;
									assign node557 = (inp[0]) ? node567 : node558;
										assign node558 = (inp[10]) ? node562 : node559;
											assign node559 = (inp[3]) ? 11'b11001110001 : 11'b01001110111;
											assign node562 = (inp[3]) ? node564 : 11'b11100110101;
												assign node564 = (inp[9]) ? 11'b01100110011 : 11'b01101110011;
										assign node567 = (inp[3]) ? 11'b01110110011 : node568;
											assign node568 = (inp[9]) ? 11'b01011100101 : 11'b01111100111;
							assign node572 = (inp[11]) ? node582 : node573;
								assign node573 = (inp[4]) ? 11'b11010110010 : node574;
									assign node574 = (inp[0]) ? node578 : node575;
										assign node575 = (inp[3]) ? 11'b01001000111 : 11'b11111000101;
										assign node578 = (inp[9]) ? 11'b01101010001 : 11'b01000000001;
								assign node582 = (inp[4]) ? node590 : node583;
									assign node583 = (inp[10]) ? node587 : node584;
										assign node584 = (inp[0]) ? 11'b01110110110 : 11'b01010110000;
										assign node587 = (inp[0]) ? 11'b01110100010 : 11'b11101000110;
									assign node590 = (inp[9]) ? node596 : node591;
										assign node591 = (inp[10]) ? 11'b11010000110 : node592;
											assign node592 = (inp[3]) ? 11'b11110010110 : 11'b01011010100;
										assign node596 = (inp[0]) ? node598 : 11'b11101000010;
											assign node598 = (inp[3]) ? 11'b01011000000 : 11'b01111000100;
						assign node601 = (inp[5]) ? node639 : node602;
							assign node602 = (inp[11]) ? node624 : node603;
								assign node603 = (inp[3]) ? node615 : node604;
									assign node604 = (inp[10]) ? 11'b01101100110 : node605;
										assign node605 = (inp[4]) ? node609 : node606;
											assign node606 = (inp[0]) ? 11'b01100000000 : 11'b01010000010;
											assign node609 = (inp[0]) ? 11'b01011010110 : node610;
												assign node610 = (inp[9]) ? 11'b01100100100 : 11'b01111100110;
									assign node615 = (inp[10]) ? node621 : node616;
										assign node616 = (inp[9]) ? 11'b01010110010 : node617;
											assign node617 = (inp[4]) ? 11'b01000110010 : 11'b01001100010;
										assign node621 = (inp[0]) ? 11'b01110100000 : 11'b01000100010;
								assign node624 = (inp[4]) ? node632 : node625;
									assign node625 = (inp[3]) ? node627 : 11'b11010010110;
										assign node627 = (inp[9]) ? node629 : 11'b01010000000;
											assign node629 = (inp[10]) ? 11'b01110010100 : 11'b01100010000;
									assign node632 = (inp[9]) ? 11'b10000111001 : node633;
										assign node633 = (inp[10]) ? node635 : 11'b00111111001;
											assign node635 = (inp[0]) ? 11'b00000101111 : 11'b00110111001;
							assign node639 = (inp[4]) ? node653 : node640;
								assign node640 = (inp[11]) ? node642 : 11'b00101011001;
									assign node642 = (inp[3]) ? node650 : node643;
										assign node643 = (inp[9]) ? node647 : node644;
											assign node644 = (inp[0]) ? 11'b00110111111 : 11'b00011111011;
											assign node647 = (inp[0]) ? 11'b00011101001 : 11'b10101101111;
										assign node650 = (inp[9]) ? 11'b00000101011 : 11'b10001101001;
								assign node653 = (inp[0]) ? node655 : 11'b10110001011;
									assign node655 = (inp[10]) ? 11'b00010001011 : 11'b00010001001;
					assign node658 = (inp[0]) ? node722 : node659;
						assign node659 = (inp[9]) ? node695 : node660;
							assign node660 = (inp[8]) ? node682 : node661;
								assign node661 = (inp[4]) ? node673 : node662;
									assign node662 = (inp[5]) ? node666 : node663;
										assign node663 = (inp[11]) ? 11'b00110101010 : 11'b10111001011;
										assign node666 = (inp[10]) ? node670 : node667;
											assign node667 = (inp[3]) ? 11'b10110111000 : 11'b00110111010;
											assign node670 = (inp[3]) ? 11'b00110001100 : 11'b10010011010;
									assign node673 = (inp[3]) ? 11'b10011011110 : node674;
										assign node674 = (inp[10]) ? node678 : node675;
											assign node675 = (inp[5]) ? 11'b00110111111 : 11'b00101001100;
											assign node678 = (inp[5]) ? 11'b10100101111 : 11'b10100111110;
								assign node682 = (inp[5]) ? node690 : node683;
									assign node683 = (inp[11]) ? 11'b00100111101 : node684;
										assign node684 = (inp[4]) ? 11'b00110001001 : node685;
											assign node685 = (inp[3]) ? 11'b10000101001 : 11'b00110101011;
									assign node690 = (inp[11]) ? node692 : 11'b00001011101;
										assign node692 = (inp[4]) ? 11'b10000011100 : 11'b10100101000;
							assign node695 = (inp[11]) ? node707 : node696;
								assign node696 = (inp[5]) ? node704 : node697;
									assign node697 = (inp[10]) ? 11'b10101101011 : node698;
										assign node698 = (inp[8]) ? node700 : 11'b00011101100;
											assign node700 = (inp[3]) ? 11'b10010001101 : 11'b00000001111;
									assign node704 = (inp[4]) ? 11'b00011101000 : 11'b00011101100;
								assign node707 = (inp[4]) ? node715 : node708;
									assign node708 = (inp[3]) ? node712 : node709;
										assign node709 = (inp[8]) ? 11'b00011111011 : 11'b00000001010;
										assign node712 = (inp[5]) ? 11'b10111111111 : 11'b00010111111;
									assign node715 = (inp[3]) ? node717 : 11'b00111011101;
										assign node717 = (inp[5]) ? node719 : 11'b00000011011;
											assign node719 = (inp[8]) ? 11'b00000001000 : 11'b00000101001;
						assign node722 = (inp[9]) ? node756 : node723;
							assign node723 = (inp[8]) ? node739 : node724;
								assign node724 = (inp[10]) ? node732 : node725;
									assign node725 = (inp[11]) ? node727 : 11'b00001001001;
										assign node727 = (inp[4]) ? node729 : 11'b00011011010;
											assign node729 = (inp[5]) ? 11'b00100111011 : 11'b00011011010;
									assign node732 = (inp[5]) ? node736 : node733;
										assign node733 = (inp[4]) ? 11'b00010001010 : 11'b00010001111;
										assign node736 = (inp[11]) ? 11'b00110001010 : 11'b00110101100;
								assign node739 = (inp[3]) ? node749 : node740;
									assign node740 = (inp[10]) ? node744 : node741;
										assign node741 = (inp[5]) ? 11'b00101001011 : 11'b00100101001;
										assign node744 = (inp[11]) ? 11'b00100111111 : node745;
											assign node745 = (inp[4]) ? 11'b00100011111 : 11'b00101001101;
									assign node749 = (inp[11]) ? node751 : 11'b00011011001;
										assign node751 = (inp[10]) ? node753 : 11'b00000101001;
											assign node753 = (inp[4]) ? 11'b00001001011 : 11'b00111101011;
							assign node756 = (inp[10]) ? node768 : node757;
								assign node757 = (inp[11]) ? node763 : node758;
									assign node758 = (inp[5]) ? node760 : 11'b00101101011;
										assign node760 = (inp[3]) ? 11'b00111111000 : 11'b00011101110;
									assign node763 = (inp[8]) ? 11'b00011011110 : node764;
										assign node764 = (inp[5]) ? 11'b00110011100 : 11'b00110011010;
								assign node768 = (inp[11]) ? node780 : node769;
									assign node769 = (inp[3]) ? node775 : node770;
										assign node770 = (inp[5]) ? 11'b00011111010 : node771;
											assign node771 = (inp[8]) ? 11'b00011111001 : 11'b00011111000;
										assign node775 = (inp[5]) ? 11'b00010101010 : node776;
											assign node776 = (inp[8]) ? 11'b00001001011 : 11'b00001101010;
									assign node780 = (inp[8]) ? node788 : node781;
										assign node781 = (inp[5]) ? node785 : node782;
											assign node782 = (inp[3]) ? 11'b00001101000 : 11'b00000001000;
											assign node785 = (inp[3]) ? 11'b00001101001 : 11'b00111101011;
										assign node788 = (inp[3]) ? 11'b00000001000 : 11'b00010001010;
				assign node791 = (inp[8]) ? node913 : node792;
					assign node792 = (inp[5]) ? node852 : node793;
						assign node793 = (inp[2]) ? node825 : node794;
							assign node794 = (inp[4]) ? node810 : node795;
								assign node795 = (inp[11]) ? node801 : node796;
									assign node796 = (inp[9]) ? 11'b00001101000 : node797;
										assign node797 = (inp[0]) ? 11'b00000101010 : 11'b00011101010;
									assign node801 = (inp[9]) ? node807 : node802;
										assign node802 = (inp[10]) ? node804 : 11'b00000001010;
											assign node804 = (inp[0]) ? 11'b00101001010 : 11'b00011011110;
										assign node807 = (inp[10]) ? 11'b00010001000 : 11'b00111011110;
								assign node810 = (inp[0]) ? node822 : node811;
									assign node811 = (inp[10]) ? node819 : node812;
										assign node812 = (inp[11]) ? node816 : node813;
											assign node813 = (inp[3]) ? 11'b10001101100 : 11'b00110101100;
											assign node816 = (inp[3]) ? 11'b10110001100 : 11'b00000001110;
										assign node819 = (inp[3]) ? 11'b00101011000 : 11'b10111001010;
									assign node822 = (inp[9]) ? 11'b00000100001 : 11'b00111110011;
							assign node825 = (inp[10]) ? node841 : node826;
								assign node826 = (inp[4]) ? node836 : node827;
									assign node827 = (inp[11]) ? node831 : node828;
										assign node828 = (inp[3]) ? 11'b10110000110 : 11'b00111000010;
										assign node831 = (inp[0]) ? 11'b00111010011 : node832;
											assign node832 = (inp[9]) ? 11'b10000100101 : 11'b10111110001;
									assign node836 = (inp[3]) ? 11'b10010110001 : node837;
										assign node837 = (inp[11]) ? 11'b00110010101 : 11'b00110110111;
								assign node841 = (inp[9]) ? node847 : node842;
									assign node842 = (inp[3]) ? 11'b00100100011 : node843;
										assign node843 = (inp[4]) ? 11'b00110000111 : 11'b00010110101;
									assign node847 = (inp[0]) ? 11'b00101110011 : node848;
										assign node848 = (inp[11]) ? 11'b00001010011 : 11'b00001110001;
						assign node852 = (inp[0]) ? node884 : node853;
							assign node853 = (inp[10]) ? node861 : node854;
								assign node854 = (inp[3]) ? node858 : node855;
									assign node855 = (inp[11]) ? 11'b00010110101 : 11'b00001010101;
									assign node858 = (inp[2]) ? 11'b10000110101 : 11'b10001110101;
								assign node861 = (inp[3]) ? node873 : node862;
									assign node862 = (inp[9]) ? node868 : node863;
										assign node863 = (inp[4]) ? node865 : 11'b10100010001;
											assign node865 = (inp[2]) ? 11'b10111000111 : 11'b10010000111;
										assign node868 = (inp[2]) ? node870 : 11'b10111100111;
											assign node870 = (inp[11]) ? 11'b10001000101 : 11'b10011100111;
									assign node873 = (inp[4]) ? node879 : node874;
										assign node874 = (inp[2]) ? 11'b00111100101 : node875;
											assign node875 = (inp[9]) ? 11'b00011000111 : 11'b00010000101;
										assign node879 = (inp[2]) ? 11'b00000100011 : node880;
											assign node880 = (inp[11]) ? 11'b00100100001 : 11'b00101000011;
							assign node884 = (inp[3]) ? node900 : node885;
								assign node885 = (inp[4]) ? node897 : node886;
									assign node886 = (inp[9]) ? node888 : 11'b00010010011;
										assign node888 = (inp[11]) ? node894 : node889;
											assign node889 = (inp[10]) ? node891 : 11'b00010100101;
												assign node891 = (inp[2]) ? 11'b00111110001 : 11'b00111010011;
											assign node894 = (inp[2]) ? 11'b00101010111 : 11'b00101110111;
									assign node897 = (inp[9]) ? 11'b00100100011 : 11'b00110110001;
								assign node900 = (inp[11]) ? node910 : node901;
									assign node901 = (inp[10]) ? 11'b00111100011 : node902;
										assign node902 = (inp[9]) ? 11'b00100110011 : node903;
											assign node903 = (inp[4]) ? 11'b00100110011 : node904;
												assign node904 = (inp[2]) ? 11'b00110000001 : 11'b00101100001;
									assign node910 = (inp[9]) ? 11'b00011100001 : 11'b00011000001;
					assign node913 = (inp[9]) ? node969 : node914;
						assign node914 = (inp[11]) ? node938 : node915;
							assign node915 = (inp[2]) ? node923 : node916;
								assign node916 = (inp[5]) ? node920 : node917;
									assign node917 = (inp[4]) ? 11'b00111000011 : 11'b00111000101;
									assign node920 = (inp[3]) ? 11'b00100000000 : 11'b00000000000;
								assign node923 = (inp[5]) ? node933 : node924;
									assign node924 = (inp[10]) ? node928 : node925;
										assign node925 = (inp[4]) ? 11'b00110100000 : 11'b10010000001;
										assign node928 = (inp[3]) ? 11'b00011100100 : node929;
											assign node929 = (inp[0]) ? 11'b00111100100 : 11'b10111100010;
									assign node933 = (inp[3]) ? 11'b10111110000 : node934;
										assign node934 = (inp[4]) ? 11'b00011110110 : 11'b00111110010;
							assign node938 = (inp[2]) ? node950 : node939;
								assign node939 = (inp[4]) ? node947 : node940;
									assign node940 = (inp[10]) ? 11'b00000110110 : node941;
										assign node941 = (inp[5]) ? node943 : 11'b10111110010;
											assign node943 = (inp[0]) ? 11'b00111100010 : 11'b10010100000;
									assign node947 = (inp[5]) ? 11'b00101000010 : 11'b00101100110;
								assign node950 = (inp[10]) ? node956 : node951;
									assign node951 = (inp[5]) ? node953 : 11'b00101010000;
										assign node953 = (inp[3]) ? 11'b00001010000 : 11'b00001010010;
									assign node956 = (inp[3]) ? node964 : node957;
										assign node957 = (inp[0]) ? node961 : node958;
											assign node958 = (inp[4]) ? 11'b10001010100 : 11'b10001000000;
											assign node961 = (inp[4]) ? 11'b00001000110 : 11'b00101010110;
										assign node964 = (inp[5]) ? 11'b00101000100 : node965;
											assign node965 = (inp[0]) ? 11'b00111000000 : 11'b00111010110;
						assign node969 = (inp[0]) ? node999 : node970;
							assign node970 = (inp[4]) ? node988 : node971;
								assign node971 = (inp[5]) ? node977 : node972;
									assign node972 = (inp[11]) ? node974 : 11'b00000110100;
										assign node974 = (inp[3]) ? 11'b00111110100 : 11'b10110010100;
									assign node977 = (inp[10]) ? node983 : node978;
										assign node978 = (inp[2]) ? node980 : 11'b00011010010;
											assign node980 = (inp[11]) ? 11'b00100000010 : 11'b00110110010;
										assign node983 = (inp[11]) ? 11'b00100100110 : node984;
											assign node984 = (inp[2]) ? 11'b10110100110 : 11'b10001000110;
								assign node988 = (inp[10]) ? node992 : node989;
									assign node989 = (inp[2]) ? 11'b00000000110 : 11'b00100000111;
									assign node992 = (inp[5]) ? node996 : node993;
										assign node993 = (inp[3]) ? 11'b00000010010 : 11'b10000010000;
										assign node996 = (inp[11]) ? 11'b00100000000 : 11'b00100100000;
							assign node999 = (inp[11]) ? node1017 : node1000;
								assign node1000 = (inp[2]) ? node1008 : node1001;
									assign node1001 = (inp[10]) ? node1003 : 11'b00101000101;
										assign node1003 = (inp[5]) ? node1005 : 11'b00010010001;
											assign node1005 = (inp[4]) ? 11'b00000100000 : 11'b00010000010;
									assign node1008 = (inp[4]) ? node1012 : node1009;
										assign node1009 = (inp[5]) ? 11'b00110110000 : 11'b00100110000;
										assign node1012 = (inp[3]) ? node1014 : 11'b00000110010;
											assign node1014 = (inp[5]) ? 11'b00000100000 : 11'b00000100010;
								assign node1017 = (inp[3]) ? node1023 : node1018;
									assign node1018 = (inp[5]) ? 11'b00000000010 : node1019;
										assign node1019 = (inp[4]) ? 11'b00000000010 : 11'b00110000010;
									assign node1023 = (inp[2]) ? node1027 : node1024;
										assign node1024 = (inp[5]) ? 11'b00010000000 : 11'b00111000000;
										assign node1027 = (inp[5]) ? 11'b00000010000 : node1028;
											assign node1028 = (inp[4]) ? 11'b00000000000 : 11'b00010000000;
		assign node1032 = (inp[7]) ? node1488 : node1033;
			assign node1033 = (inp[6]) ? node1265 : node1034;
				assign node1034 = (inp[8]) ? node1148 : node1035;
					assign node1035 = (inp[3]) ? node1093 : node1036;
						assign node1036 = (inp[11]) ? node1064 : node1037;
							assign node1037 = (inp[2]) ? node1045 : node1038;
								assign node1038 = (inp[0]) ? node1040 : 11'b00111111101;
									assign node1040 = (inp[5]) ? node1042 : 11'b00100111111;
										assign node1042 = (inp[4]) ? 11'b00100111001 : 11'b00100111011;
								assign node1045 = (inp[4]) ? node1057 : node1046;
									assign node1046 = (inp[5]) ? node1052 : node1047;
										assign node1047 = (inp[10]) ? 11'b10110011100 : node1048;
											assign node1048 = (inp[0]) ? 11'b00001001010 : 11'b00101001000;
										assign node1052 = (inp[10]) ? node1054 : 11'b00101011001;
											assign node1054 = (inp[0]) ? 11'b00101011001 : 11'b10001001111;
									assign node1057 = (inp[5]) ? node1059 : 11'b10111111101;
										assign node1059 = (inp[10]) ? 11'b00111111011 : node1060;
											assign node1060 = (inp[0]) ? 11'b00111001001 : 11'b00111011111;
							assign node1064 = (inp[2]) ? node1076 : node1065;
								assign node1065 = (inp[10]) ? node1071 : node1066;
									assign node1066 = (inp[0]) ? node1068 : 11'b00011001111;
										assign node1068 = (inp[9]) ? 11'b00111001101 : 11'b00011011011;
									assign node1071 = (inp[5]) ? node1073 : 11'b10111011111;
										assign node1073 = (inp[9]) ? 11'b10010001011 : 11'b10001001111;
								assign node1076 = (inp[10]) ? node1080 : node1077;
									assign node1077 = (inp[0]) ? 11'b00010111011 : 11'b00010101011;
									assign node1080 = (inp[0]) ? node1090 : node1081;
										assign node1081 = (inp[9]) ? node1087 : node1082;
											assign node1082 = (inp[4]) ? 11'b10111101101 : node1083;
												assign node1083 = (inp[5]) ? 11'b10001111011 : 11'b10111101011;
											assign node1087 = (inp[4]) ? 11'b10011011011 : 11'b10001111101;
										assign node1090 = (inp[5]) ? 11'b00001111101 : 11'b00100101101;
						assign node1093 = (inp[9]) ? node1111 : node1094;
							assign node1094 = (inp[2]) ? node1106 : node1095;
								assign node1095 = (inp[0]) ? node1101 : node1096;
									assign node1096 = (inp[4]) ? 11'b00101001001 : node1097;
										assign node1097 = (inp[11]) ? 11'b00011001111 : 11'b00101111111;
									assign node1101 = (inp[5]) ? 11'b00111101001 : node1102;
										assign node1102 = (inp[4]) ? 11'b00101101001 : 11'b00001101001;
								assign node1106 = (inp[5]) ? node1108 : 11'b00011001000;
									assign node1108 = (inp[4]) ? 11'b00110011001 : 11'b00110001001;
							assign node1111 = (inp[5]) ? node1131 : node1112;
								assign node1112 = (inp[11]) ? node1122 : node1113;
									assign node1113 = (inp[2]) ? 11'b10100001110 : node1114;
										assign node1114 = (inp[4]) ? node1116 : 11'b00000111101;
											assign node1116 = (inp[0]) ? 11'b00100101001 : node1117;
												assign node1117 = (inp[10]) ? 11'b00100111001 : 11'b10100111001;
									assign node1122 = (inp[10]) ? node1124 : 11'b00100011001;
										assign node1124 = (inp[0]) ? node1128 : node1125;
											assign node1125 = (inp[2]) ? 11'b00011011001 : 11'b00010011101;
											assign node1128 = (inp[2]) ? 11'b00010101011 : 11'b00010001001;
								assign node1131 = (inp[0]) ? node1139 : node1132;
									assign node1132 = (inp[11]) ? node1136 : node1133;
										assign node1133 = (inp[2]) ? 11'b00001101011 : 11'b00100101011;
										assign node1136 = (inp[10]) ? 11'b00010101001 : 11'b10001101001;
									assign node1139 = (inp[10]) ? node1145 : node1140;
										assign node1140 = (inp[2]) ? node1142 : 11'b00010011011;
											assign node1142 = (inp[11]) ? 11'b00000101011 : 11'b00010001001;
										assign node1145 = (inp[2]) ? 11'b00000101001 : 11'b00010101001;
					assign node1148 = (inp[0]) ? node1196 : node1149;
						assign node1149 = (inp[10]) ? node1173 : node1150;
							assign node1150 = (inp[3]) ? node1162 : node1151;
								assign node1151 = (inp[11]) ? node1157 : node1152;
									assign node1152 = (inp[9]) ? 11'b00010011000 : node1153;
										assign node1153 = (inp[2]) ? 11'b00100111000 : 11'b00111111100;
									assign node1157 = (inp[2]) ? node1159 : 11'b00000101000;
										assign node1159 = (inp[9]) ? 11'b00100001000 : 11'b00101001001;
								assign node1162 = (inp[9]) ? node1166 : node1163;
									assign node1163 = (inp[4]) ? 11'b10100111110 : 11'b10111111010;
									assign node1166 = (inp[4]) ? node1170 : node1167;
										assign node1167 = (inp[2]) ? 11'b10001001111 : 11'b10111101100;
										assign node1170 = (inp[11]) ? 11'b10100001000 : 11'b10001001000;
							assign node1173 = (inp[3]) ? node1189 : node1174;
								assign node1174 = (inp[5]) ? node1186 : node1175;
									assign node1175 = (inp[11]) ? node1179 : node1176;
										assign node1176 = (inp[9]) ? 11'b10101011101 : 11'b10100111100;
										assign node1179 = (inp[2]) ? node1181 : 11'b10111011010;
											assign node1181 = (inp[9]) ? node1183 : 11'b10011111100;
												assign node1183 = (inp[4]) ? 11'b10000111010 : 11'b10111111110;
									assign node1186 = (inp[11]) ? 11'b10001001100 : 11'b10001101100;
								assign node1189 = (inp[11]) ? node1193 : node1190;
									assign node1190 = (inp[2]) ? 11'b00001011011 : 11'b00100111010;
									assign node1193 = (inp[9]) ? 11'b00111001110 : 11'b00110011101;
						assign node1196 = (inp[3]) ? node1220 : node1197;
							assign node1197 = (inp[5]) ? node1209 : node1198;
								assign node1198 = (inp[4]) ? node1204 : node1199;
									assign node1199 = (inp[11]) ? 11'b00111011001 : node1200;
										assign node1200 = (inp[10]) ? 11'b00111011001 : 11'b00111001111;
									assign node1204 = (inp[11]) ? 11'b00011101100 : node1205;
										assign node1205 = (inp[10]) ? 11'b00100011111 : 11'b00001011111;
								assign node1209 = (inp[10]) ? node1217 : node1210;
									assign node1210 = (inp[4]) ? node1214 : node1211;
										assign node1211 = (inp[9]) ? 11'b00010011100 : 11'b00110011010;
										assign node1214 = (inp[2]) ? 11'b00011011100 : 11'b00001011000;
									assign node1217 = (inp[2]) ? 11'b00000111010 : 11'b00011001010;
							assign node1220 = (inp[10]) ? node1244 : node1221;
								assign node1221 = (inp[2]) ? node1227 : node1222;
									assign node1222 = (inp[5]) ? node1224 : 11'b00110011010;
										assign node1224 = (inp[11]) ? 11'b00111101000 : 11'b00100001000;
									assign node1227 = (inp[4]) ? node1235 : node1228;
										assign node1228 = (inp[5]) ? node1232 : node1229;
											assign node1229 = (inp[9]) ? 11'b00001011011 : 11'b00000001011;
											assign node1232 = (inp[11]) ? 11'b00001011010 : 11'b00110111010;
										assign node1235 = (inp[9]) ? node1239 : node1236;
											assign node1236 = (inp[5]) ? 11'b00001011000 : 11'b00101111010;
											assign node1239 = (inp[5]) ? 11'b00000001010 : node1240;
												assign node1240 = (inp[11]) ? 11'b00100101000 : 11'b00101001001;
								assign node1244 = (inp[9]) ? node1256 : node1245;
									assign node1245 = (inp[5]) ? node1253 : node1246;
										assign node1246 = (inp[2]) ? node1250 : node1247;
											assign node1247 = (inp[4]) ? 11'b00111101000 : 11'b00011101000;
											assign node1250 = (inp[4]) ? 11'b00110001001 : 11'b00011001001;
										assign node1253 = (inp[11]) ? 11'b00100101000 : 11'b00100101010;
									assign node1256 = (inp[4]) ? node1258 : 11'b00011101010;
										assign node1258 = (inp[5]) ? 11'b00001001000 : node1259;
											assign node1259 = (inp[11]) ? node1261 : 11'b00000101010;
												assign node1261 = (inp[2]) ? 11'b00000101000 : 11'b00001001000;
				assign node1265 = (inp[2]) ? node1365 : node1266;
					assign node1266 = (inp[8]) ? node1322 : node1267;
						assign node1267 = (inp[11]) ? node1295 : node1268;
							assign node1268 = (inp[5]) ? node1282 : node1269;
								assign node1269 = (inp[4]) ? node1275 : node1270;
									assign node1270 = (inp[9]) ? 11'b00000101000 : node1271;
										assign node1271 = (inp[10]) ? 11'b00011101110 : 11'b10011101000;
									assign node1275 = (inp[9]) ? node1277 : 11'b00000111000;
										assign node1277 = (inp[3]) ? node1279 : 11'b10101101010;
											assign node1279 = (inp[10]) ? 11'b00111111000 : 11'b00101101010;
								assign node1282 = (inp[0]) ? node1284 : 11'b00000001110;
									assign node1284 = (inp[4]) ? 11'b00100001000 : node1285;
										assign node1285 = (inp[10]) ? node1291 : node1286;
											assign node1286 = (inp[9]) ? 11'b00011001100 : node1287;
												assign node1287 = (inp[3]) ? 11'b00101001010 : 11'b00011001010;
											assign node1291 = (inp[3]) ? 11'b00010001000 : 11'b00110011010;
							assign node1295 = (inp[5]) ? node1309 : node1296;
								assign node1296 = (inp[0]) ? node1302 : node1297;
									assign node1297 = (inp[10]) ? 11'b10111011110 : node1298;
										assign node1298 = (inp[9]) ? 11'b00110111000 : 11'b10000111010;
									assign node1302 = (inp[10]) ? node1304 : 11'b00110001010;
										assign node1304 = (inp[3]) ? 11'b00100101010 : node1305;
											assign node1305 = (inp[4]) ? 11'b00100001010 : 11'b00001001010;
								assign node1309 = (inp[0]) ? node1317 : node1310;
									assign node1310 = (inp[3]) ? node1312 : 11'b00001110111;
										assign node1312 = (inp[10]) ? 11'b00000100101 : node1313;
											assign node1313 = (inp[9]) ? 11'b10100100011 : 11'b10101100001;
									assign node1317 = (inp[10]) ? node1319 : 11'b00111110001;
										assign node1319 = (inp[4]) ? 11'b00011100001 : 11'b00110100001;
						assign node1322 = (inp[0]) ? node1344 : node1323;
							assign node1323 = (inp[11]) ? node1339 : node1324;
								assign node1324 = (inp[5]) ? node1332 : node1325;
									assign node1325 = (inp[4]) ? node1327 : 11'b10001010111;
										assign node1327 = (inp[9]) ? 11'b10010010001 : node1328;
											assign node1328 = (inp[10]) ? 11'b10110010101 : 11'b10000000111;
									assign node1332 = (inp[9]) ? node1336 : node1333;
										assign node1333 = (inp[10]) ? 11'b10001100111 : 11'b00111110101;
										assign node1336 = (inp[10]) ? 11'b10100110011 : 11'b00000110011;
								assign node1339 = (inp[5]) ? node1341 : 11'b00011000001;
									assign node1341 = (inp[3]) ? 11'b10101010101 : 11'b10111000111;
							assign node1344 = (inp[10]) ? node1358 : node1345;
								assign node1345 = (inp[5]) ? node1355 : node1346;
									assign node1346 = (inp[11]) ? node1348 : 11'b00011010011;
										assign node1348 = (inp[9]) ? node1352 : node1349;
											assign node1349 = (inp[3]) ? 11'b00110010001 : 11'b00100010011;
											assign node1352 = (inp[4]) ? 11'b00111100011 : 11'b00100010011;
									assign node1355 = (inp[4]) ? 11'b00111110011 : 11'b00100110001;
								assign node1358 = (inp[9]) ? node1362 : node1359;
									assign node1359 = (inp[5]) ? 11'b00111110111 : 11'b00011000011;
									assign node1362 = (inp[3]) ? 11'b00001000011 : 11'b00000000001;
					assign node1365 = (inp[5]) ? node1433 : node1366;
						assign node1366 = (inp[0]) ? node1394 : node1367;
							assign node1367 = (inp[8]) ? node1383 : node1368;
								assign node1368 = (inp[11]) ? node1374 : node1369;
									assign node1369 = (inp[10]) ? 11'b00111000111 : node1370;
										assign node1370 = (inp[9]) ? 11'b10101000101 : 11'b10101000011;
									assign node1374 = (inp[4]) ? node1378 : node1375;
										assign node1375 = (inp[9]) ? 11'b00100110110 : 11'b00110110110;
										assign node1378 = (inp[10]) ? node1380 : 11'b00101110100;
											assign node1380 = (inp[3]) ? 11'b00001110010 : 11'b10011110010;
								assign node1383 = (inp[4]) ? node1387 : node1384;
									assign node1384 = (inp[10]) ? 11'b10100000000 : 11'b00110100000;
									assign node1387 = (inp[3]) ? node1389 : 11'b10110100010;
										assign node1389 = (inp[10]) ? 11'b00010110010 : node1390;
											assign node1390 = (inp[11]) ? 11'b10110110010 : 11'b10110110000;
							assign node1394 = (inp[4]) ? node1412 : node1395;
								assign node1395 = (inp[10]) ? node1399 : node1396;
									assign node1396 = (inp[8]) ? 11'b00001110000 : 11'b00001110010;
									assign node1399 = (inp[8]) ? node1405 : node1400;
										assign node1400 = (inp[3]) ? 11'b00100100010 : node1401;
											assign node1401 = (inp[11]) ? 11'b00011110100 : 11'b00001000101;
										assign node1405 = (inp[3]) ? node1407 : 11'b00111100010;
											assign node1407 = (inp[11]) ? 11'b00011100000 : node1408;
												assign node1408 = (inp[9]) ? 11'b00001100010 : 11'b00011100010;
								assign node1412 = (inp[11]) ? node1422 : node1413;
									assign node1413 = (inp[10]) ? node1419 : node1414;
										assign node1414 = (inp[8]) ? node1416 : 11'b00010000001;
											assign node1416 = (inp[3]) ? 11'b00011110000 : 11'b00111100000;
										assign node1419 = (inp[3]) ? 11'b00110100010 : 11'b00110110110;
									assign node1422 = (inp[9]) ? node1428 : node1423;
										assign node1423 = (inp[8]) ? 11'b00100110010 : node1424;
											assign node1424 = (inp[3]) ? 11'b00100110000 : 11'b00000110000;
										assign node1428 = (inp[10]) ? node1430 : 11'b00011100100;
											assign node1430 = (inp[3]) ? 11'b00000100000 : 11'b00000100010;
						assign node1433 = (inp[0]) ? node1463 : node1434;
							assign node1434 = (inp[4]) ? node1446 : node1435;
								assign node1435 = (inp[9]) ? node1439 : node1436;
									assign node1436 = (inp[8]) ? 11'b10101010010 : 11'b10000010010;
									assign node1439 = (inp[10]) ? node1441 : 11'b00111000010;
										assign node1441 = (inp[11]) ? 11'b10011000100 : node1442;
											assign node1442 = (inp[3]) ? 11'b00001000100 : 11'b10101000110;
								assign node1446 = (inp[8]) ? node1452 : node1447;
									assign node1447 = (inp[10]) ? 11'b00010000010 : node1448;
										assign node1448 = (inp[11]) ? 11'b00101010100 : 11'b10101000000;
									assign node1452 = (inp[10]) ? node1458 : node1453;
										assign node1453 = (inp[3]) ? 11'b10010000010 : node1454;
											assign node1454 = (inp[11]) ? 11'b00010000110 : 11'b00010010110;
										assign node1458 = (inp[11]) ? node1460 : 11'b00010000000;
											assign node1460 = (inp[9]) ? 11'b10010000000 : 11'b10010000100;
							assign node1463 = (inp[8]) ? node1477 : node1464;
								assign node1464 = (inp[10]) ? node1472 : node1465;
									assign node1465 = (inp[4]) ? 11'b00111010100 : node1466;
										assign node1466 = (inp[3]) ? node1468 : 11'b00000100110;
											assign node1468 = (inp[9]) ? 11'b00110110000 : 11'b00110100010;
									assign node1472 = (inp[3]) ? node1474 : 11'b00100100100;
										assign node1474 = (inp[9]) ? 11'b00000000000 : 11'b00000100000;
								assign node1477 = (inp[10]) ? 11'b00000000100 : node1478;
									assign node1478 = (inp[4]) ? node1484 : node1479;
										assign node1479 = (inp[9]) ? node1481 : 11'b00101000010;
											assign node1481 = (inp[3]) ? 11'b00001010010 : 11'b00001010110;
										assign node1484 = (inp[11]) ? 11'b00000010010 : 11'b00000000010;
			assign node1488 = (inp[6]) ? node1762 : node1489;
				assign node1489 = (inp[2]) ? node1613 : node1490;
					assign node1490 = (inp[5]) ? node1552 : node1491;
						assign node1491 = (inp[0]) ? node1509 : node1492;
							assign node1492 = (inp[4]) ? node1504 : node1493;
								assign node1493 = (inp[8]) ? node1497 : node1494;
									assign node1494 = (inp[10]) ? 11'b00011100101 : 11'b00011100011;
									assign node1497 = (inp[11]) ? node1499 : 11'b00110000101;
										assign node1499 = (inp[10]) ? 11'b10010110101 : node1500;
											assign node1500 = (inp[3]) ? 11'b10110110001 : 11'b00010100001;
								assign node1504 = (inp[9]) ? node1506 : 11'b10100100111;
									assign node1506 = (inp[3]) ? 11'b10001110001 : 11'b00000110101;
							assign node1509 = (inp[10]) ? node1529 : node1510;
								assign node1510 = (inp[8]) ? node1522 : node1511;
									assign node1511 = (inp[4]) ? node1517 : node1512;
										assign node1512 = (inp[3]) ? node1514 : 11'b00101110111;
											assign node1514 = (inp[11]) ? 11'b00101110011 : 11'b00001110011;
										assign node1517 = (inp[11]) ? 11'b00110100011 : node1518;
											assign node1518 = (inp[9]) ? 11'b00100100011 : 11'b00000100011;
									assign node1522 = (inp[11]) ? node1526 : node1523;
										assign node1523 = (inp[9]) ? 11'b00111100111 : 11'b00101100001;
										assign node1526 = (inp[4]) ? 11'b00111110001 : 11'b00100110001;
								assign node1529 = (inp[3]) ? node1537 : node1530;
									assign node1530 = (inp[8]) ? node1534 : node1531;
										assign node1531 = (inp[4]) ? 11'b00000110101 : 11'b00001100101;
										assign node1534 = (inp[9]) ? 11'b00111110001 : 11'b00101110111;
									assign node1537 = (inp[8]) ? node1545 : node1538;
										assign node1538 = (inp[4]) ? node1542 : node1539;
											assign node1539 = (inp[11]) ? 11'b00101100001 : 11'b00001100001;
											assign node1542 = (inp[9]) ? 11'b00000100001 : 11'b00010100001;
										assign node1545 = (inp[4]) ? node1549 : node1546;
											assign node1546 = (inp[11]) ? 11'b00110100011 : 11'b00010000001;
											assign node1549 = (inp[9]) ? 11'b00000100011 : 11'b00001100001;
						assign node1552 = (inp[0]) ? node1584 : node1553;
							assign node1553 = (inp[10]) ? node1561 : node1554;
								assign node1554 = (inp[9]) ? 11'b00000110001 : node1555;
									assign node1555 = (inp[3]) ? 11'b10111010101 : node1556;
										assign node1556 = (inp[4]) ? 11'b00011010111 : 11'b00011010011;
								assign node1561 = (inp[3]) ? node1573 : node1562;
									assign node1562 = (inp[8]) ? node1566 : node1563;
										assign node1563 = (inp[11]) ? 11'b10011000101 : 11'b10000000111;
										assign node1566 = (inp[11]) ? node1568 : 11'b10101010001;
											assign node1568 = (inp[4]) ? 11'b10100000101 : node1569;
												assign node1569 = (inp[9]) ? 11'b10100000111 : 11'b10001010011;
									assign node1573 = (inp[4]) ? node1577 : node1574;
										assign node1574 = (inp[9]) ? 11'b00100000111 : 11'b00001000111;
										assign node1577 = (inp[8]) ? 11'b00111000001 : node1578;
											assign node1578 = (inp[9]) ? 11'b00110000011 : node1579;
												assign node1579 = (inp[11]) ? 11'b00110000011 : 11'b00000010011;
							assign node1584 = (inp[4]) ? node1596 : node1585;
								assign node1585 = (inp[8]) ? node1593 : node1586;
									assign node1586 = (inp[3]) ? node1590 : node1587;
										assign node1587 = (inp[10]) ? 11'b00011010111 : 11'b00111010101;
										assign node1590 = (inp[10]) ? 11'b00111000011 : 11'b00101010011;
									assign node1593 = (inp[10]) ? 11'b00000000011 : 11'b00100110001;
								assign node1596 = (inp[8]) ? node1600 : node1597;
									assign node1597 = (inp[9]) ? 11'b00000000001 : 11'b00101010011;
									assign node1600 = (inp[11]) ? node1606 : node1601;
										assign node1601 = (inp[10]) ? 11'b00001010001 : node1602;
											assign node1602 = (inp[9]) ? 11'b00011000001 : 11'b00010100001;
										assign node1606 = (inp[9]) ? node1608 : 11'b00010010001;
											assign node1608 = (inp[10]) ? 11'b00010000001 : node1609;
												assign node1609 = (inp[3]) ? 11'b00010000001 : 11'b00000000111;
					assign node1613 = (inp[8]) ? node1709 : node1614;
						assign node1614 = (inp[5]) ? node1666 : node1615;
							assign node1615 = (inp[11]) ? node1639 : node1616;
								assign node1616 = (inp[4]) ? node1628 : node1617;
									assign node1617 = (inp[0]) ? node1625 : node1618;
										assign node1618 = (inp[10]) ? 11'b10101000011 : node1619;
											assign node1619 = (inp[3]) ? node1621 : 11'b00111000001;
												assign node1621 = (inp[9]) ? 11'b10111000111 : 11'b10111000011;
										assign node1625 = (inp[9]) ? 11'b00001000011 : 11'b00001000001;
									assign node1628 = (inp[3]) ? node1636 : node1629;
										assign node1629 = (inp[10]) ? node1631 : 11'b00010000111;
											assign node1631 = (inp[0]) ? node1633 : 11'b10101010101;
												assign node1633 = (inp[9]) ? 11'b00110010001 : 11'b00010010111;
										assign node1636 = (inp[0]) ? 11'b00100000011 : 11'b00010000011;
								assign node1639 = (inp[4]) ? node1657 : node1640;
									assign node1640 = (inp[9]) ? node1648 : node1641;
										assign node1641 = (inp[0]) ? node1643 : 11'b10100010011;
											assign node1643 = (inp[3]) ? node1645 : 11'b00000010111;
												assign node1645 = (inp[10]) ? 11'b00100000001 : 11'b00010000011;
										assign node1648 = (inp[0]) ? node1652 : node1649;
											assign node1649 = (inp[10]) ? 11'b10011110110 : 11'b00000010001;
											assign node1652 = (inp[10]) ? node1654 : 11'b00111110010;
												assign node1654 = (inp[3]) ? 11'b00011100010 : 11'b00001100010;
									assign node1657 = (inp[9]) ? node1663 : node1658;
										assign node1658 = (inp[3]) ? node1660 : 11'b10011110100;
											assign node1660 = (inp[10]) ? 11'b00001110000 : 11'b00101110000;
										assign node1663 = (inp[3]) ? 11'b10111110010 : 11'b10001110010;
							assign node1666 = (inp[0]) ? node1692 : node1667;
								assign node1667 = (inp[11]) ? node1681 : node1668;
									assign node1668 = (inp[3]) ? node1676 : node1669;
										assign node1669 = (inp[10]) ? node1673 : node1670;
											assign node1670 = (inp[9]) ? 11'b00110110000 : 11'b00100110110;
											assign node1673 = (inp[9]) ? 11'b10010100100 : 11'b10110100100;
										assign node1676 = (inp[10]) ? node1678 : 11'b10010110110;
											assign node1678 = (inp[4]) ? 11'b00100110000 : 11'b00010110110;
									assign node1681 = (inp[3]) ? node1685 : node1682;
										assign node1682 = (inp[4]) ? 11'b00111110100 : 11'b10011110000;
										assign node1685 = (inp[4]) ? node1687 : 11'b00101100100;
											assign node1687 = (inp[10]) ? 11'b00010100010 : node1688;
												assign node1688 = (inp[9]) ? 11'b10010100000 : 11'b10001110100;
								assign node1692 = (inp[11]) ? node1700 : node1693;
									assign node1693 = (inp[3]) ? node1697 : node1694;
										assign node1694 = (inp[9]) ? 11'b00010100100 : 11'b00001100000;
										assign node1697 = (inp[9]) ? 11'b00001100010 : 11'b00110100000;
									assign node1700 = (inp[4]) ? 11'b00101110000 : node1701;
										assign node1701 = (inp[10]) ? 11'b00111100000 : node1702;
											assign node1702 = (inp[9]) ? 11'b00001110010 : node1703;
												assign node1703 = (inp[3]) ? 11'b00111100000 : 11'b00011110000;
						assign node1709 = (inp[3]) ? node1737 : node1710;
							assign node1710 = (inp[4]) ? node1724 : node1711;
								assign node1711 = (inp[0]) ? node1717 : node1712;
									assign node1712 = (inp[9]) ? 11'b00101010010 : node1713;
										assign node1713 = (inp[11]) ? 11'b00110010010 : 11'b00110010000;
									assign node1717 = (inp[5]) ? node1721 : node1718;
										assign node1718 = (inp[9]) ? 11'b00100000010 : 11'b00101010100;
										assign node1721 = (inp[10]) ? 11'b00010000000 : 11'b00010010100;
								assign node1724 = (inp[11]) ? node1732 : node1725;
									assign node1725 = (inp[0]) ? 11'b00111010110 : node1726;
										assign node1726 = (inp[10]) ? 11'b10011010100 : node1727;
											assign node1727 = (inp[9]) ? 11'b00001000100 : 11'b00001010100;
									assign node1732 = (inp[0]) ? 11'b00010000000 : node1733;
										assign node1733 = (inp[10]) ? 11'b10000010100 : 11'b00000000100;
							assign node1737 = (inp[9]) ? node1747 : node1738;
								assign node1738 = (inp[4]) ? node1744 : node1739;
									assign node1739 = (inp[11]) ? 11'b00001000000 : node1740;
										assign node1740 = (inp[0]) ? 11'b00010100010 : 11'b10000100010;
									assign node1744 = (inp[0]) ? 11'b00101000010 : 11'b00000000010;
								assign node1747 = (inp[10]) ? node1753 : node1748;
									assign node1748 = (inp[0]) ? 11'b00110010010 : node1749;
										assign node1749 = (inp[4]) ? 11'b10000000000 : 11'b10000010100;
									assign node1753 = (inp[11]) ? node1757 : node1754;
										assign node1754 = (inp[0]) ? 11'b00001000000 : 11'b00011000000;
										assign node1757 = (inp[4]) ? 11'b00000000000 : node1758;
											assign node1758 = (inp[0]) ? 11'b00000000000 : 11'b00000000100;
				assign node1762 = (inp[2]) ? node1880 : node1763;
					assign node1763 = (inp[8]) ? node1819 : node1764;
						assign node1764 = (inp[3]) ? node1790 : node1765;
							assign node1765 = (inp[9]) ? node1779 : node1766;
								assign node1766 = (inp[10]) ? node1774 : node1767;
									assign node1767 = (inp[0]) ? node1769 : 11'b00001100000;
										assign node1769 = (inp[11]) ? 11'b00010110010 : node1770;
											assign node1770 = (inp[5]) ? 11'b00010100000 : 11'b00011100010;
									assign node1774 = (inp[4]) ? node1776 : 11'b10011100010;
										assign node1776 = (inp[0]) ? 11'b00011110110 : 11'b10011110110;
								assign node1779 = (inp[10]) ? 11'b00011110000 : node1780;
									assign node1780 = (inp[11]) ? node1786 : node1781;
										assign node1781 = (inp[0]) ? 11'b00011100110 : node1782;
											assign node1782 = (inp[5]) ? 11'b00111110110 : 11'b00111100100;
										assign node1786 = (inp[0]) ? 11'b00101110100 : 11'b00010110110;
							assign node1790 = (inp[11]) ? node1800 : node1791;
								assign node1791 = (inp[4]) ? 11'b00101100010 : node1792;
									assign node1792 = (inp[0]) ? node1796 : node1793;
										assign node1793 = (inp[5]) ? 11'b10000110000 : 11'b00001110100;
										assign node1796 = (inp[9]) ? 11'b00001100000 : 11'b00001100010;
								assign node1800 = (inp[0]) ? node1808 : node1801;
									assign node1801 = (inp[9]) ? 11'b10000110010 : node1802;
										assign node1802 = (inp[4]) ? 11'b10110100110 : node1803;
											assign node1803 = (inp[10]) ? 11'b00010110110 : 11'b10010110010;
									assign node1808 = (inp[4]) ? node1816 : node1809;
										assign node1809 = (inp[9]) ? 11'b00000100010 : node1810;
											assign node1810 = (inp[5]) ? 11'b00101100000 : node1811;
												assign node1811 = (inp[10]) ? 11'b00100100010 : 11'b00000100010;
										assign node1816 = (inp[9]) ? 11'b00110100000 : 11'b00110110010;
						assign node1819 = (inp[0]) ? node1851 : node1820;
							assign node1820 = (inp[9]) ? node1832 : node1821;
								assign node1821 = (inp[3]) ? node1825 : node1822;
									assign node1822 = (inp[10]) ? 11'b10100110100 : 11'b00110100100;
									assign node1825 = (inp[4]) ? 11'b00011000010 : node1826;
										assign node1826 = (inp[5]) ? 11'b10011010000 : node1827;
											assign node1827 = (inp[11]) ? 11'b10111010000 : 11'b10100100010;
								assign node1832 = (inp[5]) ? node1840 : node1833;
									assign node1833 = (inp[4]) ? node1837 : node1834;
										assign node1834 = (inp[3]) ? 11'b10110100100 : 11'b10001010100;
										assign node1837 = (inp[10]) ? 11'b00101010010 : 11'b00101000110;
									assign node1840 = (inp[4]) ? node1844 : node1841;
										assign node1841 = (inp[10]) ? 11'b00100000110 : 11'b00000000010;
										assign node1844 = (inp[10]) ? node1846 : 11'b00100010100;
											assign node1846 = (inp[11]) ? node1848 : 11'b10110010000;
												assign node1848 = (inp[3]) ? 11'b00100000000 : 11'b10100000000;
							assign node1851 = (inp[5]) ? node1871 : node1852;
								assign node1852 = (inp[11]) ? node1860 : node1853;
									assign node1853 = (inp[4]) ? node1855 : 11'b00100110000;
										assign node1855 = (inp[10]) ? node1857 : 11'b00000110000;
											assign node1857 = (inp[3]) ? 11'b00001000010 : 11'b00011010010;
									assign node1860 = (inp[10]) ? node1868 : node1861;
										assign node1861 = (inp[3]) ? node1863 : 11'b00101010010;
											assign node1863 = (inp[9]) ? node1865 : 11'b00011000000;
												assign node1865 = (inp[4]) ? 11'b00111000000 : 11'b00101010000;
										assign node1868 = (inp[3]) ? 11'b00011000010 : 11'b00111000010;
								assign node1871 = (inp[4]) ? node1873 : 11'b00010010010;
									assign node1873 = (inp[9]) ? node1875 : 11'b00010010000;
										assign node1875 = (inp[10]) ? node1877 : 11'b00000010100;
											assign node1877 = (inp[3]) ? 11'b00000000000 : 11'b00010010000;
					assign node1880 = (inp[8]) ? node1938 : node1881;
						assign node1881 = (inp[5]) ? node1913 : node1882;
							assign node1882 = (inp[4]) ? node1900 : node1883;
								assign node1883 = (inp[9]) ? node1891 : node1884;
									assign node1884 = (inp[10]) ? node1886 : 11'b00101000000;
										assign node1886 = (inp[0]) ? node1888 : 11'b10111000010;
											assign node1888 = (inp[3]) ? 11'b00101000010 : 11'b00011010110;
									assign node1891 = (inp[11]) ? node1897 : node1892;
										assign node1892 = (inp[10]) ? 11'b00001010010 : node1893;
											assign node1893 = (inp[3]) ? 11'b00011010010 : 11'b00011000110;
										assign node1897 = (inp[3]) ? 11'b10001000110 : 11'b10011010110;
								assign node1900 = (inp[10]) ? node1908 : node1901;
									assign node1901 = (inp[0]) ? node1905 : node1902;
										assign node1902 = (inp[3]) ? 11'b10111000100 : 11'b00111010100;
										assign node1905 = (inp[9]) ? 11'b00111000000 : 11'b00011010000;
									assign node1908 = (inp[9]) ? node1910 : 11'b00011000000;
										assign node1910 = (inp[0]) ? 11'b00001000000 : 11'b00001010000;
							assign node1913 = (inp[11]) ? node1925 : node1914;
								assign node1914 = (inp[4]) ? 11'b00110000010 : node1915;
									assign node1915 = (inp[10]) ? node1921 : node1916;
										assign node1916 = (inp[0]) ? 11'b00011000000 : node1917;
											assign node1917 = (inp[3]) ? 11'b10111010000 : 11'b00101010000;
										assign node1921 = (inp[3]) ? 11'b00001010100 : 11'b00101000100;
								assign node1925 = (inp[3]) ? node1931 : node1926;
									assign node1926 = (inp[0]) ? 11'b00100010100 : node1927;
										assign node1927 = (inp[4]) ? 11'b00110010100 : 11'b00010000000;
									assign node1931 = (inp[4]) ? 11'b00010000000 : node1932;
										assign node1932 = (inp[0]) ? node1934 : 11'b10000000010;
											assign node1934 = (inp[10]) ? 11'b00000000000 : 11'b00000010000;
						assign node1938 = (inp[5]) ? node1974 : node1939;
							assign node1939 = (inp[11]) ? node1959 : node1940;
								assign node1940 = (inp[10]) ? node1950 : node1941;
									assign node1941 = (inp[4]) ? node1945 : node1942;
										assign node1942 = (inp[0]) ? 11'b00010000010 : 11'b00100000010;
										assign node1945 = (inp[0]) ? node1947 : 11'b00010000110;
											assign node1947 = (inp[3]) ? 11'b00010010010 : 11'b00010010110;
									assign node1950 = (inp[9]) ? node1956 : node1951;
										assign node1951 = (inp[3]) ? 11'b00110000010 : node1952;
											assign node1952 = (inp[4]) ? 11'b00110010110 : 11'b00110000110;
										assign node1956 = (inp[3]) ? 11'b00000010110 : 11'b00100010010;
								assign node1959 = (inp[10]) ? node1967 : node1960;
									assign node1960 = (inp[9]) ? 11'b00110010000 : node1961;
										assign node1961 = (inp[3]) ? 11'b00000000010 : node1962;
											assign node1962 = (inp[0]) ? 11'b00100010010 : 11'b00100000010;
									assign node1967 = (inp[4]) ? node1971 : node1968;
										assign node1968 = (inp[9]) ? 11'b10110010100 : 11'b00110010100;
										assign node1971 = (inp[3]) ? 11'b00000000000 : 11'b00000000100;
							assign node1974 = (inp[4]) ? node1988 : node1975;
								assign node1975 = (inp[10]) ? node1981 : node1976;
									assign node1976 = (inp[11]) ? 11'b00100010000 : node1977;
										assign node1977 = (inp[3]) ? 11'b00110010000 : 11'b00110000100;
									assign node1981 = (inp[11]) ? 11'b00000000100 : node1982;
										assign node1982 = (inp[9]) ? node1984 : 11'b00010010100;
											assign node1984 = (inp[3]) ? 11'b00010000000 : 11'b00010010000;
								assign node1988 = (inp[9]) ? node1992 : node1989;
									assign node1989 = (inp[11]) ? 11'b10000000100 : 11'b00010010100;
									assign node1992 = (inp[10]) ? 11'b00000000000 : 11'b10000000000;

endmodule