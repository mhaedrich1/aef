module dtc_split66_bm26 (
	input  wire [15-1:0] inp,
	output wire [15-1:0] outp
);

	wire [15-1:0] node1;
	wire [15-1:0] node2;
	wire [15-1:0] node3;
	wire [15-1:0] node4;
	wire [15-1:0] node5;
	wire [15-1:0] node6;
	wire [15-1:0] node7;
	wire [15-1:0] node8;
	wire [15-1:0] node9;
	wire [15-1:0] node10;
	wire [15-1:0] node13;
	wire [15-1:0] node16;
	wire [15-1:0] node17;
	wire [15-1:0] node20;
	wire [15-1:0] node23;
	wire [15-1:0] node24;
	wire [15-1:0] node25;
	wire [15-1:0] node28;
	wire [15-1:0] node31;
	wire [15-1:0] node32;
	wire [15-1:0] node35;
	wire [15-1:0] node38;
	wire [15-1:0] node39;
	wire [15-1:0] node40;
	wire [15-1:0] node41;
	wire [15-1:0] node44;
	wire [15-1:0] node47;
	wire [15-1:0] node48;
	wire [15-1:0] node51;
	wire [15-1:0] node54;
	wire [15-1:0] node55;
	wire [15-1:0] node56;
	wire [15-1:0] node59;
	wire [15-1:0] node62;
	wire [15-1:0] node63;
	wire [15-1:0] node66;
	wire [15-1:0] node69;
	wire [15-1:0] node70;
	wire [15-1:0] node71;
	wire [15-1:0] node72;
	wire [15-1:0] node73;
	wire [15-1:0] node76;
	wire [15-1:0] node79;
	wire [15-1:0] node80;
	wire [15-1:0] node83;
	wire [15-1:0] node86;
	wire [15-1:0] node87;
	wire [15-1:0] node88;
	wire [15-1:0] node91;
	wire [15-1:0] node94;
	wire [15-1:0] node95;
	wire [15-1:0] node98;
	wire [15-1:0] node101;
	wire [15-1:0] node102;
	wire [15-1:0] node103;
	wire [15-1:0] node104;
	wire [15-1:0] node107;
	wire [15-1:0] node110;
	wire [15-1:0] node111;
	wire [15-1:0] node114;
	wire [15-1:0] node117;
	wire [15-1:0] node118;
	wire [15-1:0] node119;
	wire [15-1:0] node122;
	wire [15-1:0] node125;
	wire [15-1:0] node126;
	wire [15-1:0] node129;
	wire [15-1:0] node132;
	wire [15-1:0] node133;
	wire [15-1:0] node134;
	wire [15-1:0] node135;
	wire [15-1:0] node136;
	wire [15-1:0] node137;
	wire [15-1:0] node140;
	wire [15-1:0] node143;
	wire [15-1:0] node144;
	wire [15-1:0] node147;
	wire [15-1:0] node150;
	wire [15-1:0] node151;
	wire [15-1:0] node152;
	wire [15-1:0] node155;
	wire [15-1:0] node158;
	wire [15-1:0] node159;
	wire [15-1:0] node162;
	wire [15-1:0] node165;
	wire [15-1:0] node166;
	wire [15-1:0] node167;
	wire [15-1:0] node168;
	wire [15-1:0] node171;
	wire [15-1:0] node174;
	wire [15-1:0] node175;
	wire [15-1:0] node178;
	wire [15-1:0] node181;
	wire [15-1:0] node182;
	wire [15-1:0] node183;
	wire [15-1:0] node186;
	wire [15-1:0] node189;
	wire [15-1:0] node190;
	wire [15-1:0] node193;
	wire [15-1:0] node196;
	wire [15-1:0] node197;
	wire [15-1:0] node198;
	wire [15-1:0] node199;
	wire [15-1:0] node200;
	wire [15-1:0] node203;
	wire [15-1:0] node206;
	wire [15-1:0] node207;
	wire [15-1:0] node210;
	wire [15-1:0] node213;
	wire [15-1:0] node214;
	wire [15-1:0] node215;
	wire [15-1:0] node218;
	wire [15-1:0] node221;
	wire [15-1:0] node222;
	wire [15-1:0] node225;
	wire [15-1:0] node228;
	wire [15-1:0] node229;
	wire [15-1:0] node230;
	wire [15-1:0] node231;
	wire [15-1:0] node234;
	wire [15-1:0] node237;
	wire [15-1:0] node238;
	wire [15-1:0] node241;
	wire [15-1:0] node244;
	wire [15-1:0] node245;
	wire [15-1:0] node246;
	wire [15-1:0] node249;
	wire [15-1:0] node252;
	wire [15-1:0] node253;
	wire [15-1:0] node256;
	wire [15-1:0] node259;
	wire [15-1:0] node260;
	wire [15-1:0] node261;
	wire [15-1:0] node262;
	wire [15-1:0] node263;
	wire [15-1:0] node264;
	wire [15-1:0] node265;
	wire [15-1:0] node268;
	wire [15-1:0] node271;
	wire [15-1:0] node272;
	wire [15-1:0] node275;
	wire [15-1:0] node278;
	wire [15-1:0] node279;
	wire [15-1:0] node280;
	wire [15-1:0] node283;
	wire [15-1:0] node286;
	wire [15-1:0] node287;
	wire [15-1:0] node290;
	wire [15-1:0] node293;
	wire [15-1:0] node294;
	wire [15-1:0] node295;
	wire [15-1:0] node296;
	wire [15-1:0] node299;
	wire [15-1:0] node302;
	wire [15-1:0] node303;
	wire [15-1:0] node306;
	wire [15-1:0] node309;
	wire [15-1:0] node310;
	wire [15-1:0] node311;
	wire [15-1:0] node314;
	wire [15-1:0] node317;
	wire [15-1:0] node318;
	wire [15-1:0] node321;
	wire [15-1:0] node324;
	wire [15-1:0] node325;
	wire [15-1:0] node326;
	wire [15-1:0] node327;
	wire [15-1:0] node328;
	wire [15-1:0] node331;
	wire [15-1:0] node334;
	wire [15-1:0] node335;
	wire [15-1:0] node338;
	wire [15-1:0] node341;
	wire [15-1:0] node342;
	wire [15-1:0] node343;
	wire [15-1:0] node346;
	wire [15-1:0] node349;
	wire [15-1:0] node350;
	wire [15-1:0] node353;
	wire [15-1:0] node356;
	wire [15-1:0] node357;
	wire [15-1:0] node358;
	wire [15-1:0] node359;
	wire [15-1:0] node362;
	wire [15-1:0] node365;
	wire [15-1:0] node366;
	wire [15-1:0] node369;
	wire [15-1:0] node372;
	wire [15-1:0] node373;
	wire [15-1:0] node374;
	wire [15-1:0] node377;
	wire [15-1:0] node380;
	wire [15-1:0] node381;
	wire [15-1:0] node384;
	wire [15-1:0] node387;
	wire [15-1:0] node388;
	wire [15-1:0] node389;
	wire [15-1:0] node390;
	wire [15-1:0] node391;
	wire [15-1:0] node392;
	wire [15-1:0] node395;
	wire [15-1:0] node398;
	wire [15-1:0] node399;
	wire [15-1:0] node402;
	wire [15-1:0] node405;
	wire [15-1:0] node406;
	wire [15-1:0] node407;
	wire [15-1:0] node410;
	wire [15-1:0] node413;
	wire [15-1:0] node414;
	wire [15-1:0] node417;
	wire [15-1:0] node420;
	wire [15-1:0] node421;
	wire [15-1:0] node422;
	wire [15-1:0] node423;
	wire [15-1:0] node426;
	wire [15-1:0] node429;
	wire [15-1:0] node430;
	wire [15-1:0] node433;
	wire [15-1:0] node436;
	wire [15-1:0] node437;
	wire [15-1:0] node438;
	wire [15-1:0] node441;
	wire [15-1:0] node444;
	wire [15-1:0] node445;
	wire [15-1:0] node448;
	wire [15-1:0] node451;
	wire [15-1:0] node452;
	wire [15-1:0] node453;
	wire [15-1:0] node454;
	wire [15-1:0] node455;
	wire [15-1:0] node458;
	wire [15-1:0] node461;
	wire [15-1:0] node462;
	wire [15-1:0] node465;
	wire [15-1:0] node468;
	wire [15-1:0] node469;
	wire [15-1:0] node470;
	wire [15-1:0] node473;
	wire [15-1:0] node476;
	wire [15-1:0] node477;
	wire [15-1:0] node480;
	wire [15-1:0] node483;
	wire [15-1:0] node484;
	wire [15-1:0] node485;
	wire [15-1:0] node486;
	wire [15-1:0] node489;
	wire [15-1:0] node492;
	wire [15-1:0] node493;
	wire [15-1:0] node496;
	wire [15-1:0] node499;
	wire [15-1:0] node500;
	wire [15-1:0] node501;
	wire [15-1:0] node504;
	wire [15-1:0] node507;
	wire [15-1:0] node508;
	wire [15-1:0] node511;
	wire [15-1:0] node514;
	wire [15-1:0] node515;
	wire [15-1:0] node516;
	wire [15-1:0] node517;
	wire [15-1:0] node518;
	wire [15-1:0] node519;
	wire [15-1:0] node520;
	wire [15-1:0] node521;
	wire [15-1:0] node524;
	wire [15-1:0] node527;
	wire [15-1:0] node528;
	wire [15-1:0] node531;
	wire [15-1:0] node534;
	wire [15-1:0] node535;
	wire [15-1:0] node536;
	wire [15-1:0] node539;
	wire [15-1:0] node542;
	wire [15-1:0] node543;
	wire [15-1:0] node546;
	wire [15-1:0] node549;
	wire [15-1:0] node550;
	wire [15-1:0] node551;
	wire [15-1:0] node552;
	wire [15-1:0] node555;
	wire [15-1:0] node558;
	wire [15-1:0] node559;
	wire [15-1:0] node562;
	wire [15-1:0] node565;
	wire [15-1:0] node566;
	wire [15-1:0] node567;
	wire [15-1:0] node570;
	wire [15-1:0] node573;
	wire [15-1:0] node574;
	wire [15-1:0] node577;
	wire [15-1:0] node580;
	wire [15-1:0] node581;
	wire [15-1:0] node582;
	wire [15-1:0] node583;
	wire [15-1:0] node584;
	wire [15-1:0] node587;
	wire [15-1:0] node590;
	wire [15-1:0] node591;
	wire [15-1:0] node594;
	wire [15-1:0] node597;
	wire [15-1:0] node598;
	wire [15-1:0] node599;
	wire [15-1:0] node602;
	wire [15-1:0] node605;
	wire [15-1:0] node606;
	wire [15-1:0] node609;
	wire [15-1:0] node612;
	wire [15-1:0] node613;
	wire [15-1:0] node614;
	wire [15-1:0] node615;
	wire [15-1:0] node618;
	wire [15-1:0] node621;
	wire [15-1:0] node622;
	wire [15-1:0] node625;
	wire [15-1:0] node628;
	wire [15-1:0] node629;
	wire [15-1:0] node630;
	wire [15-1:0] node633;
	wire [15-1:0] node636;
	wire [15-1:0] node637;
	wire [15-1:0] node640;
	wire [15-1:0] node643;
	wire [15-1:0] node644;
	wire [15-1:0] node645;
	wire [15-1:0] node646;
	wire [15-1:0] node647;
	wire [15-1:0] node648;
	wire [15-1:0] node651;
	wire [15-1:0] node654;
	wire [15-1:0] node655;
	wire [15-1:0] node658;
	wire [15-1:0] node661;
	wire [15-1:0] node662;
	wire [15-1:0] node663;
	wire [15-1:0] node666;
	wire [15-1:0] node669;
	wire [15-1:0] node670;
	wire [15-1:0] node673;
	wire [15-1:0] node676;
	wire [15-1:0] node677;
	wire [15-1:0] node678;
	wire [15-1:0] node679;
	wire [15-1:0] node682;
	wire [15-1:0] node685;
	wire [15-1:0] node686;
	wire [15-1:0] node689;
	wire [15-1:0] node692;
	wire [15-1:0] node693;
	wire [15-1:0] node694;
	wire [15-1:0] node697;
	wire [15-1:0] node700;
	wire [15-1:0] node701;
	wire [15-1:0] node704;
	wire [15-1:0] node707;
	wire [15-1:0] node708;
	wire [15-1:0] node709;
	wire [15-1:0] node710;
	wire [15-1:0] node711;
	wire [15-1:0] node714;
	wire [15-1:0] node717;
	wire [15-1:0] node718;
	wire [15-1:0] node721;
	wire [15-1:0] node724;
	wire [15-1:0] node725;
	wire [15-1:0] node726;
	wire [15-1:0] node729;
	wire [15-1:0] node732;
	wire [15-1:0] node733;
	wire [15-1:0] node736;
	wire [15-1:0] node739;
	wire [15-1:0] node740;
	wire [15-1:0] node741;
	wire [15-1:0] node742;
	wire [15-1:0] node745;
	wire [15-1:0] node748;
	wire [15-1:0] node749;
	wire [15-1:0] node752;
	wire [15-1:0] node755;
	wire [15-1:0] node756;
	wire [15-1:0] node757;
	wire [15-1:0] node760;
	wire [15-1:0] node763;
	wire [15-1:0] node764;
	wire [15-1:0] node767;
	wire [15-1:0] node770;
	wire [15-1:0] node771;
	wire [15-1:0] node772;
	wire [15-1:0] node773;
	wire [15-1:0] node774;
	wire [15-1:0] node775;
	wire [15-1:0] node776;
	wire [15-1:0] node779;
	wire [15-1:0] node782;
	wire [15-1:0] node783;
	wire [15-1:0] node786;
	wire [15-1:0] node789;
	wire [15-1:0] node790;
	wire [15-1:0] node791;
	wire [15-1:0] node794;
	wire [15-1:0] node797;
	wire [15-1:0] node798;
	wire [15-1:0] node801;
	wire [15-1:0] node804;
	wire [15-1:0] node805;
	wire [15-1:0] node806;
	wire [15-1:0] node807;
	wire [15-1:0] node810;
	wire [15-1:0] node813;
	wire [15-1:0] node814;
	wire [15-1:0] node817;
	wire [15-1:0] node820;
	wire [15-1:0] node821;
	wire [15-1:0] node822;
	wire [15-1:0] node825;
	wire [15-1:0] node828;
	wire [15-1:0] node829;
	wire [15-1:0] node832;
	wire [15-1:0] node835;
	wire [15-1:0] node836;
	wire [15-1:0] node837;
	wire [15-1:0] node838;
	wire [15-1:0] node839;
	wire [15-1:0] node842;
	wire [15-1:0] node845;
	wire [15-1:0] node846;
	wire [15-1:0] node849;
	wire [15-1:0] node852;
	wire [15-1:0] node853;
	wire [15-1:0] node854;
	wire [15-1:0] node857;
	wire [15-1:0] node860;
	wire [15-1:0] node861;
	wire [15-1:0] node864;
	wire [15-1:0] node867;
	wire [15-1:0] node868;
	wire [15-1:0] node869;
	wire [15-1:0] node870;
	wire [15-1:0] node873;
	wire [15-1:0] node876;
	wire [15-1:0] node877;
	wire [15-1:0] node880;
	wire [15-1:0] node883;
	wire [15-1:0] node884;
	wire [15-1:0] node885;
	wire [15-1:0] node888;
	wire [15-1:0] node891;
	wire [15-1:0] node892;
	wire [15-1:0] node895;
	wire [15-1:0] node898;
	wire [15-1:0] node899;
	wire [15-1:0] node900;
	wire [15-1:0] node901;
	wire [15-1:0] node902;
	wire [15-1:0] node903;
	wire [15-1:0] node906;
	wire [15-1:0] node909;
	wire [15-1:0] node910;
	wire [15-1:0] node913;
	wire [15-1:0] node916;
	wire [15-1:0] node917;
	wire [15-1:0] node918;
	wire [15-1:0] node921;
	wire [15-1:0] node924;
	wire [15-1:0] node925;
	wire [15-1:0] node928;
	wire [15-1:0] node931;
	wire [15-1:0] node932;
	wire [15-1:0] node933;
	wire [15-1:0] node934;
	wire [15-1:0] node937;
	wire [15-1:0] node940;
	wire [15-1:0] node941;
	wire [15-1:0] node944;
	wire [15-1:0] node947;
	wire [15-1:0] node948;
	wire [15-1:0] node949;
	wire [15-1:0] node952;
	wire [15-1:0] node955;
	wire [15-1:0] node956;
	wire [15-1:0] node959;
	wire [15-1:0] node962;
	wire [15-1:0] node963;
	wire [15-1:0] node964;
	wire [15-1:0] node965;
	wire [15-1:0] node966;
	wire [15-1:0] node969;
	wire [15-1:0] node972;
	wire [15-1:0] node973;
	wire [15-1:0] node976;
	wire [15-1:0] node979;
	wire [15-1:0] node980;
	wire [15-1:0] node981;
	wire [15-1:0] node984;
	wire [15-1:0] node987;
	wire [15-1:0] node988;
	wire [15-1:0] node991;
	wire [15-1:0] node994;
	wire [15-1:0] node995;
	wire [15-1:0] node996;
	wire [15-1:0] node997;
	wire [15-1:0] node1000;
	wire [15-1:0] node1003;
	wire [15-1:0] node1004;
	wire [15-1:0] node1007;
	wire [15-1:0] node1010;
	wire [15-1:0] node1011;
	wire [15-1:0] node1012;
	wire [15-1:0] node1015;
	wire [15-1:0] node1018;
	wire [15-1:0] node1019;
	wire [15-1:0] node1022;
	wire [15-1:0] node1025;
	wire [15-1:0] node1026;
	wire [15-1:0] node1027;
	wire [15-1:0] node1028;
	wire [15-1:0] node1029;
	wire [15-1:0] node1030;
	wire [15-1:0] node1031;
	wire [15-1:0] node1032;
	wire [15-1:0] node1033;
	wire [15-1:0] node1036;
	wire [15-1:0] node1039;
	wire [15-1:0] node1040;
	wire [15-1:0] node1043;
	wire [15-1:0] node1046;
	wire [15-1:0] node1047;
	wire [15-1:0] node1048;
	wire [15-1:0] node1051;
	wire [15-1:0] node1054;
	wire [15-1:0] node1055;
	wire [15-1:0] node1058;
	wire [15-1:0] node1061;
	wire [15-1:0] node1062;
	wire [15-1:0] node1063;
	wire [15-1:0] node1064;
	wire [15-1:0] node1067;
	wire [15-1:0] node1070;
	wire [15-1:0] node1071;
	wire [15-1:0] node1074;
	wire [15-1:0] node1077;
	wire [15-1:0] node1078;
	wire [15-1:0] node1079;
	wire [15-1:0] node1082;
	wire [15-1:0] node1085;
	wire [15-1:0] node1086;
	wire [15-1:0] node1089;
	wire [15-1:0] node1092;
	wire [15-1:0] node1093;
	wire [15-1:0] node1094;
	wire [15-1:0] node1095;
	wire [15-1:0] node1096;
	wire [15-1:0] node1099;
	wire [15-1:0] node1102;
	wire [15-1:0] node1103;
	wire [15-1:0] node1106;
	wire [15-1:0] node1109;
	wire [15-1:0] node1110;
	wire [15-1:0] node1111;
	wire [15-1:0] node1114;
	wire [15-1:0] node1117;
	wire [15-1:0] node1118;
	wire [15-1:0] node1121;
	wire [15-1:0] node1124;
	wire [15-1:0] node1125;
	wire [15-1:0] node1126;
	wire [15-1:0] node1127;
	wire [15-1:0] node1130;
	wire [15-1:0] node1133;
	wire [15-1:0] node1134;
	wire [15-1:0] node1137;
	wire [15-1:0] node1140;
	wire [15-1:0] node1141;
	wire [15-1:0] node1142;
	wire [15-1:0] node1145;
	wire [15-1:0] node1148;
	wire [15-1:0] node1149;
	wire [15-1:0] node1152;
	wire [15-1:0] node1155;
	wire [15-1:0] node1156;
	wire [15-1:0] node1157;
	wire [15-1:0] node1158;
	wire [15-1:0] node1159;
	wire [15-1:0] node1160;
	wire [15-1:0] node1163;
	wire [15-1:0] node1166;
	wire [15-1:0] node1167;
	wire [15-1:0] node1170;
	wire [15-1:0] node1173;
	wire [15-1:0] node1174;
	wire [15-1:0] node1175;
	wire [15-1:0] node1178;
	wire [15-1:0] node1181;
	wire [15-1:0] node1182;
	wire [15-1:0] node1185;
	wire [15-1:0] node1188;
	wire [15-1:0] node1189;
	wire [15-1:0] node1190;
	wire [15-1:0] node1191;
	wire [15-1:0] node1194;
	wire [15-1:0] node1197;
	wire [15-1:0] node1198;
	wire [15-1:0] node1201;
	wire [15-1:0] node1204;
	wire [15-1:0] node1205;
	wire [15-1:0] node1206;
	wire [15-1:0] node1209;
	wire [15-1:0] node1212;
	wire [15-1:0] node1213;
	wire [15-1:0] node1216;
	wire [15-1:0] node1219;
	wire [15-1:0] node1220;
	wire [15-1:0] node1221;
	wire [15-1:0] node1222;
	wire [15-1:0] node1223;
	wire [15-1:0] node1226;
	wire [15-1:0] node1229;
	wire [15-1:0] node1230;
	wire [15-1:0] node1233;
	wire [15-1:0] node1236;
	wire [15-1:0] node1237;
	wire [15-1:0] node1238;
	wire [15-1:0] node1241;
	wire [15-1:0] node1244;
	wire [15-1:0] node1245;
	wire [15-1:0] node1248;
	wire [15-1:0] node1251;
	wire [15-1:0] node1252;
	wire [15-1:0] node1253;
	wire [15-1:0] node1254;
	wire [15-1:0] node1257;
	wire [15-1:0] node1260;
	wire [15-1:0] node1261;
	wire [15-1:0] node1264;
	wire [15-1:0] node1267;
	wire [15-1:0] node1268;
	wire [15-1:0] node1269;
	wire [15-1:0] node1272;
	wire [15-1:0] node1275;
	wire [15-1:0] node1276;
	wire [15-1:0] node1279;
	wire [15-1:0] node1282;
	wire [15-1:0] node1283;
	wire [15-1:0] node1284;
	wire [15-1:0] node1285;
	wire [15-1:0] node1286;
	wire [15-1:0] node1287;
	wire [15-1:0] node1288;
	wire [15-1:0] node1291;
	wire [15-1:0] node1294;
	wire [15-1:0] node1295;
	wire [15-1:0] node1298;
	wire [15-1:0] node1301;
	wire [15-1:0] node1302;
	wire [15-1:0] node1303;
	wire [15-1:0] node1306;
	wire [15-1:0] node1309;
	wire [15-1:0] node1310;
	wire [15-1:0] node1313;
	wire [15-1:0] node1316;
	wire [15-1:0] node1317;
	wire [15-1:0] node1318;
	wire [15-1:0] node1319;
	wire [15-1:0] node1322;
	wire [15-1:0] node1325;
	wire [15-1:0] node1326;
	wire [15-1:0] node1329;
	wire [15-1:0] node1332;
	wire [15-1:0] node1333;
	wire [15-1:0] node1334;
	wire [15-1:0] node1337;
	wire [15-1:0] node1340;
	wire [15-1:0] node1341;
	wire [15-1:0] node1344;
	wire [15-1:0] node1347;
	wire [15-1:0] node1348;
	wire [15-1:0] node1349;
	wire [15-1:0] node1350;
	wire [15-1:0] node1351;
	wire [15-1:0] node1354;
	wire [15-1:0] node1357;
	wire [15-1:0] node1358;
	wire [15-1:0] node1361;
	wire [15-1:0] node1364;
	wire [15-1:0] node1365;
	wire [15-1:0] node1366;
	wire [15-1:0] node1369;
	wire [15-1:0] node1372;
	wire [15-1:0] node1373;
	wire [15-1:0] node1376;
	wire [15-1:0] node1379;
	wire [15-1:0] node1380;
	wire [15-1:0] node1381;
	wire [15-1:0] node1382;
	wire [15-1:0] node1385;
	wire [15-1:0] node1388;
	wire [15-1:0] node1389;
	wire [15-1:0] node1392;
	wire [15-1:0] node1395;
	wire [15-1:0] node1396;
	wire [15-1:0] node1397;
	wire [15-1:0] node1400;
	wire [15-1:0] node1403;
	wire [15-1:0] node1404;
	wire [15-1:0] node1407;
	wire [15-1:0] node1410;
	wire [15-1:0] node1411;
	wire [15-1:0] node1412;
	wire [15-1:0] node1413;
	wire [15-1:0] node1414;
	wire [15-1:0] node1415;
	wire [15-1:0] node1418;
	wire [15-1:0] node1421;
	wire [15-1:0] node1422;
	wire [15-1:0] node1425;
	wire [15-1:0] node1428;
	wire [15-1:0] node1429;
	wire [15-1:0] node1430;
	wire [15-1:0] node1433;
	wire [15-1:0] node1436;
	wire [15-1:0] node1437;
	wire [15-1:0] node1440;
	wire [15-1:0] node1443;
	wire [15-1:0] node1444;
	wire [15-1:0] node1445;
	wire [15-1:0] node1446;
	wire [15-1:0] node1449;
	wire [15-1:0] node1452;
	wire [15-1:0] node1453;
	wire [15-1:0] node1456;
	wire [15-1:0] node1459;
	wire [15-1:0] node1460;
	wire [15-1:0] node1461;
	wire [15-1:0] node1464;
	wire [15-1:0] node1467;
	wire [15-1:0] node1468;
	wire [15-1:0] node1471;
	wire [15-1:0] node1474;
	wire [15-1:0] node1475;
	wire [15-1:0] node1476;
	wire [15-1:0] node1477;
	wire [15-1:0] node1478;
	wire [15-1:0] node1481;
	wire [15-1:0] node1484;
	wire [15-1:0] node1485;
	wire [15-1:0] node1488;
	wire [15-1:0] node1491;
	wire [15-1:0] node1492;
	wire [15-1:0] node1493;
	wire [15-1:0] node1496;
	wire [15-1:0] node1499;
	wire [15-1:0] node1500;
	wire [15-1:0] node1503;
	wire [15-1:0] node1506;
	wire [15-1:0] node1507;
	wire [15-1:0] node1508;
	wire [15-1:0] node1509;
	wire [15-1:0] node1512;
	wire [15-1:0] node1515;
	wire [15-1:0] node1516;
	wire [15-1:0] node1519;
	wire [15-1:0] node1522;
	wire [15-1:0] node1523;
	wire [15-1:0] node1524;
	wire [15-1:0] node1527;
	wire [15-1:0] node1530;
	wire [15-1:0] node1531;
	wire [15-1:0] node1534;
	wire [15-1:0] node1537;
	wire [15-1:0] node1538;
	wire [15-1:0] node1539;
	wire [15-1:0] node1540;
	wire [15-1:0] node1541;
	wire [15-1:0] node1542;
	wire [15-1:0] node1543;
	wire [15-1:0] node1544;
	wire [15-1:0] node1547;
	wire [15-1:0] node1550;
	wire [15-1:0] node1551;
	wire [15-1:0] node1554;
	wire [15-1:0] node1557;
	wire [15-1:0] node1558;
	wire [15-1:0] node1559;
	wire [15-1:0] node1562;
	wire [15-1:0] node1565;
	wire [15-1:0] node1566;
	wire [15-1:0] node1569;
	wire [15-1:0] node1572;
	wire [15-1:0] node1573;
	wire [15-1:0] node1574;
	wire [15-1:0] node1575;
	wire [15-1:0] node1578;
	wire [15-1:0] node1581;
	wire [15-1:0] node1582;
	wire [15-1:0] node1585;
	wire [15-1:0] node1588;
	wire [15-1:0] node1589;
	wire [15-1:0] node1590;
	wire [15-1:0] node1593;
	wire [15-1:0] node1596;
	wire [15-1:0] node1597;
	wire [15-1:0] node1600;
	wire [15-1:0] node1603;
	wire [15-1:0] node1604;
	wire [15-1:0] node1605;
	wire [15-1:0] node1606;
	wire [15-1:0] node1607;
	wire [15-1:0] node1610;
	wire [15-1:0] node1613;
	wire [15-1:0] node1614;
	wire [15-1:0] node1617;
	wire [15-1:0] node1620;
	wire [15-1:0] node1621;
	wire [15-1:0] node1622;
	wire [15-1:0] node1625;
	wire [15-1:0] node1628;
	wire [15-1:0] node1629;
	wire [15-1:0] node1632;
	wire [15-1:0] node1635;
	wire [15-1:0] node1636;
	wire [15-1:0] node1637;
	wire [15-1:0] node1638;
	wire [15-1:0] node1641;
	wire [15-1:0] node1644;
	wire [15-1:0] node1645;
	wire [15-1:0] node1648;
	wire [15-1:0] node1651;
	wire [15-1:0] node1652;
	wire [15-1:0] node1653;
	wire [15-1:0] node1656;
	wire [15-1:0] node1659;
	wire [15-1:0] node1660;
	wire [15-1:0] node1663;
	wire [15-1:0] node1666;
	wire [15-1:0] node1667;
	wire [15-1:0] node1668;
	wire [15-1:0] node1669;
	wire [15-1:0] node1670;
	wire [15-1:0] node1671;
	wire [15-1:0] node1674;
	wire [15-1:0] node1677;
	wire [15-1:0] node1678;
	wire [15-1:0] node1681;
	wire [15-1:0] node1684;
	wire [15-1:0] node1685;
	wire [15-1:0] node1686;
	wire [15-1:0] node1689;
	wire [15-1:0] node1692;
	wire [15-1:0] node1693;
	wire [15-1:0] node1696;
	wire [15-1:0] node1699;
	wire [15-1:0] node1700;
	wire [15-1:0] node1701;
	wire [15-1:0] node1702;
	wire [15-1:0] node1705;
	wire [15-1:0] node1708;
	wire [15-1:0] node1709;
	wire [15-1:0] node1712;
	wire [15-1:0] node1715;
	wire [15-1:0] node1716;
	wire [15-1:0] node1717;
	wire [15-1:0] node1720;
	wire [15-1:0] node1723;
	wire [15-1:0] node1724;
	wire [15-1:0] node1727;
	wire [15-1:0] node1730;
	wire [15-1:0] node1731;
	wire [15-1:0] node1732;
	wire [15-1:0] node1733;
	wire [15-1:0] node1734;
	wire [15-1:0] node1737;
	wire [15-1:0] node1740;
	wire [15-1:0] node1741;
	wire [15-1:0] node1744;
	wire [15-1:0] node1747;
	wire [15-1:0] node1748;
	wire [15-1:0] node1749;
	wire [15-1:0] node1752;
	wire [15-1:0] node1755;
	wire [15-1:0] node1756;
	wire [15-1:0] node1759;
	wire [15-1:0] node1762;
	wire [15-1:0] node1763;
	wire [15-1:0] node1764;
	wire [15-1:0] node1765;
	wire [15-1:0] node1768;
	wire [15-1:0] node1771;
	wire [15-1:0] node1772;
	wire [15-1:0] node1775;
	wire [15-1:0] node1778;
	wire [15-1:0] node1779;
	wire [15-1:0] node1780;
	wire [15-1:0] node1783;
	wire [15-1:0] node1786;
	wire [15-1:0] node1787;
	wire [15-1:0] node1790;
	wire [15-1:0] node1793;
	wire [15-1:0] node1794;
	wire [15-1:0] node1795;
	wire [15-1:0] node1796;
	wire [15-1:0] node1797;
	wire [15-1:0] node1798;
	wire [15-1:0] node1799;
	wire [15-1:0] node1802;
	wire [15-1:0] node1805;
	wire [15-1:0] node1806;
	wire [15-1:0] node1809;
	wire [15-1:0] node1812;
	wire [15-1:0] node1813;
	wire [15-1:0] node1814;
	wire [15-1:0] node1817;
	wire [15-1:0] node1820;
	wire [15-1:0] node1821;
	wire [15-1:0] node1824;
	wire [15-1:0] node1827;
	wire [15-1:0] node1828;
	wire [15-1:0] node1829;
	wire [15-1:0] node1830;
	wire [15-1:0] node1833;
	wire [15-1:0] node1836;
	wire [15-1:0] node1837;
	wire [15-1:0] node1840;
	wire [15-1:0] node1843;
	wire [15-1:0] node1844;
	wire [15-1:0] node1845;
	wire [15-1:0] node1848;
	wire [15-1:0] node1851;
	wire [15-1:0] node1852;
	wire [15-1:0] node1855;
	wire [15-1:0] node1858;
	wire [15-1:0] node1859;
	wire [15-1:0] node1860;
	wire [15-1:0] node1861;
	wire [15-1:0] node1862;
	wire [15-1:0] node1865;
	wire [15-1:0] node1868;
	wire [15-1:0] node1869;
	wire [15-1:0] node1872;
	wire [15-1:0] node1875;
	wire [15-1:0] node1876;
	wire [15-1:0] node1877;
	wire [15-1:0] node1880;
	wire [15-1:0] node1883;
	wire [15-1:0] node1884;
	wire [15-1:0] node1887;
	wire [15-1:0] node1890;
	wire [15-1:0] node1891;
	wire [15-1:0] node1892;
	wire [15-1:0] node1893;
	wire [15-1:0] node1896;
	wire [15-1:0] node1899;
	wire [15-1:0] node1900;
	wire [15-1:0] node1903;
	wire [15-1:0] node1906;
	wire [15-1:0] node1907;
	wire [15-1:0] node1908;
	wire [15-1:0] node1911;
	wire [15-1:0] node1914;
	wire [15-1:0] node1915;
	wire [15-1:0] node1918;
	wire [15-1:0] node1921;
	wire [15-1:0] node1922;
	wire [15-1:0] node1923;
	wire [15-1:0] node1924;
	wire [15-1:0] node1925;
	wire [15-1:0] node1926;
	wire [15-1:0] node1929;
	wire [15-1:0] node1932;
	wire [15-1:0] node1933;
	wire [15-1:0] node1936;
	wire [15-1:0] node1939;
	wire [15-1:0] node1940;
	wire [15-1:0] node1941;
	wire [15-1:0] node1944;
	wire [15-1:0] node1947;
	wire [15-1:0] node1948;
	wire [15-1:0] node1951;
	wire [15-1:0] node1954;
	wire [15-1:0] node1955;
	wire [15-1:0] node1956;
	wire [15-1:0] node1957;
	wire [15-1:0] node1960;
	wire [15-1:0] node1963;
	wire [15-1:0] node1964;
	wire [15-1:0] node1967;
	wire [15-1:0] node1970;
	wire [15-1:0] node1971;
	wire [15-1:0] node1972;
	wire [15-1:0] node1975;
	wire [15-1:0] node1978;
	wire [15-1:0] node1979;
	wire [15-1:0] node1982;
	wire [15-1:0] node1985;
	wire [15-1:0] node1986;
	wire [15-1:0] node1987;
	wire [15-1:0] node1988;
	wire [15-1:0] node1989;
	wire [15-1:0] node1992;
	wire [15-1:0] node1995;
	wire [15-1:0] node1996;
	wire [15-1:0] node1999;
	wire [15-1:0] node2002;
	wire [15-1:0] node2003;
	wire [15-1:0] node2004;
	wire [15-1:0] node2007;
	wire [15-1:0] node2010;
	wire [15-1:0] node2011;
	wire [15-1:0] node2014;
	wire [15-1:0] node2017;
	wire [15-1:0] node2018;
	wire [15-1:0] node2019;
	wire [15-1:0] node2020;
	wire [15-1:0] node2023;
	wire [15-1:0] node2026;
	wire [15-1:0] node2027;
	wire [15-1:0] node2030;
	wire [15-1:0] node2033;
	wire [15-1:0] node2034;
	wire [15-1:0] node2035;
	wire [15-1:0] node2038;
	wire [15-1:0] node2041;
	wire [15-1:0] node2042;
	wire [15-1:0] node2045;
	wire [15-1:0] node2048;
	wire [15-1:0] node2049;
	wire [15-1:0] node2050;
	wire [15-1:0] node2051;
	wire [15-1:0] node2052;
	wire [15-1:0] node2053;
	wire [15-1:0] node2054;
	wire [15-1:0] node2055;
	wire [15-1:0] node2056;
	wire [15-1:0] node2057;
	wire [15-1:0] node2060;
	wire [15-1:0] node2063;
	wire [15-1:0] node2064;
	wire [15-1:0] node2067;
	wire [15-1:0] node2070;
	wire [15-1:0] node2071;
	wire [15-1:0] node2072;
	wire [15-1:0] node2075;
	wire [15-1:0] node2078;
	wire [15-1:0] node2079;
	wire [15-1:0] node2082;
	wire [15-1:0] node2085;
	wire [15-1:0] node2086;
	wire [15-1:0] node2087;
	wire [15-1:0] node2088;
	wire [15-1:0] node2091;
	wire [15-1:0] node2094;
	wire [15-1:0] node2095;
	wire [15-1:0] node2098;
	wire [15-1:0] node2101;
	wire [15-1:0] node2102;
	wire [15-1:0] node2103;
	wire [15-1:0] node2106;
	wire [15-1:0] node2109;
	wire [15-1:0] node2110;
	wire [15-1:0] node2113;
	wire [15-1:0] node2116;
	wire [15-1:0] node2117;
	wire [15-1:0] node2118;
	wire [15-1:0] node2119;
	wire [15-1:0] node2120;
	wire [15-1:0] node2123;
	wire [15-1:0] node2126;
	wire [15-1:0] node2127;
	wire [15-1:0] node2130;
	wire [15-1:0] node2133;
	wire [15-1:0] node2134;
	wire [15-1:0] node2135;
	wire [15-1:0] node2138;
	wire [15-1:0] node2141;
	wire [15-1:0] node2142;
	wire [15-1:0] node2145;
	wire [15-1:0] node2148;
	wire [15-1:0] node2149;
	wire [15-1:0] node2150;
	wire [15-1:0] node2151;
	wire [15-1:0] node2154;
	wire [15-1:0] node2157;
	wire [15-1:0] node2158;
	wire [15-1:0] node2161;
	wire [15-1:0] node2164;
	wire [15-1:0] node2165;
	wire [15-1:0] node2166;
	wire [15-1:0] node2169;
	wire [15-1:0] node2172;
	wire [15-1:0] node2173;
	wire [15-1:0] node2176;
	wire [15-1:0] node2179;
	wire [15-1:0] node2180;
	wire [15-1:0] node2181;
	wire [15-1:0] node2182;
	wire [15-1:0] node2183;
	wire [15-1:0] node2184;
	wire [15-1:0] node2187;
	wire [15-1:0] node2190;
	wire [15-1:0] node2191;
	wire [15-1:0] node2194;
	wire [15-1:0] node2197;
	wire [15-1:0] node2198;
	wire [15-1:0] node2199;
	wire [15-1:0] node2202;
	wire [15-1:0] node2205;
	wire [15-1:0] node2206;
	wire [15-1:0] node2209;
	wire [15-1:0] node2212;
	wire [15-1:0] node2213;
	wire [15-1:0] node2214;
	wire [15-1:0] node2215;
	wire [15-1:0] node2218;
	wire [15-1:0] node2221;
	wire [15-1:0] node2222;
	wire [15-1:0] node2225;
	wire [15-1:0] node2228;
	wire [15-1:0] node2229;
	wire [15-1:0] node2230;
	wire [15-1:0] node2233;
	wire [15-1:0] node2236;
	wire [15-1:0] node2237;
	wire [15-1:0] node2240;
	wire [15-1:0] node2243;
	wire [15-1:0] node2244;
	wire [15-1:0] node2245;
	wire [15-1:0] node2246;
	wire [15-1:0] node2247;
	wire [15-1:0] node2250;
	wire [15-1:0] node2253;
	wire [15-1:0] node2254;
	wire [15-1:0] node2257;
	wire [15-1:0] node2260;
	wire [15-1:0] node2261;
	wire [15-1:0] node2262;
	wire [15-1:0] node2265;
	wire [15-1:0] node2268;
	wire [15-1:0] node2269;
	wire [15-1:0] node2272;
	wire [15-1:0] node2275;
	wire [15-1:0] node2276;
	wire [15-1:0] node2277;
	wire [15-1:0] node2278;
	wire [15-1:0] node2281;
	wire [15-1:0] node2284;
	wire [15-1:0] node2285;
	wire [15-1:0] node2288;
	wire [15-1:0] node2291;
	wire [15-1:0] node2292;
	wire [15-1:0] node2293;
	wire [15-1:0] node2296;
	wire [15-1:0] node2299;
	wire [15-1:0] node2300;
	wire [15-1:0] node2303;
	wire [15-1:0] node2306;
	wire [15-1:0] node2307;
	wire [15-1:0] node2308;
	wire [15-1:0] node2309;
	wire [15-1:0] node2310;
	wire [15-1:0] node2311;
	wire [15-1:0] node2312;
	wire [15-1:0] node2315;
	wire [15-1:0] node2318;
	wire [15-1:0] node2319;
	wire [15-1:0] node2322;
	wire [15-1:0] node2325;
	wire [15-1:0] node2326;
	wire [15-1:0] node2327;
	wire [15-1:0] node2330;
	wire [15-1:0] node2333;
	wire [15-1:0] node2334;
	wire [15-1:0] node2337;
	wire [15-1:0] node2340;
	wire [15-1:0] node2341;
	wire [15-1:0] node2342;
	wire [15-1:0] node2343;
	wire [15-1:0] node2346;
	wire [15-1:0] node2349;
	wire [15-1:0] node2350;
	wire [15-1:0] node2353;
	wire [15-1:0] node2356;
	wire [15-1:0] node2357;
	wire [15-1:0] node2358;
	wire [15-1:0] node2361;
	wire [15-1:0] node2364;
	wire [15-1:0] node2365;
	wire [15-1:0] node2368;
	wire [15-1:0] node2371;
	wire [15-1:0] node2372;
	wire [15-1:0] node2373;
	wire [15-1:0] node2374;
	wire [15-1:0] node2375;
	wire [15-1:0] node2378;
	wire [15-1:0] node2381;
	wire [15-1:0] node2382;
	wire [15-1:0] node2385;
	wire [15-1:0] node2388;
	wire [15-1:0] node2389;
	wire [15-1:0] node2390;
	wire [15-1:0] node2393;
	wire [15-1:0] node2396;
	wire [15-1:0] node2397;
	wire [15-1:0] node2400;
	wire [15-1:0] node2403;
	wire [15-1:0] node2404;
	wire [15-1:0] node2405;
	wire [15-1:0] node2406;
	wire [15-1:0] node2409;
	wire [15-1:0] node2412;
	wire [15-1:0] node2413;
	wire [15-1:0] node2416;
	wire [15-1:0] node2419;
	wire [15-1:0] node2420;
	wire [15-1:0] node2421;
	wire [15-1:0] node2424;
	wire [15-1:0] node2427;
	wire [15-1:0] node2428;
	wire [15-1:0] node2431;
	wire [15-1:0] node2434;
	wire [15-1:0] node2435;
	wire [15-1:0] node2436;
	wire [15-1:0] node2437;
	wire [15-1:0] node2438;
	wire [15-1:0] node2439;
	wire [15-1:0] node2442;
	wire [15-1:0] node2445;
	wire [15-1:0] node2446;
	wire [15-1:0] node2449;
	wire [15-1:0] node2452;
	wire [15-1:0] node2453;
	wire [15-1:0] node2454;
	wire [15-1:0] node2457;
	wire [15-1:0] node2460;
	wire [15-1:0] node2461;
	wire [15-1:0] node2464;
	wire [15-1:0] node2467;
	wire [15-1:0] node2468;
	wire [15-1:0] node2469;
	wire [15-1:0] node2470;
	wire [15-1:0] node2473;
	wire [15-1:0] node2476;
	wire [15-1:0] node2477;
	wire [15-1:0] node2480;
	wire [15-1:0] node2483;
	wire [15-1:0] node2484;
	wire [15-1:0] node2485;
	wire [15-1:0] node2488;
	wire [15-1:0] node2491;
	wire [15-1:0] node2492;
	wire [15-1:0] node2495;
	wire [15-1:0] node2498;
	wire [15-1:0] node2499;
	wire [15-1:0] node2500;
	wire [15-1:0] node2501;
	wire [15-1:0] node2502;
	wire [15-1:0] node2505;
	wire [15-1:0] node2508;
	wire [15-1:0] node2509;
	wire [15-1:0] node2512;
	wire [15-1:0] node2515;
	wire [15-1:0] node2516;
	wire [15-1:0] node2517;
	wire [15-1:0] node2520;
	wire [15-1:0] node2523;
	wire [15-1:0] node2524;
	wire [15-1:0] node2527;
	wire [15-1:0] node2530;
	wire [15-1:0] node2531;
	wire [15-1:0] node2532;
	wire [15-1:0] node2533;
	wire [15-1:0] node2536;
	wire [15-1:0] node2539;
	wire [15-1:0] node2540;
	wire [15-1:0] node2543;
	wire [15-1:0] node2546;
	wire [15-1:0] node2547;
	wire [15-1:0] node2548;
	wire [15-1:0] node2551;
	wire [15-1:0] node2554;
	wire [15-1:0] node2555;
	wire [15-1:0] node2558;
	wire [15-1:0] node2561;
	wire [15-1:0] node2562;
	wire [15-1:0] node2563;
	wire [15-1:0] node2564;
	wire [15-1:0] node2565;
	wire [15-1:0] node2566;
	wire [15-1:0] node2567;
	wire [15-1:0] node2568;
	wire [15-1:0] node2571;
	wire [15-1:0] node2574;
	wire [15-1:0] node2575;
	wire [15-1:0] node2578;
	wire [15-1:0] node2581;
	wire [15-1:0] node2582;
	wire [15-1:0] node2583;
	wire [15-1:0] node2586;
	wire [15-1:0] node2589;
	wire [15-1:0] node2590;
	wire [15-1:0] node2593;
	wire [15-1:0] node2596;
	wire [15-1:0] node2597;
	wire [15-1:0] node2598;
	wire [15-1:0] node2599;
	wire [15-1:0] node2602;
	wire [15-1:0] node2605;
	wire [15-1:0] node2606;
	wire [15-1:0] node2609;
	wire [15-1:0] node2612;
	wire [15-1:0] node2613;
	wire [15-1:0] node2614;
	wire [15-1:0] node2617;
	wire [15-1:0] node2620;
	wire [15-1:0] node2621;
	wire [15-1:0] node2624;
	wire [15-1:0] node2627;
	wire [15-1:0] node2628;
	wire [15-1:0] node2629;
	wire [15-1:0] node2630;
	wire [15-1:0] node2631;
	wire [15-1:0] node2634;
	wire [15-1:0] node2637;
	wire [15-1:0] node2638;
	wire [15-1:0] node2641;
	wire [15-1:0] node2644;
	wire [15-1:0] node2645;
	wire [15-1:0] node2646;
	wire [15-1:0] node2649;
	wire [15-1:0] node2652;
	wire [15-1:0] node2653;
	wire [15-1:0] node2656;
	wire [15-1:0] node2659;
	wire [15-1:0] node2660;
	wire [15-1:0] node2661;
	wire [15-1:0] node2662;
	wire [15-1:0] node2665;
	wire [15-1:0] node2668;
	wire [15-1:0] node2669;
	wire [15-1:0] node2672;
	wire [15-1:0] node2675;
	wire [15-1:0] node2676;
	wire [15-1:0] node2677;
	wire [15-1:0] node2680;
	wire [15-1:0] node2683;
	wire [15-1:0] node2684;
	wire [15-1:0] node2687;
	wire [15-1:0] node2690;
	wire [15-1:0] node2691;
	wire [15-1:0] node2692;
	wire [15-1:0] node2693;
	wire [15-1:0] node2694;
	wire [15-1:0] node2695;
	wire [15-1:0] node2698;
	wire [15-1:0] node2701;
	wire [15-1:0] node2702;
	wire [15-1:0] node2705;
	wire [15-1:0] node2708;
	wire [15-1:0] node2709;
	wire [15-1:0] node2710;
	wire [15-1:0] node2713;
	wire [15-1:0] node2716;
	wire [15-1:0] node2717;
	wire [15-1:0] node2720;
	wire [15-1:0] node2723;
	wire [15-1:0] node2724;
	wire [15-1:0] node2725;
	wire [15-1:0] node2726;
	wire [15-1:0] node2729;
	wire [15-1:0] node2732;
	wire [15-1:0] node2733;
	wire [15-1:0] node2736;
	wire [15-1:0] node2739;
	wire [15-1:0] node2740;
	wire [15-1:0] node2741;
	wire [15-1:0] node2744;
	wire [15-1:0] node2747;
	wire [15-1:0] node2748;
	wire [15-1:0] node2751;
	wire [15-1:0] node2754;
	wire [15-1:0] node2755;
	wire [15-1:0] node2756;
	wire [15-1:0] node2757;
	wire [15-1:0] node2758;
	wire [15-1:0] node2761;
	wire [15-1:0] node2764;
	wire [15-1:0] node2765;
	wire [15-1:0] node2768;
	wire [15-1:0] node2771;
	wire [15-1:0] node2772;
	wire [15-1:0] node2773;
	wire [15-1:0] node2776;
	wire [15-1:0] node2779;
	wire [15-1:0] node2780;
	wire [15-1:0] node2783;
	wire [15-1:0] node2786;
	wire [15-1:0] node2787;
	wire [15-1:0] node2788;
	wire [15-1:0] node2789;
	wire [15-1:0] node2792;
	wire [15-1:0] node2795;
	wire [15-1:0] node2796;
	wire [15-1:0] node2799;
	wire [15-1:0] node2802;
	wire [15-1:0] node2803;
	wire [15-1:0] node2804;
	wire [15-1:0] node2807;
	wire [15-1:0] node2810;
	wire [15-1:0] node2811;
	wire [15-1:0] node2814;
	wire [15-1:0] node2817;
	wire [15-1:0] node2818;
	wire [15-1:0] node2819;
	wire [15-1:0] node2820;
	wire [15-1:0] node2821;
	wire [15-1:0] node2822;
	wire [15-1:0] node2823;
	wire [15-1:0] node2826;
	wire [15-1:0] node2829;
	wire [15-1:0] node2830;
	wire [15-1:0] node2833;
	wire [15-1:0] node2836;
	wire [15-1:0] node2837;
	wire [15-1:0] node2838;
	wire [15-1:0] node2841;
	wire [15-1:0] node2844;
	wire [15-1:0] node2845;
	wire [15-1:0] node2848;
	wire [15-1:0] node2851;
	wire [15-1:0] node2852;
	wire [15-1:0] node2853;
	wire [15-1:0] node2854;
	wire [15-1:0] node2857;
	wire [15-1:0] node2860;
	wire [15-1:0] node2861;
	wire [15-1:0] node2864;
	wire [15-1:0] node2867;
	wire [15-1:0] node2868;
	wire [15-1:0] node2869;
	wire [15-1:0] node2872;
	wire [15-1:0] node2875;
	wire [15-1:0] node2876;
	wire [15-1:0] node2879;
	wire [15-1:0] node2882;
	wire [15-1:0] node2883;
	wire [15-1:0] node2884;
	wire [15-1:0] node2885;
	wire [15-1:0] node2886;
	wire [15-1:0] node2889;
	wire [15-1:0] node2892;
	wire [15-1:0] node2893;
	wire [15-1:0] node2896;
	wire [15-1:0] node2899;
	wire [15-1:0] node2900;
	wire [15-1:0] node2901;
	wire [15-1:0] node2904;
	wire [15-1:0] node2907;
	wire [15-1:0] node2908;
	wire [15-1:0] node2911;
	wire [15-1:0] node2914;
	wire [15-1:0] node2915;
	wire [15-1:0] node2916;
	wire [15-1:0] node2917;
	wire [15-1:0] node2920;
	wire [15-1:0] node2923;
	wire [15-1:0] node2924;
	wire [15-1:0] node2927;
	wire [15-1:0] node2930;
	wire [15-1:0] node2931;
	wire [15-1:0] node2932;
	wire [15-1:0] node2935;
	wire [15-1:0] node2938;
	wire [15-1:0] node2939;
	wire [15-1:0] node2942;
	wire [15-1:0] node2945;
	wire [15-1:0] node2946;
	wire [15-1:0] node2947;
	wire [15-1:0] node2948;
	wire [15-1:0] node2949;
	wire [15-1:0] node2950;
	wire [15-1:0] node2953;
	wire [15-1:0] node2956;
	wire [15-1:0] node2957;
	wire [15-1:0] node2960;
	wire [15-1:0] node2963;
	wire [15-1:0] node2964;
	wire [15-1:0] node2965;
	wire [15-1:0] node2968;
	wire [15-1:0] node2971;
	wire [15-1:0] node2972;
	wire [15-1:0] node2975;
	wire [15-1:0] node2978;
	wire [15-1:0] node2979;
	wire [15-1:0] node2980;
	wire [15-1:0] node2981;
	wire [15-1:0] node2984;
	wire [15-1:0] node2987;
	wire [15-1:0] node2988;
	wire [15-1:0] node2991;
	wire [15-1:0] node2994;
	wire [15-1:0] node2995;
	wire [15-1:0] node2996;
	wire [15-1:0] node2999;
	wire [15-1:0] node3002;
	wire [15-1:0] node3003;
	wire [15-1:0] node3006;
	wire [15-1:0] node3009;
	wire [15-1:0] node3010;
	wire [15-1:0] node3011;
	wire [15-1:0] node3012;
	wire [15-1:0] node3013;
	wire [15-1:0] node3016;
	wire [15-1:0] node3019;
	wire [15-1:0] node3020;
	wire [15-1:0] node3023;
	wire [15-1:0] node3026;
	wire [15-1:0] node3027;
	wire [15-1:0] node3028;
	wire [15-1:0] node3031;
	wire [15-1:0] node3034;
	wire [15-1:0] node3035;
	wire [15-1:0] node3038;
	wire [15-1:0] node3041;
	wire [15-1:0] node3042;
	wire [15-1:0] node3043;
	wire [15-1:0] node3044;
	wire [15-1:0] node3047;
	wire [15-1:0] node3050;
	wire [15-1:0] node3051;
	wire [15-1:0] node3054;
	wire [15-1:0] node3057;
	wire [15-1:0] node3058;
	wire [15-1:0] node3059;
	wire [15-1:0] node3062;
	wire [15-1:0] node3065;
	wire [15-1:0] node3066;
	wire [15-1:0] node3069;
	wire [15-1:0] node3072;
	wire [15-1:0] node3073;
	wire [15-1:0] node3074;
	wire [15-1:0] node3075;
	wire [15-1:0] node3076;
	wire [15-1:0] node3077;
	wire [15-1:0] node3078;
	wire [15-1:0] node3079;
	wire [15-1:0] node3080;
	wire [15-1:0] node3083;
	wire [15-1:0] node3086;
	wire [15-1:0] node3087;
	wire [15-1:0] node3090;
	wire [15-1:0] node3093;
	wire [15-1:0] node3094;
	wire [15-1:0] node3095;
	wire [15-1:0] node3098;
	wire [15-1:0] node3101;
	wire [15-1:0] node3102;
	wire [15-1:0] node3105;
	wire [15-1:0] node3108;
	wire [15-1:0] node3109;
	wire [15-1:0] node3110;
	wire [15-1:0] node3111;
	wire [15-1:0] node3114;
	wire [15-1:0] node3117;
	wire [15-1:0] node3118;
	wire [15-1:0] node3121;
	wire [15-1:0] node3124;
	wire [15-1:0] node3125;
	wire [15-1:0] node3126;
	wire [15-1:0] node3129;
	wire [15-1:0] node3132;
	wire [15-1:0] node3133;
	wire [15-1:0] node3136;
	wire [15-1:0] node3139;
	wire [15-1:0] node3140;
	wire [15-1:0] node3141;
	wire [15-1:0] node3142;
	wire [15-1:0] node3143;
	wire [15-1:0] node3146;
	wire [15-1:0] node3149;
	wire [15-1:0] node3150;
	wire [15-1:0] node3153;
	wire [15-1:0] node3156;
	wire [15-1:0] node3157;
	wire [15-1:0] node3158;
	wire [15-1:0] node3161;
	wire [15-1:0] node3164;
	wire [15-1:0] node3165;
	wire [15-1:0] node3168;
	wire [15-1:0] node3171;
	wire [15-1:0] node3172;
	wire [15-1:0] node3173;
	wire [15-1:0] node3174;
	wire [15-1:0] node3177;
	wire [15-1:0] node3180;
	wire [15-1:0] node3181;
	wire [15-1:0] node3184;
	wire [15-1:0] node3187;
	wire [15-1:0] node3188;
	wire [15-1:0] node3189;
	wire [15-1:0] node3192;
	wire [15-1:0] node3195;
	wire [15-1:0] node3196;
	wire [15-1:0] node3199;
	wire [15-1:0] node3202;
	wire [15-1:0] node3203;
	wire [15-1:0] node3204;
	wire [15-1:0] node3205;
	wire [15-1:0] node3206;
	wire [15-1:0] node3207;
	wire [15-1:0] node3210;
	wire [15-1:0] node3213;
	wire [15-1:0] node3214;
	wire [15-1:0] node3217;
	wire [15-1:0] node3220;
	wire [15-1:0] node3221;
	wire [15-1:0] node3222;
	wire [15-1:0] node3225;
	wire [15-1:0] node3228;
	wire [15-1:0] node3229;
	wire [15-1:0] node3232;
	wire [15-1:0] node3235;
	wire [15-1:0] node3236;
	wire [15-1:0] node3237;
	wire [15-1:0] node3238;
	wire [15-1:0] node3241;
	wire [15-1:0] node3244;
	wire [15-1:0] node3245;
	wire [15-1:0] node3248;
	wire [15-1:0] node3251;
	wire [15-1:0] node3252;
	wire [15-1:0] node3253;
	wire [15-1:0] node3256;
	wire [15-1:0] node3259;
	wire [15-1:0] node3260;
	wire [15-1:0] node3263;
	wire [15-1:0] node3266;
	wire [15-1:0] node3267;
	wire [15-1:0] node3268;
	wire [15-1:0] node3269;
	wire [15-1:0] node3270;
	wire [15-1:0] node3273;
	wire [15-1:0] node3276;
	wire [15-1:0] node3277;
	wire [15-1:0] node3280;
	wire [15-1:0] node3283;
	wire [15-1:0] node3284;
	wire [15-1:0] node3285;
	wire [15-1:0] node3288;
	wire [15-1:0] node3291;
	wire [15-1:0] node3292;
	wire [15-1:0] node3295;
	wire [15-1:0] node3298;
	wire [15-1:0] node3299;
	wire [15-1:0] node3300;
	wire [15-1:0] node3301;
	wire [15-1:0] node3304;
	wire [15-1:0] node3307;
	wire [15-1:0] node3308;
	wire [15-1:0] node3311;
	wire [15-1:0] node3314;
	wire [15-1:0] node3315;
	wire [15-1:0] node3316;
	wire [15-1:0] node3319;
	wire [15-1:0] node3322;
	wire [15-1:0] node3323;
	wire [15-1:0] node3326;
	wire [15-1:0] node3329;
	wire [15-1:0] node3330;
	wire [15-1:0] node3331;
	wire [15-1:0] node3332;
	wire [15-1:0] node3333;
	wire [15-1:0] node3334;
	wire [15-1:0] node3335;
	wire [15-1:0] node3338;
	wire [15-1:0] node3341;
	wire [15-1:0] node3342;
	wire [15-1:0] node3345;
	wire [15-1:0] node3348;
	wire [15-1:0] node3349;
	wire [15-1:0] node3350;
	wire [15-1:0] node3353;
	wire [15-1:0] node3356;
	wire [15-1:0] node3357;
	wire [15-1:0] node3360;
	wire [15-1:0] node3363;
	wire [15-1:0] node3364;
	wire [15-1:0] node3365;
	wire [15-1:0] node3366;
	wire [15-1:0] node3369;
	wire [15-1:0] node3372;
	wire [15-1:0] node3373;
	wire [15-1:0] node3376;
	wire [15-1:0] node3379;
	wire [15-1:0] node3380;
	wire [15-1:0] node3381;
	wire [15-1:0] node3384;
	wire [15-1:0] node3387;
	wire [15-1:0] node3388;
	wire [15-1:0] node3391;
	wire [15-1:0] node3394;
	wire [15-1:0] node3395;
	wire [15-1:0] node3396;
	wire [15-1:0] node3397;
	wire [15-1:0] node3398;
	wire [15-1:0] node3401;
	wire [15-1:0] node3404;
	wire [15-1:0] node3405;
	wire [15-1:0] node3408;
	wire [15-1:0] node3411;
	wire [15-1:0] node3412;
	wire [15-1:0] node3413;
	wire [15-1:0] node3416;
	wire [15-1:0] node3419;
	wire [15-1:0] node3420;
	wire [15-1:0] node3423;
	wire [15-1:0] node3426;
	wire [15-1:0] node3427;
	wire [15-1:0] node3428;
	wire [15-1:0] node3429;
	wire [15-1:0] node3432;
	wire [15-1:0] node3435;
	wire [15-1:0] node3436;
	wire [15-1:0] node3439;
	wire [15-1:0] node3442;
	wire [15-1:0] node3443;
	wire [15-1:0] node3444;
	wire [15-1:0] node3447;
	wire [15-1:0] node3450;
	wire [15-1:0] node3451;
	wire [15-1:0] node3454;
	wire [15-1:0] node3457;
	wire [15-1:0] node3458;
	wire [15-1:0] node3459;
	wire [15-1:0] node3460;
	wire [15-1:0] node3461;
	wire [15-1:0] node3462;
	wire [15-1:0] node3465;
	wire [15-1:0] node3468;
	wire [15-1:0] node3469;
	wire [15-1:0] node3472;
	wire [15-1:0] node3475;
	wire [15-1:0] node3476;
	wire [15-1:0] node3477;
	wire [15-1:0] node3480;
	wire [15-1:0] node3483;
	wire [15-1:0] node3484;
	wire [15-1:0] node3487;
	wire [15-1:0] node3490;
	wire [15-1:0] node3491;
	wire [15-1:0] node3492;
	wire [15-1:0] node3493;
	wire [15-1:0] node3496;
	wire [15-1:0] node3499;
	wire [15-1:0] node3500;
	wire [15-1:0] node3503;
	wire [15-1:0] node3506;
	wire [15-1:0] node3507;
	wire [15-1:0] node3508;
	wire [15-1:0] node3511;
	wire [15-1:0] node3514;
	wire [15-1:0] node3515;
	wire [15-1:0] node3518;
	wire [15-1:0] node3521;
	wire [15-1:0] node3522;
	wire [15-1:0] node3523;
	wire [15-1:0] node3524;
	wire [15-1:0] node3525;
	wire [15-1:0] node3528;
	wire [15-1:0] node3531;
	wire [15-1:0] node3532;
	wire [15-1:0] node3535;
	wire [15-1:0] node3538;
	wire [15-1:0] node3539;
	wire [15-1:0] node3540;
	wire [15-1:0] node3543;
	wire [15-1:0] node3546;
	wire [15-1:0] node3547;
	wire [15-1:0] node3550;
	wire [15-1:0] node3553;
	wire [15-1:0] node3554;
	wire [15-1:0] node3555;
	wire [15-1:0] node3556;
	wire [15-1:0] node3559;
	wire [15-1:0] node3562;
	wire [15-1:0] node3563;
	wire [15-1:0] node3566;
	wire [15-1:0] node3569;
	wire [15-1:0] node3570;
	wire [15-1:0] node3571;
	wire [15-1:0] node3574;
	wire [15-1:0] node3577;
	wire [15-1:0] node3578;
	wire [15-1:0] node3581;
	wire [15-1:0] node3584;
	wire [15-1:0] node3585;
	wire [15-1:0] node3586;
	wire [15-1:0] node3587;
	wire [15-1:0] node3588;
	wire [15-1:0] node3589;
	wire [15-1:0] node3590;
	wire [15-1:0] node3591;
	wire [15-1:0] node3594;
	wire [15-1:0] node3597;
	wire [15-1:0] node3598;
	wire [15-1:0] node3601;
	wire [15-1:0] node3604;
	wire [15-1:0] node3605;
	wire [15-1:0] node3606;
	wire [15-1:0] node3609;
	wire [15-1:0] node3612;
	wire [15-1:0] node3613;
	wire [15-1:0] node3616;
	wire [15-1:0] node3619;
	wire [15-1:0] node3620;
	wire [15-1:0] node3621;
	wire [15-1:0] node3622;
	wire [15-1:0] node3625;
	wire [15-1:0] node3628;
	wire [15-1:0] node3629;
	wire [15-1:0] node3632;
	wire [15-1:0] node3635;
	wire [15-1:0] node3636;
	wire [15-1:0] node3637;
	wire [15-1:0] node3640;
	wire [15-1:0] node3643;
	wire [15-1:0] node3644;
	wire [15-1:0] node3647;
	wire [15-1:0] node3650;
	wire [15-1:0] node3651;
	wire [15-1:0] node3652;
	wire [15-1:0] node3653;
	wire [15-1:0] node3654;
	wire [15-1:0] node3657;
	wire [15-1:0] node3660;
	wire [15-1:0] node3661;
	wire [15-1:0] node3664;
	wire [15-1:0] node3667;
	wire [15-1:0] node3668;
	wire [15-1:0] node3669;
	wire [15-1:0] node3672;
	wire [15-1:0] node3675;
	wire [15-1:0] node3676;
	wire [15-1:0] node3679;
	wire [15-1:0] node3682;
	wire [15-1:0] node3683;
	wire [15-1:0] node3684;
	wire [15-1:0] node3685;
	wire [15-1:0] node3688;
	wire [15-1:0] node3691;
	wire [15-1:0] node3692;
	wire [15-1:0] node3695;
	wire [15-1:0] node3698;
	wire [15-1:0] node3699;
	wire [15-1:0] node3700;
	wire [15-1:0] node3703;
	wire [15-1:0] node3706;
	wire [15-1:0] node3707;
	wire [15-1:0] node3710;
	wire [15-1:0] node3713;
	wire [15-1:0] node3714;
	wire [15-1:0] node3715;
	wire [15-1:0] node3716;
	wire [15-1:0] node3717;
	wire [15-1:0] node3718;
	wire [15-1:0] node3721;
	wire [15-1:0] node3724;
	wire [15-1:0] node3725;
	wire [15-1:0] node3728;
	wire [15-1:0] node3731;
	wire [15-1:0] node3732;
	wire [15-1:0] node3733;
	wire [15-1:0] node3736;
	wire [15-1:0] node3739;
	wire [15-1:0] node3740;
	wire [15-1:0] node3743;
	wire [15-1:0] node3746;
	wire [15-1:0] node3747;
	wire [15-1:0] node3748;
	wire [15-1:0] node3749;
	wire [15-1:0] node3752;
	wire [15-1:0] node3755;
	wire [15-1:0] node3756;
	wire [15-1:0] node3759;
	wire [15-1:0] node3762;
	wire [15-1:0] node3763;
	wire [15-1:0] node3764;
	wire [15-1:0] node3767;
	wire [15-1:0] node3770;
	wire [15-1:0] node3771;
	wire [15-1:0] node3774;
	wire [15-1:0] node3777;
	wire [15-1:0] node3778;
	wire [15-1:0] node3779;
	wire [15-1:0] node3780;
	wire [15-1:0] node3781;
	wire [15-1:0] node3784;
	wire [15-1:0] node3787;
	wire [15-1:0] node3788;
	wire [15-1:0] node3791;
	wire [15-1:0] node3794;
	wire [15-1:0] node3795;
	wire [15-1:0] node3796;
	wire [15-1:0] node3799;
	wire [15-1:0] node3802;
	wire [15-1:0] node3803;
	wire [15-1:0] node3806;
	wire [15-1:0] node3809;
	wire [15-1:0] node3810;
	wire [15-1:0] node3811;
	wire [15-1:0] node3812;
	wire [15-1:0] node3815;
	wire [15-1:0] node3818;
	wire [15-1:0] node3819;
	wire [15-1:0] node3822;
	wire [15-1:0] node3825;
	wire [15-1:0] node3826;
	wire [15-1:0] node3827;
	wire [15-1:0] node3830;
	wire [15-1:0] node3833;
	wire [15-1:0] node3834;
	wire [15-1:0] node3837;
	wire [15-1:0] node3840;
	wire [15-1:0] node3841;
	wire [15-1:0] node3842;
	wire [15-1:0] node3843;
	wire [15-1:0] node3844;
	wire [15-1:0] node3845;
	wire [15-1:0] node3846;
	wire [15-1:0] node3849;
	wire [15-1:0] node3852;
	wire [15-1:0] node3853;
	wire [15-1:0] node3856;
	wire [15-1:0] node3859;
	wire [15-1:0] node3860;
	wire [15-1:0] node3861;
	wire [15-1:0] node3864;
	wire [15-1:0] node3867;
	wire [15-1:0] node3868;
	wire [15-1:0] node3871;
	wire [15-1:0] node3874;
	wire [15-1:0] node3875;
	wire [15-1:0] node3876;
	wire [15-1:0] node3877;
	wire [15-1:0] node3880;
	wire [15-1:0] node3883;
	wire [15-1:0] node3884;
	wire [15-1:0] node3887;
	wire [15-1:0] node3890;
	wire [15-1:0] node3891;
	wire [15-1:0] node3892;
	wire [15-1:0] node3895;
	wire [15-1:0] node3898;
	wire [15-1:0] node3899;
	wire [15-1:0] node3902;
	wire [15-1:0] node3905;
	wire [15-1:0] node3906;
	wire [15-1:0] node3907;
	wire [15-1:0] node3908;
	wire [15-1:0] node3909;
	wire [15-1:0] node3912;
	wire [15-1:0] node3915;
	wire [15-1:0] node3916;
	wire [15-1:0] node3919;
	wire [15-1:0] node3922;
	wire [15-1:0] node3923;
	wire [15-1:0] node3924;
	wire [15-1:0] node3927;
	wire [15-1:0] node3930;
	wire [15-1:0] node3931;
	wire [15-1:0] node3934;
	wire [15-1:0] node3937;
	wire [15-1:0] node3938;
	wire [15-1:0] node3939;
	wire [15-1:0] node3940;
	wire [15-1:0] node3943;
	wire [15-1:0] node3946;
	wire [15-1:0] node3947;
	wire [15-1:0] node3950;
	wire [15-1:0] node3953;
	wire [15-1:0] node3954;
	wire [15-1:0] node3955;
	wire [15-1:0] node3958;
	wire [15-1:0] node3961;
	wire [15-1:0] node3962;
	wire [15-1:0] node3965;
	wire [15-1:0] node3968;
	wire [15-1:0] node3969;
	wire [15-1:0] node3970;
	wire [15-1:0] node3971;
	wire [15-1:0] node3972;
	wire [15-1:0] node3973;
	wire [15-1:0] node3976;
	wire [15-1:0] node3979;
	wire [15-1:0] node3980;
	wire [15-1:0] node3983;
	wire [15-1:0] node3986;
	wire [15-1:0] node3987;
	wire [15-1:0] node3988;
	wire [15-1:0] node3991;
	wire [15-1:0] node3994;
	wire [15-1:0] node3995;
	wire [15-1:0] node3998;
	wire [15-1:0] node4001;
	wire [15-1:0] node4002;
	wire [15-1:0] node4003;
	wire [15-1:0] node4004;
	wire [15-1:0] node4007;
	wire [15-1:0] node4010;
	wire [15-1:0] node4011;
	wire [15-1:0] node4014;
	wire [15-1:0] node4017;
	wire [15-1:0] node4018;
	wire [15-1:0] node4019;
	wire [15-1:0] node4022;
	wire [15-1:0] node4025;
	wire [15-1:0] node4026;
	wire [15-1:0] node4029;
	wire [15-1:0] node4032;
	wire [15-1:0] node4033;
	wire [15-1:0] node4034;
	wire [15-1:0] node4035;
	wire [15-1:0] node4036;
	wire [15-1:0] node4039;
	wire [15-1:0] node4042;
	wire [15-1:0] node4043;
	wire [15-1:0] node4046;
	wire [15-1:0] node4049;
	wire [15-1:0] node4050;
	wire [15-1:0] node4051;
	wire [15-1:0] node4054;
	wire [15-1:0] node4057;
	wire [15-1:0] node4058;
	wire [15-1:0] node4061;
	wire [15-1:0] node4064;
	wire [15-1:0] node4065;
	wire [15-1:0] node4066;
	wire [15-1:0] node4067;
	wire [15-1:0] node4070;
	wire [15-1:0] node4073;
	wire [15-1:0] node4074;
	wire [15-1:0] node4077;
	wire [15-1:0] node4080;
	wire [15-1:0] node4081;
	wire [15-1:0] node4082;
	wire [15-1:0] node4085;
	wire [15-1:0] node4088;
	wire [15-1:0] node4089;
	wire [15-1:0] node4092;

	assign outp = (inp[9]) ? node2048 : node1;
		assign node1 = (inp[12]) ? node1025 : node2;
			assign node2 = (inp[0]) ? node514 : node3;
				assign node3 = (inp[7]) ? node259 : node4;
					assign node4 = (inp[10]) ? node132 : node5;
						assign node5 = (inp[3]) ? node69 : node6;
							assign node6 = (inp[14]) ? node38 : node7;
								assign node7 = (inp[8]) ? node23 : node8;
									assign node8 = (inp[6]) ? node16 : node9;
										assign node9 = (inp[11]) ? node13 : node10;
											assign node10 = (inp[5]) ? 15'b000111111111111 : 15'b001111111111111;
											assign node13 = (inp[5]) ? 15'b000011111111111 : 15'b000111111111111;
										assign node16 = (inp[5]) ? node20 : node17;
											assign node17 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node20 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
									assign node23 = (inp[1]) ? node31 : node24;
										assign node24 = (inp[13]) ? node28 : node25;
											assign node25 = (inp[5]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node28 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node31 = (inp[4]) ? node35 : node32;
											assign node32 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node35 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node38 = (inp[5]) ? node54 : node39;
									assign node39 = (inp[8]) ? node47 : node40;
										assign node40 = (inp[4]) ? node44 : node41;
											assign node41 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node44 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node47 = (inp[6]) ? node51 : node48;
											assign node48 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node51 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node54 = (inp[13]) ? node62 : node55;
										assign node55 = (inp[1]) ? node59 : node56;
											assign node56 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node59 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node62 = (inp[11]) ? node66 : node63;
											assign node63 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node66 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node69 = (inp[6]) ? node101 : node70;
								assign node70 = (inp[14]) ? node86 : node71;
									assign node71 = (inp[5]) ? node79 : node72;
										assign node72 = (inp[8]) ? node76 : node73;
											assign node73 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node76 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node79 = (inp[1]) ? node83 : node80;
											assign node80 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node83 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node86 = (inp[4]) ? node94 : node87;
										assign node87 = (inp[8]) ? node91 : node88;
											assign node88 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node91 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node94 = (inp[5]) ? node98 : node95;
											assign node95 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node98 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node101 = (inp[1]) ? node117 : node102;
									assign node102 = (inp[5]) ? node110 : node103;
										assign node103 = (inp[4]) ? node107 : node104;
											assign node104 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node107 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node110 = (inp[13]) ? node114 : node111;
											assign node111 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node114 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node117 = (inp[2]) ? node125 : node118;
										assign node118 = (inp[14]) ? node122 : node119;
											assign node119 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node122 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node125 = (inp[13]) ? node129 : node126;
											assign node126 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node129 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
						assign node132 = (inp[5]) ? node196 : node133;
							assign node133 = (inp[1]) ? node165 : node134;
								assign node134 = (inp[6]) ? node150 : node135;
									assign node135 = (inp[8]) ? node143 : node136;
										assign node136 = (inp[11]) ? node140 : node137;
											assign node137 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node140 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node143 = (inp[13]) ? node147 : node144;
											assign node144 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node147 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node150 = (inp[3]) ? node158 : node151;
										assign node151 = (inp[8]) ? node155 : node152;
											assign node152 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node155 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node158 = (inp[4]) ? node162 : node159;
											assign node159 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node162 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node165 = (inp[4]) ? node181 : node166;
									assign node166 = (inp[3]) ? node174 : node167;
										assign node167 = (inp[11]) ? node171 : node168;
											assign node168 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node171 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node174 = (inp[14]) ? node178 : node175;
											assign node175 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node178 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node181 = (inp[14]) ? node189 : node182;
										assign node182 = (inp[11]) ? node186 : node183;
											assign node183 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node186 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node189 = (inp[3]) ? node193 : node190;
											assign node190 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node193 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node196 = (inp[14]) ? node228 : node197;
								assign node197 = (inp[11]) ? node213 : node198;
									assign node198 = (inp[8]) ? node206 : node199;
										assign node199 = (inp[13]) ? node203 : node200;
											assign node200 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node203 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node206 = (inp[1]) ? node210 : node207;
											assign node207 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node210 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node213 = (inp[1]) ? node221 : node214;
										assign node214 = (inp[6]) ? node218 : node215;
											assign node215 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node218 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node221 = (inp[2]) ? node225 : node222;
											assign node222 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node225 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node228 = (inp[3]) ? node244 : node229;
									assign node229 = (inp[8]) ? node237 : node230;
										assign node230 = (inp[4]) ? node234 : node231;
											assign node231 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node234 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node237 = (inp[2]) ? node241 : node238;
											assign node238 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node241 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node244 = (inp[6]) ? node252 : node245;
										assign node245 = (inp[2]) ? node249 : node246;
											assign node246 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node249 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node252 = (inp[2]) ? node256 : node253;
											assign node253 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node256 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
					assign node259 = (inp[2]) ? node387 : node260;
						assign node260 = (inp[4]) ? node324 : node261;
							assign node261 = (inp[13]) ? node293 : node262;
								assign node262 = (inp[8]) ? node278 : node263;
									assign node263 = (inp[3]) ? node271 : node264;
										assign node264 = (inp[10]) ? node268 : node265;
											assign node265 = (inp[11]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node268 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node271 = (inp[14]) ? node275 : node272;
											assign node272 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node275 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node278 = (inp[5]) ? node286 : node279;
										assign node279 = (inp[10]) ? node283 : node280;
											assign node280 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node283 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node286 = (inp[3]) ? node290 : node287;
											assign node287 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node290 = (inp[6]) ? 15'b000000001111111 : 15'b000000111111111;
								assign node293 = (inp[8]) ? node309 : node294;
									assign node294 = (inp[14]) ? node302 : node295;
										assign node295 = (inp[6]) ? node299 : node296;
											assign node296 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node299 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node302 = (inp[5]) ? node306 : node303;
											assign node303 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node306 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node309 = (inp[11]) ? node317 : node310;
										assign node310 = (inp[10]) ? node314 : node311;
											assign node311 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node314 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node317 = (inp[5]) ? node321 : node318;
											assign node318 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node321 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node324 = (inp[1]) ? node356 : node325;
								assign node325 = (inp[11]) ? node341 : node326;
									assign node326 = (inp[8]) ? node334 : node327;
										assign node327 = (inp[10]) ? node331 : node328;
											assign node328 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node331 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node334 = (inp[6]) ? node338 : node335;
											assign node335 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node338 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node341 = (inp[5]) ? node349 : node342;
										assign node342 = (inp[3]) ? node346 : node343;
											assign node343 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node346 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node349 = (inp[10]) ? node353 : node350;
											assign node350 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node353 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node356 = (inp[5]) ? node372 : node357;
									assign node357 = (inp[13]) ? node365 : node358;
										assign node358 = (inp[6]) ? node362 : node359;
											assign node359 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node362 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node365 = (inp[11]) ? node369 : node366;
											assign node366 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node369 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node372 = (inp[8]) ? node380 : node373;
										assign node373 = (inp[3]) ? node377 : node374;
											assign node374 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node377 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node380 = (inp[14]) ? node384 : node381;
											assign node381 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node384 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node387 = (inp[8]) ? node451 : node388;
							assign node388 = (inp[10]) ? node420 : node389;
								assign node389 = (inp[5]) ? node405 : node390;
									assign node390 = (inp[11]) ? node398 : node391;
										assign node391 = (inp[3]) ? node395 : node392;
											assign node392 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node395 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node398 = (inp[4]) ? node402 : node399;
											assign node399 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node402 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node405 = (inp[3]) ? node413 : node406;
										assign node406 = (inp[11]) ? node410 : node407;
											assign node407 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node410 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node413 = (inp[14]) ? node417 : node414;
											assign node414 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node417 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node420 = (inp[13]) ? node436 : node421;
									assign node421 = (inp[4]) ? node429 : node422;
										assign node422 = (inp[6]) ? node426 : node423;
											assign node423 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node426 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node429 = (inp[14]) ? node433 : node430;
											assign node430 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node433 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node436 = (inp[14]) ? node444 : node437;
										assign node437 = (inp[4]) ? node441 : node438;
											assign node438 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node441 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node444 = (inp[5]) ? node448 : node445;
											assign node445 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node448 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node451 = (inp[1]) ? node483 : node452;
								assign node452 = (inp[11]) ? node468 : node453;
									assign node453 = (inp[4]) ? node461 : node454;
										assign node454 = (inp[3]) ? node458 : node455;
											assign node455 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node458 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node461 = (inp[13]) ? node465 : node462;
											assign node462 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node465 = (inp[5]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node468 = (inp[10]) ? node476 : node469;
										assign node469 = (inp[6]) ? node473 : node470;
											assign node470 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node473 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node476 = (inp[6]) ? node480 : node477;
											assign node477 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node480 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node483 = (inp[14]) ? node499 : node484;
									assign node484 = (inp[11]) ? node492 : node485;
										assign node485 = (inp[5]) ? node489 : node486;
											assign node486 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node489 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node492 = (inp[6]) ? node496 : node493;
											assign node493 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node496 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node499 = (inp[6]) ? node507 : node500;
										assign node500 = (inp[4]) ? node504 : node501;
											assign node501 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node504 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node507 = (inp[11]) ? node511 : node508;
											assign node508 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node511 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
				assign node514 = (inp[6]) ? node770 : node515;
					assign node515 = (inp[10]) ? node643 : node516;
						assign node516 = (inp[13]) ? node580 : node517;
							assign node517 = (inp[2]) ? node549 : node518;
								assign node518 = (inp[8]) ? node534 : node519;
									assign node519 = (inp[7]) ? node527 : node520;
										assign node520 = (inp[3]) ? node524 : node521;
											assign node521 = (inp[11]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node524 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node527 = (inp[3]) ? node531 : node528;
											assign node528 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node531 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node534 = (inp[3]) ? node542 : node535;
										assign node535 = (inp[1]) ? node539 : node536;
											assign node536 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node539 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node542 = (inp[4]) ? node546 : node543;
											assign node543 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node546 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node549 = (inp[3]) ? node565 : node550;
									assign node550 = (inp[7]) ? node558 : node551;
										assign node551 = (inp[11]) ? node555 : node552;
											assign node552 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node555 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node558 = (inp[5]) ? node562 : node559;
											assign node559 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node562 = (inp[8]) ? 15'b000000001111111 : 15'b000000111111111;
									assign node565 = (inp[5]) ? node573 : node566;
										assign node566 = (inp[8]) ? node570 : node567;
											assign node567 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node570 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node573 = (inp[7]) ? node577 : node574;
											assign node574 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node577 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node580 = (inp[1]) ? node612 : node581;
								assign node581 = (inp[4]) ? node597 : node582;
									assign node582 = (inp[11]) ? node590 : node583;
										assign node583 = (inp[5]) ? node587 : node584;
											assign node584 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node587 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node590 = (inp[7]) ? node594 : node591;
											assign node591 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node594 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node597 = (inp[5]) ? node605 : node598;
										assign node598 = (inp[11]) ? node602 : node599;
											assign node599 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node602 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node605 = (inp[8]) ? node609 : node606;
											assign node606 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node609 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node612 = (inp[8]) ? node628 : node613;
									assign node613 = (inp[11]) ? node621 : node614;
										assign node614 = (inp[5]) ? node618 : node615;
											assign node615 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node618 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node621 = (inp[4]) ? node625 : node622;
											assign node622 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node625 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node628 = (inp[5]) ? node636 : node629;
										assign node629 = (inp[11]) ? node633 : node630;
											assign node630 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node633 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node636 = (inp[3]) ? node640 : node637;
											assign node637 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node640 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node643 = (inp[11]) ? node707 : node644;
							assign node644 = (inp[7]) ? node676 : node645;
								assign node645 = (inp[8]) ? node661 : node646;
									assign node646 = (inp[5]) ? node654 : node647;
										assign node647 = (inp[14]) ? node651 : node648;
											assign node648 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node651 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node654 = (inp[2]) ? node658 : node655;
											assign node655 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node658 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node661 = (inp[13]) ? node669 : node662;
										assign node662 = (inp[1]) ? node666 : node663;
											assign node663 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node666 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node669 = (inp[14]) ? node673 : node670;
											assign node670 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node673 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node676 = (inp[13]) ? node692 : node677;
									assign node677 = (inp[5]) ? node685 : node678;
										assign node678 = (inp[1]) ? node682 : node679;
											assign node679 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node682 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node685 = (inp[2]) ? node689 : node686;
											assign node686 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node689 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node692 = (inp[2]) ? node700 : node693;
										assign node693 = (inp[14]) ? node697 : node694;
											assign node694 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node697 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node700 = (inp[4]) ? node704 : node701;
											assign node701 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node704 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node707 = (inp[4]) ? node739 : node708;
								assign node708 = (inp[13]) ? node724 : node709;
									assign node709 = (inp[1]) ? node717 : node710;
										assign node710 = (inp[3]) ? node714 : node711;
											assign node711 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node714 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node717 = (inp[2]) ? node721 : node718;
											assign node718 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node721 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node724 = (inp[3]) ? node732 : node725;
										assign node725 = (inp[14]) ? node729 : node726;
											assign node726 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node729 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node732 = (inp[5]) ? node736 : node733;
											assign node733 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node736 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node739 = (inp[7]) ? node755 : node740;
									assign node740 = (inp[1]) ? node748 : node741;
										assign node741 = (inp[14]) ? node745 : node742;
											assign node742 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node745 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node748 = (inp[14]) ? node752 : node749;
											assign node749 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node752 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node755 = (inp[14]) ? node763 : node756;
										assign node756 = (inp[8]) ? node760 : node757;
											assign node757 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node760 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node763 = (inp[13]) ? node767 : node764;
											assign node764 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node767 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
					assign node770 = (inp[2]) ? node898 : node771;
						assign node771 = (inp[11]) ? node835 : node772;
							assign node772 = (inp[13]) ? node804 : node773;
								assign node773 = (inp[3]) ? node789 : node774;
									assign node774 = (inp[4]) ? node782 : node775;
										assign node775 = (inp[5]) ? node779 : node776;
											assign node776 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node779 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node782 = (inp[8]) ? node786 : node783;
											assign node783 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node786 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node789 = (inp[1]) ? node797 : node790;
										assign node790 = (inp[14]) ? node794 : node791;
											assign node791 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node794 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node797 = (inp[7]) ? node801 : node798;
											assign node798 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node801 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node804 = (inp[7]) ? node820 : node805;
									assign node805 = (inp[10]) ? node813 : node806;
										assign node806 = (inp[1]) ? node810 : node807;
											assign node807 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node810 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node813 = (inp[8]) ? node817 : node814;
											assign node814 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node817 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node820 = (inp[14]) ? node828 : node821;
										assign node821 = (inp[3]) ? node825 : node822;
											assign node822 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node825 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node828 = (inp[10]) ? node832 : node829;
											assign node829 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node832 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node835 = (inp[1]) ? node867 : node836;
								assign node836 = (inp[5]) ? node852 : node837;
									assign node837 = (inp[13]) ? node845 : node838;
										assign node838 = (inp[14]) ? node842 : node839;
											assign node839 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node842 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node845 = (inp[14]) ? node849 : node846;
											assign node846 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node849 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node852 = (inp[10]) ? node860 : node853;
										assign node853 = (inp[3]) ? node857 : node854;
											assign node854 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node857 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node860 = (inp[4]) ? node864 : node861;
											assign node861 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node864 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node867 = (inp[14]) ? node883 : node868;
									assign node868 = (inp[5]) ? node876 : node869;
										assign node869 = (inp[8]) ? node873 : node870;
											assign node870 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node873 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node876 = (inp[10]) ? node880 : node877;
											assign node877 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node880 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node883 = (inp[5]) ? node891 : node884;
										assign node884 = (inp[3]) ? node888 : node885;
											assign node885 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node888 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node891 = (inp[7]) ? node895 : node892;
											assign node892 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node895 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node898 = (inp[5]) ? node962 : node899;
							assign node899 = (inp[7]) ? node931 : node900;
								assign node900 = (inp[13]) ? node916 : node901;
									assign node901 = (inp[3]) ? node909 : node902;
										assign node902 = (inp[14]) ? node906 : node903;
											assign node903 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node906 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node909 = (inp[1]) ? node913 : node910;
											assign node910 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node913 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node916 = (inp[10]) ? node924 : node917;
										assign node917 = (inp[1]) ? node921 : node918;
											assign node918 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node921 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node924 = (inp[14]) ? node928 : node925;
											assign node925 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node928 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node931 = (inp[14]) ? node947 : node932;
									assign node932 = (inp[8]) ? node940 : node933;
										assign node933 = (inp[10]) ? node937 : node934;
											assign node934 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node937 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node940 = (inp[10]) ? node944 : node941;
											assign node941 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node944 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node947 = (inp[13]) ? node955 : node948;
										assign node948 = (inp[3]) ? node952 : node949;
											assign node949 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node952 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node955 = (inp[11]) ? node959 : node956;
											assign node956 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node959 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node962 = (inp[10]) ? node994 : node963;
								assign node963 = (inp[11]) ? node979 : node964;
									assign node964 = (inp[7]) ? node972 : node965;
										assign node965 = (inp[8]) ? node969 : node966;
											assign node966 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node969 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node972 = (inp[3]) ? node976 : node973;
											assign node973 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node976 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node979 = (inp[4]) ? node987 : node980;
										assign node980 = (inp[3]) ? node984 : node981;
											assign node981 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node984 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node987 = (inp[1]) ? node991 : node988;
											assign node988 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node991 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node994 = (inp[1]) ? node1010 : node995;
									assign node995 = (inp[13]) ? node1003 : node996;
										assign node996 = (inp[4]) ? node1000 : node997;
											assign node997 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1000 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1003 = (inp[14]) ? node1007 : node1004;
											assign node1004 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1007 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node1010 = (inp[3]) ? node1018 : node1011;
										assign node1011 = (inp[4]) ? node1015 : node1012;
											assign node1012 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1015 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node1018 = (inp[13]) ? node1022 : node1019;
											assign node1019 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node1022 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
			assign node1025 = (inp[3]) ? node1537 : node1026;
				assign node1026 = (inp[2]) ? node1282 : node1027;
					assign node1027 = (inp[5]) ? node1155 : node1028;
						assign node1028 = (inp[0]) ? node1092 : node1029;
							assign node1029 = (inp[10]) ? node1061 : node1030;
								assign node1030 = (inp[14]) ? node1046 : node1031;
									assign node1031 = (inp[6]) ? node1039 : node1032;
										assign node1032 = (inp[1]) ? node1036 : node1033;
											assign node1033 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node1036 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node1039 = (inp[4]) ? node1043 : node1040;
											assign node1040 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1043 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node1046 = (inp[13]) ? node1054 : node1047;
										assign node1047 = (inp[4]) ? node1051 : node1048;
											assign node1048 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1051 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1054 = (inp[7]) ? node1058 : node1055;
											assign node1055 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1058 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node1061 = (inp[1]) ? node1077 : node1062;
									assign node1062 = (inp[7]) ? node1070 : node1063;
										assign node1063 = (inp[4]) ? node1067 : node1064;
											assign node1064 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1067 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1070 = (inp[6]) ? node1074 : node1071;
											assign node1071 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1074 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1077 = (inp[11]) ? node1085 : node1078;
										assign node1078 = (inp[4]) ? node1082 : node1079;
											assign node1079 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1082 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1085 = (inp[4]) ? node1089 : node1086;
											assign node1086 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1089 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node1092 = (inp[6]) ? node1124 : node1093;
								assign node1093 = (inp[10]) ? node1109 : node1094;
									assign node1094 = (inp[13]) ? node1102 : node1095;
										assign node1095 = (inp[1]) ? node1099 : node1096;
											assign node1096 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1099 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1102 = (inp[8]) ? node1106 : node1103;
											assign node1103 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1106 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1109 = (inp[14]) ? node1117 : node1110;
										assign node1110 = (inp[11]) ? node1114 : node1111;
											assign node1111 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1114 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1117 = (inp[4]) ? node1121 : node1118;
											assign node1118 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1121 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node1124 = (inp[7]) ? node1140 : node1125;
									assign node1125 = (inp[14]) ? node1133 : node1126;
										assign node1126 = (inp[1]) ? node1130 : node1127;
											assign node1127 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1130 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1133 = (inp[4]) ? node1137 : node1134;
											assign node1134 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1137 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1140 = (inp[13]) ? node1148 : node1141;
										assign node1141 = (inp[8]) ? node1145 : node1142;
											assign node1142 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1145 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1148 = (inp[10]) ? node1152 : node1149;
											assign node1149 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1152 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node1155 = (inp[13]) ? node1219 : node1156;
							assign node1156 = (inp[14]) ? node1188 : node1157;
								assign node1157 = (inp[1]) ? node1173 : node1158;
									assign node1158 = (inp[0]) ? node1166 : node1159;
										assign node1159 = (inp[7]) ? node1163 : node1160;
											assign node1160 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1163 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1166 = (inp[4]) ? node1170 : node1167;
											assign node1167 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1170 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1173 = (inp[7]) ? node1181 : node1174;
										assign node1174 = (inp[0]) ? node1178 : node1175;
											assign node1175 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1178 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1181 = (inp[8]) ? node1185 : node1182;
											assign node1182 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1185 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node1188 = (inp[0]) ? node1204 : node1189;
									assign node1189 = (inp[1]) ? node1197 : node1190;
										assign node1190 = (inp[8]) ? node1194 : node1191;
											assign node1191 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1194 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1197 = (inp[4]) ? node1201 : node1198;
											assign node1198 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1201 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1204 = (inp[8]) ? node1212 : node1205;
										assign node1205 = (inp[11]) ? node1209 : node1206;
											assign node1206 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1209 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1212 = (inp[10]) ? node1216 : node1213;
											assign node1213 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1216 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node1219 = (inp[8]) ? node1251 : node1220;
								assign node1220 = (inp[4]) ? node1236 : node1221;
									assign node1221 = (inp[7]) ? node1229 : node1222;
										assign node1222 = (inp[1]) ? node1226 : node1223;
											assign node1223 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1226 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1229 = (inp[6]) ? node1233 : node1230;
											assign node1230 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1233 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1236 = (inp[14]) ? node1244 : node1237;
										assign node1237 = (inp[10]) ? node1241 : node1238;
											assign node1238 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1241 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1244 = (inp[6]) ? node1248 : node1245;
											assign node1245 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1248 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1251 = (inp[0]) ? node1267 : node1252;
									assign node1252 = (inp[1]) ? node1260 : node1253;
										assign node1253 = (inp[7]) ? node1257 : node1254;
											assign node1254 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1257 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1260 = (inp[11]) ? node1264 : node1261;
											assign node1261 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1264 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1267 = (inp[14]) ? node1275 : node1268;
										assign node1268 = (inp[10]) ? node1272 : node1269;
											assign node1269 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1272 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1275 = (inp[4]) ? node1279 : node1276;
											assign node1276 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1279 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
					assign node1282 = (inp[6]) ? node1410 : node1283;
						assign node1283 = (inp[11]) ? node1347 : node1284;
							assign node1284 = (inp[8]) ? node1316 : node1285;
								assign node1285 = (inp[10]) ? node1301 : node1286;
									assign node1286 = (inp[1]) ? node1294 : node1287;
										assign node1287 = (inp[4]) ? node1291 : node1288;
											assign node1288 = (inp[7]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1291 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1294 = (inp[0]) ? node1298 : node1295;
											assign node1295 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1298 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1301 = (inp[4]) ? node1309 : node1302;
										assign node1302 = (inp[14]) ? node1306 : node1303;
											assign node1303 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1306 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1309 = (inp[1]) ? node1313 : node1310;
											assign node1310 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1313 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node1316 = (inp[13]) ? node1332 : node1317;
									assign node1317 = (inp[7]) ? node1325 : node1318;
										assign node1318 = (inp[4]) ? node1322 : node1319;
											assign node1319 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1322 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1325 = (inp[10]) ? node1329 : node1326;
											assign node1326 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1329 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1332 = (inp[4]) ? node1340 : node1333;
										assign node1333 = (inp[14]) ? node1337 : node1334;
											assign node1334 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1337 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1340 = (inp[7]) ? node1344 : node1341;
											assign node1341 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1344 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node1347 = (inp[0]) ? node1379 : node1348;
								assign node1348 = (inp[7]) ? node1364 : node1349;
									assign node1349 = (inp[4]) ? node1357 : node1350;
										assign node1350 = (inp[8]) ? node1354 : node1351;
											assign node1351 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1354 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1357 = (inp[13]) ? node1361 : node1358;
											assign node1358 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1361 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1364 = (inp[13]) ? node1372 : node1365;
										assign node1365 = (inp[1]) ? node1369 : node1366;
											assign node1366 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1369 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1372 = (inp[1]) ? node1376 : node1373;
											assign node1373 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1376 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1379 = (inp[4]) ? node1395 : node1380;
									assign node1380 = (inp[13]) ? node1388 : node1381;
										assign node1381 = (inp[8]) ? node1385 : node1382;
											assign node1382 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1385 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1388 = (inp[5]) ? node1392 : node1389;
											assign node1389 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1392 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1395 = (inp[10]) ? node1403 : node1396;
										assign node1396 = (inp[7]) ? node1400 : node1397;
											assign node1397 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1400 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1403 = (inp[1]) ? node1407 : node1404;
											assign node1404 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1407 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node1410 = (inp[8]) ? node1474 : node1411;
							assign node1411 = (inp[0]) ? node1443 : node1412;
								assign node1412 = (inp[10]) ? node1428 : node1413;
									assign node1413 = (inp[1]) ? node1421 : node1414;
										assign node1414 = (inp[7]) ? node1418 : node1415;
											assign node1415 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1418 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1421 = (inp[5]) ? node1425 : node1422;
											assign node1422 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1425 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1428 = (inp[13]) ? node1436 : node1429;
										assign node1429 = (inp[1]) ? node1433 : node1430;
											assign node1430 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1433 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1436 = (inp[11]) ? node1440 : node1437;
											assign node1437 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1440 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1443 = (inp[14]) ? node1459 : node1444;
									assign node1444 = (inp[11]) ? node1452 : node1445;
										assign node1445 = (inp[1]) ? node1449 : node1446;
											assign node1446 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1449 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1452 = (inp[4]) ? node1456 : node1453;
											assign node1453 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1456 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1459 = (inp[4]) ? node1467 : node1460;
										assign node1460 = (inp[7]) ? node1464 : node1461;
											assign node1461 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1464 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1467 = (inp[1]) ? node1471 : node1468;
											assign node1468 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1471 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node1474 = (inp[10]) ? node1506 : node1475;
								assign node1475 = (inp[7]) ? node1491 : node1476;
									assign node1476 = (inp[1]) ? node1484 : node1477;
										assign node1477 = (inp[11]) ? node1481 : node1478;
											assign node1478 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1481 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1484 = (inp[13]) ? node1488 : node1485;
											assign node1485 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1488 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1491 = (inp[4]) ? node1499 : node1492;
										assign node1492 = (inp[1]) ? node1496 : node1493;
											assign node1493 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1496 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1499 = (inp[13]) ? node1503 : node1500;
											assign node1500 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1503 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node1506 = (inp[4]) ? node1522 : node1507;
									assign node1507 = (inp[1]) ? node1515 : node1508;
										assign node1508 = (inp[5]) ? node1512 : node1509;
											assign node1509 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1512 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1515 = (inp[14]) ? node1519 : node1516;
											assign node1516 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1519 = (inp[0]) ? 15'b000000000011111 : 15'b000000000011111;
									assign node1522 = (inp[11]) ? node1530 : node1523;
										assign node1523 = (inp[7]) ? node1527 : node1524;
											assign node1524 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1527 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node1530 = (inp[0]) ? node1534 : node1531;
											assign node1531 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node1534 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
				assign node1537 = (inp[13]) ? node1793 : node1538;
					assign node1538 = (inp[8]) ? node1666 : node1539;
						assign node1539 = (inp[4]) ? node1603 : node1540;
							assign node1540 = (inp[1]) ? node1572 : node1541;
								assign node1541 = (inp[10]) ? node1557 : node1542;
									assign node1542 = (inp[6]) ? node1550 : node1543;
										assign node1543 = (inp[0]) ? node1547 : node1544;
											assign node1544 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1547 = (inp[7]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1550 = (inp[7]) ? node1554 : node1551;
											assign node1551 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1554 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1557 = (inp[14]) ? node1565 : node1558;
										assign node1558 = (inp[11]) ? node1562 : node1559;
											assign node1559 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1562 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1565 = (inp[2]) ? node1569 : node1566;
											assign node1566 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1569 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node1572 = (inp[6]) ? node1588 : node1573;
									assign node1573 = (inp[11]) ? node1581 : node1574;
										assign node1574 = (inp[10]) ? node1578 : node1575;
											assign node1575 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1578 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1581 = (inp[5]) ? node1585 : node1582;
											assign node1582 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1585 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1588 = (inp[7]) ? node1596 : node1589;
										assign node1589 = (inp[0]) ? node1593 : node1590;
											assign node1590 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1593 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1596 = (inp[2]) ? node1600 : node1597;
											assign node1597 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1600 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node1603 = (inp[14]) ? node1635 : node1604;
								assign node1604 = (inp[6]) ? node1620 : node1605;
									assign node1605 = (inp[1]) ? node1613 : node1606;
										assign node1606 = (inp[5]) ? node1610 : node1607;
											assign node1607 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1610 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1613 = (inp[2]) ? node1617 : node1614;
											assign node1614 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1617 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1620 = (inp[2]) ? node1628 : node1621;
										assign node1621 = (inp[5]) ? node1625 : node1622;
											assign node1622 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1625 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1628 = (inp[11]) ? node1632 : node1629;
											assign node1629 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1632 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1635 = (inp[1]) ? node1651 : node1636;
									assign node1636 = (inp[11]) ? node1644 : node1637;
										assign node1637 = (inp[0]) ? node1641 : node1638;
											assign node1638 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1641 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1644 = (inp[7]) ? node1648 : node1645;
											assign node1645 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1648 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1651 = (inp[2]) ? node1659 : node1652;
										assign node1652 = (inp[0]) ? node1656 : node1653;
											assign node1653 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1656 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1659 = (inp[10]) ? node1663 : node1660;
											assign node1660 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1663 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node1666 = (inp[5]) ? node1730 : node1667;
							assign node1667 = (inp[6]) ? node1699 : node1668;
								assign node1668 = (inp[14]) ? node1684 : node1669;
									assign node1669 = (inp[1]) ? node1677 : node1670;
										assign node1670 = (inp[2]) ? node1674 : node1671;
											assign node1671 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1674 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1677 = (inp[10]) ? node1681 : node1678;
											assign node1678 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1681 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1684 = (inp[7]) ? node1692 : node1685;
										assign node1685 = (inp[10]) ? node1689 : node1686;
											assign node1686 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1689 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1692 = (inp[0]) ? node1696 : node1693;
											assign node1693 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1696 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1699 = (inp[1]) ? node1715 : node1700;
									assign node1700 = (inp[7]) ? node1708 : node1701;
										assign node1701 = (inp[10]) ? node1705 : node1702;
											assign node1702 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1705 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1708 = (inp[2]) ? node1712 : node1709;
											assign node1709 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1712 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1715 = (inp[11]) ? node1723 : node1716;
										assign node1716 = (inp[0]) ? node1720 : node1717;
											assign node1717 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1720 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1723 = (inp[10]) ? node1727 : node1724;
											assign node1724 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1727 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node1730 = (inp[0]) ? node1762 : node1731;
								assign node1731 = (inp[2]) ? node1747 : node1732;
									assign node1732 = (inp[4]) ? node1740 : node1733;
										assign node1733 = (inp[7]) ? node1737 : node1734;
											assign node1734 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1737 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1740 = (inp[14]) ? node1744 : node1741;
											assign node1741 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1744 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1747 = (inp[11]) ? node1755 : node1748;
										assign node1748 = (inp[1]) ? node1752 : node1749;
											assign node1749 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1752 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1755 = (inp[6]) ? node1759 : node1756;
											assign node1756 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1759 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node1762 = (inp[11]) ? node1778 : node1763;
									assign node1763 = (inp[14]) ? node1771 : node1764;
										assign node1764 = (inp[1]) ? node1768 : node1765;
											assign node1765 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1768 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1771 = (inp[10]) ? node1775 : node1772;
											assign node1772 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1775 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node1778 = (inp[4]) ? node1786 : node1779;
										assign node1779 = (inp[10]) ? node1783 : node1780;
											assign node1780 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1783 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node1786 = (inp[7]) ? node1790 : node1787;
											assign node1787 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node1790 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
					assign node1793 = (inp[11]) ? node1921 : node1794;
						assign node1794 = (inp[10]) ? node1858 : node1795;
							assign node1795 = (inp[14]) ? node1827 : node1796;
								assign node1796 = (inp[7]) ? node1812 : node1797;
									assign node1797 = (inp[5]) ? node1805 : node1798;
										assign node1798 = (inp[6]) ? node1802 : node1799;
											assign node1799 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1802 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1805 = (inp[4]) ? node1809 : node1806;
											assign node1806 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1809 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1812 = (inp[5]) ? node1820 : node1813;
										assign node1813 = (inp[8]) ? node1817 : node1814;
											assign node1814 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1817 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1820 = (inp[0]) ? node1824 : node1821;
											assign node1821 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1824 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node1827 = (inp[1]) ? node1843 : node1828;
									assign node1828 = (inp[6]) ? node1836 : node1829;
										assign node1829 = (inp[8]) ? node1833 : node1830;
											assign node1830 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1833 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1836 = (inp[5]) ? node1840 : node1837;
											assign node1837 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1840 = (inp[4]) ? 15'b000000000011111 : 15'b000000001111111;
									assign node1843 = (inp[4]) ? node1851 : node1844;
										assign node1844 = (inp[2]) ? node1848 : node1845;
											assign node1845 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1848 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1851 = (inp[2]) ? node1855 : node1852;
											assign node1852 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1855 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node1858 = (inp[0]) ? node1890 : node1859;
								assign node1859 = (inp[6]) ? node1875 : node1860;
									assign node1860 = (inp[1]) ? node1868 : node1861;
										assign node1861 = (inp[5]) ? node1865 : node1862;
											assign node1862 = (inp[7]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1865 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1868 = (inp[8]) ? node1872 : node1869;
											assign node1869 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1872 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1875 = (inp[8]) ? node1883 : node1876;
										assign node1876 = (inp[2]) ? node1880 : node1877;
											assign node1877 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1880 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1883 = (inp[4]) ? node1887 : node1884;
											assign node1884 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1887 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node1890 = (inp[8]) ? node1906 : node1891;
									assign node1891 = (inp[2]) ? node1899 : node1892;
										assign node1892 = (inp[1]) ? node1896 : node1893;
											assign node1893 = (inp[7]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1896 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1899 = (inp[6]) ? node1903 : node1900;
											assign node1900 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1903 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node1906 = (inp[7]) ? node1914 : node1907;
										assign node1907 = (inp[4]) ? node1911 : node1908;
											assign node1908 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1911 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node1914 = (inp[1]) ? node1918 : node1915;
											assign node1915 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node1918 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node1921 = (inp[14]) ? node1985 : node1922;
							assign node1922 = (inp[1]) ? node1954 : node1923;
								assign node1923 = (inp[4]) ? node1939 : node1924;
									assign node1924 = (inp[6]) ? node1932 : node1925;
										assign node1925 = (inp[7]) ? node1929 : node1926;
											assign node1926 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1929 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1932 = (inp[5]) ? node1936 : node1933;
											assign node1933 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1936 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1939 = (inp[10]) ? node1947 : node1940;
										assign node1940 = (inp[5]) ? node1944 : node1941;
											assign node1941 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1944 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1947 = (inp[0]) ? node1951 : node1948;
											assign node1948 = (inp[7]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1951 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node1954 = (inp[10]) ? node1970 : node1955;
									assign node1955 = (inp[2]) ? node1963 : node1956;
										assign node1956 = (inp[0]) ? node1960 : node1957;
											assign node1957 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1960 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1963 = (inp[7]) ? node1967 : node1964;
											assign node1964 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1967 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node1970 = (inp[5]) ? node1978 : node1971;
										assign node1971 = (inp[7]) ? node1975 : node1972;
											assign node1972 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1975 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node1978 = (inp[4]) ? node1982 : node1979;
											assign node1979 = (inp[7]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node1982 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node1985 = (inp[2]) ? node2017 : node1986;
								assign node1986 = (inp[0]) ? node2002 : node1987;
									assign node1987 = (inp[5]) ? node1995 : node1988;
										assign node1988 = (inp[4]) ? node1992 : node1989;
											assign node1989 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1992 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1995 = (inp[10]) ? node1999 : node1996;
											assign node1996 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1999 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2002 = (inp[7]) ? node2010 : node2003;
										assign node2003 = (inp[8]) ? node2007 : node2004;
											assign node2004 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2007 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2010 = (inp[8]) ? node2014 : node2011;
											assign node2011 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2014 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node2017 = (inp[4]) ? node2033 : node2018;
									assign node2018 = (inp[1]) ? node2026 : node2019;
										assign node2019 = (inp[0]) ? node2023 : node2020;
											assign node2020 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2023 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2026 = (inp[7]) ? node2030 : node2027;
											assign node2027 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2030 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node2033 = (inp[5]) ? node2041 : node2034;
										assign node2034 = (inp[7]) ? node2038 : node2035;
											assign node2035 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2038 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node2041 = (inp[6]) ? node2045 : node2042;
											assign node2042 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node2045 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
		assign node2048 = (inp[7]) ? node3072 : node2049;
			assign node2049 = (inp[11]) ? node2561 : node2050;
				assign node2050 = (inp[14]) ? node2306 : node2051;
					assign node2051 = (inp[2]) ? node2179 : node2052;
						assign node2052 = (inp[12]) ? node2116 : node2053;
							assign node2053 = (inp[1]) ? node2085 : node2054;
								assign node2054 = (inp[5]) ? node2070 : node2055;
									assign node2055 = (inp[4]) ? node2063 : node2056;
										assign node2056 = (inp[3]) ? node2060 : node2057;
											assign node2057 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node2060 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node2063 = (inp[6]) ? node2067 : node2064;
											assign node2064 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2067 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node2070 = (inp[6]) ? node2078 : node2071;
										assign node2071 = (inp[13]) ? node2075 : node2072;
											assign node2072 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2075 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2078 = (inp[4]) ? node2082 : node2079;
											assign node2079 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2082 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node2085 = (inp[0]) ? node2101 : node2086;
									assign node2086 = (inp[10]) ? node2094 : node2087;
										assign node2087 = (inp[4]) ? node2091 : node2088;
											assign node2088 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2091 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2094 = (inp[5]) ? node2098 : node2095;
											assign node2095 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2098 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node2101 = (inp[6]) ? node2109 : node2102;
										assign node2102 = (inp[10]) ? node2106 : node2103;
											assign node2103 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2106 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2109 = (inp[5]) ? node2113 : node2110;
											assign node2110 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2113 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node2116 = (inp[13]) ? node2148 : node2117;
								assign node2117 = (inp[10]) ? node2133 : node2118;
									assign node2118 = (inp[8]) ? node2126 : node2119;
										assign node2119 = (inp[1]) ? node2123 : node2120;
											assign node2120 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2123 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2126 = (inp[5]) ? node2130 : node2127;
											assign node2127 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2130 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node2133 = (inp[5]) ? node2141 : node2134;
										assign node2134 = (inp[4]) ? node2138 : node2135;
											assign node2135 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2138 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2141 = (inp[1]) ? node2145 : node2142;
											assign node2142 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2145 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node2148 = (inp[10]) ? node2164 : node2149;
									assign node2149 = (inp[3]) ? node2157 : node2150;
										assign node2150 = (inp[0]) ? node2154 : node2151;
											assign node2151 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2154 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2157 = (inp[4]) ? node2161 : node2158;
											assign node2158 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2161 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2164 = (inp[5]) ? node2172 : node2165;
										assign node2165 = (inp[8]) ? node2169 : node2166;
											assign node2166 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2169 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2172 = (inp[6]) ? node2176 : node2173;
											assign node2173 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2176 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
						assign node2179 = (inp[10]) ? node2243 : node2180;
							assign node2180 = (inp[3]) ? node2212 : node2181;
								assign node2181 = (inp[5]) ? node2197 : node2182;
									assign node2182 = (inp[0]) ? node2190 : node2183;
										assign node2183 = (inp[8]) ? node2187 : node2184;
											assign node2184 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2187 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2190 = (inp[12]) ? node2194 : node2191;
											assign node2191 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2194 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node2197 = (inp[13]) ? node2205 : node2198;
										assign node2198 = (inp[8]) ? node2202 : node2199;
											assign node2199 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2202 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2205 = (inp[0]) ? node2209 : node2206;
											assign node2206 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2209 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node2212 = (inp[0]) ? node2228 : node2213;
									assign node2213 = (inp[1]) ? node2221 : node2214;
										assign node2214 = (inp[13]) ? node2218 : node2215;
											assign node2215 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2218 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2221 = (inp[6]) ? node2225 : node2222;
											assign node2222 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2225 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2228 = (inp[1]) ? node2236 : node2229;
										assign node2229 = (inp[6]) ? node2233 : node2230;
											assign node2230 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2233 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2236 = (inp[12]) ? node2240 : node2237;
											assign node2237 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2240 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node2243 = (inp[1]) ? node2275 : node2244;
								assign node2244 = (inp[8]) ? node2260 : node2245;
									assign node2245 = (inp[5]) ? node2253 : node2246;
										assign node2246 = (inp[13]) ? node2250 : node2247;
											assign node2247 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2250 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2253 = (inp[3]) ? node2257 : node2254;
											assign node2254 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2257 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2260 = (inp[0]) ? node2268 : node2261;
										assign node2261 = (inp[5]) ? node2265 : node2262;
											assign node2262 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2265 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2268 = (inp[12]) ? node2272 : node2269;
											assign node2269 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2272 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node2275 = (inp[8]) ? node2291 : node2276;
									assign node2276 = (inp[13]) ? node2284 : node2277;
										assign node2277 = (inp[6]) ? node2281 : node2278;
											assign node2278 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2281 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2284 = (inp[0]) ? node2288 : node2285;
											assign node2285 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2288 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2291 = (inp[5]) ? node2299 : node2292;
										assign node2292 = (inp[13]) ? node2296 : node2293;
											assign node2293 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2296 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2299 = (inp[13]) ? node2303 : node2300;
											assign node2300 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2303 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
					assign node2306 = (inp[6]) ? node2434 : node2307;
						assign node2307 = (inp[1]) ? node2371 : node2308;
							assign node2308 = (inp[2]) ? node2340 : node2309;
								assign node2309 = (inp[13]) ? node2325 : node2310;
									assign node2310 = (inp[3]) ? node2318 : node2311;
										assign node2311 = (inp[0]) ? node2315 : node2312;
											assign node2312 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2315 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2318 = (inp[10]) ? node2322 : node2319;
											assign node2319 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2322 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node2325 = (inp[12]) ? node2333 : node2326;
										assign node2326 = (inp[4]) ? node2330 : node2327;
											assign node2327 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2330 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2333 = (inp[8]) ? node2337 : node2334;
											assign node2334 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2337 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node2340 = (inp[4]) ? node2356 : node2341;
									assign node2341 = (inp[12]) ? node2349 : node2342;
										assign node2342 = (inp[13]) ? node2346 : node2343;
											assign node2343 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2346 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2349 = (inp[8]) ? node2353 : node2350;
											assign node2350 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2353 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2356 = (inp[3]) ? node2364 : node2357;
										assign node2357 = (inp[8]) ? node2361 : node2358;
											assign node2358 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2361 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2364 = (inp[12]) ? node2368 : node2365;
											assign node2365 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2368 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node2371 = (inp[13]) ? node2403 : node2372;
								assign node2372 = (inp[4]) ? node2388 : node2373;
									assign node2373 = (inp[0]) ? node2381 : node2374;
										assign node2374 = (inp[2]) ? node2378 : node2375;
											assign node2375 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2378 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2381 = (inp[8]) ? node2385 : node2382;
											assign node2382 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2385 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2388 = (inp[0]) ? node2396 : node2389;
										assign node2389 = (inp[12]) ? node2393 : node2390;
											assign node2390 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2393 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2396 = (inp[10]) ? node2400 : node2397;
											assign node2397 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2400 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node2403 = (inp[3]) ? node2419 : node2404;
									assign node2404 = (inp[5]) ? node2412 : node2405;
										assign node2405 = (inp[10]) ? node2409 : node2406;
											assign node2406 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2409 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2412 = (inp[12]) ? node2416 : node2413;
											assign node2413 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2416 = (inp[2]) ? 15'b000000000011111 : 15'b000000001111111;
									assign node2419 = (inp[4]) ? node2427 : node2420;
										assign node2420 = (inp[5]) ? node2424 : node2421;
											assign node2421 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2424 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2427 = (inp[2]) ? node2431 : node2428;
											assign node2428 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2431 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node2434 = (inp[3]) ? node2498 : node2435;
							assign node2435 = (inp[0]) ? node2467 : node2436;
								assign node2436 = (inp[2]) ? node2452 : node2437;
									assign node2437 = (inp[5]) ? node2445 : node2438;
										assign node2438 = (inp[8]) ? node2442 : node2439;
											assign node2439 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2442 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2445 = (inp[13]) ? node2449 : node2446;
											assign node2446 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2449 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2452 = (inp[10]) ? node2460 : node2453;
										assign node2453 = (inp[4]) ? node2457 : node2454;
											assign node2454 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2457 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2460 = (inp[5]) ? node2464 : node2461;
											assign node2461 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2464 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node2467 = (inp[13]) ? node2483 : node2468;
									assign node2468 = (inp[2]) ? node2476 : node2469;
										assign node2469 = (inp[8]) ? node2473 : node2470;
											assign node2470 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2473 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2476 = (inp[4]) ? node2480 : node2477;
											assign node2477 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2480 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2483 = (inp[4]) ? node2491 : node2484;
										assign node2484 = (inp[1]) ? node2488 : node2485;
											assign node2485 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2488 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2491 = (inp[12]) ? node2495 : node2492;
											assign node2492 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2495 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node2498 = (inp[12]) ? node2530 : node2499;
								assign node2499 = (inp[5]) ? node2515 : node2500;
									assign node2500 = (inp[4]) ? node2508 : node2501;
										assign node2501 = (inp[8]) ? node2505 : node2502;
											assign node2502 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2505 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2508 = (inp[1]) ? node2512 : node2509;
											assign node2509 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2512 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2515 = (inp[8]) ? node2523 : node2516;
										assign node2516 = (inp[0]) ? node2520 : node2517;
											assign node2517 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2520 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2523 = (inp[1]) ? node2527 : node2524;
											assign node2524 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2527 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node2530 = (inp[1]) ? node2546 : node2531;
									assign node2531 = (inp[0]) ? node2539 : node2532;
										assign node2532 = (inp[5]) ? node2536 : node2533;
											assign node2533 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2536 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2539 = (inp[13]) ? node2543 : node2540;
											assign node2540 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2543 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2546 = (inp[5]) ? node2554 : node2547;
										assign node2547 = (inp[8]) ? node2551 : node2548;
											assign node2548 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2551 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2554 = (inp[8]) ? node2558 : node2555;
											assign node2555 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2558 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
				assign node2561 = (inp[0]) ? node2817 : node2562;
					assign node2562 = (inp[12]) ? node2690 : node2563;
						assign node2563 = (inp[4]) ? node2627 : node2564;
							assign node2564 = (inp[10]) ? node2596 : node2565;
								assign node2565 = (inp[13]) ? node2581 : node2566;
									assign node2566 = (inp[14]) ? node2574 : node2567;
										assign node2567 = (inp[6]) ? node2571 : node2568;
											assign node2568 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2571 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2574 = (inp[8]) ? node2578 : node2575;
											assign node2575 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2578 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node2581 = (inp[2]) ? node2589 : node2582;
										assign node2582 = (inp[6]) ? node2586 : node2583;
											assign node2583 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2586 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2589 = (inp[1]) ? node2593 : node2590;
											assign node2590 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2593 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node2596 = (inp[6]) ? node2612 : node2597;
									assign node2597 = (inp[8]) ? node2605 : node2598;
										assign node2598 = (inp[14]) ? node2602 : node2599;
											assign node2599 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2602 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2605 = (inp[2]) ? node2609 : node2606;
											assign node2606 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2609 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2612 = (inp[8]) ? node2620 : node2613;
										assign node2613 = (inp[2]) ? node2617 : node2614;
											assign node2614 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2617 = (inp[1]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node2620 = (inp[13]) ? node2624 : node2621;
											assign node2621 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2624 = (inp[3]) ? 15'b000000000111111 : 15'b000000000111111;
							assign node2627 = (inp[13]) ? node2659 : node2628;
								assign node2628 = (inp[1]) ? node2644 : node2629;
									assign node2629 = (inp[14]) ? node2637 : node2630;
										assign node2630 = (inp[3]) ? node2634 : node2631;
											assign node2631 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2634 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2637 = (inp[8]) ? node2641 : node2638;
											assign node2638 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2641 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2644 = (inp[8]) ? node2652 : node2645;
										assign node2645 = (inp[14]) ? node2649 : node2646;
											assign node2646 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2649 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2652 = (inp[3]) ? node2656 : node2653;
											assign node2653 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2656 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node2659 = (inp[3]) ? node2675 : node2660;
									assign node2660 = (inp[2]) ? node2668 : node2661;
										assign node2661 = (inp[8]) ? node2665 : node2662;
											assign node2662 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2665 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2668 = (inp[10]) ? node2672 : node2669;
											assign node2669 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2672 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2675 = (inp[14]) ? node2683 : node2676;
										assign node2676 = (inp[6]) ? node2680 : node2677;
											assign node2677 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2680 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2683 = (inp[5]) ? node2687 : node2684;
											assign node2684 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2687 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node2690 = (inp[5]) ? node2754 : node2691;
							assign node2691 = (inp[3]) ? node2723 : node2692;
								assign node2692 = (inp[8]) ? node2708 : node2693;
									assign node2693 = (inp[10]) ? node2701 : node2694;
										assign node2694 = (inp[1]) ? node2698 : node2695;
											assign node2695 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2698 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2701 = (inp[6]) ? node2705 : node2702;
											assign node2702 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2705 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2708 = (inp[2]) ? node2716 : node2709;
										assign node2709 = (inp[6]) ? node2713 : node2710;
											assign node2710 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2713 = (inp[13]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node2716 = (inp[6]) ? node2720 : node2717;
											assign node2717 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2720 = (inp[13]) ? 15'b000000000011111 : 15'b000000001111111;
								assign node2723 = (inp[1]) ? node2739 : node2724;
									assign node2724 = (inp[14]) ? node2732 : node2725;
										assign node2725 = (inp[10]) ? node2729 : node2726;
											assign node2726 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2729 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2732 = (inp[8]) ? node2736 : node2733;
											assign node2733 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2736 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2739 = (inp[6]) ? node2747 : node2740;
										assign node2740 = (inp[13]) ? node2744 : node2741;
											assign node2741 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2744 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2747 = (inp[4]) ? node2751 : node2748;
											assign node2748 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2751 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node2754 = (inp[1]) ? node2786 : node2755;
								assign node2755 = (inp[6]) ? node2771 : node2756;
									assign node2756 = (inp[2]) ? node2764 : node2757;
										assign node2757 = (inp[3]) ? node2761 : node2758;
											assign node2758 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2761 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2764 = (inp[10]) ? node2768 : node2765;
											assign node2765 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2768 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2771 = (inp[13]) ? node2779 : node2772;
										assign node2772 = (inp[10]) ? node2776 : node2773;
											assign node2773 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2776 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2779 = (inp[14]) ? node2783 : node2780;
											assign node2780 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2783 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node2786 = (inp[14]) ? node2802 : node2787;
									assign node2787 = (inp[10]) ? node2795 : node2788;
										assign node2788 = (inp[8]) ? node2792 : node2789;
											assign node2789 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2792 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2795 = (inp[6]) ? node2799 : node2796;
											assign node2796 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2799 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2802 = (inp[6]) ? node2810 : node2803;
										assign node2803 = (inp[3]) ? node2807 : node2804;
											assign node2804 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2807 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2810 = (inp[10]) ? node2814 : node2811;
											assign node2811 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2814 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
					assign node2817 = (inp[13]) ? node2945 : node2818;
						assign node2818 = (inp[14]) ? node2882 : node2819;
							assign node2819 = (inp[1]) ? node2851 : node2820;
								assign node2820 = (inp[8]) ? node2836 : node2821;
									assign node2821 = (inp[4]) ? node2829 : node2822;
										assign node2822 = (inp[6]) ? node2826 : node2823;
											assign node2823 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2826 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2829 = (inp[2]) ? node2833 : node2830;
											assign node2830 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2833 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2836 = (inp[2]) ? node2844 : node2837;
										assign node2837 = (inp[3]) ? node2841 : node2838;
											assign node2838 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2841 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2844 = (inp[12]) ? node2848 : node2845;
											assign node2845 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2848 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node2851 = (inp[12]) ? node2867 : node2852;
									assign node2852 = (inp[4]) ? node2860 : node2853;
										assign node2853 = (inp[3]) ? node2857 : node2854;
											assign node2854 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2857 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2860 = (inp[6]) ? node2864 : node2861;
											assign node2861 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2864 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2867 = (inp[4]) ? node2875 : node2868;
										assign node2868 = (inp[5]) ? node2872 : node2869;
											assign node2869 = (inp[3]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node2872 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2875 = (inp[5]) ? node2879 : node2876;
											assign node2876 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2879 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node2882 = (inp[5]) ? node2914 : node2883;
								assign node2883 = (inp[12]) ? node2899 : node2884;
									assign node2884 = (inp[1]) ? node2892 : node2885;
										assign node2885 = (inp[2]) ? node2889 : node2886;
											assign node2886 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2889 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2892 = (inp[8]) ? node2896 : node2893;
											assign node2893 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2896 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2899 = (inp[2]) ? node2907 : node2900;
										assign node2900 = (inp[4]) ? node2904 : node2901;
											assign node2901 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2904 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2907 = (inp[3]) ? node2911 : node2908;
											assign node2908 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2911 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node2914 = (inp[4]) ? node2930 : node2915;
									assign node2915 = (inp[8]) ? node2923 : node2916;
										assign node2916 = (inp[6]) ? node2920 : node2917;
											assign node2917 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2920 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2923 = (inp[12]) ? node2927 : node2924;
											assign node2924 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2927 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2930 = (inp[6]) ? node2938 : node2931;
										assign node2931 = (inp[2]) ? node2935 : node2932;
											assign node2932 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2935 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2938 = (inp[12]) ? node2942 : node2939;
											assign node2939 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2942 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node2945 = (inp[8]) ? node3009 : node2946;
							assign node2946 = (inp[10]) ? node2978 : node2947;
								assign node2947 = (inp[3]) ? node2963 : node2948;
									assign node2948 = (inp[4]) ? node2956 : node2949;
										assign node2949 = (inp[2]) ? node2953 : node2950;
											assign node2950 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2953 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2956 = (inp[1]) ? node2960 : node2957;
											assign node2957 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2960 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2963 = (inp[2]) ? node2971 : node2964;
										assign node2964 = (inp[1]) ? node2968 : node2965;
											assign node2965 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2968 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2971 = (inp[4]) ? node2975 : node2972;
											assign node2972 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2975 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node2978 = (inp[1]) ? node2994 : node2979;
									assign node2979 = (inp[3]) ? node2987 : node2980;
										assign node2980 = (inp[14]) ? node2984 : node2981;
											assign node2981 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2984 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2987 = (inp[5]) ? node2991 : node2988;
											assign node2988 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2991 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node2994 = (inp[6]) ? node3002 : node2995;
										assign node2995 = (inp[2]) ? node2999 : node2996;
											assign node2996 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2999 = (inp[5]) ? 15'b000000000001111 : 15'b000000000111111;
										assign node3002 = (inp[2]) ? node3006 : node3003;
											assign node3003 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3006 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node3009 = (inp[6]) ? node3041 : node3010;
								assign node3010 = (inp[14]) ? node3026 : node3011;
									assign node3011 = (inp[3]) ? node3019 : node3012;
										assign node3012 = (inp[1]) ? node3016 : node3013;
											assign node3013 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3016 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3019 = (inp[10]) ? node3023 : node3020;
											assign node3020 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3023 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3026 = (inp[3]) ? node3034 : node3027;
										assign node3027 = (inp[4]) ? node3031 : node3028;
											assign node3028 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3031 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3034 = (inp[2]) ? node3038 : node3035;
											assign node3035 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3038 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node3041 = (inp[2]) ? node3057 : node3042;
									assign node3042 = (inp[12]) ? node3050 : node3043;
										assign node3043 = (inp[14]) ? node3047 : node3044;
											assign node3044 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3047 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3050 = (inp[10]) ? node3054 : node3051;
											assign node3051 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3054 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node3057 = (inp[5]) ? node3065 : node3058;
										assign node3058 = (inp[3]) ? node3062 : node3059;
											assign node3059 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3062 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node3065 = (inp[4]) ? node3069 : node3066;
											assign node3066 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node3069 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
			assign node3072 = (inp[4]) ? node3584 : node3073;
				assign node3073 = (inp[10]) ? node3329 : node3074;
					assign node3074 = (inp[2]) ? node3202 : node3075;
						assign node3075 = (inp[14]) ? node3139 : node3076;
							assign node3076 = (inp[13]) ? node3108 : node3077;
								assign node3077 = (inp[12]) ? node3093 : node3078;
									assign node3078 = (inp[3]) ? node3086 : node3079;
										assign node3079 = (inp[0]) ? node3083 : node3080;
											assign node3080 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node3083 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node3086 = (inp[11]) ? node3090 : node3087;
											assign node3087 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3090 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node3093 = (inp[0]) ? node3101 : node3094;
										assign node3094 = (inp[5]) ? node3098 : node3095;
											assign node3095 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3098 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3101 = (inp[6]) ? node3105 : node3102;
											assign node3102 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3105 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node3108 = (inp[6]) ? node3124 : node3109;
									assign node3109 = (inp[0]) ? node3117 : node3110;
										assign node3110 = (inp[8]) ? node3114 : node3111;
											assign node3111 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3114 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3117 = (inp[3]) ? node3121 : node3118;
											assign node3118 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3121 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node3124 = (inp[5]) ? node3132 : node3125;
										assign node3125 = (inp[11]) ? node3129 : node3126;
											assign node3126 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3129 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3132 = (inp[8]) ? node3136 : node3133;
											assign node3133 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3136 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node3139 = (inp[0]) ? node3171 : node3140;
								assign node3140 = (inp[1]) ? node3156 : node3141;
									assign node3141 = (inp[11]) ? node3149 : node3142;
										assign node3142 = (inp[5]) ? node3146 : node3143;
											assign node3143 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3146 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3149 = (inp[13]) ? node3153 : node3150;
											assign node3150 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3153 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node3156 = (inp[8]) ? node3164 : node3157;
										assign node3157 = (inp[12]) ? node3161 : node3158;
											assign node3158 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3161 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3164 = (inp[6]) ? node3168 : node3165;
											assign node3165 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3168 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node3171 = (inp[3]) ? node3187 : node3172;
									assign node3172 = (inp[11]) ? node3180 : node3173;
										assign node3173 = (inp[8]) ? node3177 : node3174;
											assign node3174 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3177 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3180 = (inp[5]) ? node3184 : node3181;
											assign node3181 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3184 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3187 = (inp[8]) ? node3195 : node3188;
										assign node3188 = (inp[1]) ? node3192 : node3189;
											assign node3189 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3192 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3195 = (inp[6]) ? node3199 : node3196;
											assign node3196 = (inp[12]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node3199 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node3202 = (inp[8]) ? node3266 : node3203;
							assign node3203 = (inp[1]) ? node3235 : node3204;
								assign node3204 = (inp[5]) ? node3220 : node3205;
									assign node3205 = (inp[3]) ? node3213 : node3206;
										assign node3206 = (inp[12]) ? node3210 : node3207;
											assign node3207 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3210 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3213 = (inp[13]) ? node3217 : node3214;
											assign node3214 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3217 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node3220 = (inp[6]) ? node3228 : node3221;
										assign node3221 = (inp[3]) ? node3225 : node3222;
											assign node3222 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3225 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3228 = (inp[11]) ? node3232 : node3229;
											assign node3229 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3232 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node3235 = (inp[13]) ? node3251 : node3236;
									assign node3236 = (inp[5]) ? node3244 : node3237;
										assign node3237 = (inp[11]) ? node3241 : node3238;
											assign node3238 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3241 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3244 = (inp[14]) ? node3248 : node3245;
											assign node3245 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3248 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3251 = (inp[3]) ? node3259 : node3252;
										assign node3252 = (inp[11]) ? node3256 : node3253;
											assign node3253 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3256 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3259 = (inp[5]) ? node3263 : node3260;
											assign node3260 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3263 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node3266 = (inp[6]) ? node3298 : node3267;
								assign node3267 = (inp[5]) ? node3283 : node3268;
									assign node3268 = (inp[3]) ? node3276 : node3269;
										assign node3269 = (inp[11]) ? node3273 : node3270;
											assign node3270 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3273 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3276 = (inp[13]) ? node3280 : node3277;
											assign node3277 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3280 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3283 = (inp[14]) ? node3291 : node3284;
										assign node3284 = (inp[12]) ? node3288 : node3285;
											assign node3285 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3288 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3291 = (inp[13]) ? node3295 : node3292;
											assign node3292 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3295 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node3298 = (inp[11]) ? node3314 : node3299;
									assign node3299 = (inp[0]) ? node3307 : node3300;
										assign node3300 = (inp[13]) ? node3304 : node3301;
											assign node3301 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3304 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3307 = (inp[1]) ? node3311 : node3308;
											assign node3308 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3311 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3314 = (inp[1]) ? node3322 : node3315;
										assign node3315 = (inp[12]) ? node3319 : node3316;
											assign node3316 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3319 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3322 = (inp[13]) ? node3326 : node3323;
											assign node3323 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3326 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
					assign node3329 = (inp[3]) ? node3457 : node3330;
						assign node3330 = (inp[12]) ? node3394 : node3331;
							assign node3331 = (inp[14]) ? node3363 : node3332;
								assign node3332 = (inp[0]) ? node3348 : node3333;
									assign node3333 = (inp[11]) ? node3341 : node3334;
										assign node3334 = (inp[1]) ? node3338 : node3335;
											assign node3335 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3338 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3341 = (inp[5]) ? node3345 : node3342;
											assign node3342 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3345 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node3348 = (inp[2]) ? node3356 : node3349;
										assign node3349 = (inp[8]) ? node3353 : node3350;
											assign node3350 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3353 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3356 = (inp[11]) ? node3360 : node3357;
											assign node3357 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3360 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node3363 = (inp[2]) ? node3379 : node3364;
									assign node3364 = (inp[8]) ? node3372 : node3365;
										assign node3365 = (inp[13]) ? node3369 : node3366;
											assign node3366 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3369 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3372 = (inp[13]) ? node3376 : node3373;
											assign node3373 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3376 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3379 = (inp[5]) ? node3387 : node3380;
										assign node3380 = (inp[6]) ? node3384 : node3381;
											assign node3381 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3384 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3387 = (inp[13]) ? node3391 : node3388;
											assign node3388 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3391 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node3394 = (inp[13]) ? node3426 : node3395;
								assign node3395 = (inp[8]) ? node3411 : node3396;
									assign node3396 = (inp[14]) ? node3404 : node3397;
										assign node3397 = (inp[0]) ? node3401 : node3398;
											assign node3398 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3401 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3404 = (inp[2]) ? node3408 : node3405;
											assign node3405 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3408 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3411 = (inp[5]) ? node3419 : node3412;
										assign node3412 = (inp[14]) ? node3416 : node3413;
											assign node3413 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3416 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3419 = (inp[6]) ? node3423 : node3420;
											assign node3420 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3423 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node3426 = (inp[0]) ? node3442 : node3427;
									assign node3427 = (inp[8]) ? node3435 : node3428;
										assign node3428 = (inp[11]) ? node3432 : node3429;
											assign node3429 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3432 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3435 = (inp[2]) ? node3439 : node3436;
											assign node3436 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3439 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3442 = (inp[1]) ? node3450 : node3443;
										assign node3443 = (inp[5]) ? node3447 : node3444;
											assign node3444 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3447 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3450 = (inp[14]) ? node3454 : node3451;
											assign node3451 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3454 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node3457 = (inp[12]) ? node3521 : node3458;
							assign node3458 = (inp[5]) ? node3490 : node3459;
								assign node3459 = (inp[14]) ? node3475 : node3460;
									assign node3460 = (inp[1]) ? node3468 : node3461;
										assign node3461 = (inp[11]) ? node3465 : node3462;
											assign node3462 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3465 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3468 = (inp[6]) ? node3472 : node3469;
											assign node3469 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3472 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3475 = (inp[1]) ? node3483 : node3476;
										assign node3476 = (inp[8]) ? node3480 : node3477;
											assign node3477 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3480 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3483 = (inp[6]) ? node3487 : node3484;
											assign node3484 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3487 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node3490 = (inp[8]) ? node3506 : node3491;
									assign node3491 = (inp[14]) ? node3499 : node3492;
										assign node3492 = (inp[11]) ? node3496 : node3493;
											assign node3493 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3496 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3499 = (inp[1]) ? node3503 : node3500;
											assign node3500 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3503 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3506 = (inp[11]) ? node3514 : node3507;
										assign node3507 = (inp[6]) ? node3511 : node3508;
											assign node3508 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3511 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3514 = (inp[13]) ? node3518 : node3515;
											assign node3515 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3518 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node3521 = (inp[6]) ? node3553 : node3522;
								assign node3522 = (inp[14]) ? node3538 : node3523;
									assign node3523 = (inp[11]) ? node3531 : node3524;
										assign node3524 = (inp[1]) ? node3528 : node3525;
											assign node3525 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3528 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3531 = (inp[13]) ? node3535 : node3532;
											assign node3532 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3535 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3538 = (inp[1]) ? node3546 : node3539;
										assign node3539 = (inp[0]) ? node3543 : node3540;
											assign node3540 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3543 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3546 = (inp[2]) ? node3550 : node3547;
											assign node3547 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3550 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node3553 = (inp[13]) ? node3569 : node3554;
									assign node3554 = (inp[14]) ? node3562 : node3555;
										assign node3555 = (inp[5]) ? node3559 : node3556;
											assign node3556 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3559 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3562 = (inp[11]) ? node3566 : node3563;
											assign node3563 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3566 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node3569 = (inp[0]) ? node3577 : node3570;
										assign node3570 = (inp[5]) ? node3574 : node3571;
											assign node3571 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3574 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node3577 = (inp[14]) ? node3581 : node3578;
											assign node3578 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node3581 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
				assign node3584 = (inp[11]) ? node3840 : node3585;
					assign node3585 = (inp[14]) ? node3713 : node3586;
						assign node3586 = (inp[12]) ? node3650 : node3587;
							assign node3587 = (inp[0]) ? node3619 : node3588;
								assign node3588 = (inp[8]) ? node3604 : node3589;
									assign node3589 = (inp[3]) ? node3597 : node3590;
										assign node3590 = (inp[2]) ? node3594 : node3591;
											assign node3591 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3594 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3597 = (inp[1]) ? node3601 : node3598;
											assign node3598 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3601 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node3604 = (inp[5]) ? node3612 : node3605;
										assign node3605 = (inp[13]) ? node3609 : node3606;
											assign node3606 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3609 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3612 = (inp[2]) ? node3616 : node3613;
											assign node3613 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3616 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node3619 = (inp[6]) ? node3635 : node3620;
									assign node3620 = (inp[3]) ? node3628 : node3621;
										assign node3621 = (inp[1]) ? node3625 : node3622;
											assign node3622 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3625 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3628 = (inp[5]) ? node3632 : node3629;
											assign node3629 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3632 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3635 = (inp[2]) ? node3643 : node3636;
										assign node3636 = (inp[5]) ? node3640 : node3637;
											assign node3637 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3640 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3643 = (inp[1]) ? node3647 : node3644;
											assign node3644 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3647 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node3650 = (inp[3]) ? node3682 : node3651;
								assign node3651 = (inp[8]) ? node3667 : node3652;
									assign node3652 = (inp[5]) ? node3660 : node3653;
										assign node3653 = (inp[1]) ? node3657 : node3654;
											assign node3654 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3657 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3660 = (inp[13]) ? node3664 : node3661;
											assign node3661 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3664 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3667 = (inp[10]) ? node3675 : node3668;
										assign node3668 = (inp[2]) ? node3672 : node3669;
											assign node3669 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3672 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3675 = (inp[13]) ? node3679 : node3676;
											assign node3676 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3679 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node3682 = (inp[8]) ? node3698 : node3683;
									assign node3683 = (inp[1]) ? node3691 : node3684;
										assign node3684 = (inp[2]) ? node3688 : node3685;
											assign node3685 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3688 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3691 = (inp[13]) ? node3695 : node3692;
											assign node3692 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3695 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3698 = (inp[5]) ? node3706 : node3699;
										assign node3699 = (inp[6]) ? node3703 : node3700;
											assign node3700 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3703 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3706 = (inp[10]) ? node3710 : node3707;
											assign node3707 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3710 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node3713 = (inp[0]) ? node3777 : node3714;
							assign node3714 = (inp[10]) ? node3746 : node3715;
								assign node3715 = (inp[6]) ? node3731 : node3716;
									assign node3716 = (inp[13]) ? node3724 : node3717;
										assign node3717 = (inp[5]) ? node3721 : node3718;
											assign node3718 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3721 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3724 = (inp[2]) ? node3728 : node3725;
											assign node3725 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3728 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3731 = (inp[3]) ? node3739 : node3732;
										assign node3732 = (inp[5]) ? node3736 : node3733;
											assign node3733 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3736 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3739 = (inp[5]) ? node3743 : node3740;
											assign node3740 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3743 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node3746 = (inp[3]) ? node3762 : node3747;
									assign node3747 = (inp[13]) ? node3755 : node3748;
										assign node3748 = (inp[1]) ? node3752 : node3749;
											assign node3749 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3752 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3755 = (inp[2]) ? node3759 : node3756;
											assign node3756 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3759 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3762 = (inp[2]) ? node3770 : node3763;
										assign node3763 = (inp[8]) ? node3767 : node3764;
											assign node3764 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3767 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3770 = (inp[12]) ? node3774 : node3771;
											assign node3771 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3774 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node3777 = (inp[8]) ? node3809 : node3778;
								assign node3778 = (inp[5]) ? node3794 : node3779;
									assign node3779 = (inp[10]) ? node3787 : node3780;
										assign node3780 = (inp[3]) ? node3784 : node3781;
											assign node3781 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3784 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3787 = (inp[12]) ? node3791 : node3788;
											assign node3788 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3791 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3794 = (inp[2]) ? node3802 : node3795;
										assign node3795 = (inp[6]) ? node3799 : node3796;
											assign node3796 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3799 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3802 = (inp[13]) ? node3806 : node3803;
											assign node3803 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3806 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node3809 = (inp[10]) ? node3825 : node3810;
									assign node3810 = (inp[12]) ? node3818 : node3811;
										assign node3811 = (inp[5]) ? node3815 : node3812;
											assign node3812 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3815 = (inp[2]) ? 15'b000000000001111 : 15'b000000000111111;
										assign node3818 = (inp[1]) ? node3822 : node3819;
											assign node3819 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3822 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node3825 = (inp[5]) ? node3833 : node3826;
										assign node3826 = (inp[6]) ? node3830 : node3827;
											assign node3827 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3830 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node3833 = (inp[6]) ? node3837 : node3834;
											assign node3834 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node3837 = (inp[12]) ? 15'b000000000000111 : 15'b000000000001111;
					assign node3840 = (inp[0]) ? node3968 : node3841;
						assign node3841 = (inp[1]) ? node3905 : node3842;
							assign node3842 = (inp[14]) ? node3874 : node3843;
								assign node3843 = (inp[2]) ? node3859 : node3844;
									assign node3844 = (inp[3]) ? node3852 : node3845;
										assign node3845 = (inp[6]) ? node3849 : node3846;
											assign node3846 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3849 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3852 = (inp[8]) ? node3856 : node3853;
											assign node3853 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3856 = (inp[6]) ? 15'b000000000011111 : 15'b000000001111111;
									assign node3859 = (inp[12]) ? node3867 : node3860;
										assign node3860 = (inp[6]) ? node3864 : node3861;
											assign node3861 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3864 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3867 = (inp[3]) ? node3871 : node3868;
											assign node3868 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3871 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node3874 = (inp[5]) ? node3890 : node3875;
									assign node3875 = (inp[10]) ? node3883 : node3876;
										assign node3876 = (inp[2]) ? node3880 : node3877;
											assign node3877 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3880 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3883 = (inp[12]) ? node3887 : node3884;
											assign node3884 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3887 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3890 = (inp[3]) ? node3898 : node3891;
										assign node3891 = (inp[2]) ? node3895 : node3892;
											assign node3892 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3895 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3898 = (inp[13]) ? node3902 : node3899;
											assign node3899 = (inp[12]) ? 15'b000000000001111 : 15'b000000000111111;
											assign node3902 = (inp[2]) ? 15'b000000000000111 : 15'b000000000011111;
							assign node3905 = (inp[2]) ? node3937 : node3906;
								assign node3906 = (inp[6]) ? node3922 : node3907;
									assign node3907 = (inp[12]) ? node3915 : node3908;
										assign node3908 = (inp[13]) ? node3912 : node3909;
											assign node3909 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3912 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3915 = (inp[10]) ? node3919 : node3916;
											assign node3916 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3919 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3922 = (inp[12]) ? node3930 : node3923;
										assign node3923 = (inp[14]) ? node3927 : node3924;
											assign node3924 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3927 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3930 = (inp[3]) ? node3934 : node3931;
											assign node3931 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3934 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node3937 = (inp[8]) ? node3953 : node3938;
									assign node3938 = (inp[5]) ? node3946 : node3939;
										assign node3939 = (inp[14]) ? node3943 : node3940;
											assign node3940 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3943 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3946 = (inp[10]) ? node3950 : node3947;
											assign node3947 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3950 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node3953 = (inp[6]) ? node3961 : node3954;
										assign node3954 = (inp[10]) ? node3958 : node3955;
											assign node3955 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3958 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node3961 = (inp[12]) ? node3965 : node3962;
											assign node3962 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node3965 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node3968 = (inp[10]) ? node4032 : node3969;
							assign node3969 = (inp[1]) ? node4001 : node3970;
								assign node3970 = (inp[8]) ? node3986 : node3971;
									assign node3971 = (inp[5]) ? node3979 : node3972;
										assign node3972 = (inp[13]) ? node3976 : node3973;
											assign node3973 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3976 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3979 = (inp[2]) ? node3983 : node3980;
											assign node3980 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3983 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3986 = (inp[13]) ? node3994 : node3987;
										assign node3987 = (inp[2]) ? node3991 : node3988;
											assign node3988 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3991 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node3994 = (inp[2]) ? node3998 : node3995;
											assign node3995 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3998 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node4001 = (inp[3]) ? node4017 : node4002;
									assign node4002 = (inp[13]) ? node4010 : node4003;
										assign node4003 = (inp[2]) ? node4007 : node4004;
											assign node4004 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4007 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node4010 = (inp[6]) ? node4014 : node4011;
											assign node4011 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4014 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node4017 = (inp[8]) ? node4025 : node4018;
										assign node4018 = (inp[6]) ? node4022 : node4019;
											assign node4019 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4022 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node4025 = (inp[14]) ? node4029 : node4026;
											assign node4026 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node4029 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
							assign node4032 = (inp[12]) ? node4064 : node4033;
								assign node4033 = (inp[13]) ? node4049 : node4034;
									assign node4034 = (inp[1]) ? node4042 : node4035;
										assign node4035 = (inp[8]) ? node4039 : node4036;
											assign node4036 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4039 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node4042 = (inp[6]) ? node4046 : node4043;
											assign node4043 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4046 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node4049 = (inp[5]) ? node4057 : node4050;
										assign node4050 = (inp[3]) ? node4054 : node4051;
											assign node4051 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4054 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node4057 = (inp[6]) ? node4061 : node4058;
											assign node4058 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node4061 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node4064 = (inp[8]) ? node4080 : node4065;
									assign node4065 = (inp[13]) ? node4073 : node4066;
										assign node4066 = (inp[3]) ? node4070 : node4067;
											assign node4067 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4070 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node4073 = (inp[2]) ? node4077 : node4074;
											assign node4074 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node4077 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node4080 = (inp[14]) ? node4088 : node4081;
										assign node4081 = (inp[2]) ? node4085 : node4082;
											assign node4082 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node4085 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node4088 = (inp[2]) ? node4092 : node4089;
											assign node4089 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node4092 = (inp[6]) ? 15'b000000000000011 : 15'b000000000000111;

endmodule