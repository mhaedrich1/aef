module dtc_split66_bm45 (
	input  wire [16-1:0] inp,
	output wire [46-1:0] outp
);

	wire [46-1:0] node1;
	wire [46-1:0] node2;
	wire [46-1:0] node4;
	wire [46-1:0] node5;
	wire [46-1:0] node7;
	wire [46-1:0] node9;
	wire [46-1:0] node11;
	wire [46-1:0] node13;
	wire [46-1:0] node14;
	wire [46-1:0] node15;
	wire [46-1:0] node17;
	wire [46-1:0] node22;
	wire [46-1:0] node24;
	wire [46-1:0] node26;
	wire [46-1:0] node27;
	wire [46-1:0] node29;
	wire [46-1:0] node31;
	wire [46-1:0] node33;
	wire [46-1:0] node34;
	wire [46-1:0] node36;
	wire [46-1:0] node38;
	wire [46-1:0] node41;
	wire [46-1:0] node42;
	wire [46-1:0] node44;
	wire [46-1:0] node48;
	wire [46-1:0] node50;
	wire [46-1:0] node52;
	wire [46-1:0] node54;
	wire [46-1:0] node56;
	wire [46-1:0] node58;
	wire [46-1:0] node60;
	wire [46-1:0] node63;
	wire [46-1:0] node65;
	wire [46-1:0] node66;
	wire [46-1:0] node67;
	wire [46-1:0] node68;
	wire [46-1:0] node69;
	wire [46-1:0] node72;
	wire [46-1:0] node74;
	wire [46-1:0] node76;
	wire [46-1:0] node78;
	wire [46-1:0] node79;
	wire [46-1:0] node81;
	wire [46-1:0] node82;
	wire [46-1:0] node85;
	wire [46-1:0] node89;
	wire [46-1:0] node90;
	wire [46-1:0] node92;
	wire [46-1:0] node94;
	wire [46-1:0] node96;
	wire [46-1:0] node98;
	wire [46-1:0] node99;
	wire [46-1:0] node101;
	wire [46-1:0] node104;
	wire [46-1:0] node105;
	wire [46-1:0] node108;
	wire [46-1:0] node112;
	wire [46-1:0] node113;
	wire [46-1:0] node114;
	wire [46-1:0] node118;
	wire [46-1:0] node119;
	wire [46-1:0] node122;
	wire [46-1:0] node125;
	wire [46-1:0] node126;
	wire [46-1:0] node127;
	wire [46-1:0] node128;
	wire [46-1:0] node131;
	wire [46-1:0] node133;
	wire [46-1:0] node135;
	wire [46-1:0] node136;
	wire [46-1:0] node138;
	wire [46-1:0] node140;
	wire [46-1:0] node142;
	wire [46-1:0] node145;
	wire [46-1:0] node146;
	wire [46-1:0] node148;
	wire [46-1:0] node150;
	wire [46-1:0] node153;
	wire [46-1:0] node154;
	wire [46-1:0] node156;
	wire [46-1:0] node159;
	wire [46-1:0] node160;
	wire [46-1:0] node164;
	wire [46-1:0] node165;
	wire [46-1:0] node167;
	wire [46-1:0] node169;
	wire [46-1:0] node171;
	wire [46-1:0] node172;
	wire [46-1:0] node174;
	wire [46-1:0] node175;
	wire [46-1:0] node178;
	wire [46-1:0] node182;
	wire [46-1:0] node184;
	wire [46-1:0] node186;
	wire [46-1:0] node188;
	wire [46-1:0] node189;
	wire [46-1:0] node191;
	wire [46-1:0] node193;
	wire [46-1:0] node196;
	wire [46-1:0] node197;
	wire [46-1:0] node199;
	wire [46-1:0] node202;
	wire [46-1:0] node203;
	wire [46-1:0] node206;
	wire [46-1:0] node209;
	wire [46-1:0] node211;
	wire [46-1:0] node213;
	wire [46-1:0] node215;
	wire [46-1:0] node216;
	wire [46-1:0] node218;
	wire [46-1:0] node220;
	wire [46-1:0] node222;
	wire [46-1:0] node224;
	wire [46-1:0] node227;
	wire [46-1:0] node228;
	wire [46-1:0] node230;
	wire [46-1:0] node232;
	wire [46-1:0] node233;
	wire [46-1:0] node236;
	wire [46-1:0] node239;
	wire [46-1:0] node240;
	wire [46-1:0] node241;
	wire [46-1:0] node242;
	wire [46-1:0] node245;
	wire [46-1:0] node249;
	wire [46-1:0] node250;
	wire [46-1:0] node251;
	wire [46-1:0] node254;
	wire [46-1:0] node257;
	wire [46-1:0] node258;
	wire [46-1:0] node262;
	wire [46-1:0] node263;
	wire [46-1:0] node264;
	wire [46-1:0] node267;
	wire [46-1:0] node268;
	wire [46-1:0] node269;
	wire [46-1:0] node270;
	wire [46-1:0] node271;
	wire [46-1:0] node274;
	wire [46-1:0] node277;
	wire [46-1:0] node278;
	wire [46-1:0] node281;
	wire [46-1:0] node284;
	wire [46-1:0] node285;
	wire [46-1:0] node286;
	wire [46-1:0] node289;
	wire [46-1:0] node292;
	wire [46-1:0] node293;
	wire [46-1:0] node296;
	wire [46-1:0] node299;
	wire [46-1:0] node300;
	wire [46-1:0] node301;
	wire [46-1:0] node302;
	wire [46-1:0] node305;
	wire [46-1:0] node308;
	wire [46-1:0] node309;
	wire [46-1:0] node312;
	wire [46-1:0] node315;
	wire [46-1:0] node316;
	wire [46-1:0] node317;
	wire [46-1:0] node320;
	wire [46-1:0] node323;
	wire [46-1:0] node324;
	wire [46-1:0] node327;
	wire [46-1:0] node330;
	wire [46-1:0] node331;
	wire [46-1:0] node334;
	wire [46-1:0] node336;
	wire [46-1:0] node337;
	wire [46-1:0] node338;
	wire [46-1:0] node339;
	wire [46-1:0] node340;
	wire [46-1:0] node341;
	wire [46-1:0] node342;
	wire [46-1:0] node343;
	wire [46-1:0] node344;
	wire [46-1:0] node345;
	wire [46-1:0] node348;
	wire [46-1:0] node351;
	wire [46-1:0] node352;
	wire [46-1:0] node355;
	wire [46-1:0] node358;
	wire [46-1:0] node359;
	wire [46-1:0] node360;
	wire [46-1:0] node363;
	wire [46-1:0] node366;
	wire [46-1:0] node367;
	wire [46-1:0] node370;
	wire [46-1:0] node373;
	wire [46-1:0] node374;
	wire [46-1:0] node375;
	wire [46-1:0] node376;
	wire [46-1:0] node379;
	wire [46-1:0] node382;
	wire [46-1:0] node383;
	wire [46-1:0] node386;
	wire [46-1:0] node389;
	wire [46-1:0] node390;
	wire [46-1:0] node391;
	wire [46-1:0] node394;
	wire [46-1:0] node397;
	wire [46-1:0] node398;
	wire [46-1:0] node401;
	wire [46-1:0] node404;
	wire [46-1:0] node405;
	wire [46-1:0] node406;
	wire [46-1:0] node407;
	wire [46-1:0] node408;
	wire [46-1:0] node411;
	wire [46-1:0] node414;
	wire [46-1:0] node415;
	wire [46-1:0] node419;
	wire [46-1:0] node420;
	wire [46-1:0] node421;
	wire [46-1:0] node424;
	wire [46-1:0] node427;
	wire [46-1:0] node428;
	wire [46-1:0] node431;
	wire [46-1:0] node434;
	wire [46-1:0] node435;
	wire [46-1:0] node436;
	wire [46-1:0] node437;
	wire [46-1:0] node440;
	wire [46-1:0] node443;
	wire [46-1:0] node444;
	wire [46-1:0] node447;
	wire [46-1:0] node450;
	wire [46-1:0] node451;
	wire [46-1:0] node452;
	wire [46-1:0] node455;
	wire [46-1:0] node458;
	wire [46-1:0] node459;
	wire [46-1:0] node462;
	wire [46-1:0] node465;
	wire [46-1:0] node466;
	wire [46-1:0] node467;
	wire [46-1:0] node468;
	wire [46-1:0] node469;
	wire [46-1:0] node470;
	wire [46-1:0] node473;
	wire [46-1:0] node476;
	wire [46-1:0] node477;
	wire [46-1:0] node480;
	wire [46-1:0] node483;
	wire [46-1:0] node484;
	wire [46-1:0] node485;
	wire [46-1:0] node488;
	wire [46-1:0] node491;
	wire [46-1:0] node492;
	wire [46-1:0] node495;
	wire [46-1:0] node498;
	wire [46-1:0] node499;
	wire [46-1:0] node500;
	wire [46-1:0] node501;
	wire [46-1:0] node504;
	wire [46-1:0] node507;
	wire [46-1:0] node508;
	wire [46-1:0] node511;
	wire [46-1:0] node514;
	wire [46-1:0] node515;
	wire [46-1:0] node516;
	wire [46-1:0] node519;
	wire [46-1:0] node522;
	wire [46-1:0] node523;
	wire [46-1:0] node526;
	wire [46-1:0] node529;
	wire [46-1:0] node530;
	wire [46-1:0] node531;
	wire [46-1:0] node532;
	wire [46-1:0] node533;
	wire [46-1:0] node536;
	wire [46-1:0] node539;
	wire [46-1:0] node540;
	wire [46-1:0] node543;
	wire [46-1:0] node546;
	wire [46-1:0] node547;
	wire [46-1:0] node548;
	wire [46-1:0] node551;
	wire [46-1:0] node554;
	wire [46-1:0] node555;
	wire [46-1:0] node558;
	wire [46-1:0] node561;
	wire [46-1:0] node562;
	wire [46-1:0] node563;
	wire [46-1:0] node564;
	wire [46-1:0] node567;
	wire [46-1:0] node570;
	wire [46-1:0] node571;
	wire [46-1:0] node574;
	wire [46-1:0] node577;
	wire [46-1:0] node578;
	wire [46-1:0] node579;
	wire [46-1:0] node582;
	wire [46-1:0] node585;
	wire [46-1:0] node586;
	wire [46-1:0] node589;
	wire [46-1:0] node592;
	wire [46-1:0] node593;
	wire [46-1:0] node594;
	wire [46-1:0] node595;
	wire [46-1:0] node597;
	wire [46-1:0] node598;
	wire [46-1:0] node600;
	wire [46-1:0] node603;
	wire [46-1:0] node604;
	wire [46-1:0] node607;
	wire [46-1:0] node610;
	wire [46-1:0] node611;
	wire [46-1:0] node612;
	wire [46-1:0] node613;
	wire [46-1:0] node616;
	wire [46-1:0] node619;
	wire [46-1:0] node620;
	wire [46-1:0] node625;
	wire [46-1:0] node626;
	wire [46-1:0] node627;
	wire [46-1:0] node628;
	wire [46-1:0] node630;
	wire [46-1:0] node634;
	wire [46-1:0] node636;
	wire [46-1:0] node637;
	wire [46-1:0] node643;
	wire [46-1:0] node644;
	wire [46-1:0] node645;
	wire [46-1:0] node647;
	wire [46-1:0] node649;
	wire [46-1:0] node650;
	wire [46-1:0] node652;
	wire [46-1:0] node653;
	wire [46-1:0] node656;
	wire [46-1:0] node659;
	wire [46-1:0] node660;
	wire [46-1:0] node661;
	wire [46-1:0] node664;
	wire [46-1:0] node668;
	wire [46-1:0] node669;
	wire [46-1:0] node670;
	wire [46-1:0] node671;
	wire [46-1:0] node672;
	wire [46-1:0] node673;
	wire [46-1:0] node676;
	wire [46-1:0] node679;
	wire [46-1:0] node680;
	wire [46-1:0] node683;
	wire [46-1:0] node686;
	wire [46-1:0] node687;
	wire [46-1:0] node688;
	wire [46-1:0] node691;
	wire [46-1:0] node694;
	wire [46-1:0] node695;
	wire [46-1:0] node698;
	wire [46-1:0] node701;
	wire [46-1:0] node702;
	wire [46-1:0] node703;
	wire [46-1:0] node704;
	wire [46-1:0] node707;
	wire [46-1:0] node710;
	wire [46-1:0] node711;
	wire [46-1:0] node714;
	wire [46-1:0] node717;
	wire [46-1:0] node718;
	wire [46-1:0] node719;
	wire [46-1:0] node722;
	wire [46-1:0] node725;
	wire [46-1:0] node726;
	wire [46-1:0] node729;
	wire [46-1:0] node732;
	wire [46-1:0] node733;
	wire [46-1:0] node734;
	wire [46-1:0] node735;
	wire [46-1:0] node736;
	wire [46-1:0] node739;
	wire [46-1:0] node742;
	wire [46-1:0] node743;
	wire [46-1:0] node746;
	wire [46-1:0] node749;
	wire [46-1:0] node750;
	wire [46-1:0] node751;
	wire [46-1:0] node754;
	wire [46-1:0] node757;
	wire [46-1:0] node758;
	wire [46-1:0] node761;
	wire [46-1:0] node764;
	wire [46-1:0] node765;
	wire [46-1:0] node766;
	wire [46-1:0] node767;
	wire [46-1:0] node770;
	wire [46-1:0] node773;
	wire [46-1:0] node774;
	wire [46-1:0] node777;
	wire [46-1:0] node780;
	wire [46-1:0] node781;
	wire [46-1:0] node782;
	wire [46-1:0] node785;
	wire [46-1:0] node788;
	wire [46-1:0] node789;
	wire [46-1:0] node792;
	wire [46-1:0] node795;
	wire [46-1:0] node796;
	wire [46-1:0] node797;
	wire [46-1:0] node798;
	wire [46-1:0] node799;
	wire [46-1:0] node800;
	wire [46-1:0] node801;
	wire [46-1:0] node804;
	wire [46-1:0] node807;
	wire [46-1:0] node808;
	wire [46-1:0] node811;
	wire [46-1:0] node814;
	wire [46-1:0] node815;
	wire [46-1:0] node816;
	wire [46-1:0] node819;
	wire [46-1:0] node822;
	wire [46-1:0] node823;
	wire [46-1:0] node826;
	wire [46-1:0] node829;
	wire [46-1:0] node830;
	wire [46-1:0] node831;
	wire [46-1:0] node832;
	wire [46-1:0] node835;
	wire [46-1:0] node838;
	wire [46-1:0] node839;
	wire [46-1:0] node842;
	wire [46-1:0] node845;
	wire [46-1:0] node846;
	wire [46-1:0] node847;
	wire [46-1:0] node850;
	wire [46-1:0] node853;
	wire [46-1:0] node854;
	wire [46-1:0] node857;
	wire [46-1:0] node860;
	wire [46-1:0] node861;
	wire [46-1:0] node862;
	wire [46-1:0] node863;
	wire [46-1:0] node864;
	wire [46-1:0] node867;
	wire [46-1:0] node870;
	wire [46-1:0] node871;
	wire [46-1:0] node874;
	wire [46-1:0] node877;
	wire [46-1:0] node878;
	wire [46-1:0] node879;
	wire [46-1:0] node882;
	wire [46-1:0] node885;
	wire [46-1:0] node886;
	wire [46-1:0] node889;
	wire [46-1:0] node892;
	wire [46-1:0] node893;
	wire [46-1:0] node894;
	wire [46-1:0] node895;
	wire [46-1:0] node898;
	wire [46-1:0] node901;
	wire [46-1:0] node902;
	wire [46-1:0] node905;
	wire [46-1:0] node908;
	wire [46-1:0] node909;
	wire [46-1:0] node910;
	wire [46-1:0] node913;
	wire [46-1:0] node916;
	wire [46-1:0] node917;
	wire [46-1:0] node920;
	wire [46-1:0] node923;
	wire [46-1:0] node924;
	wire [46-1:0] node925;
	wire [46-1:0] node926;
	wire [46-1:0] node927;
	wire [46-1:0] node928;
	wire [46-1:0] node931;
	wire [46-1:0] node934;
	wire [46-1:0] node935;
	wire [46-1:0] node938;
	wire [46-1:0] node941;
	wire [46-1:0] node942;
	wire [46-1:0] node943;
	wire [46-1:0] node946;
	wire [46-1:0] node949;
	wire [46-1:0] node950;
	wire [46-1:0] node953;
	wire [46-1:0] node956;
	wire [46-1:0] node957;
	wire [46-1:0] node958;
	wire [46-1:0] node959;
	wire [46-1:0] node962;
	wire [46-1:0] node965;
	wire [46-1:0] node966;
	wire [46-1:0] node969;
	wire [46-1:0] node972;
	wire [46-1:0] node973;
	wire [46-1:0] node974;
	wire [46-1:0] node977;
	wire [46-1:0] node980;
	wire [46-1:0] node981;
	wire [46-1:0] node984;
	wire [46-1:0] node987;
	wire [46-1:0] node988;
	wire [46-1:0] node989;
	wire [46-1:0] node990;
	wire [46-1:0] node991;
	wire [46-1:0] node994;
	wire [46-1:0] node997;
	wire [46-1:0] node998;
	wire [46-1:0] node1001;
	wire [46-1:0] node1004;
	wire [46-1:0] node1005;
	wire [46-1:0] node1006;
	wire [46-1:0] node1009;
	wire [46-1:0] node1012;
	wire [46-1:0] node1013;
	wire [46-1:0] node1017;
	wire [46-1:0] node1018;
	wire [46-1:0] node1019;
	wire [46-1:0] node1020;
	wire [46-1:0] node1023;
	wire [46-1:0] node1026;
	wire [46-1:0] node1027;
	wire [46-1:0] node1030;
	wire [46-1:0] node1033;
	wire [46-1:0] node1034;
	wire [46-1:0] node1035;
	wire [46-1:0] node1038;
	wire [46-1:0] node1041;
	wire [46-1:0] node1042;
	wire [46-1:0] node1045;
	wire [46-1:0] node1048;
	wire [46-1:0] node1049;
	wire [46-1:0] node1050;
	wire [46-1:0] node1051;
	wire [46-1:0] node1053;
	wire [46-1:0] node1055;
	wire [46-1:0] node1057;
	wire [46-1:0] node1059;
	wire [46-1:0] node1060;
	wire [46-1:0] node1063;
	wire [46-1:0] node1066;
	wire [46-1:0] node1067;
	wire [46-1:0] node1069;
	wire [46-1:0] node1071;
	wire [46-1:0] node1073;
	wire [46-1:0] node1074;
	wire [46-1:0] node1077;
	wire [46-1:0] node1080;
	wire [46-1:0] node1081;
	wire [46-1:0] node1082;
	wire [46-1:0] node1083;
	wire [46-1:0] node1084;
	wire [46-1:0] node1087;
	wire [46-1:0] node1090;
	wire [46-1:0] node1091;
	wire [46-1:0] node1094;
	wire [46-1:0] node1097;
	wire [46-1:0] node1098;
	wire [46-1:0] node1099;
	wire [46-1:0] node1102;
	wire [46-1:0] node1105;
	wire [46-1:0] node1106;
	wire [46-1:0] node1109;
	wire [46-1:0] node1112;
	wire [46-1:0] node1113;
	wire [46-1:0] node1115;
	wire [46-1:0] node1116;
	wire [46-1:0] node1119;
	wire [46-1:0] node1122;
	wire [46-1:0] node1123;
	wire [46-1:0] node1124;
	wire [46-1:0] node1127;
	wire [46-1:0] node1131;
	wire [46-1:0] node1132;
	wire [46-1:0] node1133;
	wire [46-1:0] node1134;
	wire [46-1:0] node1135;
	wire [46-1:0] node1136;
	wire [46-1:0] node1137;
	wire [46-1:0] node1140;
	wire [46-1:0] node1143;
	wire [46-1:0] node1144;
	wire [46-1:0] node1147;
	wire [46-1:0] node1150;
	wire [46-1:0] node1151;
	wire [46-1:0] node1152;
	wire [46-1:0] node1155;
	wire [46-1:0] node1158;
	wire [46-1:0] node1159;
	wire [46-1:0] node1162;
	wire [46-1:0] node1165;
	wire [46-1:0] node1166;
	wire [46-1:0] node1167;
	wire [46-1:0] node1168;
	wire [46-1:0] node1171;
	wire [46-1:0] node1174;
	wire [46-1:0] node1175;
	wire [46-1:0] node1178;
	wire [46-1:0] node1181;
	wire [46-1:0] node1182;
	wire [46-1:0] node1183;
	wire [46-1:0] node1186;
	wire [46-1:0] node1189;
	wire [46-1:0] node1190;
	wire [46-1:0] node1193;
	wire [46-1:0] node1196;
	wire [46-1:0] node1197;
	wire [46-1:0] node1198;
	wire [46-1:0] node1199;
	wire [46-1:0] node1200;
	wire [46-1:0] node1203;
	wire [46-1:0] node1206;
	wire [46-1:0] node1207;
	wire [46-1:0] node1210;
	wire [46-1:0] node1213;
	wire [46-1:0] node1214;
	wire [46-1:0] node1215;
	wire [46-1:0] node1218;
	wire [46-1:0] node1221;
	wire [46-1:0] node1222;
	wire [46-1:0] node1225;
	wire [46-1:0] node1228;
	wire [46-1:0] node1229;
	wire [46-1:0] node1230;
	wire [46-1:0] node1231;
	wire [46-1:0] node1234;
	wire [46-1:0] node1237;
	wire [46-1:0] node1238;
	wire [46-1:0] node1241;
	wire [46-1:0] node1244;
	wire [46-1:0] node1245;
	wire [46-1:0] node1246;
	wire [46-1:0] node1249;
	wire [46-1:0] node1252;
	wire [46-1:0] node1253;
	wire [46-1:0] node1256;
	wire [46-1:0] node1259;
	wire [46-1:0] node1260;
	wire [46-1:0] node1261;
	wire [46-1:0] node1262;
	wire [46-1:0] node1263;
	wire [46-1:0] node1264;
	wire [46-1:0] node1267;
	wire [46-1:0] node1270;
	wire [46-1:0] node1271;
	wire [46-1:0] node1274;
	wire [46-1:0] node1277;
	wire [46-1:0] node1278;
	wire [46-1:0] node1279;
	wire [46-1:0] node1282;
	wire [46-1:0] node1285;
	wire [46-1:0] node1286;
	wire [46-1:0] node1289;
	wire [46-1:0] node1292;
	wire [46-1:0] node1293;
	wire [46-1:0] node1294;
	wire [46-1:0] node1295;
	wire [46-1:0] node1298;
	wire [46-1:0] node1301;
	wire [46-1:0] node1302;
	wire [46-1:0] node1305;
	wire [46-1:0] node1308;
	wire [46-1:0] node1309;
	wire [46-1:0] node1310;
	wire [46-1:0] node1313;
	wire [46-1:0] node1316;
	wire [46-1:0] node1317;
	wire [46-1:0] node1320;
	wire [46-1:0] node1323;
	wire [46-1:0] node1324;
	wire [46-1:0] node1325;
	wire [46-1:0] node1326;
	wire [46-1:0] node1327;
	wire [46-1:0] node1330;
	wire [46-1:0] node1333;
	wire [46-1:0] node1334;
	wire [46-1:0] node1337;
	wire [46-1:0] node1340;
	wire [46-1:0] node1341;
	wire [46-1:0] node1342;
	wire [46-1:0] node1345;
	wire [46-1:0] node1348;
	wire [46-1:0] node1349;
	wire [46-1:0] node1352;
	wire [46-1:0] node1355;
	wire [46-1:0] node1356;
	wire [46-1:0] node1357;
	wire [46-1:0] node1358;
	wire [46-1:0] node1361;
	wire [46-1:0] node1364;
	wire [46-1:0] node1365;
	wire [46-1:0] node1368;
	wire [46-1:0] node1371;
	wire [46-1:0] node1372;
	wire [46-1:0] node1373;
	wire [46-1:0] node1376;
	wire [46-1:0] node1379;
	wire [46-1:0] node1380;
	wire [46-1:0] node1383;
	wire [46-1:0] node1386;
	wire [46-1:0] node1387;
	wire [46-1:0] node1388;
	wire [46-1:0] node1389;
	wire [46-1:0] node1390;
	wire [46-1:0] node1391;
	wire [46-1:0] node1394;
	wire [46-1:0] node1399;
	wire [46-1:0] node1400;
	wire [46-1:0] node1401;
	wire [46-1:0] node1402;
	wire [46-1:0] node1405;
	wire [46-1:0] node1408;
	wire [46-1:0] node1409;
	wire [46-1:0] node1412;
	wire [46-1:0] node1415;
	wire [46-1:0] node1416;
	wire [46-1:0] node1417;
	wire [46-1:0] node1420;
	wire [46-1:0] node1424;
	wire [46-1:0] node1425;
	wire [46-1:0] node1426;
	wire [46-1:0] node1427;
	wire [46-1:0] node1428;
	wire [46-1:0] node1431;
	wire [46-1:0] node1434;
	wire [46-1:0] node1435;
	wire [46-1:0] node1438;
	wire [46-1:0] node1441;
	wire [46-1:0] node1442;
	wire [46-1:0] node1443;
	wire [46-1:0] node1446;
	wire [46-1:0] node1450;
	wire [46-1:0] node1451;
	wire [46-1:0] node1452;
	wire [46-1:0] node1453;
	wire [46-1:0] node1456;

	assign outp = (inp[1]) ? node262 : node1;
		assign node1 = (inp[15]) ? node63 : node2;
			assign node2 = (inp[12]) ? node4 : 46'b0000000000000000000000000000000000000000000000;
				assign node4 = (inp[0]) ? node22 : node5;
					assign node5 = (inp[5]) ? node7 : 46'b0000000000000000000000000000000000000000000000;
						assign node7 = (inp[3]) ? node9 : 46'b0000000000000000000000000000000000000000000000;
							assign node9 = (inp[2]) ? node11 : 46'b0000000000000000000000000000000000000000000000;
								assign node11 = (inp[6]) ? node13 : 46'b0000000000000000000000000000000000000000000000;
									assign node13 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : node14;
										assign node14 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node15;
											assign node15 = (inp[13]) ? node17 : 46'b0000000000000000000000000000000000000000000000;
												assign node17 = (inp[7]) ? 46'b0000000000000000000000000000000000000100000000 : 46'b0000000000000000000000000000000000000000000000;
					assign node22 = (inp[7]) ? node24 : 46'b0000000000000000000000000000000000000000000000;
						assign node24 = (inp[6]) ? node26 : 46'b0000000000000000000000000000000000000000000000;
							assign node26 = (inp[13]) ? node48 : node27;
								assign node27 = (inp[4]) ? node29 : 46'b0000000000000000000000000000000000000000000000;
									assign node29 = (inp[9]) ? node31 : 46'b0000000000000000000000000000000000000000000000;
										assign node31 = (inp[10]) ? node33 : 46'b0000000000000000000000000000000000000000000000;
											assign node33 = (inp[11]) ? node41 : node34;
												assign node34 = (inp[8]) ? node36 : 46'b0000000000000000000000000000000000000000000000;
													assign node36 = (inp[14]) ? node38 : 46'b0000000000000000000000000000000000000000000000;
														assign node38 = (inp[3]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
												assign node41 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node42;
													assign node42 = (inp[8]) ? node44 : 46'b0000000000000000000000000000000000000000000000;
														assign node44 = (inp[14]) ? 46'b0000000000000000100000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
								assign node48 = (inp[2]) ? node50 : 46'b0000000000000000000000000000000000000000000000;
									assign node50 = (inp[3]) ? node52 : 46'b0000000000000000000000000000000000000000000000;
										assign node52 = (inp[10]) ? node54 : 46'b0000000000000000000000000000000000000000000000;
											assign node54 = (inp[14]) ? node56 : 46'b0000000000000000000000000000000000000000000000;
												assign node56 = (inp[4]) ? node58 : 46'b0000000000000000000000000000000000000000000000;
													assign node58 = (inp[8]) ? node60 : 46'b0000000000000000000000000000000000000000000000;
														assign node60 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000001000000000000000000000000000000000000;
			assign node63 = (inp[3]) ? node65 : 46'b0000000000000000000000000000001000000000000000;
				assign node65 = (inp[9]) ? node125 : node66;
					assign node66 = (inp[11]) ? node112 : node67;
						assign node67 = (inp[2]) ? node89 : node68;
							assign node68 = (inp[13]) ? node72 : node69;
								assign node69 = (inp[0]) ? 46'b0000000000001000000000000010000000000000000000 : 46'b0000001000001000000000000000000000000000000000;
								assign node72 = (inp[14]) ? node74 : 46'b0000000000000000000000000000000000000000000000;
									assign node74 = (inp[6]) ? node76 : 46'b0000000000000000000000000000000000000000000000;
										assign node76 = (inp[5]) ? node78 : 46'b0000000000000000000000000000000000000000000000;
											assign node78 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node79;
												assign node79 = (inp[10]) ? node81 : 46'b0000000000000000000000000000000000000000000000;
													assign node81 = (inp[12]) ? node85 : node82;
														assign node82 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
														assign node85 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000010000000000010100000000000000000000010000;
							assign node89 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node90;
								assign node90 = (inp[14]) ? node92 : 46'b0000000000000000000000000000000000000000000000;
									assign node92 = (inp[13]) ? node94 : 46'b0000000000000000000000000000000000000000000000;
										assign node94 = (inp[6]) ? node96 : 46'b0000000000000000000000000000000000000000000000;
											assign node96 = (inp[5]) ? node98 : 46'b0000000000000000000000000000000000000000000000;
												assign node98 = (inp[10]) ? node104 : node99;
													assign node99 = (inp[4]) ? node101 : 46'b0000000000000000000000000000000000000000000000;
														assign node101 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
													assign node104 = (inp[7]) ? node108 : node105;
														assign node105 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
														assign node108 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000001000010000000000000001000010000000;
						assign node112 = (inp[13]) ? node118 : node113;
							assign node113 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node114;
								assign node114 = (inp[0]) ? 46'b0000010000000000000000000010000000000000000000 : 46'b0000011000000000000000000000000000000000000000;
							assign node118 = (inp[2]) ? node122 : node119;
								assign node119 = (inp[0]) ? 46'b0000001000000000011000000100000000000000010000 : 46'b0000001000000000010000000100000000000000010010;
								assign node122 = (inp[0]) ? 46'b0000001000000000010010000000010000000010000000 : 46'b0000001000000000010010100000000000000010000000;
					assign node125 = (inp[2]) ? node209 : node126;
						assign node126 = (inp[0]) ? node164 : node127;
							assign node127 = (inp[13]) ? node131 : node128;
								assign node128 = (inp[11]) ? 46'b0000010100000000000000000000000000000000000000 : 46'b0000000100001000000000000000000000000000000000;
								assign node131 = (inp[5]) ? node133 : 46'b0000000000000000000000000000000000000000000000;
									assign node133 = (inp[14]) ? node135 : 46'b0000000000000000000000000000000000000000000000;
										assign node135 = (inp[6]) ? node145 : node136;
											assign node136 = (inp[4]) ? node138 : 46'b0000000000000000000000000000000000000000000000;
												assign node138 = (inp[10]) ? node140 : 46'b0000000000000000000000000000000000000000000000;
													assign node140 = (inp[8]) ? node142 : 46'b0000000000000000000000000000000000000000000000;
														assign node142 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
											assign node145 = (inp[10]) ? node153 : node146;
												assign node146 = (inp[4]) ? node148 : 46'b0000000000000000000000000000000000000000000000;
													assign node148 = (inp[8]) ? node150 : 46'b0000000000000000000000000000000000000000000000;
														assign node150 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000100000000010000;
												assign node153 = (inp[4]) ? node159 : node154;
													assign node154 = (inp[8]) ? node156 : 46'b0000000000000000000000000000000000000000000000;
														assign node156 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000010000000000010000010100000000000000010010;
													assign node159 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : node160;
														assign node160 = (inp[7]) ? 46'b0000000000011000010000000000000000000000010000 : 46'b0010000000010000000000000100000000000000010010;
							assign node164 = (inp[11]) ? node182 : node165;
								assign node165 = (inp[13]) ? node167 : 46'b0010001000000000000000000000000000000000010000;
									assign node167 = (inp[14]) ? node169 : 46'b0000000000000000000000000000000000000000000000;
										assign node169 = (inp[6]) ? node171 : 46'b0000000000000000000000000000000000000000000000;
											assign node171 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node172;
												assign node172 = (inp[5]) ? node174 : 46'b0000000000000000000000000000000000000000000000;
													assign node174 = (inp[7]) ? node178 : node175;
														assign node175 = (inp[10]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
														assign node178 = (inp[8]) ? 46'b0000000000001000010000000000000000000000010100 : 46'b0000000000000000000000000000000000000000000000;
								assign node182 = (inp[14]) ? node184 : 46'b0000000000000000000000000000000000000000000000;
									assign node184 = (inp[13]) ? node186 : 46'b0000000000000000000000000000000000000000000000;
										assign node186 = (inp[5]) ? node188 : 46'b0000000000000000000000000000000000000000000000;
											assign node188 = (inp[6]) ? node196 : node189;
												assign node189 = (inp[10]) ? node191 : 46'b0000000000000000000000000000000000000000000000;
													assign node191 = (inp[8]) ? node193 : 46'b0000000000000000000000000000000000000000000000;
														assign node193 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
												assign node196 = (inp[4]) ? node202 : node197;
													assign node197 = (inp[10]) ? node199 : 46'b0000000000000000000000000000000000000000000000;
														assign node199 = (inp[8]) ? 46'b0010000000000000001000010100000000000000010000 : 46'b0000000000000000000000000000000000000000000000;
													assign node202 = (inp[7]) ? node206 : node203;
														assign node203 = (inp[12]) ? 46'b0000010000000000011000000100000000000000010000 : 46'b0000000000000000000000000000000000000000000000;
														assign node206 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
						assign node209 = (inp[13]) ? node211 : 46'b0000000000000000000000000000000000000000000000;
							assign node211 = (inp[5]) ? node213 : 46'b0000000000000000000000000000000000000000000000;
								assign node213 = (inp[14]) ? node215 : 46'b0000000000000000000000000000000000000000000000;
									assign node215 = (inp[6]) ? node227 : node216;
										assign node216 = (inp[10]) ? node218 : 46'b0000000000000000000000000000000000000000000000;
											assign node218 = (inp[11]) ? node220 : 46'b0000000000000000000000000000000000000000000000;
												assign node220 = (inp[4]) ? node222 : 46'b0000000000000000000000000000000000000000000000;
													assign node222 = (inp[8]) ? node224 : 46'b0000000000000000000000000000000000000000000000;
														assign node224 = (inp[7]) ? 46'b0000000000000000000010000000010000000000000000 : 46'b0000000000000000000000000000000000000000000000;
										assign node227 = (inp[10]) ? node239 : node228;
											assign node228 = (inp[4]) ? node230 : 46'b0000000000000000000000000000000000000000000000;
												assign node230 = (inp[8]) ? node232 : 46'b0000000000000000000000000000000000000000000000;
													assign node232 = (inp[0]) ? node236 : node233;
														assign node233 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000001000010000000000000100000010000000;
														assign node236 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
											assign node239 = (inp[11]) ? node249 : node240;
												assign node240 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node241;
													assign node241 = (inp[8]) ? node245 : node242;
														assign node242 = (inp[4]) ? 46'b0000000000010000010000000000000000000010000000 : 46'b0000000000000000000000000000000000000000000000;
														assign node245 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000010000000000000010000000;
												assign node249 = (inp[12]) ? node257 : node250;
													assign node250 = (inp[7]) ? node254 : node251;
														assign node251 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0010000000000000000010100000000000000010000000;
														assign node254 = (inp[4]) ? 46'b0000000000011000010010000000000000000010000000 : 46'b0000000000001000010010010000000000000010000000;
													assign node257 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node258;
														assign node258 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
		assign node262 = (inp[15]) ? node330 : node263;
			assign node263 = (inp[13]) ? node267 : node264;
				assign node264 = (inp[3]) ? 46'b0000100000000000000000000000001000000000000000 : 46'b0000100000000000000000000000000000000000000000;
				assign node267 = (inp[2]) ? node299 : node268;
					assign node268 = (inp[9]) ? node284 : node269;
						assign node269 = (inp[11]) ? node277 : node270;
							assign node270 = (inp[0]) ? node274 : node271;
								assign node271 = (inp[3]) ? 46'b0000100000001000010000010100001000000000010010 : 46'b0000100000001000010000010100000000000000010010;
								assign node274 = (inp[3]) ? 46'b0000100000001000010000000100001100000000010010 : 46'b0000100000001000010000000100000100000000010010;
							assign node277 = (inp[0]) ? node281 : node278;
								assign node278 = (inp[3]) ? 46'b0000100000001000011000010100001000000000010000 : 46'b0000100000001000011000010100000000000000010000;
								assign node281 = (inp[3]) ? 46'b0000100000001000011000000100001100000000010000 : 46'b0000100000001000011000000100000100000000010000;
						assign node284 = (inp[11]) ? node292 : node285;
							assign node285 = (inp[0]) ? node289 : node286;
								assign node286 = (inp[3]) ? 46'b0000110000000000010000010100001000000000010010 : 46'b0000110000000000010000010100000000000000010010;
								assign node289 = (inp[3]) ? 46'b0000110000000000010000000100001100000000010010 : 46'b0000110000000000010000000100000100000000010010;
							assign node292 = (inp[0]) ? node296 : node293;
								assign node293 = (inp[3]) ? 46'b0000110000000000011000010100001000000000010000 : 46'b0000110000000000011000010100000000000000010000;
								assign node296 = (inp[3]) ? 46'b0000110000000000011000000100001100000000010000 : 46'b0000110000000000011000000100000100000000010000;
					assign node299 = (inp[9]) ? node315 : node300;
						assign node300 = (inp[0]) ? node308 : node301;
							assign node301 = (inp[11]) ? node305 : node302;
								assign node302 = (inp[3]) ? 46'b0000100000001000010010110000001000000010000000 : 46'b0000100000001000010010110000000000000010000000;
								assign node305 = (inp[3]) ? 46'b0000100000001000010010010000011000000010000000 : 46'b0000100000001000010010010000010000000010000000;
							assign node308 = (inp[11]) ? node312 : node309;
								assign node309 = (inp[3]) ? 46'b0000100000001000010010100000001100000010000000 : 46'b0000100000001000010010100000000100000010000000;
								assign node312 = (inp[3]) ? 46'b0000100000001000010010000000011100000010000000 : 46'b0000100000001000010010000000010100000010000000;
						assign node315 = (inp[0]) ? node323 : node316;
							assign node316 = (inp[11]) ? node320 : node317;
								assign node317 = (inp[3]) ? 46'b0000110000000000010010110000001000000010000000 : 46'b0000110000000000010010110000000000000010000000;
								assign node320 = (inp[3]) ? 46'b0000110000000000010010010000011000000010000000 : 46'b0000110000000000010010010000010000000010000000;
							assign node323 = (inp[11]) ? node327 : node324;
								assign node324 = (inp[3]) ? 46'b0000110000000000010010100000001100000010000000 : 46'b0000110000000000010010100000000100000010000000;
								assign node327 = (inp[3]) ? 46'b0000110000000000010010000000011100000010000000 : 46'b0000110000000000010010000000010100000010000000;
			assign node330 = (inp[13]) ? node334 : node331;
				assign node331 = (inp[3]) ? 46'b0000000000000000000000000000000000000000001000 : 46'b0000000000000000000000000000001000000000001000;
				assign node334 = (inp[3]) ? node336 : 46'b0000000000000000000000000000001000000000000000;
					assign node336 = (inp[2]) ? node1048 : node337;
						assign node337 = (inp[11]) ? node643 : node338;
							assign node338 = (inp[9]) ? node592 : node339;
								assign node339 = (inp[0]) ? node465 : node340;
									assign node340 = (inp[7]) ? node404 : node341;
										assign node341 = (inp[12]) ? node373 : node342;
											assign node342 = (inp[6]) ? node358 : node343;
												assign node343 = (inp[5]) ? node351 : node344;
													assign node344 = (inp[8]) ? node348 : node345;
														assign node345 = (inp[14]) ? 46'b0011000000000000001000010001100010110001010000 : 46'b0011000000000100000000010000100010110001010000;
														assign node348 = (inp[14]) ? 46'b0011000000000010000000010000100010110001010000 : 46'b0011000000000000000000010001100010110001010010;
													assign node351 = (inp[14]) ? node355 : node352;
														assign node352 = (inp[8]) ? 46'b0010000000000000000000010001100010110001010010 : 46'b0010000000000100000000010000100010110001010000;
														assign node355 = (inp[4]) ? 46'b0010000000000010001000010001100010110001010000 : 46'b0010000000000110000000010000100010110001010000;
												assign node358 = (inp[10]) ? node366 : node359;
													assign node359 = (inp[4]) ? node363 : node360;
														assign node360 = (inp[5]) ? 46'b0010000000000100000000010000100010010001010000 : 46'b0011000000000100000000010000100010010001010000;
														assign node363 = (inp[5]) ? 46'b0010000000000000001000010001100010010001010000 : 46'b0011000000000000001000010001100010010001010000;
													assign node366 = (inp[5]) ? node370 : node367;
														assign node367 = (inp[8]) ? 46'b0011000000000010000000010001100010010001010010 : 46'b0011000000000010001000010001100010010001010000;
														assign node370 = (inp[8]) ? 46'b0010000000000010000000010001100010010001010010 : 46'b0010000000000110000000010000100010010001010000;
											assign node373 = (inp[5]) ? node389 : node374;
												assign node374 = (inp[14]) ? node382 : node375;
													assign node375 = (inp[6]) ? node379 : node376;
														assign node376 = (inp[4]) ? 46'b0011000000000100000000010000100000110001010000 : 46'b0011000000000100000000010001100000110001010010;
														assign node379 = (inp[8]) ? 46'b0011000000000100000000010001100000010001010010 : 46'b0011000000000100000000010000100000010001010000;
													assign node382 = (inp[6]) ? node386 : node383;
														assign node383 = (inp[4]) ? 46'b0011000000000010001000010001100000110001010000 : 46'b0011000000000010000000010000100000110001010000;
														assign node386 = (inp[8]) ? 46'b0011000000000010000000010000100000010001010000 : 46'b0011000000000000001000010001100000010001010010;
												assign node389 = (inp[6]) ? node397 : node390;
													assign node390 = (inp[4]) ? node394 : node391;
														assign node391 = (inp[14]) ? 46'b0010000000000000001000010001100000110001010010 : 46'b0010000000000100000000010001100000110001010010;
														assign node394 = (inp[10]) ? 46'b0010000000000010000000010000100000110001010000 : 46'b0010000000000000001000010001100000110001010000;
													assign node397 = (inp[8]) ? node401 : node398;
														assign node398 = (inp[10]) ? 46'b0010000000000100000000010001100000010001010010 : 46'b0010000000000100001000010001100000010001010000;
														assign node401 = (inp[10]) ? 46'b0010000000000010000000010001100000010001010010 : 46'b0010000000000010000000010000100000010001010000;
										assign node404 = (inp[5]) ? node434 : node405;
											assign node405 = (inp[6]) ? node419 : node406;
												assign node406 = (inp[12]) ? node414 : node407;
													assign node407 = (inp[14]) ? node411 : node408;
														assign node408 = (inp[4]) ? 46'b0011000000000110000000010000000010110001010000 : 46'b0011000000000100000000010001000010110001010010;
														assign node411 = (inp[8]) ? 46'b0011000000000010000000010000000010110001010000 : 46'b0011000000000000001000010001000010110001010000;
													assign node414 = (inp[8]) ? 46'b0011000000000010000000010001000000110001010010 : node415;
														assign node415 = (inp[14]) ? 46'b0011000000000000001000010001000000110001010000 : 46'b0011000000000100000000010000000000110001010000;
												assign node419 = (inp[12]) ? node427 : node420;
													assign node420 = (inp[8]) ? node424 : node421;
														assign node421 = (inp[14]) ? 46'b0011000000000000001000010001000010010001010000 : 46'b0011000000000100000000010000000010010001010000;
														assign node424 = (inp[10]) ? 46'b0011000000000010000000010001000010010001010010 : 46'b0011000000000010000000010000000010010001010000;
													assign node427 = (inp[4]) ? node431 : node428;
														assign node428 = (inp[14]) ? 46'b0011000000000100001000010001000000010001010000 : 46'b0011000000000100000000010001000000010001010010;
														assign node431 = (inp[10]) ? 46'b0011000000000010000000010000000000010001010000 : 46'b0011000000000000001000010001000000010001010000;
											assign node434 = (inp[12]) ? node450 : node435;
												assign node435 = (inp[6]) ? node443 : node436;
													assign node436 = (inp[8]) ? node440 : node437;
														assign node437 = (inp[14]) ? 46'b0010000000000000001000010001000010110001010000 : 46'b0010000000000100000000010000000010110001010000;
														assign node440 = (inp[14]) ? 46'b0010000000000010000000010001000010110001010000 : 46'b0010000000000000000000010001000010110001010010;
													assign node443 = (inp[10]) ? node447 : node444;
														assign node444 = (inp[8]) ? 46'b0010000000000000000000010001000010010001010010 : 46'b0010000000000100001000010001000010010001010000;
														assign node447 = (inp[4]) ? 46'b0010000000000010000000010000000010010001010000 : 46'b0010000000000000000000010001000010010001010010;
												assign node450 = (inp[6]) ? node458 : node451;
													assign node451 = (inp[10]) ? node455 : node452;
														assign node452 = (inp[4]) ? 46'b0010000000000000001000010001000000110001010000 : 46'b0010000000000100000000010000000000110001010000;
														assign node455 = (inp[14]) ? 46'b0010000000000010000000010001000000110001010000 : 46'b0010000000000000000000010001000000110001010010;
													assign node458 = (inp[4]) ? node462 : node459;
														assign node459 = (inp[14]) ? 46'b0010000000000110000000010000000000010001010000 : 46'b0010000000000100000000010001000000010001010010;
														assign node462 = (inp[10]) ? 46'b0010000000000010000000010000000000010001010000 : 46'b0010000000000000001000010001000000010001010000;
									assign node465 = (inp[6]) ? node529 : node466;
										assign node466 = (inp[12]) ? node498 : node467;
											assign node467 = (inp[5]) ? node483 : node468;
												assign node468 = (inp[7]) ? node476 : node469;
													assign node469 = (inp[10]) ? node473 : node470;
														assign node470 = (inp[4]) ? 46'b0011000000000000001000010001100010110000010000 : 46'b0011000000000100000000010000100010110000010000;
														assign node473 = (inp[14]) ? 46'b0011000000000000001000010001100010110000010010 : 46'b0011000000000000000000010001100010110000010010;
													assign node476 = (inp[14]) ? node480 : node477;
														assign node477 = (inp[8]) ? 46'b0011000000000000000000010001000010110000010010 : 46'b0011000000000100000000010000000010110000010000;
														assign node480 = (inp[8]) ? 46'b0011000000000010000000010000000010110000010000 : 46'b0011000000000000001000010001000010110000010000;
												assign node483 = (inp[7]) ? node491 : node484;
													assign node484 = (inp[14]) ? node488 : node485;
														assign node485 = (inp[4]) ? 46'b0010000000000000001000010001100010110000010000 : 46'b0010000000000100000000010001100010110000010010;
														assign node488 = (inp[8]) ? 46'b0010000000000010000000010000100010110000010000 : 46'b0010000000000000001000010001100010110000010000;
													assign node491 = (inp[10]) ? node495 : node492;
														assign node492 = (inp[4]) ? 46'b0010000000000000001000010001000010110000010000 : 46'b0010000000000100000000010000000010110000010000;
														assign node495 = (inp[4]) ? 46'b0010000000000010000000010000000010110000010000 : 46'b0010000000000000000000010001000010110000010010;
											assign node498 = (inp[7]) ? node514 : node499;
												assign node499 = (inp[5]) ? node507 : node500;
													assign node500 = (inp[14]) ? node504 : node501;
														assign node501 = (inp[4]) ? 46'b0011000000000010000000010000100000110000010000 : 46'b0011000000000100000000010001100000110000010010;
														assign node504 = (inp[8]) ? 46'b0011000000000010000000010000100000110000010000 : 46'b0011000000000000001000010001100000110000010000;
													assign node507 = (inp[8]) ? node511 : node508;
														assign node508 = (inp[10]) ? 46'b0010000000000000001000010001100000110000010010 : 46'b0010000000000100001000010001100000110000010000;
														assign node511 = (inp[14]) ? 46'b0010000000000010000000010000100000110000010000 : 46'b0010000000000000000000010001100000110000010010;
												assign node514 = (inp[5]) ? node522 : node515;
													assign node515 = (inp[8]) ? node519 : node516;
														assign node516 = (inp[14]) ? 46'b0011000000000000001000010001000000110000010000 : 46'b0011000000000100000000010000000000110000010000;
														assign node519 = (inp[14]) ? 46'b0011000000000010000000010000000000110000010000 : 46'b0011000000000100000000010001000000110000010010;
													assign node522 = (inp[8]) ? node526 : node523;
														assign node523 = (inp[14]) ? 46'b0010000000000000001000010001000000110000010000 : 46'b0010000000000100000000010000000000110000010000;
														assign node526 = (inp[14]) ? 46'b0010000000000010000000010000000000110000010000 : 46'b0010000000000000000000010001000000110000010010;
										assign node529 = (inp[12]) ? node561 : node530;
											assign node530 = (inp[5]) ? node546 : node531;
												assign node531 = (inp[7]) ? node539 : node532;
													assign node532 = (inp[8]) ? node536 : node533;
														assign node533 = (inp[14]) ? 46'b0011000000000000001000010001100010010000010000 : 46'b0011000000000100000000010000100010010000010000;
														assign node536 = (inp[14]) ? 46'b0011000000000010000000010001100010010000010000 : 46'b0011000000000000000000010001100010010000010010;
													assign node539 = (inp[8]) ? node543 : node540;
														assign node540 = (inp[14]) ? 46'b0011000000000000001000010001000010010000010000 : 46'b0011000000000100000000010000000010010000010000;
														assign node543 = (inp[10]) ? 46'b0011000000000010000000010001000010010000010010 : 46'b0011000000000010000000010000000010010000010000;
												assign node546 = (inp[7]) ? node554 : node547;
													assign node547 = (inp[4]) ? node551 : node548;
														assign node548 = (inp[10]) ? 46'b0010000000000000000000010001100010010000010010 : 46'b0010000000000100000000010000100010010000010000;
														assign node551 = (inp[10]) ? 46'b0010000000000010000000010000100010010000010000 : 46'b0010000000000000001000010001100010010000010000;
													assign node554 = (inp[10]) ? node558 : node555;
														assign node555 = (inp[4]) ? 46'b0010000000000000001000010001000010010000010010 : 46'b0010000000000100000000010000000010010000010000;
														assign node558 = (inp[4]) ? 46'b0010000000000010000000010000000010010000010000 : 46'b0010000000000000000000010001000010010000010010;
											assign node561 = (inp[5]) ? node577 : node562;
												assign node562 = (inp[7]) ? node570 : node563;
													assign node563 = (inp[4]) ? node567 : node564;
														assign node564 = (inp[10]) ? 46'b0011000000000000000000010001100000010000010010 : 46'b0011000000000100000000010000100000010000010000;
														assign node567 = (inp[10]) ? 46'b0011000000000010000000010001100000010000010010 : 46'b0011000000000000001000010001100000010000010000;
													assign node570 = (inp[4]) ? node574 : node571;
														assign node571 = (inp[10]) ? 46'b0011000000000000000000010001000000010000010010 : 46'b0011000000000100000000010000000000010000010000;
														assign node574 = (inp[10]) ? 46'b0011000000000010000000010001000000010000010000 : 46'b0011000000000000001000010001000000010000010000;
												assign node577 = (inp[7]) ? node585 : node578;
													assign node578 = (inp[14]) ? node582 : node579;
														assign node579 = (inp[8]) ? 46'b0010000000000000000000010001100000010000010010 : 46'b0010000000000100000000010001100000010000010000;
														assign node582 = (inp[4]) ? 46'b0010000000000010001000010001100000010000010000 : 46'b0010000000000100001000010001100000010000010000;
													assign node585 = (inp[4]) ? node589 : node586;
														assign node586 = (inp[8]) ? 46'b0010000000000100000000010000000000010000010000 : 46'b0010000000000100000000010000000000010000010000;
														assign node589 = (inp[10]) ? 46'b0010000000000010000000010001000000010000010000 : 46'b0010000000000000001000010001000000010000010000;
								assign node592 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node593;
									assign node593 = (inp[4]) ? node625 : node594;
										assign node594 = (inp[7]) ? node610 : node595;
											assign node595 = (inp[5]) ? node597 : 46'b0000000000000000000000000000000000000000000000;
												assign node597 = (inp[10]) ? node603 : node598;
													assign node598 = (inp[8]) ? node600 : 46'b0000000000000000000000000000000000000000000000;
														assign node600 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000100000000001001100000000000000010;
													assign node603 = (inp[6]) ? node607 : node604;
														assign node604 = (inp[8]) ? 46'b0000000000000010000000001001100000100000000010 : 46'b0000000000000100000000001001100000100000000010;
														assign node607 = (inp[12]) ? 46'b0000000000000000000000001001100000000000000010 : 46'b0000000000000000000000001001100010000000000010;
											assign node610 = (inp[5]) ? 46'b0000000000000000000000000000000000000000000000 : node611;
												assign node611 = (inp[10]) ? node619 : node612;
													assign node612 = (inp[6]) ? node616 : node613;
														assign node613 = (inp[12]) ? 46'b0001000000000100000000001000000000100000000000 : 46'b0001000000000100000000001000000010100000000000;
														assign node616 = (inp[12]) ? 46'b0001000000000100000000001001000000000000000000 : 46'b0001000000000100000000001001000010000000000000;
													assign node619 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : node620;
														assign node620 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000000100000000001001000000000000000010;
										assign node625 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : node626;
											assign node626 = (inp[8]) ? node634 : node627;
												assign node627 = (inp[5]) ? 46'b0000000000000000000000000000000000000000000000 : node628;
													assign node628 = (inp[7]) ? node630 : 46'b0000000000000000000000000000000000000000000000;
														assign node630 = (inp[10]) ? 46'b0001000000000110000000001000000000000000000000 : 46'b0001000000000100001000001001000000000000000000;
												assign node634 = (inp[5]) ? node636 : 46'b0000000000000000000000000000000000000000000000;
													assign node636 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node637;
														assign node637 = (inp[10]) ? 46'b0000000000000010000000001001100000100000000010 : 46'b0000000000000000001000001001100010000000000010;
							assign node643 = (inp[9]) ? node795 : node644;
								assign node644 = (inp[0]) ? node668 : node645;
									assign node645 = (inp[5]) ? node647 : 46'b0000000000000000000000000000000000000000000000;
										assign node647 = (inp[7]) ? node649 : 46'b0000000000000000000000000000000000000000000000;
											assign node649 = (inp[12]) ? node659 : node650;
												assign node650 = (inp[6]) ? node652 : 46'b0000000000000000000000000000000000000000000000;
													assign node652 = (inp[8]) ? node656 : node653;
														assign node653 = (inp[14]) ? 46'b0000000000000010001001000001000010000000000000 : 46'b0000000000000100000001000000000010000000000000;
														assign node656 = (inp[14]) ? 46'b0000000000000010000001000001000010000000000000 : 46'b0000000000000000000001000001000010000000000010;
												assign node659 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : node660;
													assign node660 = (inp[10]) ? node664 : node661;
														assign node661 = (inp[4]) ? 46'b0000000000000000001001000001000000100000000000 : 46'b0000000000000100000001000000000000100000000000;
														assign node664 = (inp[4]) ? 46'b0000000000000010000001000000000000100000000000 : 46'b0000000000000000000001000001000000100000000010;
									assign node668 = (inp[12]) ? node732 : node669;
										assign node669 = (inp[6]) ? node701 : node670;
											assign node670 = (inp[7]) ? node686 : node671;
												assign node671 = (inp[5]) ? node679 : node672;
													assign node672 = (inp[8]) ? node676 : node673;
														assign node673 = (inp[14]) ? 46'b0101000000000000001000000001100010100000000000 : 46'b0101000000000100000000000000100010100000000000;
														assign node676 = (inp[10]) ? 46'b0101000000000010000000000001100010100000000010 : 46'b0101000000000100000000000000100010100000000000;
													assign node679 = (inp[14]) ? node683 : node680;
														assign node680 = (inp[4]) ? 46'b0100000000000000001000000001100010100000000000 : 46'b0100000000000100000000000001100010100000000010;
														assign node683 = (inp[4]) ? 46'b0100000000000010001000000001100010100000000000 : 46'b0100000000000000000000000001100010100000000010;
												assign node686 = (inp[5]) ? node694 : node687;
													assign node687 = (inp[10]) ? node691 : node688;
														assign node688 = (inp[14]) ? 46'b0101000000000100000000000000000010100000000000 : 46'b0101000000000100000000000000000010100000000000;
														assign node691 = (inp[8]) ? 46'b0101000000000010000000000001000010100000000010 : 46'b0101000000000010000000000000000010100000000000;
													assign node694 = (inp[10]) ? node698 : node695;
														assign node695 = (inp[4]) ? 46'b0100000000000000001000000001000010100000000000 : 46'b0100000000000100000000000000000010100000000000;
														assign node698 = (inp[4]) ? 46'b0100000000000010000000000000000010100000000000 : 46'b0100000000000000000000000001000010100000000010;
											assign node701 = (inp[7]) ? node717 : node702;
												assign node702 = (inp[5]) ? node710 : node703;
													assign node703 = (inp[4]) ? node707 : node704;
														assign node704 = (inp[10]) ? 46'b0101000000000000000000000001100010000000000010 : 46'b0101000000000100000000000000100010000000000000;
														assign node707 = (inp[10]) ? 46'b0101000000000010000000000000100010000000000000 : 46'b0101000000000000001000000001100010000000000000;
													assign node710 = (inp[4]) ? node714 : node711;
														assign node711 = (inp[10]) ? 46'b0100000000000000000000000001100010000000000010 : 46'b0100000000000100000000000000100010000000000000;
														assign node714 = (inp[10]) ? 46'b0100000000000010000000000000100010000000000000 : 46'b0100000000000000001000000001100010000000000000;
												assign node717 = (inp[5]) ? node725 : node718;
													assign node718 = (inp[4]) ? node722 : node719;
														assign node719 = (inp[10]) ? 46'b0101000000000000000000000001000010000000000010 : 46'b0101000000000100000000000000000010000000000000;
														assign node722 = (inp[10]) ? 46'b0101000000000010000000000000000010000000000000 : 46'b0101000000000000001000000001000010000000000000;
													assign node725 = (inp[8]) ? node729 : node726;
														assign node726 = (inp[14]) ? 46'b0100000000000000001000000001000010000000000000 : 46'b0100000000000100000000000000000010000000000000;
														assign node729 = (inp[10]) ? 46'b0100000000000010000000000001000010000000000010 : 46'b0100000000000100000000000001000010000000000010;
										assign node732 = (inp[5]) ? node764 : node733;
											assign node733 = (inp[7]) ? node749 : node734;
												assign node734 = (inp[6]) ? node742 : node735;
													assign node735 = (inp[10]) ? node739 : node736;
														assign node736 = (inp[8]) ? 46'b0101000000000110000000000000100000100000000000 : 46'b0101000000000100000000000000100000100000000000;
														assign node739 = (inp[8]) ? 46'b0101000000000010000000000001100000100000000010 : 46'b0101000000000000001000000001100000100000000010;
													assign node742 = (inp[8]) ? node746 : node743;
														assign node743 = (inp[14]) ? 46'b0101000000000000001000000001100000000000000000 : 46'b0101000000000100000000000000100000000000000000;
														assign node746 = (inp[14]) ? 46'b0101000000000010000000000001100000000000000000 : 46'b0101000000000000000000000001100000000000000010;
												assign node749 = (inp[6]) ? node757 : node750;
													assign node750 = (inp[8]) ? node754 : node751;
														assign node751 = (inp[14]) ? 46'b0101000000000000001000000001000000100000000000 : 46'b0101000000000100000000000000000000100000000000;
														assign node754 = (inp[10]) ? 46'b0101000000000010000000000001000000100000000010 : 46'b0101000000000000000000000001000000100000000010;
													assign node757 = (inp[8]) ? node761 : node758;
														assign node758 = (inp[14]) ? 46'b0101000000000000001000000001000000000000000000 : 46'b0101000000000100000000000001000000000000000000;
														assign node761 = (inp[14]) ? 46'b0101000000000010000000000000000000000000000000 : 46'b0101000000000000000000000001000000000000000010;
											assign node764 = (inp[7]) ? node780 : node765;
												assign node765 = (inp[6]) ? node773 : node766;
													assign node766 = (inp[8]) ? node770 : node767;
														assign node767 = (inp[14]) ? 46'b0100000000000000001000000001100000100000000000 : 46'b0100000000000100000000000000100000100000000000;
														assign node770 = (inp[14]) ? 46'b0100000000000010000000000001100000100000000000 : 46'b0100000000000000000000000001100000100000000010;
													assign node773 = (inp[10]) ? node777 : node774;
														assign node774 = (inp[4]) ? 46'b0100000000000000001000000001100000000000000000 : 46'b0100000000000100000000000001100000000000000000;
														assign node777 = (inp[8]) ? 46'b0100000000000010000000000001100000000000000010 : 46'b0100000000000100000000000000100000000000000000;
												assign node780 = (inp[6]) ? node788 : node781;
													assign node781 = (inp[10]) ? node785 : node782;
														assign node782 = (inp[4]) ? 46'b0100000000000000001000000001000000100000000000 : 46'b0100000000000100000000000000000000100000000000;
														assign node785 = (inp[4]) ? 46'b0100000000000010000000000000000000100000000000 : 46'b0100000000000000000000000001000000100000000010;
													assign node788 = (inp[4]) ? node792 : node789;
														assign node789 = (inp[10]) ? 46'b0100000000000000000000000001000000000000000010 : 46'b0100000000000100000000000001000000000000000000;
														assign node792 = (inp[14]) ? 46'b0100000000000010000000000000000000000000000000 : 46'b0100000000000110000000000000000000000000000000;
								assign node795 = (inp[0]) ? node923 : node796;
									assign node796 = (inp[7]) ? node860 : node797;
										assign node797 = (inp[6]) ? node829 : node798;
											assign node798 = (inp[5]) ? node814 : node799;
												assign node799 = (inp[12]) ? node807 : node800;
													assign node800 = (inp[10]) ? node804 : node801;
														assign node801 = (inp[8]) ? 46'b1001000000000000001000000001100010100000000010 : 46'b1001000000000100001000000001100010100000000000;
														assign node804 = (inp[14]) ? 46'b1001000000000000001000000001100010100000000000 : 46'b1001000000000000000000000001100010100000000010;
													assign node807 = (inp[10]) ? node811 : node808;
														assign node808 = (inp[4]) ? 46'b1001000000000000001000000001100000100000000000 : 46'b1001000000000100000000000000100000100000000000;
														assign node811 = (inp[4]) ? 46'b1001000000000010000000000000100000100000000000 : 46'b1001000000000000000000000001100000100000000010;
												assign node814 = (inp[12]) ? node822 : node815;
													assign node815 = (inp[8]) ? node819 : node816;
														assign node816 = (inp[10]) ? 46'b1000000000000000001000000001100010100000000010 : 46'b1000000000000100001000000001100010100000000000;
														assign node819 = (inp[10]) ? 46'b1000000000000000000000000001100010100000000010 : 46'b1000000000000000000000000001100010100000000010;
													assign node822 = (inp[8]) ? node826 : node823;
														assign node823 = (inp[10]) ? 46'b1000000000000000001000000001100000100000000000 : 46'b1000000000000100001000000001100000100000000000;
														assign node826 = (inp[10]) ? 46'b1000000000000010000000000001100000100000000010 : 46'b1000000000000000001000000001100000100000000000;
											assign node829 = (inp[5]) ? node845 : node830;
												assign node830 = (inp[8]) ? node838 : node831;
													assign node831 = (inp[12]) ? node835 : node832;
														assign node832 = (inp[14]) ? 46'b1001000000000000001000000001100010000000000000 : 46'b1001000000000100001000000001100010000000000000;
														assign node835 = (inp[14]) ? 46'b1001000000000000001000000001100000000000000000 : 46'b1001000000000100000000000000100000000000000000;
													assign node838 = (inp[14]) ? node842 : node839;
														assign node839 = (inp[4]) ? 46'b1001000000000010000000000001100000000000000010 : 46'b1001000000000100000000000001100010000000000010;
														assign node842 = (inp[12]) ? 46'b1001000000000010000000000000100000000000000000 : 46'b1001000000000010000000000000100010000000000000;
												assign node845 = (inp[12]) ? node853 : node846;
													assign node846 = (inp[8]) ? node850 : node847;
														assign node847 = (inp[14]) ? 46'b1000000000000000001000000001100010000000000000 : 46'b1000000000000100000000000000100010000000000000;
														assign node850 = (inp[14]) ? 46'b1000000000000010000000000000100010000000000000 : 46'b1000000000000000000000000001100010000000000010;
													assign node853 = (inp[8]) ? node857 : node854;
														assign node854 = (inp[14]) ? 46'b1000000000000000001000000001100000000000000000 : 46'b1000000000000100000000000000100000000000000000;
														assign node857 = (inp[14]) ? 46'b1000000000000010000000000000100000000000000000 : 46'b1000000000000000000000000001100000000000000010;
										assign node860 = (inp[12]) ? node892 : node861;
											assign node861 = (inp[6]) ? node877 : node862;
												assign node862 = (inp[5]) ? node870 : node863;
													assign node863 = (inp[8]) ? node867 : node864;
														assign node864 = (inp[14]) ? 46'b1001000000000000001000000001000010100000000000 : 46'b1001000000000100000000000000000010100000000000;
														assign node867 = (inp[14]) ? 46'b1001000000000010000000000000000010100000000000 : 46'b1001000000000000000000000001000010100000000010;
													assign node870 = (inp[14]) ? node874 : node871;
														assign node871 = (inp[8]) ? 46'b1000000000000000000000000001000010100000000010 : 46'b1000000000000100000000000001000010100000000000;
														assign node874 = (inp[4]) ? 46'b1000000000000010001000000001000010100000000000 : 46'b1000000000000010000000000000000010100000000000;
												assign node877 = (inp[5]) ? node885 : node878;
													assign node878 = (inp[14]) ? node882 : node879;
														assign node879 = (inp[8]) ? 46'b1001000000000000000000000001000010000000000010 : 46'b1001000000000100000000000001000010000000000000;
														assign node882 = (inp[8]) ? 46'b1001000000000010000000000000000010000000000000 : 46'b1001000000000000001000000001000010000000000000;
													assign node885 = (inp[8]) ? node889 : node886;
														assign node886 = (inp[10]) ? 46'b1000000000000000001000000001000010000000000000 : 46'b1000000000000100001000000001000010000000000000;
														assign node889 = (inp[14]) ? 46'b1000000000000010000000000000000010000000000000 : 46'b1000000000000000000000000001000010000000000010;
											assign node892 = (inp[5]) ? node908 : node893;
												assign node893 = (inp[6]) ? node901 : node894;
													assign node894 = (inp[8]) ? node898 : node895;
														assign node895 = (inp[14]) ? 46'b1001000000000000001000000001000000100000000000 : 46'b1001000000000100000000000000000000100000000000;
														assign node898 = (inp[14]) ? 46'b1001000000000010000000000000000000100000000000 : 46'b1001000000000000000000000001000000100000000010;
													assign node901 = (inp[4]) ? node905 : node902;
														assign node902 = (inp[10]) ? 46'b1001000000000000000000000001000000000000000010 : 46'b1001000000000100000000000000000000000000000000;
														assign node905 = (inp[10]) ? 46'b1001000000000010000000000000000000000000000000 : 46'b1001000000000000001000000001000000000000000000;
												assign node908 = (inp[6]) ? node916 : node909;
													assign node909 = (inp[8]) ? node913 : node910;
														assign node910 = (inp[14]) ? 46'b1000000000000000001000000001000000100000000010 : 46'b1000000000000100000000000000000000100000000000;
														assign node913 = (inp[14]) ? 46'b1000000000000010000000000001000000100000000000 : 46'b1000000000000000000000000001000000100000000010;
													assign node916 = (inp[8]) ? node920 : node917;
														assign node917 = (inp[14]) ? 46'b1000000000000000001000000001000000000000000000 : 46'b1000000000000100000000000000000000000000000000;
														assign node920 = (inp[4]) ? 46'b1000000000000010000000000001000000000000000000 : 46'b1000000000000000000000000001000000000000000010;
									assign node923 = (inp[6]) ? node987 : node924;
										assign node924 = (inp[5]) ? node956 : node925;
											assign node925 = (inp[7]) ? node941 : node926;
												assign node926 = (inp[12]) ? node934 : node927;
													assign node927 = (inp[10]) ? node931 : node928;
														assign node928 = (inp[4]) ? 46'b0001000000000000001000000001100010101000000000 : 46'b0001000000000100000000000000100010101000000000;
														assign node931 = (inp[8]) ? 46'b0001000000000010000000000001100010101000000010 : 46'b0001000000000110000000000000100010101000000000;
													assign node934 = (inp[4]) ? node938 : node935;
														assign node935 = (inp[10]) ? 46'b0001000000000100000000000001100000101000000010 : 46'b0001000000000100000000000000100000101000000000;
														assign node938 = (inp[10]) ? 46'b0001000000000010000000000000100000101000000000 : 46'b0001000000000000001000000001100000101000000000;
												assign node941 = (inp[12]) ? node949 : node942;
													assign node942 = (inp[10]) ? node946 : node943;
														assign node943 = (inp[4]) ? 46'b0001000000000000001000000001000010101000000000 : 46'b0001000000000100000000000000000010101000000000;
														assign node946 = (inp[4]) ? 46'b0001000000000010000000000000000010101000000000 : 46'b0001000000000000000000000001000010101000000010;
													assign node949 = (inp[4]) ? node953 : node950;
														assign node950 = (inp[10]) ? 46'b0001000000000000000000000001000000101000000010 : 46'b0001000000000100000000000000000000101000000000;
														assign node953 = (inp[14]) ? 46'b0001000000000010001000000001000000101000000000 : 46'b0001000000000000001000000001000000101000000010;
											assign node956 = (inp[7]) ? node972 : node957;
												assign node957 = (inp[12]) ? node965 : node958;
													assign node958 = (inp[10]) ? node962 : node959;
														assign node959 = (inp[4]) ? 46'b0000000000000000001000000001100010101000000000 : 46'b0000000000000100000000000000100010101000000000;
														assign node962 = (inp[8]) ? 46'b0000000000000010000000000001100010101000000010 : 46'b0000000000000000001000000001100010101000000000;
													assign node965 = (inp[14]) ? node969 : node966;
														assign node966 = (inp[8]) ? 46'b0000000000000000000000000001100000101000000010 : 46'b0000000000000100001000000001100000101000000000;
														assign node969 = (inp[8]) ? 46'b0000000000000010000000000000100000101000000000 : 46'b0000000000000000001000000001100000101000000000;
												assign node972 = (inp[12]) ? node980 : node973;
													assign node973 = (inp[4]) ? node977 : node974;
														assign node974 = (inp[8]) ? 46'b0000000000000000000000000001000010101000000010 : 46'b0000000000000100000000000000000010101000000000;
														assign node977 = (inp[10]) ? 46'b0000000000000010000000000000000010101000000000 : 46'b0000000000000000001000000001000010101000000000;
													assign node980 = (inp[4]) ? node984 : node981;
														assign node981 = (inp[10]) ? 46'b0000000000000000000000000001000000101000000010 : 46'b0000000000000100000000000000000000101000000000;
														assign node984 = (inp[10]) ? 46'b0000000000000010000000000000000000101000000000 : 46'b0000000000000000001000000001000000101000000000;
										assign node987 = (inp[12]) ? node1017 : node988;
											assign node988 = (inp[5]) ? node1004 : node989;
												assign node989 = (inp[7]) ? node997 : node990;
													assign node990 = (inp[14]) ? node994 : node991;
														assign node991 = (inp[8]) ? 46'b0001000000000000000000000001100010001000000010 : 46'b0001000000000100000000000000100010001000000000;
														assign node994 = (inp[8]) ? 46'b0001000000000010000000000000100010001000000000 : 46'b0001000000000000001000000001100010001000000000;
													assign node997 = (inp[10]) ? node1001 : node998;
														assign node998 = (inp[4]) ? 46'b0001000000000000001000000001000010001000000000 : 46'b0001000000000100000000000001000010001000000000;
														assign node1001 = (inp[8]) ? 46'b0001000000000010000000000001000010001000000010 : 46'b0001000000000110000000000000000010001000000000;
												assign node1004 = (inp[7]) ? node1012 : node1005;
													assign node1005 = (inp[8]) ? node1009 : node1006;
														assign node1006 = (inp[10]) ? 46'b0000000000000000000000000001100010001000000010 : 46'b0000000000000100001000000001100010001000000000;
														assign node1009 = (inp[14]) ? 46'b0000000000000010000000000000100010001000000000 : 46'b0000000000000000000000000001100010001000000010;
													assign node1012 = (inp[10]) ? 46'b0000000000000000000000000001000010001000000010 : node1013;
														assign node1013 = (inp[4]) ? 46'b0000000000000000001000000001000010001000000000 : 46'b0000000000000100000000000000000010001000000000;
											assign node1017 = (inp[7]) ? node1033 : node1018;
												assign node1018 = (inp[5]) ? node1026 : node1019;
													assign node1019 = (inp[4]) ? node1023 : node1020;
														assign node1020 = (inp[14]) ? 46'b0001000000000000001000000001100000001000000000 : 46'b0001000000000100000000000001100000001000000010;
														assign node1023 = (inp[10]) ? 46'b0001000000000010000000000000100000001000000000 : 46'b0001000000000000001000000001100000001000000000;
													assign node1026 = (inp[8]) ? node1030 : node1027;
														assign node1027 = (inp[14]) ? 46'b0000000000000000001000000001100000001000000000 : 46'b0000000000000100001000000001100000001000000000;
														assign node1030 = (inp[14]) ? 46'b0000000000000010000000000000100000001000000000 : 46'b0000000000000000000000000001100000001000000010;
												assign node1033 = (inp[5]) ? node1041 : node1034;
													assign node1034 = (inp[14]) ? node1038 : node1035;
														assign node1035 = (inp[8]) ? 46'b0001000000000000001000000001000000001000000010 : 46'b0001000000000100000000000000000000001000000000;
														assign node1038 = (inp[4]) ? 46'b0001000000000010001000000001000000001000000000 : 46'b0001000000000000001000000001000000001000000010;
													assign node1041 = (inp[4]) ? node1045 : node1042;
														assign node1042 = (inp[10]) ? 46'b0000000000000000000000000001000000001000000010 : 46'b0000000000000100000000000000000000001000000000;
														assign node1045 = (inp[14]) ? 46'b0000000000000010001000000001000000001000000000 : 46'b0000000000000000000000000001000000001000000010;
						assign node1048 = (inp[11]) ? node1386 : node1049;
							assign node1049 = (inp[9]) ? node1131 : node1050;
								assign node1050 = (inp[7]) ? node1066 : node1051;
									assign node1051 = (inp[12]) ? node1053 : 46'b0000000000000000000000000000000000000000000000;
										assign node1053 = (inp[5]) ? node1055 : 46'b0000000000000000000000000000000000000000000000;
											assign node1055 = (inp[0]) ? node1057 : 46'b0000000000000000000000000000000000000000000000;
												assign node1057 = (inp[6]) ? node1059 : 46'b0000000000000000000000000000000000000000000000;
													assign node1059 = (inp[10]) ? node1063 : node1060;
														assign node1060 = (inp[8]) ? 46'b0000000000000111000000000000100000000000100000 : 46'b0000000000000101001000000001100000000000100000;
														assign node1063 = (inp[8]) ? 46'b0000000000000001000000000001100000000000100010 : 46'b0000000000000011000000000000100000000000100000;
									assign node1066 = (inp[5]) ? node1080 : node1067;
										assign node1067 = (inp[12]) ? node1069 : 46'b0000000000000000000000000000000000000000000000;
											assign node1069 = (inp[6]) ? node1071 : 46'b0000000000000000000000000000000000000000000000;
												assign node1071 = (inp[0]) ? node1073 : 46'b0000000000000000000000000000000000000000000000;
													assign node1073 = (inp[14]) ? node1077 : node1074;
														assign node1074 = (inp[8]) ? 46'b0001000000000001000000000001000000000000100010 : 46'b0001000000000101000000000000000000000000100000;
														assign node1077 = (inp[4]) ? 46'b0001000000000011001000000001000000000000100000 : 46'b0001000000000001001000000001000000000000100010;
										assign node1080 = (inp[0]) ? node1112 : node1081;
											assign node1081 = (inp[12]) ? node1097 : node1082;
												assign node1082 = (inp[6]) ? node1090 : node1083;
													assign node1083 = (inp[4]) ? node1087 : node1084;
														assign node1084 = (inp[10]) ? 46'b0000000000100000000001000001000010100000000010 : 46'b0000000000100100000001000000000010100000000000;
														assign node1087 = (inp[10]) ? 46'b0000000000100010000001000001000010100000000000 : 46'b0000000000100000001001000001000010100000000000;
													assign node1090 = (inp[10]) ? node1094 : node1091;
														assign node1091 = (inp[4]) ? 46'b0000000000100000001001000001000010000000000000 : 46'b0000000000100100000001000000000010000000000000;
														assign node1094 = (inp[4]) ? 46'b0000000000100010000001000001000010000000000000 : 46'b0000000000100000000001000001000010000000000010;
												assign node1097 = (inp[6]) ? node1105 : node1098;
													assign node1098 = (inp[4]) ? node1102 : node1099;
														assign node1099 = (inp[14]) ? 46'b0000000000100100000001000000000000100000000000 : 46'b0000000000100100000001000001000000100000000010;
														assign node1102 = (inp[10]) ? 46'b0000000000100010000001000000000000100000000000 : 46'b0000000000100000001001000001000000100000000000;
													assign node1105 = (inp[14]) ? node1109 : node1106;
														assign node1106 = (inp[8]) ? 46'b0000000000100000000001000001000000000000000010 : 46'b0000000000100100000001000000000000000000000000;
														assign node1109 = (inp[8]) ? 46'b0000000000100010000001000000000000000000000000 : 46'b0000000000100010001001000001000000000000000000;
											assign node1112 = (inp[12]) ? node1122 : node1113;
												assign node1113 = (inp[6]) ? node1115 : 46'b0000000000000000000000000000000000000000000000;
													assign node1115 = (inp[10]) ? node1119 : node1116;
														assign node1116 = (inp[4]) ? 46'b0000000000000001001000000001000010000000100000 : 46'b0000000000000101000000000001000010000000100000;
														assign node1119 = (inp[4]) ? 46'b0000000000000011000000000000000010000000100000 : 46'b0000000000000011000000000001000010000000100010;
												assign node1122 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : node1123;
													assign node1123 = (inp[14]) ? node1127 : node1124;
														assign node1124 = (inp[8]) ? 46'b0000000000000001000000000001000000100000100010 : 46'b0000000000000101000000000000000000100000100000;
														assign node1127 = (inp[8]) ? 46'b0000000000000011000000000001000000100000100000 : 46'b0000000000000001001000000001000000100000100000;
								assign node1131 = (inp[5]) ? node1259 : node1132;
									assign node1132 = (inp[7]) ? node1196 : node1133;
										assign node1133 = (inp[12]) ? node1165 : node1134;
											assign node1134 = (inp[0]) ? node1150 : node1135;
												assign node1135 = (inp[14]) ? node1143 : node1136;
													assign node1136 = (inp[4]) ? node1140 : node1137;
														assign node1137 = (inp[6]) ? 46'b0001000000100100000000000001100010000000100010 : 46'b0001000000100100000000000001100010100000100010;
														assign node1140 = (inp[10]) ? 46'b0001000000100010000000000001100010000000100010 : 46'b0001000000100000001000000001100010000000100010;
													assign node1143 = (inp[6]) ? node1147 : node1144;
														assign node1144 = (inp[4]) ? 46'b0001000000100010001000000001100010100000100000 : 46'b0001000000100000001000000001100010100000100000;
														assign node1147 = (inp[8]) ? 46'b0001000000100010000000000000100010000000100000 : 46'b0001000000100000001000000001100010000000100000;
												assign node1150 = (inp[6]) ? node1158 : node1151;
													assign node1151 = (inp[14]) ? node1155 : node1152;
														assign node1152 = (inp[4]) ? 46'b0001000000000100000000000000100010100000100000 : 46'b0001000000000100000000000001100010100000100010;
														assign node1155 = (inp[8]) ? 46'b0001000000000010000000000001100010100000100000 : 46'b0001000000000000001000000001100010100000100000;
													assign node1158 = (inp[10]) ? node1162 : node1159;
														assign node1159 = (inp[4]) ? 46'b0001000000000000001000000001100010000000100000 : 46'b0001000000000100000000000000100010000000100000;
														assign node1162 = (inp[14]) ? 46'b0001000000000000001000000001100010000000100000 : 46'b0001000000000000000000000001100010000000100010;
											assign node1165 = (inp[0]) ? node1181 : node1166;
												assign node1166 = (inp[8]) ? node1174 : node1167;
													assign node1167 = (inp[14]) ? node1171 : node1168;
														assign node1168 = (inp[6]) ? 46'b0001000000100100000000000000100000000000100000 : 46'b0001000000100100000000000000100000100000100000;
														assign node1171 = (inp[10]) ? 46'b0001000000100000001000000001100000000000100010 : 46'b0001000000100100001000000001100000000000100000;
													assign node1174 = (inp[4]) ? node1178 : node1175;
														assign node1175 = (inp[14]) ? 46'b0001000000100010000000000001100000000000100010 : 46'b0001000000100000000000000001100000000000100010;
														assign node1178 = (inp[14]) ? 46'b0001000000100010000000000000100000000000100000 : 46'b0001000000100010000000000001100000000000100010;
												assign node1181 = (inp[4]) ? node1189 : node1182;
													assign node1182 = (inp[10]) ? node1186 : node1183;
														assign node1183 = (inp[6]) ? 46'b0001000000000100000000000000100000000000100000 : 46'b0001000000000100000000000000100000100000100000;
														assign node1186 = (inp[6]) ? 46'b0001000000000000000000000001100000000000100010 : 46'b0001000000000000000000000001100000100000100010;
													assign node1189 = (inp[10]) ? node1193 : node1190;
														assign node1190 = (inp[8]) ? 46'b0001000000000010001000000001100000000000100000 : 46'b0001000000000000001000000001100000000000100000;
														assign node1193 = (inp[14]) ? 46'b0001000000000010000000000000100000000000100000 : 46'b0001000000000010000000000000100000000000100000;
										assign node1196 = (inp[6]) ? node1228 : node1197;
											assign node1197 = (inp[0]) ? node1213 : node1198;
												assign node1198 = (inp[12]) ? node1206 : node1199;
													assign node1199 = (inp[8]) ? node1203 : node1200;
														assign node1200 = (inp[14]) ? 46'b0001000000100000001000000001000010100000100000 : 46'b0001000000100100000000000000000010100000100000;
														assign node1203 = (inp[10]) ? 46'b0001000000100010000000000001000010100000100010 : 46'b0001000000100100000000000000000010100000100000;
													assign node1206 = (inp[8]) ? node1210 : node1207;
														assign node1207 = (inp[4]) ? 46'b0001000000100000001000000001000000100000100000 : 46'b0001000000100100000000000001000000100000100000;
														assign node1210 = (inp[14]) ? 46'b0001000000100010000000000000000000100000100000 : 46'b0001000000100000001000000001000000100000100010;
												assign node1213 = (inp[12]) ? node1221 : node1214;
													assign node1214 = (inp[8]) ? node1218 : node1215;
														assign node1215 = (inp[14]) ? 46'b0001000000000000001000000001000010100000100000 : 46'b0001000000000100000000000000000010100000100000;
														assign node1218 = (inp[14]) ? 46'b0001000000000010000000000000000010100000100000 : 46'b0001000000000000001000000001000010100000100010;
													assign node1221 = (inp[8]) ? node1225 : node1222;
														assign node1222 = (inp[10]) ? 46'b0001000000000000001000000001000000100000100010 : 46'b0001000000000100001000000001000000100000100000;
														assign node1225 = (inp[14]) ? 46'b0001000000000010000000000000000000100000100000 : 46'b0001000000000000000000000001000000100000100010;
											assign node1228 = (inp[12]) ? node1244 : node1229;
												assign node1229 = (inp[0]) ? node1237 : node1230;
													assign node1230 = (inp[4]) ? node1234 : node1231;
														assign node1231 = (inp[10]) ? 46'b0001000000100000000000000001000010000000100010 : 46'b0001000000100100000000000000000010000000100000;
														assign node1234 = (inp[14]) ? 46'b0001000000100010001000000001000010000000100000 : 46'b0001000000100010000000000001000010000000100010;
													assign node1237 = (inp[4]) ? node1241 : node1238;
														assign node1238 = (inp[10]) ? 46'b0001000000000010000000000001000010000000100010 : 46'b0001000000000100000000000001000010000000100000;
														assign node1241 = (inp[14]) ? 46'b0001000000000010001000000001000010000000100000 : 46'b0001000000000000001000000001000010000000100010;
												assign node1244 = (inp[0]) ? node1252 : node1245;
													assign node1245 = (inp[14]) ? node1249 : node1246;
														assign node1246 = (inp[4]) ? 46'b0001000000100000001000000001000000000000100010 : 46'b0001000000100100000000000001000000000000100010;
														assign node1249 = (inp[4]) ? 46'b0001000000100010001000000001000000000000100000 : 46'b0001000000100000001000000001000000000000100010;
													assign node1252 = (inp[8]) ? node1256 : node1253;
														assign node1253 = (inp[10]) ? 46'b0001000000000000001000000001000000000000100000 : 46'b0001000000000100001000000001000000000000100000;
														assign node1256 = (inp[14]) ? 46'b0001000000000010000000000000000000000000100000 : 46'b0001000000000000000000000001000000000000100010;
									assign node1259 = (inp[6]) ? node1323 : node1260;
										assign node1260 = (inp[7]) ? node1292 : node1261;
											assign node1261 = (inp[12]) ? node1277 : node1262;
												assign node1262 = (inp[4]) ? node1270 : node1263;
													assign node1263 = (inp[10]) ? node1267 : node1264;
														assign node1264 = (inp[14]) ? 46'b0000000000000110000000000000100010100000100000 : 46'b0000000000000100000000000000100010100000100000;
														assign node1267 = (inp[14]) ? 46'b0000000000000000001000000001100010100000100010 : 46'b0000000000000000000000000001100010100000100010;
													assign node1270 = (inp[10]) ? node1274 : node1271;
														assign node1271 = (inp[14]) ? 46'b0000000000100010001000000001100010100000100000 : 46'b0000000000000000001000000001100010100000100010;
														assign node1274 = (inp[0]) ? 46'b0000000000000010000000000000100010100000100000 : 46'b0000000000100010000000000000100010100000100000;
												assign node1277 = (inp[0]) ? node1285 : node1278;
													assign node1278 = (inp[4]) ? node1282 : node1279;
														assign node1279 = (inp[10]) ? 46'b0000000000100000000000000001100000100000100010 : 46'b0000000000100100000000000000100000100000100000;
														assign node1282 = (inp[10]) ? 46'b0000000000100010000000000000100000100000100000 : 46'b0000000000100010001000000001100000100000100000;
													assign node1285 = (inp[10]) ? node1289 : node1286;
														assign node1286 = (inp[4]) ? 46'b0000000000000000001000000001100000100000100000 : 46'b0000000000000100000000000000100000100000100000;
														assign node1289 = (inp[4]) ? 46'b0000000000000010000000000000100000100000100000 : 46'b0000000000000000000000000001100000100000100010;
											assign node1292 = (inp[0]) ? node1308 : node1293;
												assign node1293 = (inp[12]) ? node1301 : node1294;
													assign node1294 = (inp[10]) ? node1298 : node1295;
														assign node1295 = (inp[8]) ? 46'b0000000000100110000000000000000010100000100000 : 46'b0000000000100100001000000001000010100000100000;
														assign node1298 = (inp[4]) ? 46'b0000000000100010000000000000000010100000100000 : 46'b0000000000100000000000000001000010100000100010;
													assign node1301 = (inp[10]) ? node1305 : node1302;
														assign node1302 = (inp[4]) ? 46'b0000000000100000001000000001000000100000100000 : 46'b0000000000100100000000000000000000100000100000;
														assign node1305 = (inp[4]) ? 46'b0000000000100010000000000000000000100000100000 : 46'b0000000000100000000000000001000000100000100010;
												assign node1308 = (inp[8]) ? node1316 : node1309;
													assign node1309 = (inp[14]) ? node1313 : node1310;
														assign node1310 = (inp[10]) ? 46'b0000000000000110000000000000000000100000100000 : 46'b0000000000000100001000000001000000100000100000;
														assign node1313 = (inp[12]) ? 46'b0000000000000000001000000001000000100000100000 : 46'b0000000000000000001000000001000010100000100000;
													assign node1316 = (inp[14]) ? node1320 : node1317;
														assign node1317 = (inp[4]) ? 46'b0000000000000010000000000001000000100000100010 : 46'b0000000000000000000000000001000000100000100010;
														assign node1320 = (inp[12]) ? 46'b0000000000000010000000000000000000100000100000 : 46'b0000000000000010000000000000000010100000100000;
										assign node1323 = (inp[12]) ? node1355 : node1324;
											assign node1324 = (inp[7]) ? node1340 : node1325;
												assign node1325 = (inp[0]) ? node1333 : node1326;
													assign node1326 = (inp[4]) ? node1330 : node1327;
														assign node1327 = (inp[10]) ? 46'b0000000000100000000000000001100010000000100010 : 46'b0000000000100100000000000000100010000000100000;
														assign node1330 = (inp[10]) ? 46'b0000000000100010000000000001100010000000100000 : 46'b0000000000100000001000000001100010000000100000;
													assign node1333 = (inp[8]) ? node1337 : node1334;
														assign node1334 = (inp[10]) ? 46'b0000000000000010001000000001100010000000100000 : 46'b0000000000000100001000000001100010000000100000;
														assign node1337 = (inp[10]) ? 46'b0000000000000010000000000001100010000000100010 : 46'b0000000000000000000000000001100010000000100010;
												assign node1340 = (inp[0]) ? node1348 : node1341;
													assign node1341 = (inp[8]) ? node1345 : node1342;
														assign node1342 = (inp[14]) ? 46'b0000000000100000001000000001000010000000100000 : 46'b0000000000100100000000000000000010000000100000;
														assign node1345 = (inp[10]) ? 46'b0000000000100010000000000001000010000000100010 : 46'b0000000000100010000000000000000010000000100000;
													assign node1348 = (inp[4]) ? node1352 : node1349;
														assign node1349 = (inp[14]) ? 46'b0000000000000000001000000001000010000000100000 : 46'b0000000000000100000000000001000010000000100010;
														assign node1352 = (inp[10]) ? 46'b0000000000000010000000000000000010000000100000 : 46'b0000000000000000001000000001000010000000100000;
											assign node1355 = (inp[7]) ? node1371 : node1356;
												assign node1356 = (inp[0]) ? node1364 : node1357;
													assign node1357 = (inp[14]) ? node1361 : node1358;
														assign node1358 = (inp[8]) ? 46'b0000000000100000000000000001100000000000100010 : 46'b0000000000100100000000000000100000000000100000;
														assign node1361 = (inp[8]) ? 46'b0000000000100010000000000000100000000000100000 : 46'b0000000000100000001000000001100000000000100000;
													assign node1364 = (inp[8]) ? node1368 : node1365;
														assign node1365 = (inp[10]) ? 46'b0000000000000100000000000000100000000000100000 : 46'b0000000000000100000000000000100000000000100000;
														assign node1368 = (inp[4]) ? 46'b0000000000000000001000000001100000000000100000 : 46'b0000000000000010000000000000100000000000100000;
												assign node1371 = (inp[0]) ? node1379 : node1372;
													assign node1372 = (inp[10]) ? node1376 : node1373;
														assign node1373 = (inp[4]) ? 46'b0000000000100000001000000001000000000000100000 : 46'b0000000000100100000000000000000000000000100000;
														assign node1376 = (inp[4]) ? 46'b0000000000100010000000000000000000000000100000 : 46'b0000000000100000000000000001000000000000100010;
													assign node1379 = (inp[10]) ? node1383 : node1380;
														assign node1380 = (inp[4]) ? 46'b0000000000000000001000000001000000000000100000 : 46'b0000000000000100000000000000000000000000100000;
														assign node1383 = (inp[4]) ? 46'b0000000000000010000000000001000000000000100000 : 46'b0000000000000000000000000001000000000000100010;
							assign node1386 = (inp[7]) ? node1424 : node1387;
								assign node1387 = (inp[5]) ? node1399 : node1388;
									assign node1388 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1389;
										assign node1389 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1390;
											assign node1390 = (inp[6]) ? node1394 : node1391;
												assign node1391 = (inp[12]) ? 46'b0001000000100000001000000001100000100000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1394 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000100010000000000000100010000000100000;
									assign node1399 = (inp[9]) ? node1415 : node1400;
										assign node1400 = (inp[0]) ? node1408 : node1401;
											assign node1401 = (inp[12]) ? node1405 : node1402;
												assign node1402 = (inp[6]) ? 46'b0000000000100010000000000000100010000000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1405 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000100000001000000001100000100000100000;
											assign node1408 = (inp[6]) ? node1412 : node1409;
												assign node1409 = (inp[12]) ? 46'b0000000010000000000000000001100000100000000010 : 46'b0000000010000000000000000001100010100000000010;
												assign node1412 = (inp[12]) ? 46'b0000000010000000000000000001100000000000000010 : 46'b0000000010000000000000000001100010000000000010;
										assign node1415 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1416;
											assign node1416 = (inp[12]) ? node1420 : node1417;
												assign node1417 = (inp[6]) ? 46'b0000000010000000000000000001100010000001000010 : 46'b0000000010000000000000000001100010100001000010;
												assign node1420 = (inp[6]) ? 46'b0000000010000000000000000001100000000001000010 : 46'b0000000010000000000000000001100000100001000010;
								assign node1424 = (inp[5]) ? node1450 : node1425;
									assign node1425 = (inp[0]) ? node1441 : node1426;
										assign node1426 = (inp[9]) ? node1434 : node1427;
											assign node1427 = (inp[6]) ? node1431 : node1428;
												assign node1428 = (inp[12]) ? 46'b0001000000100000001000000001000000100000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1431 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000100010000000000000000010000000100000;
											assign node1434 = (inp[12]) ? node1438 : node1435;
												assign node1435 = (inp[6]) ? 46'b0001000010000100000000000000000010000001000000 : 46'b0001000010000100000000000000000010100001000000;
												assign node1438 = (inp[6]) ? 46'b0001000010000100000000000000000000000001000000 : 46'b0001000010000100000000000000000000100001000000;
										assign node1441 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1442;
											assign node1442 = (inp[12]) ? node1446 : node1443;
												assign node1443 = (inp[6]) ? 46'b0001000010000100000000000000000010000000000000 : 46'b0001000010000100000000000000000010100000000000;
												assign node1446 = (inp[6]) ? 46'b0001000010000100000000000000000000000000000000 : 46'b0001000010000100000000000000000000100000000000;
									assign node1450 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1451;
										assign node1451 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1452;
											assign node1452 = (inp[12]) ? node1456 : node1453;
												assign node1453 = (inp[6]) ? 46'b0000000000100010000000000000000010000000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1456 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000100000001000000001000000100000100000;

endmodule