module dtc_split5_bm96 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node15;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node170;
	wire [3-1:0] node172;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node198;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node205;

	assign outp = (inp[6]) ? node2 : 3'b000;
		assign node2 = (inp[7]) ? node20 : node3;
			assign node3 = (inp[3]) ? node5 : 3'b000;
				assign node5 = (inp[1]) ? node7 : 3'b000;
					assign node7 = (inp[5]) ? 3'b000 : node8;
						assign node8 = (inp[10]) ? 3'b000 : node9;
							assign node9 = (inp[2]) ? node11 : 3'b000;
								assign node11 = (inp[8]) ? node13 : 3'b000;
									assign node13 = (inp[4]) ? node15 : 3'b000;
										assign node15 = (inp[9]) ? 3'b000 : 3'b100;
			assign node20 = (inp[3]) ? node104 : node21;
				assign node21 = (inp[4]) ? node33 : node22;
					assign node22 = (inp[9]) ? node24 : 3'b011;
						assign node24 = (inp[1]) ? 3'b011 : node25;
							assign node25 = (inp[10]) ? node29 : node26;
								assign node26 = (inp[5]) ? 3'b011 : 3'b111;
								assign node29 = (inp[5]) ? 3'b101 : 3'b011;
					assign node33 = (inp[0]) ? node81 : node34;
						assign node34 = (inp[1]) ? node72 : node35;
							assign node35 = (inp[5]) ? node53 : node36;
								assign node36 = (inp[10]) ? node48 : node37;
									assign node37 = (inp[11]) ? node43 : node38;
										assign node38 = (inp[9]) ? 3'b010 : node39;
											assign node39 = (inp[8]) ? 3'b010 : 3'b001;
										assign node43 = (inp[9]) ? 3'b001 : node44;
											assign node44 = (inp[2]) ? 3'b001 : 3'b010;
									assign node48 = (inp[9]) ? 3'b001 : node49;
										assign node49 = (inp[8]) ? 3'b001 : 3'b010;
								assign node53 = (inp[10]) ? node67 : node54;
									assign node54 = (inp[8]) ? node60 : node55;
										assign node55 = (inp[11]) ? node57 : 3'b001;
											assign node57 = (inp[9]) ? 3'b001 : 3'b010;
										assign node60 = (inp[11]) ? node62 : 3'b010;
											assign node62 = (inp[9]) ? 3'b001 : node63;
												assign node63 = (inp[2]) ? 3'b001 : 3'b010;
									assign node67 = (inp[11]) ? 3'b010 : node68;
										assign node68 = (inp[2]) ? 3'b010 : 3'b001;
							assign node72 = (inp[9]) ? node74 : 3'b010;
								assign node74 = (inp[8]) ? node76 : 3'b010;
									assign node76 = (inp[5]) ? node78 : 3'b010;
										assign node78 = (inp[10]) ? 3'b001 : 3'b010;
						assign node81 = (inp[9]) ? node89 : node82;
							assign node82 = (inp[11]) ? 3'b001 : node83;
								assign node83 = (inp[1]) ? node85 : 3'b001;
									assign node85 = (inp[8]) ? 3'b001 : 3'b010;
							assign node89 = (inp[1]) ? 3'b010 : node90;
								assign node90 = (inp[11]) ? node96 : node91;
									assign node91 = (inp[10]) ? node93 : 3'b110;
										assign node93 = (inp[5]) ? 3'b001 : 3'b101;
									assign node96 = (inp[10]) ? node98 : 3'b001;
										assign node98 = (inp[5]) ? node100 : 3'b001;
											assign node100 = (inp[8]) ? 3'b110 : 3'b010;
				assign node104 = (inp[1]) ? node166 : node105;
					assign node105 = (inp[4]) ? node127 : node106;
						assign node106 = (inp[9]) ? node112 : node107;
							assign node107 = (inp[10]) ? node109 : 3'b111;
								assign node109 = (inp[0]) ? 3'b111 : 3'b110;
							assign node112 = (inp[0]) ? node120 : node113;
								assign node113 = (inp[10]) ? node117 : node114;
									assign node114 = (inp[11]) ? 3'b111 : 3'b110;
									assign node117 = (inp[5]) ? 3'b011 : 3'b111;
								assign node120 = (inp[10]) ? node124 : node121;
									assign node121 = (inp[11]) ? 3'b110 : 3'b111;
									assign node124 = (inp[5]) ? 3'b010 : 3'b110;
						assign node127 = (inp[0]) ? node149 : node128;
							assign node128 = (inp[9]) ? node140 : node129;
								assign node129 = (inp[10]) ? node135 : node130;
									assign node130 = (inp[11]) ? node132 : 3'b111;
										assign node132 = (inp[8]) ? 3'b111 : 3'b011;
									assign node135 = (inp[11]) ? 3'b001 : node136;
										assign node136 = (inp[8]) ? 3'b101 : 3'b001;
								assign node140 = (inp[10]) ? node144 : node141;
									assign node141 = (inp[11]) ? 3'b110 : 3'b001;
									assign node144 = (inp[11]) ? node146 : 3'b110;
										assign node146 = (inp[5]) ? 3'b010 : 3'b110;
							assign node149 = (inp[9]) ? node157 : node150;
								assign node150 = (inp[8]) ? node152 : 3'b110;
									assign node152 = (inp[2]) ? 3'b110 : node153;
										assign node153 = (inp[5]) ? 3'b010 : 3'b110;
								assign node157 = (inp[11]) ? node161 : node158;
									assign node158 = (inp[10]) ? 3'b100 : 3'b010;
									assign node161 = (inp[5]) ? node163 : 3'b100;
										assign node163 = (inp[10]) ? 3'b000 : 3'b100;
					assign node166 = (inp[4]) ? node186 : node167;
						assign node167 = (inp[0]) ? node177 : node168;
							assign node168 = (inp[9]) ? node170 : 3'b100;
								assign node170 = (inp[5]) ? node172 : 3'b101;
									assign node172 = (inp[11]) ? node174 : 3'b101;
										assign node174 = (inp[10]) ? 3'b100 : 3'b101;
							assign node177 = (inp[9]) ? 3'b100 : node178;
								assign node178 = (inp[11]) ? 3'b100 : node179;
									assign node179 = (inp[10]) ? node181 : 3'b101;
										assign node181 = (inp[8]) ? 3'b101 : 3'b100;
						assign node186 = (inp[0]) ? node190 : node187;
							assign node187 = (inp[9]) ? 3'b010 : 3'b001;
							assign node190 = (inp[9]) ? node202 : node191;
								assign node191 = (inp[11]) ? 3'b100 : node192;
									assign node192 = (inp[5]) ? node198 : node193;
										assign node193 = (inp[10]) ? 3'b010 : node194;
											assign node194 = (inp[8]) ? 3'b110 : 3'b010;
										assign node198 = (inp[10]) ? 3'b100 : 3'b010;
								assign node202 = (inp[8]) ? node204 : 3'b000;
									assign node204 = (inp[10]) ? 3'b000 : node205;
										assign node205 = (inp[11]) ? 3'b000 : 3'b100;

endmodule