module dtc_split5_bm25 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node5;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node10;
	wire [14-1:0] node11;
	wire [14-1:0] node15;
	wire [14-1:0] node16;
	wire [14-1:0] node19;
	wire [14-1:0] node22;
	wire [14-1:0] node23;
	wire [14-1:0] node24;
	wire [14-1:0] node27;
	wire [14-1:0] node30;
	wire [14-1:0] node31;
	wire [14-1:0] node34;
	wire [14-1:0] node37;
	wire [14-1:0] node38;
	wire [14-1:0] node39;
	wire [14-1:0] node40;
	wire [14-1:0] node43;
	wire [14-1:0] node46;
	wire [14-1:0] node47;
	wire [14-1:0] node50;
	wire [14-1:0] node53;
	wire [14-1:0] node54;
	wire [14-1:0] node55;
	wire [14-1:0] node58;
	wire [14-1:0] node61;
	wire [14-1:0] node63;
	wire [14-1:0] node66;
	wire [14-1:0] node67;
	wire [14-1:0] node68;
	wire [14-1:0] node69;
	wire [14-1:0] node70;
	wire [14-1:0] node73;
	wire [14-1:0] node76;
	wire [14-1:0] node77;
	wire [14-1:0] node80;
	wire [14-1:0] node83;
	wire [14-1:0] node84;
	wire [14-1:0] node85;
	wire [14-1:0] node88;
	wire [14-1:0] node91;
	wire [14-1:0] node93;
	wire [14-1:0] node96;
	wire [14-1:0] node97;
	wire [14-1:0] node98;
	wire [14-1:0] node99;
	wire [14-1:0] node102;
	wire [14-1:0] node105;
	wire [14-1:0] node106;
	wire [14-1:0] node109;
	wire [14-1:0] node112;
	wire [14-1:0] node113;
	wire [14-1:0] node114;
	wire [14-1:0] node117;
	wire [14-1:0] node120;
	wire [14-1:0] node121;
	wire [14-1:0] node124;
	wire [14-1:0] node127;
	wire [14-1:0] node128;
	wire [14-1:0] node129;
	wire [14-1:0] node130;
	wire [14-1:0] node131;
	wire [14-1:0] node132;
	wire [14-1:0] node135;
	wire [14-1:0] node138;
	wire [14-1:0] node139;
	wire [14-1:0] node142;
	wire [14-1:0] node145;
	wire [14-1:0] node146;
	wire [14-1:0] node147;
	wire [14-1:0] node150;
	wire [14-1:0] node153;
	wire [14-1:0] node155;
	wire [14-1:0] node158;
	wire [14-1:0] node159;
	wire [14-1:0] node160;
	wire [14-1:0] node161;
	wire [14-1:0] node164;
	wire [14-1:0] node167;
	wire [14-1:0] node168;
	wire [14-1:0] node171;
	wire [14-1:0] node174;
	wire [14-1:0] node175;
	wire [14-1:0] node176;
	wire [14-1:0] node179;
	wire [14-1:0] node182;
	wire [14-1:0] node183;
	wire [14-1:0] node186;
	wire [14-1:0] node189;
	wire [14-1:0] node190;
	wire [14-1:0] node191;
	wire [14-1:0] node192;
	wire [14-1:0] node193;
	wire [14-1:0] node196;
	wire [14-1:0] node199;
	wire [14-1:0] node200;
	wire [14-1:0] node203;
	wire [14-1:0] node206;
	wire [14-1:0] node207;
	wire [14-1:0] node208;
	wire [14-1:0] node211;
	wire [14-1:0] node214;
	wire [14-1:0] node215;
	wire [14-1:0] node218;
	wire [14-1:0] node221;
	wire [14-1:0] node222;
	wire [14-1:0] node223;
	wire [14-1:0] node225;
	wire [14-1:0] node228;
	wire [14-1:0] node229;
	wire [14-1:0] node232;
	wire [14-1:0] node235;
	wire [14-1:0] node236;
	wire [14-1:0] node238;
	wire [14-1:0] node241;
	wire [14-1:0] node242;
	wire [14-1:0] node245;
	wire [14-1:0] node248;
	wire [14-1:0] node249;
	wire [14-1:0] node250;
	wire [14-1:0] node251;
	wire [14-1:0] node252;
	wire [14-1:0] node253;
	wire [14-1:0] node255;
	wire [14-1:0] node258;
	wire [14-1:0] node259;
	wire [14-1:0] node262;
	wire [14-1:0] node265;
	wire [14-1:0] node266;
	wire [14-1:0] node267;
	wire [14-1:0] node270;
	wire [14-1:0] node273;
	wire [14-1:0] node274;
	wire [14-1:0] node278;
	wire [14-1:0] node279;
	wire [14-1:0] node280;
	wire [14-1:0] node281;
	wire [14-1:0] node284;
	wire [14-1:0] node287;
	wire [14-1:0] node288;
	wire [14-1:0] node291;
	wire [14-1:0] node294;
	wire [14-1:0] node295;
	wire [14-1:0] node296;
	wire [14-1:0] node300;
	wire [14-1:0] node301;
	wire [14-1:0] node304;
	wire [14-1:0] node307;
	wire [14-1:0] node308;
	wire [14-1:0] node309;
	wire [14-1:0] node310;
	wire [14-1:0] node311;
	wire [14-1:0] node314;
	wire [14-1:0] node317;
	wire [14-1:0] node318;
	wire [14-1:0] node321;
	wire [14-1:0] node324;
	wire [14-1:0] node325;
	wire [14-1:0] node326;
	wire [14-1:0] node329;
	wire [14-1:0] node332;
	wire [14-1:0] node333;
	wire [14-1:0] node336;
	wire [14-1:0] node339;
	wire [14-1:0] node340;
	wire [14-1:0] node341;
	wire [14-1:0] node342;
	wire [14-1:0] node345;
	wire [14-1:0] node348;
	wire [14-1:0] node349;
	wire [14-1:0] node352;
	wire [14-1:0] node355;
	wire [14-1:0] node356;
	wire [14-1:0] node357;
	wire [14-1:0] node360;
	wire [14-1:0] node363;
	wire [14-1:0] node365;
	wire [14-1:0] node368;
	wire [14-1:0] node369;
	wire [14-1:0] node370;
	wire [14-1:0] node371;
	wire [14-1:0] node372;
	wire [14-1:0] node373;
	wire [14-1:0] node376;
	wire [14-1:0] node379;
	wire [14-1:0] node380;
	wire [14-1:0] node383;
	wire [14-1:0] node386;
	wire [14-1:0] node387;
	wire [14-1:0] node388;
	wire [14-1:0] node391;
	wire [14-1:0] node394;
	wire [14-1:0] node395;
	wire [14-1:0] node398;
	wire [14-1:0] node401;
	wire [14-1:0] node402;
	wire [14-1:0] node403;
	wire [14-1:0] node404;
	wire [14-1:0] node407;
	wire [14-1:0] node410;
	wire [14-1:0] node411;
	wire [14-1:0] node414;
	wire [14-1:0] node417;
	wire [14-1:0] node418;
	wire [14-1:0] node419;
	wire [14-1:0] node422;
	wire [14-1:0] node425;
	wire [14-1:0] node426;
	wire [14-1:0] node429;
	wire [14-1:0] node432;
	wire [14-1:0] node433;
	wire [14-1:0] node434;
	wire [14-1:0] node435;
	wire [14-1:0] node436;
	wire [14-1:0] node439;
	wire [14-1:0] node442;
	wire [14-1:0] node443;
	wire [14-1:0] node446;
	wire [14-1:0] node449;
	wire [14-1:0] node450;
	wire [14-1:0] node451;
	wire [14-1:0] node454;
	wire [14-1:0] node457;
	wire [14-1:0] node458;
	wire [14-1:0] node461;
	wire [14-1:0] node464;
	wire [14-1:0] node465;
	wire [14-1:0] node466;
	wire [14-1:0] node467;
	wire [14-1:0] node470;
	wire [14-1:0] node473;
	wire [14-1:0] node474;
	wire [14-1:0] node477;
	wire [14-1:0] node480;
	wire [14-1:0] node481;
	wire [14-1:0] node482;
	wire [14-1:0] node485;
	wire [14-1:0] node488;
	wire [14-1:0] node490;
	wire [14-1:0] node493;
	wire [14-1:0] node494;
	wire [14-1:0] node495;
	wire [14-1:0] node496;
	wire [14-1:0] node497;
	wire [14-1:0] node498;
	wire [14-1:0] node499;
	wire [14-1:0] node500;
	wire [14-1:0] node503;
	wire [14-1:0] node506;
	wire [14-1:0] node507;
	wire [14-1:0] node510;
	wire [14-1:0] node513;
	wire [14-1:0] node514;
	wire [14-1:0] node515;
	wire [14-1:0] node518;
	wire [14-1:0] node521;
	wire [14-1:0] node522;
	wire [14-1:0] node525;
	wire [14-1:0] node528;
	wire [14-1:0] node529;
	wire [14-1:0] node530;
	wire [14-1:0] node531;
	wire [14-1:0] node534;
	wire [14-1:0] node537;
	wire [14-1:0] node538;
	wire [14-1:0] node541;
	wire [14-1:0] node544;
	wire [14-1:0] node545;
	wire [14-1:0] node546;
	wire [14-1:0] node549;
	wire [14-1:0] node552;
	wire [14-1:0] node553;
	wire [14-1:0] node556;
	wire [14-1:0] node559;
	wire [14-1:0] node560;
	wire [14-1:0] node561;
	wire [14-1:0] node562;
	wire [14-1:0] node563;
	wire [14-1:0] node566;
	wire [14-1:0] node569;
	wire [14-1:0] node570;
	wire [14-1:0] node573;
	wire [14-1:0] node576;
	wire [14-1:0] node577;
	wire [14-1:0] node578;
	wire [14-1:0] node581;
	wire [14-1:0] node584;
	wire [14-1:0] node585;
	wire [14-1:0] node588;
	wire [14-1:0] node591;
	wire [14-1:0] node592;
	wire [14-1:0] node593;
	wire [14-1:0] node594;
	wire [14-1:0] node597;
	wire [14-1:0] node600;
	wire [14-1:0] node601;
	wire [14-1:0] node604;
	wire [14-1:0] node607;
	wire [14-1:0] node608;
	wire [14-1:0] node609;
	wire [14-1:0] node612;
	wire [14-1:0] node615;
	wire [14-1:0] node616;
	wire [14-1:0] node620;
	wire [14-1:0] node621;
	wire [14-1:0] node622;
	wire [14-1:0] node623;
	wire [14-1:0] node624;
	wire [14-1:0] node625;
	wire [14-1:0] node628;
	wire [14-1:0] node631;
	wire [14-1:0] node633;
	wire [14-1:0] node636;
	wire [14-1:0] node637;
	wire [14-1:0] node638;
	wire [14-1:0] node641;
	wire [14-1:0] node644;
	wire [14-1:0] node645;
	wire [14-1:0] node649;
	wire [14-1:0] node650;
	wire [14-1:0] node651;
	wire [14-1:0] node652;
	wire [14-1:0] node655;
	wire [14-1:0] node658;
	wire [14-1:0] node659;
	wire [14-1:0] node662;
	wire [14-1:0] node665;
	wire [14-1:0] node666;
	wire [14-1:0] node667;
	wire [14-1:0] node670;
	wire [14-1:0] node673;
	wire [14-1:0] node675;
	wire [14-1:0] node678;
	wire [14-1:0] node679;
	wire [14-1:0] node680;
	wire [14-1:0] node681;
	wire [14-1:0] node682;
	wire [14-1:0] node685;
	wire [14-1:0] node688;
	wire [14-1:0] node689;
	wire [14-1:0] node692;
	wire [14-1:0] node695;
	wire [14-1:0] node696;
	wire [14-1:0] node697;
	wire [14-1:0] node700;
	wire [14-1:0] node703;
	wire [14-1:0] node704;
	wire [14-1:0] node707;
	wire [14-1:0] node710;
	wire [14-1:0] node711;
	wire [14-1:0] node712;
	wire [14-1:0] node713;
	wire [14-1:0] node716;
	wire [14-1:0] node719;
	wire [14-1:0] node720;
	wire [14-1:0] node723;
	wire [14-1:0] node726;
	wire [14-1:0] node727;
	wire [14-1:0] node728;
	wire [14-1:0] node731;
	wire [14-1:0] node734;
	wire [14-1:0] node735;
	wire [14-1:0] node738;
	wire [14-1:0] node741;
	wire [14-1:0] node742;
	wire [14-1:0] node743;
	wire [14-1:0] node744;
	wire [14-1:0] node745;
	wire [14-1:0] node746;
	wire [14-1:0] node747;
	wire [14-1:0] node751;
	wire [14-1:0] node752;
	wire [14-1:0] node755;
	wire [14-1:0] node758;
	wire [14-1:0] node759;
	wire [14-1:0] node761;
	wire [14-1:0] node764;
	wire [14-1:0] node765;
	wire [14-1:0] node768;
	wire [14-1:0] node771;
	wire [14-1:0] node772;
	wire [14-1:0] node773;
	wire [14-1:0] node774;
	wire [14-1:0] node777;
	wire [14-1:0] node780;
	wire [14-1:0] node781;
	wire [14-1:0] node784;
	wire [14-1:0] node787;
	wire [14-1:0] node788;
	wire [14-1:0] node789;
	wire [14-1:0] node792;
	wire [14-1:0] node796;
	wire [14-1:0] node797;
	wire [14-1:0] node798;
	wire [14-1:0] node799;
	wire [14-1:0] node800;
	wire [14-1:0] node803;
	wire [14-1:0] node806;
	wire [14-1:0] node807;
	wire [14-1:0] node810;
	wire [14-1:0] node813;
	wire [14-1:0] node814;
	wire [14-1:0] node815;
	wire [14-1:0] node818;
	wire [14-1:0] node821;
	wire [14-1:0] node822;
	wire [14-1:0] node825;
	wire [14-1:0] node828;
	wire [14-1:0] node829;
	wire [14-1:0] node830;
	wire [14-1:0] node831;
	wire [14-1:0] node834;
	wire [14-1:0] node837;
	wire [14-1:0] node838;
	wire [14-1:0] node842;
	wire [14-1:0] node843;
	wire [14-1:0] node844;
	wire [14-1:0] node847;
	wire [14-1:0] node850;
	wire [14-1:0] node851;
	wire [14-1:0] node854;
	wire [14-1:0] node857;
	wire [14-1:0] node858;
	wire [14-1:0] node859;
	wire [14-1:0] node860;
	wire [14-1:0] node861;
	wire [14-1:0] node862;
	wire [14-1:0] node865;
	wire [14-1:0] node868;
	wire [14-1:0] node869;
	wire [14-1:0] node872;
	wire [14-1:0] node875;
	wire [14-1:0] node876;
	wire [14-1:0] node877;
	wire [14-1:0] node880;
	wire [14-1:0] node883;
	wire [14-1:0] node884;
	wire [14-1:0] node887;
	wire [14-1:0] node890;
	wire [14-1:0] node891;
	wire [14-1:0] node892;
	wire [14-1:0] node893;
	wire [14-1:0] node896;
	wire [14-1:0] node899;
	wire [14-1:0] node900;
	wire [14-1:0] node903;
	wire [14-1:0] node906;
	wire [14-1:0] node907;
	wire [14-1:0] node909;
	wire [14-1:0] node912;
	wire [14-1:0] node913;
	wire [14-1:0] node916;
	wire [14-1:0] node919;
	wire [14-1:0] node920;
	wire [14-1:0] node921;
	wire [14-1:0] node922;
	wire [14-1:0] node923;
	wire [14-1:0] node926;
	wire [14-1:0] node929;
	wire [14-1:0] node930;
	wire [14-1:0] node933;
	wire [14-1:0] node936;
	wire [14-1:0] node937;
	wire [14-1:0] node938;
	wire [14-1:0] node941;
	wire [14-1:0] node944;
	wire [14-1:0] node945;
	wire [14-1:0] node948;
	wire [14-1:0] node951;
	wire [14-1:0] node952;
	wire [14-1:0] node953;
	wire [14-1:0] node954;
	wire [14-1:0] node957;
	wire [14-1:0] node960;
	wire [14-1:0] node961;
	wire [14-1:0] node964;
	wire [14-1:0] node967;
	wire [14-1:0] node968;
	wire [14-1:0] node969;
	wire [14-1:0] node973;
	wire [14-1:0] node975;
	wire [14-1:0] node978;
	wire [14-1:0] node979;
	wire [14-1:0] node980;
	wire [14-1:0] node981;
	wire [14-1:0] node982;
	wire [14-1:0] node983;
	wire [14-1:0] node984;
	wire [14-1:0] node985;
	wire [14-1:0] node986;
	wire [14-1:0] node990;
	wire [14-1:0] node991;
	wire [14-1:0] node994;
	wire [14-1:0] node997;
	wire [14-1:0] node998;
	wire [14-1:0] node999;
	wire [14-1:0] node1002;
	wire [14-1:0] node1005;
	wire [14-1:0] node1006;
	wire [14-1:0] node1009;
	wire [14-1:0] node1012;
	wire [14-1:0] node1013;
	wire [14-1:0] node1014;
	wire [14-1:0] node1015;
	wire [14-1:0] node1019;
	wire [14-1:0] node1020;
	wire [14-1:0] node1023;
	wire [14-1:0] node1026;
	wire [14-1:0] node1027;
	wire [14-1:0] node1028;
	wire [14-1:0] node1031;
	wire [14-1:0] node1034;
	wire [14-1:0] node1035;
	wire [14-1:0] node1038;
	wire [14-1:0] node1041;
	wire [14-1:0] node1042;
	wire [14-1:0] node1043;
	wire [14-1:0] node1044;
	wire [14-1:0] node1045;
	wire [14-1:0] node1049;
	wire [14-1:0] node1050;
	wire [14-1:0] node1053;
	wire [14-1:0] node1056;
	wire [14-1:0] node1057;
	wire [14-1:0] node1059;
	wire [14-1:0] node1062;
	wire [14-1:0] node1063;
	wire [14-1:0] node1066;
	wire [14-1:0] node1069;
	wire [14-1:0] node1070;
	wire [14-1:0] node1071;
	wire [14-1:0] node1072;
	wire [14-1:0] node1075;
	wire [14-1:0] node1078;
	wire [14-1:0] node1079;
	wire [14-1:0] node1082;
	wire [14-1:0] node1085;
	wire [14-1:0] node1086;
	wire [14-1:0] node1087;
	wire [14-1:0] node1090;
	wire [14-1:0] node1093;
	wire [14-1:0] node1094;
	wire [14-1:0] node1097;
	wire [14-1:0] node1100;
	wire [14-1:0] node1101;
	wire [14-1:0] node1102;
	wire [14-1:0] node1103;
	wire [14-1:0] node1104;
	wire [14-1:0] node1105;
	wire [14-1:0] node1108;
	wire [14-1:0] node1111;
	wire [14-1:0] node1112;
	wire [14-1:0] node1116;
	wire [14-1:0] node1117;
	wire [14-1:0] node1118;
	wire [14-1:0] node1121;
	wire [14-1:0] node1124;
	wire [14-1:0] node1125;
	wire [14-1:0] node1128;
	wire [14-1:0] node1131;
	wire [14-1:0] node1132;
	wire [14-1:0] node1133;
	wire [14-1:0] node1135;
	wire [14-1:0] node1138;
	wire [14-1:0] node1139;
	wire [14-1:0] node1143;
	wire [14-1:0] node1144;
	wire [14-1:0] node1145;
	wire [14-1:0] node1148;
	wire [14-1:0] node1151;
	wire [14-1:0] node1152;
	wire [14-1:0] node1155;
	wire [14-1:0] node1158;
	wire [14-1:0] node1159;
	wire [14-1:0] node1160;
	wire [14-1:0] node1161;
	wire [14-1:0] node1162;
	wire [14-1:0] node1165;
	wire [14-1:0] node1168;
	wire [14-1:0] node1169;
	wire [14-1:0] node1172;
	wire [14-1:0] node1175;
	wire [14-1:0] node1176;
	wire [14-1:0] node1177;
	wire [14-1:0] node1180;
	wire [14-1:0] node1183;
	wire [14-1:0] node1184;
	wire [14-1:0] node1187;
	wire [14-1:0] node1190;
	wire [14-1:0] node1191;
	wire [14-1:0] node1192;
	wire [14-1:0] node1193;
	wire [14-1:0] node1196;
	wire [14-1:0] node1199;
	wire [14-1:0] node1200;
	wire [14-1:0] node1203;
	wire [14-1:0] node1206;
	wire [14-1:0] node1207;
	wire [14-1:0] node1208;
	wire [14-1:0] node1211;
	wire [14-1:0] node1214;
	wire [14-1:0] node1215;
	wire [14-1:0] node1219;
	wire [14-1:0] node1220;
	wire [14-1:0] node1221;
	wire [14-1:0] node1222;
	wire [14-1:0] node1223;
	wire [14-1:0] node1224;
	wire [14-1:0] node1225;
	wire [14-1:0] node1228;
	wire [14-1:0] node1231;
	wire [14-1:0] node1232;
	wire [14-1:0] node1236;
	wire [14-1:0] node1237;
	wire [14-1:0] node1238;
	wire [14-1:0] node1241;
	wire [14-1:0] node1244;
	wire [14-1:0] node1245;
	wire [14-1:0] node1248;
	wire [14-1:0] node1251;
	wire [14-1:0] node1252;
	wire [14-1:0] node1253;
	wire [14-1:0] node1254;
	wire [14-1:0] node1257;
	wire [14-1:0] node1260;
	wire [14-1:0] node1261;
	wire [14-1:0] node1264;
	wire [14-1:0] node1267;
	wire [14-1:0] node1268;
	wire [14-1:0] node1269;
	wire [14-1:0] node1272;
	wire [14-1:0] node1275;
	wire [14-1:0] node1276;
	wire [14-1:0] node1279;
	wire [14-1:0] node1282;
	wire [14-1:0] node1283;
	wire [14-1:0] node1284;
	wire [14-1:0] node1285;
	wire [14-1:0] node1286;
	wire [14-1:0] node1289;
	wire [14-1:0] node1292;
	wire [14-1:0] node1293;
	wire [14-1:0] node1297;
	wire [14-1:0] node1298;
	wire [14-1:0] node1299;
	wire [14-1:0] node1302;
	wire [14-1:0] node1305;
	wire [14-1:0] node1306;
	wire [14-1:0] node1309;
	wire [14-1:0] node1312;
	wire [14-1:0] node1313;
	wire [14-1:0] node1314;
	wire [14-1:0] node1315;
	wire [14-1:0] node1318;
	wire [14-1:0] node1321;
	wire [14-1:0] node1323;
	wire [14-1:0] node1326;
	wire [14-1:0] node1327;
	wire [14-1:0] node1328;
	wire [14-1:0] node1331;
	wire [14-1:0] node1334;
	wire [14-1:0] node1335;
	wire [14-1:0] node1338;
	wire [14-1:0] node1341;
	wire [14-1:0] node1342;
	wire [14-1:0] node1343;
	wire [14-1:0] node1344;
	wire [14-1:0] node1345;
	wire [14-1:0] node1346;
	wire [14-1:0] node1350;
	wire [14-1:0] node1351;
	wire [14-1:0] node1354;
	wire [14-1:0] node1357;
	wire [14-1:0] node1358;
	wire [14-1:0] node1360;
	wire [14-1:0] node1363;
	wire [14-1:0] node1364;
	wire [14-1:0] node1367;
	wire [14-1:0] node1370;
	wire [14-1:0] node1371;
	wire [14-1:0] node1372;
	wire [14-1:0] node1373;
	wire [14-1:0] node1376;
	wire [14-1:0] node1379;
	wire [14-1:0] node1380;
	wire [14-1:0] node1383;
	wire [14-1:0] node1386;
	wire [14-1:0] node1387;
	wire [14-1:0] node1388;
	wire [14-1:0] node1391;
	wire [14-1:0] node1394;
	wire [14-1:0] node1395;
	wire [14-1:0] node1398;
	wire [14-1:0] node1401;
	wire [14-1:0] node1402;
	wire [14-1:0] node1403;
	wire [14-1:0] node1404;
	wire [14-1:0] node1406;
	wire [14-1:0] node1409;
	wire [14-1:0] node1410;
	wire [14-1:0] node1413;
	wire [14-1:0] node1416;
	wire [14-1:0] node1417;
	wire [14-1:0] node1418;
	wire [14-1:0] node1422;
	wire [14-1:0] node1425;
	wire [14-1:0] node1426;
	wire [14-1:0] node1427;
	wire [14-1:0] node1429;
	wire [14-1:0] node1432;
	wire [14-1:0] node1433;
	wire [14-1:0] node1436;
	wire [14-1:0] node1439;
	wire [14-1:0] node1440;
	wire [14-1:0] node1441;
	wire [14-1:0] node1444;
	wire [14-1:0] node1447;
	wire [14-1:0] node1448;
	wire [14-1:0] node1451;
	wire [14-1:0] node1454;
	wire [14-1:0] node1455;
	wire [14-1:0] node1456;
	wire [14-1:0] node1457;
	wire [14-1:0] node1458;
	wire [14-1:0] node1459;
	wire [14-1:0] node1460;
	wire [14-1:0] node1461;
	wire [14-1:0] node1464;
	wire [14-1:0] node1467;
	wire [14-1:0] node1468;
	wire [14-1:0] node1472;
	wire [14-1:0] node1473;
	wire [14-1:0] node1474;
	wire [14-1:0] node1477;
	wire [14-1:0] node1480;
	wire [14-1:0] node1481;
	wire [14-1:0] node1484;
	wire [14-1:0] node1487;
	wire [14-1:0] node1488;
	wire [14-1:0] node1489;
	wire [14-1:0] node1490;
	wire [14-1:0] node1493;
	wire [14-1:0] node1496;
	wire [14-1:0] node1497;
	wire [14-1:0] node1500;
	wire [14-1:0] node1503;
	wire [14-1:0] node1504;
	wire [14-1:0] node1505;
	wire [14-1:0] node1508;
	wire [14-1:0] node1511;
	wire [14-1:0] node1512;
	wire [14-1:0] node1515;
	wire [14-1:0] node1518;
	wire [14-1:0] node1519;
	wire [14-1:0] node1520;
	wire [14-1:0] node1521;
	wire [14-1:0] node1522;
	wire [14-1:0] node1526;
	wire [14-1:0] node1527;
	wire [14-1:0] node1530;
	wire [14-1:0] node1533;
	wire [14-1:0] node1534;
	wire [14-1:0] node1535;
	wire [14-1:0] node1538;
	wire [14-1:0] node1541;
	wire [14-1:0] node1542;
	wire [14-1:0] node1545;
	wire [14-1:0] node1548;
	wire [14-1:0] node1549;
	wire [14-1:0] node1550;
	wire [14-1:0] node1551;
	wire [14-1:0] node1554;
	wire [14-1:0] node1557;
	wire [14-1:0] node1558;
	wire [14-1:0] node1561;
	wire [14-1:0] node1564;
	wire [14-1:0] node1565;
	wire [14-1:0] node1567;
	wire [14-1:0] node1570;
	wire [14-1:0] node1571;
	wire [14-1:0] node1574;
	wire [14-1:0] node1577;
	wire [14-1:0] node1578;
	wire [14-1:0] node1579;
	wire [14-1:0] node1580;
	wire [14-1:0] node1581;
	wire [14-1:0] node1582;
	wire [14-1:0] node1585;
	wire [14-1:0] node1588;
	wire [14-1:0] node1589;
	wire [14-1:0] node1592;
	wire [14-1:0] node1595;
	wire [14-1:0] node1596;
	wire [14-1:0] node1599;
	wire [14-1:0] node1600;
	wire [14-1:0] node1603;
	wire [14-1:0] node1606;
	wire [14-1:0] node1607;
	wire [14-1:0] node1608;
	wire [14-1:0] node1609;
	wire [14-1:0] node1612;
	wire [14-1:0] node1615;
	wire [14-1:0] node1616;
	wire [14-1:0] node1619;
	wire [14-1:0] node1622;
	wire [14-1:0] node1623;
	wire [14-1:0] node1624;
	wire [14-1:0] node1627;
	wire [14-1:0] node1630;
	wire [14-1:0] node1631;
	wire [14-1:0] node1634;
	wire [14-1:0] node1637;
	wire [14-1:0] node1638;
	wire [14-1:0] node1639;
	wire [14-1:0] node1640;
	wire [14-1:0] node1641;
	wire [14-1:0] node1644;
	wire [14-1:0] node1647;
	wire [14-1:0] node1648;
	wire [14-1:0] node1651;
	wire [14-1:0] node1654;
	wire [14-1:0] node1655;
	wire [14-1:0] node1657;
	wire [14-1:0] node1660;
	wire [14-1:0] node1661;
	wire [14-1:0] node1664;
	wire [14-1:0] node1667;
	wire [14-1:0] node1668;
	wire [14-1:0] node1669;
	wire [14-1:0] node1670;
	wire [14-1:0] node1673;
	wire [14-1:0] node1676;
	wire [14-1:0] node1677;
	wire [14-1:0] node1680;
	wire [14-1:0] node1683;
	wire [14-1:0] node1684;
	wire [14-1:0] node1685;
	wire [14-1:0] node1688;
	wire [14-1:0] node1691;
	wire [14-1:0] node1692;
	wire [14-1:0] node1695;
	wire [14-1:0] node1698;
	wire [14-1:0] node1699;
	wire [14-1:0] node1700;
	wire [14-1:0] node1701;
	wire [14-1:0] node1702;
	wire [14-1:0] node1703;
	wire [14-1:0] node1704;
	wire [14-1:0] node1708;
	wire [14-1:0] node1709;
	wire [14-1:0] node1712;
	wire [14-1:0] node1715;
	wire [14-1:0] node1716;
	wire [14-1:0] node1717;
	wire [14-1:0] node1720;
	wire [14-1:0] node1723;
	wire [14-1:0] node1724;
	wire [14-1:0] node1727;
	wire [14-1:0] node1730;
	wire [14-1:0] node1731;
	wire [14-1:0] node1732;
	wire [14-1:0] node1733;
	wire [14-1:0] node1736;
	wire [14-1:0] node1739;
	wire [14-1:0] node1740;
	wire [14-1:0] node1743;
	wire [14-1:0] node1746;
	wire [14-1:0] node1747;
	wire [14-1:0] node1748;
	wire [14-1:0] node1751;
	wire [14-1:0] node1754;
	wire [14-1:0] node1755;
	wire [14-1:0] node1758;
	wire [14-1:0] node1761;
	wire [14-1:0] node1762;
	wire [14-1:0] node1763;
	wire [14-1:0] node1764;
	wire [14-1:0] node1765;
	wire [14-1:0] node1768;
	wire [14-1:0] node1771;
	wire [14-1:0] node1772;
	wire [14-1:0] node1775;
	wire [14-1:0] node1778;
	wire [14-1:0] node1779;
	wire [14-1:0] node1781;
	wire [14-1:0] node1784;
	wire [14-1:0] node1785;
	wire [14-1:0] node1789;
	wire [14-1:0] node1790;
	wire [14-1:0] node1791;
	wire [14-1:0] node1792;
	wire [14-1:0] node1795;
	wire [14-1:0] node1798;
	wire [14-1:0] node1799;
	wire [14-1:0] node1802;
	wire [14-1:0] node1805;
	wire [14-1:0] node1806;
	wire [14-1:0] node1807;
	wire [14-1:0] node1810;
	wire [14-1:0] node1813;
	wire [14-1:0] node1814;
	wire [14-1:0] node1818;
	wire [14-1:0] node1819;
	wire [14-1:0] node1820;
	wire [14-1:0] node1821;
	wire [14-1:0] node1822;
	wire [14-1:0] node1823;
	wire [14-1:0] node1826;
	wire [14-1:0] node1829;
	wire [14-1:0] node1830;
	wire [14-1:0] node1833;
	wire [14-1:0] node1836;
	wire [14-1:0] node1837;
	wire [14-1:0] node1838;
	wire [14-1:0] node1841;
	wire [14-1:0] node1844;
	wire [14-1:0] node1845;
	wire [14-1:0] node1848;
	wire [14-1:0] node1851;
	wire [14-1:0] node1852;
	wire [14-1:0] node1853;
	wire [14-1:0] node1854;
	wire [14-1:0] node1858;
	wire [14-1:0] node1859;
	wire [14-1:0] node1862;
	wire [14-1:0] node1865;
	wire [14-1:0] node1866;
	wire [14-1:0] node1867;
	wire [14-1:0] node1870;
	wire [14-1:0] node1873;
	wire [14-1:0] node1874;
	wire [14-1:0] node1877;
	wire [14-1:0] node1880;
	wire [14-1:0] node1881;
	wire [14-1:0] node1882;
	wire [14-1:0] node1883;
	wire [14-1:0] node1884;
	wire [14-1:0] node1887;
	wire [14-1:0] node1890;
	wire [14-1:0] node1891;
	wire [14-1:0] node1895;
	wire [14-1:0] node1896;
	wire [14-1:0] node1897;
	wire [14-1:0] node1900;
	wire [14-1:0] node1903;
	wire [14-1:0] node1904;
	wire [14-1:0] node1907;
	wire [14-1:0] node1910;
	wire [14-1:0] node1911;
	wire [14-1:0] node1912;
	wire [14-1:0] node1913;
	wire [14-1:0] node1916;
	wire [14-1:0] node1919;
	wire [14-1:0] node1920;
	wire [14-1:0] node1923;
	wire [14-1:0] node1926;
	wire [14-1:0] node1927;
	wire [14-1:0] node1928;
	wire [14-1:0] node1931;
	wire [14-1:0] node1934;
	wire [14-1:0] node1935;
	wire [14-1:0] node1938;
	wire [14-1:0] node1941;
	wire [14-1:0] node1942;
	wire [14-1:0] node1943;
	wire [14-1:0] node1944;
	wire [14-1:0] node1945;
	wire [14-1:0] node1946;
	wire [14-1:0] node1947;
	wire [14-1:0] node1948;
	wire [14-1:0] node1949;
	wire [14-1:0] node1950;
	wire [14-1:0] node1953;
	wire [14-1:0] node1956;
	wire [14-1:0] node1957;
	wire [14-1:0] node1961;
	wire [14-1:0] node1962;
	wire [14-1:0] node1963;
	wire [14-1:0] node1966;
	wire [14-1:0] node1969;
	wire [14-1:0] node1970;
	wire [14-1:0] node1973;
	wire [14-1:0] node1976;
	wire [14-1:0] node1977;
	wire [14-1:0] node1978;
	wire [14-1:0] node1979;
	wire [14-1:0] node1982;
	wire [14-1:0] node1985;
	wire [14-1:0] node1986;
	wire [14-1:0] node1989;
	wire [14-1:0] node1992;
	wire [14-1:0] node1993;
	wire [14-1:0] node1995;
	wire [14-1:0] node1998;
	wire [14-1:0] node1999;
	wire [14-1:0] node2002;
	wire [14-1:0] node2005;
	wire [14-1:0] node2006;
	wire [14-1:0] node2007;
	wire [14-1:0] node2008;
	wire [14-1:0] node2009;
	wire [14-1:0] node2012;
	wire [14-1:0] node2015;
	wire [14-1:0] node2016;
	wire [14-1:0] node2019;
	wire [14-1:0] node2022;
	wire [14-1:0] node2023;
	wire [14-1:0] node2024;
	wire [14-1:0] node2027;
	wire [14-1:0] node2030;
	wire [14-1:0] node2031;
	wire [14-1:0] node2034;
	wire [14-1:0] node2037;
	wire [14-1:0] node2038;
	wire [14-1:0] node2039;
	wire [14-1:0] node2040;
	wire [14-1:0] node2043;
	wire [14-1:0] node2046;
	wire [14-1:0] node2047;
	wire [14-1:0] node2050;
	wire [14-1:0] node2053;
	wire [14-1:0] node2054;
	wire [14-1:0] node2055;
	wire [14-1:0] node2058;
	wire [14-1:0] node2061;
	wire [14-1:0] node2062;
	wire [14-1:0] node2065;
	wire [14-1:0] node2068;
	wire [14-1:0] node2069;
	wire [14-1:0] node2070;
	wire [14-1:0] node2071;
	wire [14-1:0] node2072;
	wire [14-1:0] node2073;
	wire [14-1:0] node2076;
	wire [14-1:0] node2079;
	wire [14-1:0] node2080;
	wire [14-1:0] node2083;
	wire [14-1:0] node2086;
	wire [14-1:0] node2087;
	wire [14-1:0] node2088;
	wire [14-1:0] node2091;
	wire [14-1:0] node2094;
	wire [14-1:0] node2095;
	wire [14-1:0] node2098;
	wire [14-1:0] node2101;
	wire [14-1:0] node2102;
	wire [14-1:0] node2103;
	wire [14-1:0] node2104;
	wire [14-1:0] node2107;
	wire [14-1:0] node2110;
	wire [14-1:0] node2111;
	wire [14-1:0] node2114;
	wire [14-1:0] node2117;
	wire [14-1:0] node2118;
	wire [14-1:0] node2119;
	wire [14-1:0] node2122;
	wire [14-1:0] node2125;
	wire [14-1:0] node2126;
	wire [14-1:0] node2129;
	wire [14-1:0] node2132;
	wire [14-1:0] node2133;
	wire [14-1:0] node2134;
	wire [14-1:0] node2135;
	wire [14-1:0] node2136;
	wire [14-1:0] node2139;
	wire [14-1:0] node2142;
	wire [14-1:0] node2143;
	wire [14-1:0] node2146;
	wire [14-1:0] node2149;
	wire [14-1:0] node2150;
	wire [14-1:0] node2151;
	wire [14-1:0] node2154;
	wire [14-1:0] node2157;
	wire [14-1:0] node2158;
	wire [14-1:0] node2162;
	wire [14-1:0] node2163;
	wire [14-1:0] node2164;
	wire [14-1:0] node2165;
	wire [14-1:0] node2168;
	wire [14-1:0] node2171;
	wire [14-1:0] node2172;
	wire [14-1:0] node2176;
	wire [14-1:0] node2177;
	wire [14-1:0] node2178;
	wire [14-1:0] node2181;
	wire [14-1:0] node2184;
	wire [14-1:0] node2185;
	wire [14-1:0] node2188;
	wire [14-1:0] node2191;
	wire [14-1:0] node2192;
	wire [14-1:0] node2193;
	wire [14-1:0] node2194;
	wire [14-1:0] node2195;
	wire [14-1:0] node2196;
	wire [14-1:0] node2197;
	wire [14-1:0] node2200;
	wire [14-1:0] node2203;
	wire [14-1:0] node2204;
	wire [14-1:0] node2207;
	wire [14-1:0] node2210;
	wire [14-1:0] node2211;
	wire [14-1:0] node2212;
	wire [14-1:0] node2215;
	wire [14-1:0] node2218;
	wire [14-1:0] node2219;
	wire [14-1:0] node2222;
	wire [14-1:0] node2225;
	wire [14-1:0] node2226;
	wire [14-1:0] node2227;
	wire [14-1:0] node2228;
	wire [14-1:0] node2232;
	wire [14-1:0] node2233;
	wire [14-1:0] node2236;
	wire [14-1:0] node2239;
	wire [14-1:0] node2240;
	wire [14-1:0] node2241;
	wire [14-1:0] node2244;
	wire [14-1:0] node2247;
	wire [14-1:0] node2248;
	wire [14-1:0] node2251;
	wire [14-1:0] node2254;
	wire [14-1:0] node2255;
	wire [14-1:0] node2256;
	wire [14-1:0] node2257;
	wire [14-1:0] node2258;
	wire [14-1:0] node2261;
	wire [14-1:0] node2264;
	wire [14-1:0] node2265;
	wire [14-1:0] node2268;
	wire [14-1:0] node2271;
	wire [14-1:0] node2272;
	wire [14-1:0] node2273;
	wire [14-1:0] node2276;
	wire [14-1:0] node2279;
	wire [14-1:0] node2280;
	wire [14-1:0] node2283;
	wire [14-1:0] node2286;
	wire [14-1:0] node2287;
	wire [14-1:0] node2288;
	wire [14-1:0] node2289;
	wire [14-1:0] node2292;
	wire [14-1:0] node2296;
	wire [14-1:0] node2297;
	wire [14-1:0] node2298;
	wire [14-1:0] node2302;
	wire [14-1:0] node2303;
	wire [14-1:0] node2306;
	wire [14-1:0] node2309;
	wire [14-1:0] node2310;
	wire [14-1:0] node2311;
	wire [14-1:0] node2312;
	wire [14-1:0] node2313;
	wire [14-1:0] node2314;
	wire [14-1:0] node2317;
	wire [14-1:0] node2320;
	wire [14-1:0] node2321;
	wire [14-1:0] node2324;
	wire [14-1:0] node2327;
	wire [14-1:0] node2328;
	wire [14-1:0] node2330;
	wire [14-1:0] node2333;
	wire [14-1:0] node2334;
	wire [14-1:0] node2337;
	wire [14-1:0] node2340;
	wire [14-1:0] node2341;
	wire [14-1:0] node2342;
	wire [14-1:0] node2343;
	wire [14-1:0] node2346;
	wire [14-1:0] node2349;
	wire [14-1:0] node2350;
	wire [14-1:0] node2353;
	wire [14-1:0] node2356;
	wire [14-1:0] node2357;
	wire [14-1:0] node2358;
	wire [14-1:0] node2361;
	wire [14-1:0] node2364;
	wire [14-1:0] node2365;
	wire [14-1:0] node2368;
	wire [14-1:0] node2371;
	wire [14-1:0] node2372;
	wire [14-1:0] node2373;
	wire [14-1:0] node2374;
	wire [14-1:0] node2375;
	wire [14-1:0] node2378;
	wire [14-1:0] node2381;
	wire [14-1:0] node2382;
	wire [14-1:0] node2385;
	wire [14-1:0] node2388;
	wire [14-1:0] node2389;
	wire [14-1:0] node2391;
	wire [14-1:0] node2394;
	wire [14-1:0] node2395;
	wire [14-1:0] node2398;
	wire [14-1:0] node2401;
	wire [14-1:0] node2402;
	wire [14-1:0] node2403;
	wire [14-1:0] node2405;
	wire [14-1:0] node2408;
	wire [14-1:0] node2409;
	wire [14-1:0] node2412;
	wire [14-1:0] node2415;
	wire [14-1:0] node2416;
	wire [14-1:0] node2417;
	wire [14-1:0] node2420;
	wire [14-1:0] node2423;
	wire [14-1:0] node2424;
	wire [14-1:0] node2427;
	wire [14-1:0] node2430;
	wire [14-1:0] node2431;
	wire [14-1:0] node2432;
	wire [14-1:0] node2433;
	wire [14-1:0] node2434;
	wire [14-1:0] node2435;
	wire [14-1:0] node2436;
	wire [14-1:0] node2437;
	wire [14-1:0] node2440;
	wire [14-1:0] node2443;
	wire [14-1:0] node2444;
	wire [14-1:0] node2447;
	wire [14-1:0] node2450;
	wire [14-1:0] node2451;
	wire [14-1:0] node2452;
	wire [14-1:0] node2456;
	wire [14-1:0] node2457;
	wire [14-1:0] node2461;
	wire [14-1:0] node2462;
	wire [14-1:0] node2463;
	wire [14-1:0] node2464;
	wire [14-1:0] node2467;
	wire [14-1:0] node2470;
	wire [14-1:0] node2471;
	wire [14-1:0] node2474;
	wire [14-1:0] node2477;
	wire [14-1:0] node2478;
	wire [14-1:0] node2479;
	wire [14-1:0] node2482;
	wire [14-1:0] node2485;
	wire [14-1:0] node2487;
	wire [14-1:0] node2490;
	wire [14-1:0] node2491;
	wire [14-1:0] node2492;
	wire [14-1:0] node2493;
	wire [14-1:0] node2494;
	wire [14-1:0] node2497;
	wire [14-1:0] node2500;
	wire [14-1:0] node2501;
	wire [14-1:0] node2504;
	wire [14-1:0] node2507;
	wire [14-1:0] node2509;
	wire [14-1:0] node2510;
	wire [14-1:0] node2513;
	wire [14-1:0] node2516;
	wire [14-1:0] node2517;
	wire [14-1:0] node2518;
	wire [14-1:0] node2519;
	wire [14-1:0] node2522;
	wire [14-1:0] node2525;
	wire [14-1:0] node2526;
	wire [14-1:0] node2529;
	wire [14-1:0] node2532;
	wire [14-1:0] node2533;
	wire [14-1:0] node2534;
	wire [14-1:0] node2537;
	wire [14-1:0] node2540;
	wire [14-1:0] node2541;
	wire [14-1:0] node2544;
	wire [14-1:0] node2547;
	wire [14-1:0] node2548;
	wire [14-1:0] node2549;
	wire [14-1:0] node2550;
	wire [14-1:0] node2551;
	wire [14-1:0] node2552;
	wire [14-1:0] node2555;
	wire [14-1:0] node2558;
	wire [14-1:0] node2559;
	wire [14-1:0] node2562;
	wire [14-1:0] node2565;
	wire [14-1:0] node2566;
	wire [14-1:0] node2568;
	wire [14-1:0] node2571;
	wire [14-1:0] node2572;
	wire [14-1:0] node2575;
	wire [14-1:0] node2578;
	wire [14-1:0] node2579;
	wire [14-1:0] node2580;
	wire [14-1:0] node2581;
	wire [14-1:0] node2584;
	wire [14-1:0] node2587;
	wire [14-1:0] node2588;
	wire [14-1:0] node2591;
	wire [14-1:0] node2594;
	wire [14-1:0] node2595;
	wire [14-1:0] node2597;
	wire [14-1:0] node2600;
	wire [14-1:0] node2601;
	wire [14-1:0] node2604;
	wire [14-1:0] node2607;
	wire [14-1:0] node2608;
	wire [14-1:0] node2609;
	wire [14-1:0] node2610;
	wire [14-1:0] node2611;
	wire [14-1:0] node2614;
	wire [14-1:0] node2617;
	wire [14-1:0] node2618;
	wire [14-1:0] node2621;
	wire [14-1:0] node2624;
	wire [14-1:0] node2625;
	wire [14-1:0] node2626;
	wire [14-1:0] node2629;
	wire [14-1:0] node2632;
	wire [14-1:0] node2633;
	wire [14-1:0] node2636;
	wire [14-1:0] node2639;
	wire [14-1:0] node2640;
	wire [14-1:0] node2641;
	wire [14-1:0] node2642;
	wire [14-1:0] node2645;
	wire [14-1:0] node2648;
	wire [14-1:0] node2649;
	wire [14-1:0] node2652;
	wire [14-1:0] node2655;
	wire [14-1:0] node2656;
	wire [14-1:0] node2657;
	wire [14-1:0] node2660;
	wire [14-1:0] node2663;
	wire [14-1:0] node2664;
	wire [14-1:0] node2667;
	wire [14-1:0] node2670;
	wire [14-1:0] node2671;
	wire [14-1:0] node2672;
	wire [14-1:0] node2673;
	wire [14-1:0] node2674;
	wire [14-1:0] node2675;
	wire [14-1:0] node2676;
	wire [14-1:0] node2679;
	wire [14-1:0] node2682;
	wire [14-1:0] node2683;
	wire [14-1:0] node2686;
	wire [14-1:0] node2689;
	wire [14-1:0] node2690;
	wire [14-1:0] node2691;
	wire [14-1:0] node2694;
	wire [14-1:0] node2697;
	wire [14-1:0] node2698;
	wire [14-1:0] node2701;
	wire [14-1:0] node2704;
	wire [14-1:0] node2705;
	wire [14-1:0] node2706;
	wire [14-1:0] node2707;
	wire [14-1:0] node2710;
	wire [14-1:0] node2713;
	wire [14-1:0] node2714;
	wire [14-1:0] node2717;
	wire [14-1:0] node2720;
	wire [14-1:0] node2721;
	wire [14-1:0] node2722;
	wire [14-1:0] node2725;
	wire [14-1:0] node2728;
	wire [14-1:0] node2729;
	wire [14-1:0] node2732;
	wire [14-1:0] node2735;
	wire [14-1:0] node2736;
	wire [14-1:0] node2737;
	wire [14-1:0] node2738;
	wire [14-1:0] node2740;
	wire [14-1:0] node2743;
	wire [14-1:0] node2744;
	wire [14-1:0] node2748;
	wire [14-1:0] node2749;
	wire [14-1:0] node2750;
	wire [14-1:0] node2753;
	wire [14-1:0] node2756;
	wire [14-1:0] node2757;
	wire [14-1:0] node2761;
	wire [14-1:0] node2762;
	wire [14-1:0] node2763;
	wire [14-1:0] node2764;
	wire [14-1:0] node2767;
	wire [14-1:0] node2770;
	wire [14-1:0] node2771;
	wire [14-1:0] node2774;
	wire [14-1:0] node2777;
	wire [14-1:0] node2778;
	wire [14-1:0] node2779;
	wire [14-1:0] node2782;
	wire [14-1:0] node2785;
	wire [14-1:0] node2786;
	wire [14-1:0] node2789;
	wire [14-1:0] node2792;
	wire [14-1:0] node2793;
	wire [14-1:0] node2794;
	wire [14-1:0] node2795;
	wire [14-1:0] node2796;
	wire [14-1:0] node2797;
	wire [14-1:0] node2800;
	wire [14-1:0] node2803;
	wire [14-1:0] node2804;
	wire [14-1:0] node2807;
	wire [14-1:0] node2810;
	wire [14-1:0] node2811;
	wire [14-1:0] node2812;
	wire [14-1:0] node2815;
	wire [14-1:0] node2818;
	wire [14-1:0] node2819;
	wire [14-1:0] node2822;
	wire [14-1:0] node2825;
	wire [14-1:0] node2826;
	wire [14-1:0] node2827;
	wire [14-1:0] node2828;
	wire [14-1:0] node2831;
	wire [14-1:0] node2834;
	wire [14-1:0] node2835;
	wire [14-1:0] node2838;
	wire [14-1:0] node2841;
	wire [14-1:0] node2842;
	wire [14-1:0] node2843;
	wire [14-1:0] node2846;
	wire [14-1:0] node2849;
	wire [14-1:0] node2851;
	wire [14-1:0] node2854;
	wire [14-1:0] node2855;
	wire [14-1:0] node2856;
	wire [14-1:0] node2857;
	wire [14-1:0] node2858;
	wire [14-1:0] node2861;
	wire [14-1:0] node2864;
	wire [14-1:0] node2865;
	wire [14-1:0] node2868;
	wire [14-1:0] node2871;
	wire [14-1:0] node2872;
	wire [14-1:0] node2873;
	wire [14-1:0] node2876;
	wire [14-1:0] node2879;
	wire [14-1:0] node2880;
	wire [14-1:0] node2883;
	wire [14-1:0] node2886;
	wire [14-1:0] node2887;
	wire [14-1:0] node2888;
	wire [14-1:0] node2890;
	wire [14-1:0] node2893;
	wire [14-1:0] node2894;
	wire [14-1:0] node2897;
	wire [14-1:0] node2900;
	wire [14-1:0] node2901;
	wire [14-1:0] node2902;
	wire [14-1:0] node2905;
	wire [14-1:0] node2908;
	wire [14-1:0] node2909;
	wire [14-1:0] node2912;
	wire [14-1:0] node2915;
	wire [14-1:0] node2916;
	wire [14-1:0] node2917;
	wire [14-1:0] node2918;
	wire [14-1:0] node2919;
	wire [14-1:0] node2920;
	wire [14-1:0] node2921;
	wire [14-1:0] node2922;
	wire [14-1:0] node2923;
	wire [14-1:0] node2926;
	wire [14-1:0] node2929;
	wire [14-1:0] node2930;
	wire [14-1:0] node2933;
	wire [14-1:0] node2936;
	wire [14-1:0] node2937;
	wire [14-1:0] node2938;
	wire [14-1:0] node2941;
	wire [14-1:0] node2944;
	wire [14-1:0] node2945;
	wire [14-1:0] node2948;
	wire [14-1:0] node2951;
	wire [14-1:0] node2952;
	wire [14-1:0] node2953;
	wire [14-1:0] node2954;
	wire [14-1:0] node2957;
	wire [14-1:0] node2960;
	wire [14-1:0] node2961;
	wire [14-1:0] node2964;
	wire [14-1:0] node2967;
	wire [14-1:0] node2968;
	wire [14-1:0] node2969;
	wire [14-1:0] node2972;
	wire [14-1:0] node2975;
	wire [14-1:0] node2976;
	wire [14-1:0] node2979;
	wire [14-1:0] node2982;
	wire [14-1:0] node2983;
	wire [14-1:0] node2984;
	wire [14-1:0] node2985;
	wire [14-1:0] node2986;
	wire [14-1:0] node2989;
	wire [14-1:0] node2992;
	wire [14-1:0] node2994;
	wire [14-1:0] node2997;
	wire [14-1:0] node2998;
	wire [14-1:0] node2999;
	wire [14-1:0] node3002;
	wire [14-1:0] node3005;
	wire [14-1:0] node3006;
	wire [14-1:0] node3009;
	wire [14-1:0] node3012;
	wire [14-1:0] node3013;
	wire [14-1:0] node3014;
	wire [14-1:0] node3016;
	wire [14-1:0] node3019;
	wire [14-1:0] node3020;
	wire [14-1:0] node3023;
	wire [14-1:0] node3026;
	wire [14-1:0] node3027;
	wire [14-1:0] node3028;
	wire [14-1:0] node3031;
	wire [14-1:0] node3034;
	wire [14-1:0] node3035;
	wire [14-1:0] node3038;
	wire [14-1:0] node3041;
	wire [14-1:0] node3042;
	wire [14-1:0] node3043;
	wire [14-1:0] node3044;
	wire [14-1:0] node3045;
	wire [14-1:0] node3046;
	wire [14-1:0] node3050;
	wire [14-1:0] node3051;
	wire [14-1:0] node3055;
	wire [14-1:0] node3056;
	wire [14-1:0] node3057;
	wire [14-1:0] node3060;
	wire [14-1:0] node3063;
	wire [14-1:0] node3064;
	wire [14-1:0] node3068;
	wire [14-1:0] node3069;
	wire [14-1:0] node3070;
	wire [14-1:0] node3071;
	wire [14-1:0] node3074;
	wire [14-1:0] node3077;
	wire [14-1:0] node3078;
	wire [14-1:0] node3081;
	wire [14-1:0] node3084;
	wire [14-1:0] node3085;
	wire [14-1:0] node3086;
	wire [14-1:0] node3089;
	wire [14-1:0] node3092;
	wire [14-1:0] node3093;
	wire [14-1:0] node3096;
	wire [14-1:0] node3099;
	wire [14-1:0] node3100;
	wire [14-1:0] node3101;
	wire [14-1:0] node3102;
	wire [14-1:0] node3103;
	wire [14-1:0] node3107;
	wire [14-1:0] node3108;
	wire [14-1:0] node3111;
	wire [14-1:0] node3114;
	wire [14-1:0] node3115;
	wire [14-1:0] node3116;
	wire [14-1:0] node3120;
	wire [14-1:0] node3121;
	wire [14-1:0] node3124;
	wire [14-1:0] node3127;
	wire [14-1:0] node3128;
	wire [14-1:0] node3129;
	wire [14-1:0] node3130;
	wire [14-1:0] node3133;
	wire [14-1:0] node3136;
	wire [14-1:0] node3137;
	wire [14-1:0] node3140;
	wire [14-1:0] node3143;
	wire [14-1:0] node3144;
	wire [14-1:0] node3145;
	wire [14-1:0] node3148;
	wire [14-1:0] node3151;
	wire [14-1:0] node3152;
	wire [14-1:0] node3155;
	wire [14-1:0] node3158;
	wire [14-1:0] node3159;
	wire [14-1:0] node3160;
	wire [14-1:0] node3161;
	wire [14-1:0] node3162;
	wire [14-1:0] node3163;
	wire [14-1:0] node3165;
	wire [14-1:0] node3168;
	wire [14-1:0] node3169;
	wire [14-1:0] node3173;
	wire [14-1:0] node3174;
	wire [14-1:0] node3175;
	wire [14-1:0] node3178;
	wire [14-1:0] node3181;
	wire [14-1:0] node3182;
	wire [14-1:0] node3185;
	wire [14-1:0] node3188;
	wire [14-1:0] node3189;
	wire [14-1:0] node3190;
	wire [14-1:0] node3191;
	wire [14-1:0] node3194;
	wire [14-1:0] node3197;
	wire [14-1:0] node3198;
	wire [14-1:0] node3201;
	wire [14-1:0] node3204;
	wire [14-1:0] node3205;
	wire [14-1:0] node3206;
	wire [14-1:0] node3209;
	wire [14-1:0] node3212;
	wire [14-1:0] node3213;
	wire [14-1:0] node3216;
	wire [14-1:0] node3219;
	wire [14-1:0] node3220;
	wire [14-1:0] node3221;
	wire [14-1:0] node3222;
	wire [14-1:0] node3223;
	wire [14-1:0] node3227;
	wire [14-1:0] node3228;
	wire [14-1:0] node3231;
	wire [14-1:0] node3234;
	wire [14-1:0] node3235;
	wire [14-1:0] node3236;
	wire [14-1:0] node3239;
	wire [14-1:0] node3242;
	wire [14-1:0] node3243;
	wire [14-1:0] node3246;
	wire [14-1:0] node3249;
	wire [14-1:0] node3250;
	wire [14-1:0] node3251;
	wire [14-1:0] node3252;
	wire [14-1:0] node3255;
	wire [14-1:0] node3258;
	wire [14-1:0] node3260;
	wire [14-1:0] node3263;
	wire [14-1:0] node3264;
	wire [14-1:0] node3266;
	wire [14-1:0] node3269;
	wire [14-1:0] node3270;
	wire [14-1:0] node3273;
	wire [14-1:0] node3276;
	wire [14-1:0] node3277;
	wire [14-1:0] node3278;
	wire [14-1:0] node3279;
	wire [14-1:0] node3280;
	wire [14-1:0] node3281;
	wire [14-1:0] node3284;
	wire [14-1:0] node3287;
	wire [14-1:0] node3288;
	wire [14-1:0] node3291;
	wire [14-1:0] node3294;
	wire [14-1:0] node3295;
	wire [14-1:0] node3296;
	wire [14-1:0] node3299;
	wire [14-1:0] node3302;
	wire [14-1:0] node3304;
	wire [14-1:0] node3307;
	wire [14-1:0] node3308;
	wire [14-1:0] node3309;
	wire [14-1:0] node3310;
	wire [14-1:0] node3313;
	wire [14-1:0] node3316;
	wire [14-1:0] node3317;
	wire [14-1:0] node3321;
	wire [14-1:0] node3322;
	wire [14-1:0] node3323;
	wire [14-1:0] node3326;
	wire [14-1:0] node3329;
	wire [14-1:0] node3330;
	wire [14-1:0] node3333;
	wire [14-1:0] node3336;
	wire [14-1:0] node3337;
	wire [14-1:0] node3338;
	wire [14-1:0] node3339;
	wire [14-1:0] node3340;
	wire [14-1:0] node3343;
	wire [14-1:0] node3346;
	wire [14-1:0] node3347;
	wire [14-1:0] node3350;
	wire [14-1:0] node3353;
	wire [14-1:0] node3354;
	wire [14-1:0] node3355;
	wire [14-1:0] node3358;
	wire [14-1:0] node3361;
	wire [14-1:0] node3362;
	wire [14-1:0] node3365;
	wire [14-1:0] node3368;
	wire [14-1:0] node3369;
	wire [14-1:0] node3370;
	wire [14-1:0] node3371;
	wire [14-1:0] node3374;
	wire [14-1:0] node3377;
	wire [14-1:0] node3378;
	wire [14-1:0] node3381;
	wire [14-1:0] node3384;
	wire [14-1:0] node3385;
	wire [14-1:0] node3386;
	wire [14-1:0] node3389;
	wire [14-1:0] node3392;
	wire [14-1:0] node3394;
	wire [14-1:0] node3397;
	wire [14-1:0] node3398;
	wire [14-1:0] node3399;
	wire [14-1:0] node3400;
	wire [14-1:0] node3401;
	wire [14-1:0] node3402;
	wire [14-1:0] node3403;
	wire [14-1:0] node3405;
	wire [14-1:0] node3408;
	wire [14-1:0] node3409;
	wire [14-1:0] node3413;
	wire [14-1:0] node3414;
	wire [14-1:0] node3415;
	wire [14-1:0] node3418;
	wire [14-1:0] node3421;
	wire [14-1:0] node3422;
	wire [14-1:0] node3425;
	wire [14-1:0] node3428;
	wire [14-1:0] node3429;
	wire [14-1:0] node3430;
	wire [14-1:0] node3431;
	wire [14-1:0] node3434;
	wire [14-1:0] node3437;
	wire [14-1:0] node3438;
	wire [14-1:0] node3441;
	wire [14-1:0] node3444;
	wire [14-1:0] node3445;
	wire [14-1:0] node3446;
	wire [14-1:0] node3449;
	wire [14-1:0] node3452;
	wire [14-1:0] node3453;
	wire [14-1:0] node3456;
	wire [14-1:0] node3459;
	wire [14-1:0] node3460;
	wire [14-1:0] node3461;
	wire [14-1:0] node3462;
	wire [14-1:0] node3463;
	wire [14-1:0] node3466;
	wire [14-1:0] node3469;
	wire [14-1:0] node3470;
	wire [14-1:0] node3473;
	wire [14-1:0] node3476;
	wire [14-1:0] node3477;
	wire [14-1:0] node3478;
	wire [14-1:0] node3481;
	wire [14-1:0] node3484;
	wire [14-1:0] node3485;
	wire [14-1:0] node3488;
	wire [14-1:0] node3491;
	wire [14-1:0] node3492;
	wire [14-1:0] node3493;
	wire [14-1:0] node3495;
	wire [14-1:0] node3498;
	wire [14-1:0] node3499;
	wire [14-1:0] node3502;
	wire [14-1:0] node3505;
	wire [14-1:0] node3506;
	wire [14-1:0] node3507;
	wire [14-1:0] node3510;
	wire [14-1:0] node3513;
	wire [14-1:0] node3514;
	wire [14-1:0] node3517;
	wire [14-1:0] node3520;
	wire [14-1:0] node3521;
	wire [14-1:0] node3522;
	wire [14-1:0] node3523;
	wire [14-1:0] node3524;
	wire [14-1:0] node3525;
	wire [14-1:0] node3528;
	wire [14-1:0] node3531;
	wire [14-1:0] node3532;
	wire [14-1:0] node3536;
	wire [14-1:0] node3537;
	wire [14-1:0] node3538;
	wire [14-1:0] node3541;
	wire [14-1:0] node3544;
	wire [14-1:0] node3545;
	wire [14-1:0] node3548;
	wire [14-1:0] node3551;
	wire [14-1:0] node3552;
	wire [14-1:0] node3553;
	wire [14-1:0] node3555;
	wire [14-1:0] node3558;
	wire [14-1:0] node3559;
	wire [14-1:0] node3562;
	wire [14-1:0] node3565;
	wire [14-1:0] node3566;
	wire [14-1:0] node3567;
	wire [14-1:0] node3570;
	wire [14-1:0] node3573;
	wire [14-1:0] node3574;
	wire [14-1:0] node3577;
	wire [14-1:0] node3580;
	wire [14-1:0] node3581;
	wire [14-1:0] node3582;
	wire [14-1:0] node3583;
	wire [14-1:0] node3584;
	wire [14-1:0] node3588;
	wire [14-1:0] node3590;
	wire [14-1:0] node3593;
	wire [14-1:0] node3594;
	wire [14-1:0] node3595;
	wire [14-1:0] node3598;
	wire [14-1:0] node3601;
	wire [14-1:0] node3602;
	wire [14-1:0] node3605;
	wire [14-1:0] node3608;
	wire [14-1:0] node3609;
	wire [14-1:0] node3610;
	wire [14-1:0] node3611;
	wire [14-1:0] node3614;
	wire [14-1:0] node3617;
	wire [14-1:0] node3618;
	wire [14-1:0] node3621;
	wire [14-1:0] node3624;
	wire [14-1:0] node3625;
	wire [14-1:0] node3626;
	wire [14-1:0] node3629;
	wire [14-1:0] node3632;
	wire [14-1:0] node3633;
	wire [14-1:0] node3636;
	wire [14-1:0] node3639;
	wire [14-1:0] node3640;
	wire [14-1:0] node3641;
	wire [14-1:0] node3642;
	wire [14-1:0] node3643;
	wire [14-1:0] node3644;
	wire [14-1:0] node3645;
	wire [14-1:0] node3648;
	wire [14-1:0] node3651;
	wire [14-1:0] node3652;
	wire [14-1:0] node3655;
	wire [14-1:0] node3658;
	wire [14-1:0] node3659;
	wire [14-1:0] node3660;
	wire [14-1:0] node3663;
	wire [14-1:0] node3666;
	wire [14-1:0] node3667;
	wire [14-1:0] node3670;
	wire [14-1:0] node3673;
	wire [14-1:0] node3674;
	wire [14-1:0] node3675;
	wire [14-1:0] node3676;
	wire [14-1:0] node3679;
	wire [14-1:0] node3682;
	wire [14-1:0] node3683;
	wire [14-1:0] node3686;
	wire [14-1:0] node3689;
	wire [14-1:0] node3690;
	wire [14-1:0] node3692;
	wire [14-1:0] node3695;
	wire [14-1:0] node3696;
	wire [14-1:0] node3699;
	wire [14-1:0] node3702;
	wire [14-1:0] node3703;
	wire [14-1:0] node3704;
	wire [14-1:0] node3705;
	wire [14-1:0] node3706;
	wire [14-1:0] node3709;
	wire [14-1:0] node3712;
	wire [14-1:0] node3713;
	wire [14-1:0] node3716;
	wire [14-1:0] node3719;
	wire [14-1:0] node3720;
	wire [14-1:0] node3722;
	wire [14-1:0] node3725;
	wire [14-1:0] node3726;
	wire [14-1:0] node3729;
	wire [14-1:0] node3732;
	wire [14-1:0] node3733;
	wire [14-1:0] node3734;
	wire [14-1:0] node3736;
	wire [14-1:0] node3739;
	wire [14-1:0] node3741;
	wire [14-1:0] node3744;
	wire [14-1:0] node3745;
	wire [14-1:0] node3746;
	wire [14-1:0] node3749;
	wire [14-1:0] node3752;
	wire [14-1:0] node3753;
	wire [14-1:0] node3756;
	wire [14-1:0] node3759;
	wire [14-1:0] node3760;
	wire [14-1:0] node3761;
	wire [14-1:0] node3762;
	wire [14-1:0] node3763;
	wire [14-1:0] node3764;
	wire [14-1:0] node3767;
	wire [14-1:0] node3770;
	wire [14-1:0] node3771;
	wire [14-1:0] node3774;
	wire [14-1:0] node3777;
	wire [14-1:0] node3778;
	wire [14-1:0] node3779;
	wire [14-1:0] node3782;
	wire [14-1:0] node3785;
	wire [14-1:0] node3786;
	wire [14-1:0] node3789;
	wire [14-1:0] node3792;
	wire [14-1:0] node3793;
	wire [14-1:0] node3794;
	wire [14-1:0] node3796;
	wire [14-1:0] node3799;
	wire [14-1:0] node3800;
	wire [14-1:0] node3803;
	wire [14-1:0] node3806;
	wire [14-1:0] node3807;
	wire [14-1:0] node3808;
	wire [14-1:0] node3811;
	wire [14-1:0] node3814;
	wire [14-1:0] node3815;
	wire [14-1:0] node3818;
	wire [14-1:0] node3821;
	wire [14-1:0] node3822;
	wire [14-1:0] node3823;
	wire [14-1:0] node3824;
	wire [14-1:0] node3825;
	wire [14-1:0] node3828;
	wire [14-1:0] node3831;
	wire [14-1:0] node3832;
	wire [14-1:0] node3835;
	wire [14-1:0] node3838;
	wire [14-1:0] node3839;
	wire [14-1:0] node3840;
	wire [14-1:0] node3843;
	wire [14-1:0] node3846;
	wire [14-1:0] node3847;
	wire [14-1:0] node3850;
	wire [14-1:0] node3853;
	wire [14-1:0] node3854;
	wire [14-1:0] node3855;
	wire [14-1:0] node3856;
	wire [14-1:0] node3859;
	wire [14-1:0] node3862;
	wire [14-1:0] node3864;
	wire [14-1:0] node3867;
	wire [14-1:0] node3868;
	wire [14-1:0] node3869;
	wire [14-1:0] node3872;
	wire [14-1:0] node3875;
	wire [14-1:0] node3876;
	wire [14-1:0] node3879;
	wire [14-1:0] node3882;
	wire [14-1:0] node3883;
	wire [14-1:0] node3884;
	wire [14-1:0] node3885;
	wire [14-1:0] node3886;
	wire [14-1:0] node3887;
	wire [14-1:0] node3888;
	wire [14-1:0] node3889;
	wire [14-1:0] node3890;
	wire [14-1:0] node3891;
	wire [14-1:0] node3892;
	wire [14-1:0] node3895;
	wire [14-1:0] node3898;
	wire [14-1:0] node3899;
	wire [14-1:0] node3902;
	wire [14-1:0] node3905;
	wire [14-1:0] node3906;
	wire [14-1:0] node3907;
	wire [14-1:0] node3910;
	wire [14-1:0] node3913;
	wire [14-1:0] node3914;
	wire [14-1:0] node3917;
	wire [14-1:0] node3920;
	wire [14-1:0] node3921;
	wire [14-1:0] node3922;
	wire [14-1:0] node3923;
	wire [14-1:0] node3927;
	wire [14-1:0] node3928;
	wire [14-1:0] node3932;
	wire [14-1:0] node3933;
	wire [14-1:0] node3934;
	wire [14-1:0] node3937;
	wire [14-1:0] node3940;
	wire [14-1:0] node3941;
	wire [14-1:0] node3944;
	wire [14-1:0] node3947;
	wire [14-1:0] node3948;
	wire [14-1:0] node3949;
	wire [14-1:0] node3950;
	wire [14-1:0] node3951;
	wire [14-1:0] node3954;
	wire [14-1:0] node3957;
	wire [14-1:0] node3958;
	wire [14-1:0] node3961;
	wire [14-1:0] node3964;
	wire [14-1:0] node3965;
	wire [14-1:0] node3966;
	wire [14-1:0] node3969;
	wire [14-1:0] node3972;
	wire [14-1:0] node3973;
	wire [14-1:0] node3976;
	wire [14-1:0] node3979;
	wire [14-1:0] node3980;
	wire [14-1:0] node3981;
	wire [14-1:0] node3982;
	wire [14-1:0] node3985;
	wire [14-1:0] node3988;
	wire [14-1:0] node3989;
	wire [14-1:0] node3992;
	wire [14-1:0] node3995;
	wire [14-1:0] node3996;
	wire [14-1:0] node3997;
	wire [14-1:0] node4000;
	wire [14-1:0] node4003;
	wire [14-1:0] node4004;
	wire [14-1:0] node4007;
	wire [14-1:0] node4010;
	wire [14-1:0] node4011;
	wire [14-1:0] node4012;
	wire [14-1:0] node4013;
	wire [14-1:0] node4014;
	wire [14-1:0] node4015;
	wire [14-1:0] node4018;
	wire [14-1:0] node4021;
	wire [14-1:0] node4024;
	wire [14-1:0] node4026;
	wire [14-1:0] node4027;
	wire [14-1:0] node4030;
	wire [14-1:0] node4033;
	wire [14-1:0] node4034;
	wire [14-1:0] node4035;
	wire [14-1:0] node4036;
	wire [14-1:0] node4039;
	wire [14-1:0] node4042;
	wire [14-1:0] node4043;
	wire [14-1:0] node4046;
	wire [14-1:0] node4049;
	wire [14-1:0] node4050;
	wire [14-1:0] node4051;
	wire [14-1:0] node4054;
	wire [14-1:0] node4057;
	wire [14-1:0] node4058;
	wire [14-1:0] node4061;
	wire [14-1:0] node4064;
	wire [14-1:0] node4065;
	wire [14-1:0] node4066;
	wire [14-1:0] node4067;
	wire [14-1:0] node4068;
	wire [14-1:0] node4071;
	wire [14-1:0] node4074;
	wire [14-1:0] node4075;
	wire [14-1:0] node4078;
	wire [14-1:0] node4081;
	wire [14-1:0] node4082;
	wire [14-1:0] node4083;
	wire [14-1:0] node4086;
	wire [14-1:0] node4089;
	wire [14-1:0] node4091;
	wire [14-1:0] node4094;
	wire [14-1:0] node4095;
	wire [14-1:0] node4096;
	wire [14-1:0] node4097;
	wire [14-1:0] node4100;
	wire [14-1:0] node4103;
	wire [14-1:0] node4104;
	wire [14-1:0] node4107;
	wire [14-1:0] node4110;
	wire [14-1:0] node4111;
	wire [14-1:0] node4112;
	wire [14-1:0] node4115;
	wire [14-1:0] node4118;
	wire [14-1:0] node4119;
	wire [14-1:0] node4123;
	wire [14-1:0] node4124;
	wire [14-1:0] node4125;
	wire [14-1:0] node4126;
	wire [14-1:0] node4127;
	wire [14-1:0] node4128;
	wire [14-1:0] node4129;
	wire [14-1:0] node4132;
	wire [14-1:0] node4135;
	wire [14-1:0] node4136;
	wire [14-1:0] node4139;
	wire [14-1:0] node4142;
	wire [14-1:0] node4143;
	wire [14-1:0] node4144;
	wire [14-1:0] node4147;
	wire [14-1:0] node4150;
	wire [14-1:0] node4151;
	wire [14-1:0] node4154;
	wire [14-1:0] node4157;
	wire [14-1:0] node4158;
	wire [14-1:0] node4159;
	wire [14-1:0] node4160;
	wire [14-1:0] node4163;
	wire [14-1:0] node4166;
	wire [14-1:0] node4167;
	wire [14-1:0] node4170;
	wire [14-1:0] node4173;
	wire [14-1:0] node4174;
	wire [14-1:0] node4175;
	wire [14-1:0] node4178;
	wire [14-1:0] node4181;
	wire [14-1:0] node4183;
	wire [14-1:0] node4186;
	wire [14-1:0] node4187;
	wire [14-1:0] node4188;
	wire [14-1:0] node4189;
	wire [14-1:0] node4190;
	wire [14-1:0] node4193;
	wire [14-1:0] node4196;
	wire [14-1:0] node4197;
	wire [14-1:0] node4201;
	wire [14-1:0] node4202;
	wire [14-1:0] node4203;
	wire [14-1:0] node4206;
	wire [14-1:0] node4209;
	wire [14-1:0] node4210;
	wire [14-1:0] node4213;
	wire [14-1:0] node4216;
	wire [14-1:0] node4217;
	wire [14-1:0] node4218;
	wire [14-1:0] node4219;
	wire [14-1:0] node4222;
	wire [14-1:0] node4225;
	wire [14-1:0] node4226;
	wire [14-1:0] node4229;
	wire [14-1:0] node4232;
	wire [14-1:0] node4233;
	wire [14-1:0] node4235;
	wire [14-1:0] node4238;
	wire [14-1:0] node4239;
	wire [14-1:0] node4242;
	wire [14-1:0] node4245;
	wire [14-1:0] node4246;
	wire [14-1:0] node4247;
	wire [14-1:0] node4248;
	wire [14-1:0] node4249;
	wire [14-1:0] node4250;
	wire [14-1:0] node4253;
	wire [14-1:0] node4256;
	wire [14-1:0] node4257;
	wire [14-1:0] node4260;
	wire [14-1:0] node4263;
	wire [14-1:0] node4264;
	wire [14-1:0] node4265;
	wire [14-1:0] node4268;
	wire [14-1:0] node4271;
	wire [14-1:0] node4272;
	wire [14-1:0] node4275;
	wire [14-1:0] node4278;
	wire [14-1:0] node4279;
	wire [14-1:0] node4280;
	wire [14-1:0] node4281;
	wire [14-1:0] node4284;
	wire [14-1:0] node4287;
	wire [14-1:0] node4288;
	wire [14-1:0] node4291;
	wire [14-1:0] node4294;
	wire [14-1:0] node4295;
	wire [14-1:0] node4297;
	wire [14-1:0] node4300;
	wire [14-1:0] node4301;
	wire [14-1:0] node4304;
	wire [14-1:0] node4307;
	wire [14-1:0] node4308;
	wire [14-1:0] node4309;
	wire [14-1:0] node4310;
	wire [14-1:0] node4311;
	wire [14-1:0] node4315;
	wire [14-1:0] node4316;
	wire [14-1:0] node4319;
	wire [14-1:0] node4322;
	wire [14-1:0] node4323;
	wire [14-1:0] node4324;
	wire [14-1:0] node4327;
	wire [14-1:0] node4330;
	wire [14-1:0] node4332;
	wire [14-1:0] node4335;
	wire [14-1:0] node4336;
	wire [14-1:0] node4337;
	wire [14-1:0] node4338;
	wire [14-1:0] node4341;
	wire [14-1:0] node4344;
	wire [14-1:0] node4345;
	wire [14-1:0] node4348;
	wire [14-1:0] node4351;
	wire [14-1:0] node4352;
	wire [14-1:0] node4353;
	wire [14-1:0] node4356;
	wire [14-1:0] node4359;
	wire [14-1:0] node4360;
	wire [14-1:0] node4363;
	wire [14-1:0] node4366;
	wire [14-1:0] node4367;
	wire [14-1:0] node4368;
	wire [14-1:0] node4369;
	wire [14-1:0] node4370;
	wire [14-1:0] node4371;
	wire [14-1:0] node4372;
	wire [14-1:0] node4373;
	wire [14-1:0] node4376;
	wire [14-1:0] node4379;
	wire [14-1:0] node4380;
	wire [14-1:0] node4383;
	wire [14-1:0] node4386;
	wire [14-1:0] node4387;
	wire [14-1:0] node4388;
	wire [14-1:0] node4391;
	wire [14-1:0] node4394;
	wire [14-1:0] node4395;
	wire [14-1:0] node4398;
	wire [14-1:0] node4401;
	wire [14-1:0] node4402;
	wire [14-1:0] node4403;
	wire [14-1:0] node4405;
	wire [14-1:0] node4408;
	wire [14-1:0] node4409;
	wire [14-1:0] node4413;
	wire [14-1:0] node4414;
	wire [14-1:0] node4416;
	wire [14-1:0] node4419;
	wire [14-1:0] node4421;
	wire [14-1:0] node4424;
	wire [14-1:0] node4425;
	wire [14-1:0] node4426;
	wire [14-1:0] node4427;
	wire [14-1:0] node4428;
	wire [14-1:0] node4431;
	wire [14-1:0] node4434;
	wire [14-1:0] node4435;
	wire [14-1:0] node4439;
	wire [14-1:0] node4440;
	wire [14-1:0] node4441;
	wire [14-1:0] node4444;
	wire [14-1:0] node4447;
	wire [14-1:0] node4448;
	wire [14-1:0] node4451;
	wire [14-1:0] node4454;
	wire [14-1:0] node4455;
	wire [14-1:0] node4456;
	wire [14-1:0] node4457;
	wire [14-1:0] node4460;
	wire [14-1:0] node4464;
	wire [14-1:0] node4465;
	wire [14-1:0] node4466;
	wire [14-1:0] node4469;
	wire [14-1:0] node4472;
	wire [14-1:0] node4473;
	wire [14-1:0] node4476;
	wire [14-1:0] node4479;
	wire [14-1:0] node4480;
	wire [14-1:0] node4481;
	wire [14-1:0] node4482;
	wire [14-1:0] node4483;
	wire [14-1:0] node4484;
	wire [14-1:0] node4487;
	wire [14-1:0] node4490;
	wire [14-1:0] node4491;
	wire [14-1:0] node4494;
	wire [14-1:0] node4497;
	wire [14-1:0] node4498;
	wire [14-1:0] node4499;
	wire [14-1:0] node4502;
	wire [14-1:0] node4505;
	wire [14-1:0] node4506;
	wire [14-1:0] node4510;
	wire [14-1:0] node4511;
	wire [14-1:0] node4512;
	wire [14-1:0] node4513;
	wire [14-1:0] node4516;
	wire [14-1:0] node4519;
	wire [14-1:0] node4520;
	wire [14-1:0] node4523;
	wire [14-1:0] node4526;
	wire [14-1:0] node4527;
	wire [14-1:0] node4528;
	wire [14-1:0] node4531;
	wire [14-1:0] node4534;
	wire [14-1:0] node4535;
	wire [14-1:0] node4538;
	wire [14-1:0] node4541;
	wire [14-1:0] node4542;
	wire [14-1:0] node4543;
	wire [14-1:0] node4544;
	wire [14-1:0] node4545;
	wire [14-1:0] node4548;
	wire [14-1:0] node4551;
	wire [14-1:0] node4552;
	wire [14-1:0] node4555;
	wire [14-1:0] node4558;
	wire [14-1:0] node4559;
	wire [14-1:0] node4560;
	wire [14-1:0] node4563;
	wire [14-1:0] node4566;
	wire [14-1:0] node4567;
	wire [14-1:0] node4570;
	wire [14-1:0] node4573;
	wire [14-1:0] node4574;
	wire [14-1:0] node4575;
	wire [14-1:0] node4576;
	wire [14-1:0] node4579;
	wire [14-1:0] node4582;
	wire [14-1:0] node4583;
	wire [14-1:0] node4586;
	wire [14-1:0] node4589;
	wire [14-1:0] node4590;
	wire [14-1:0] node4591;
	wire [14-1:0] node4595;
	wire [14-1:0] node4596;
	wire [14-1:0] node4599;
	wire [14-1:0] node4602;
	wire [14-1:0] node4603;
	wire [14-1:0] node4604;
	wire [14-1:0] node4605;
	wire [14-1:0] node4606;
	wire [14-1:0] node4607;
	wire [14-1:0] node4608;
	wire [14-1:0] node4611;
	wire [14-1:0] node4614;
	wire [14-1:0] node4615;
	wire [14-1:0] node4618;
	wire [14-1:0] node4621;
	wire [14-1:0] node4622;
	wire [14-1:0] node4623;
	wire [14-1:0] node4626;
	wire [14-1:0] node4629;
	wire [14-1:0] node4630;
	wire [14-1:0] node4633;
	wire [14-1:0] node4636;
	wire [14-1:0] node4637;
	wire [14-1:0] node4638;
	wire [14-1:0] node4639;
	wire [14-1:0] node4642;
	wire [14-1:0] node4645;
	wire [14-1:0] node4646;
	wire [14-1:0] node4649;
	wire [14-1:0] node4652;
	wire [14-1:0] node4653;
	wire [14-1:0] node4654;
	wire [14-1:0] node4657;
	wire [14-1:0] node4660;
	wire [14-1:0] node4661;
	wire [14-1:0] node4664;
	wire [14-1:0] node4667;
	wire [14-1:0] node4668;
	wire [14-1:0] node4669;
	wire [14-1:0] node4670;
	wire [14-1:0] node4671;
	wire [14-1:0] node4674;
	wire [14-1:0] node4677;
	wire [14-1:0] node4678;
	wire [14-1:0] node4681;
	wire [14-1:0] node4684;
	wire [14-1:0] node4685;
	wire [14-1:0] node4686;
	wire [14-1:0] node4689;
	wire [14-1:0] node4692;
	wire [14-1:0] node4693;
	wire [14-1:0] node4696;
	wire [14-1:0] node4699;
	wire [14-1:0] node4700;
	wire [14-1:0] node4701;
	wire [14-1:0] node4702;
	wire [14-1:0] node4705;
	wire [14-1:0] node4708;
	wire [14-1:0] node4709;
	wire [14-1:0] node4712;
	wire [14-1:0] node4715;
	wire [14-1:0] node4716;
	wire [14-1:0] node4717;
	wire [14-1:0] node4720;
	wire [14-1:0] node4723;
	wire [14-1:0] node4724;
	wire [14-1:0] node4727;
	wire [14-1:0] node4730;
	wire [14-1:0] node4731;
	wire [14-1:0] node4732;
	wire [14-1:0] node4733;
	wire [14-1:0] node4734;
	wire [14-1:0] node4735;
	wire [14-1:0] node4738;
	wire [14-1:0] node4741;
	wire [14-1:0] node4742;
	wire [14-1:0] node4746;
	wire [14-1:0] node4747;
	wire [14-1:0] node4748;
	wire [14-1:0] node4751;
	wire [14-1:0] node4754;
	wire [14-1:0] node4755;
	wire [14-1:0] node4758;
	wire [14-1:0] node4761;
	wire [14-1:0] node4762;
	wire [14-1:0] node4763;
	wire [14-1:0] node4764;
	wire [14-1:0] node4767;
	wire [14-1:0] node4770;
	wire [14-1:0] node4771;
	wire [14-1:0] node4774;
	wire [14-1:0] node4777;
	wire [14-1:0] node4778;
	wire [14-1:0] node4779;
	wire [14-1:0] node4782;
	wire [14-1:0] node4785;
	wire [14-1:0] node4786;
	wire [14-1:0] node4789;
	wire [14-1:0] node4792;
	wire [14-1:0] node4793;
	wire [14-1:0] node4794;
	wire [14-1:0] node4795;
	wire [14-1:0] node4796;
	wire [14-1:0] node4799;
	wire [14-1:0] node4802;
	wire [14-1:0] node4803;
	wire [14-1:0] node4806;
	wire [14-1:0] node4809;
	wire [14-1:0] node4811;
	wire [14-1:0] node4812;
	wire [14-1:0] node4815;
	wire [14-1:0] node4818;
	wire [14-1:0] node4819;
	wire [14-1:0] node4820;
	wire [14-1:0] node4821;
	wire [14-1:0] node4824;
	wire [14-1:0] node4827;
	wire [14-1:0] node4828;
	wire [14-1:0] node4831;
	wire [14-1:0] node4834;
	wire [14-1:0] node4835;
	wire [14-1:0] node4836;
	wire [14-1:0] node4839;
	wire [14-1:0] node4842;
	wire [14-1:0] node4843;
	wire [14-1:0] node4846;
	wire [14-1:0] node4849;
	wire [14-1:0] node4850;
	wire [14-1:0] node4851;
	wire [14-1:0] node4852;
	wire [14-1:0] node4853;
	wire [14-1:0] node4854;
	wire [14-1:0] node4855;
	wire [14-1:0] node4856;
	wire [14-1:0] node4857;
	wire [14-1:0] node4860;
	wire [14-1:0] node4863;
	wire [14-1:0] node4864;
	wire [14-1:0] node4867;
	wire [14-1:0] node4870;
	wire [14-1:0] node4871;
	wire [14-1:0] node4872;
	wire [14-1:0] node4875;
	wire [14-1:0] node4878;
	wire [14-1:0] node4879;
	wire [14-1:0] node4882;
	wire [14-1:0] node4885;
	wire [14-1:0] node4886;
	wire [14-1:0] node4887;
	wire [14-1:0] node4888;
	wire [14-1:0] node4891;
	wire [14-1:0] node4894;
	wire [14-1:0] node4896;
	wire [14-1:0] node4899;
	wire [14-1:0] node4900;
	wire [14-1:0] node4901;
	wire [14-1:0] node4904;
	wire [14-1:0] node4907;
	wire [14-1:0] node4908;
	wire [14-1:0] node4911;
	wire [14-1:0] node4914;
	wire [14-1:0] node4915;
	wire [14-1:0] node4916;
	wire [14-1:0] node4917;
	wire [14-1:0] node4919;
	wire [14-1:0] node4922;
	wire [14-1:0] node4923;
	wire [14-1:0] node4926;
	wire [14-1:0] node4929;
	wire [14-1:0] node4930;
	wire [14-1:0] node4931;
	wire [14-1:0] node4934;
	wire [14-1:0] node4937;
	wire [14-1:0] node4938;
	wire [14-1:0] node4942;
	wire [14-1:0] node4943;
	wire [14-1:0] node4944;
	wire [14-1:0] node4945;
	wire [14-1:0] node4948;
	wire [14-1:0] node4951;
	wire [14-1:0] node4952;
	wire [14-1:0] node4955;
	wire [14-1:0] node4958;
	wire [14-1:0] node4959;
	wire [14-1:0] node4960;
	wire [14-1:0] node4963;
	wire [14-1:0] node4966;
	wire [14-1:0] node4967;
	wire [14-1:0] node4970;
	wire [14-1:0] node4973;
	wire [14-1:0] node4974;
	wire [14-1:0] node4975;
	wire [14-1:0] node4976;
	wire [14-1:0] node4977;
	wire [14-1:0] node4978;
	wire [14-1:0] node4981;
	wire [14-1:0] node4984;
	wire [14-1:0] node4985;
	wire [14-1:0] node4988;
	wire [14-1:0] node4991;
	wire [14-1:0] node4992;
	wire [14-1:0] node4993;
	wire [14-1:0] node4996;
	wire [14-1:0] node4999;
	wire [14-1:0] node5000;
	wire [14-1:0] node5003;
	wire [14-1:0] node5006;
	wire [14-1:0] node5007;
	wire [14-1:0] node5008;
	wire [14-1:0] node5009;
	wire [14-1:0] node5012;
	wire [14-1:0] node5015;
	wire [14-1:0] node5016;
	wire [14-1:0] node5019;
	wire [14-1:0] node5022;
	wire [14-1:0] node5023;
	wire [14-1:0] node5024;
	wire [14-1:0] node5027;
	wire [14-1:0] node5030;
	wire [14-1:0] node5032;
	wire [14-1:0] node5035;
	wire [14-1:0] node5036;
	wire [14-1:0] node5037;
	wire [14-1:0] node5038;
	wire [14-1:0] node5039;
	wire [14-1:0] node5042;
	wire [14-1:0] node5045;
	wire [14-1:0] node5047;
	wire [14-1:0] node5050;
	wire [14-1:0] node5051;
	wire [14-1:0] node5053;
	wire [14-1:0] node5056;
	wire [14-1:0] node5057;
	wire [14-1:0] node5061;
	wire [14-1:0] node5062;
	wire [14-1:0] node5063;
	wire [14-1:0] node5064;
	wire [14-1:0] node5067;
	wire [14-1:0] node5070;
	wire [14-1:0] node5072;
	wire [14-1:0] node5075;
	wire [14-1:0] node5076;
	wire [14-1:0] node5077;
	wire [14-1:0] node5080;
	wire [14-1:0] node5083;
	wire [14-1:0] node5084;
	wire [14-1:0] node5087;
	wire [14-1:0] node5090;
	wire [14-1:0] node5091;
	wire [14-1:0] node5092;
	wire [14-1:0] node5093;
	wire [14-1:0] node5094;
	wire [14-1:0] node5095;
	wire [14-1:0] node5096;
	wire [14-1:0] node5099;
	wire [14-1:0] node5102;
	wire [14-1:0] node5103;
	wire [14-1:0] node5107;
	wire [14-1:0] node5108;
	wire [14-1:0] node5109;
	wire [14-1:0] node5112;
	wire [14-1:0] node5115;
	wire [14-1:0] node5116;
	wire [14-1:0] node5119;
	wire [14-1:0] node5122;
	wire [14-1:0] node5123;
	wire [14-1:0] node5124;
	wire [14-1:0] node5125;
	wire [14-1:0] node5128;
	wire [14-1:0] node5131;
	wire [14-1:0] node5132;
	wire [14-1:0] node5136;
	wire [14-1:0] node5137;
	wire [14-1:0] node5138;
	wire [14-1:0] node5141;
	wire [14-1:0] node5144;
	wire [14-1:0] node5146;
	wire [14-1:0] node5149;
	wire [14-1:0] node5150;
	wire [14-1:0] node5151;
	wire [14-1:0] node5152;
	wire [14-1:0] node5153;
	wire [14-1:0] node5156;
	wire [14-1:0] node5159;
	wire [14-1:0] node5160;
	wire [14-1:0] node5163;
	wire [14-1:0] node5166;
	wire [14-1:0] node5167;
	wire [14-1:0] node5168;
	wire [14-1:0] node5171;
	wire [14-1:0] node5174;
	wire [14-1:0] node5175;
	wire [14-1:0] node5178;
	wire [14-1:0] node5181;
	wire [14-1:0] node5182;
	wire [14-1:0] node5183;
	wire [14-1:0] node5184;
	wire [14-1:0] node5187;
	wire [14-1:0] node5190;
	wire [14-1:0] node5191;
	wire [14-1:0] node5194;
	wire [14-1:0] node5197;
	wire [14-1:0] node5198;
	wire [14-1:0] node5199;
	wire [14-1:0] node5202;
	wire [14-1:0] node5205;
	wire [14-1:0] node5206;
	wire [14-1:0] node5209;
	wire [14-1:0] node5212;
	wire [14-1:0] node5213;
	wire [14-1:0] node5214;
	wire [14-1:0] node5215;
	wire [14-1:0] node5216;
	wire [14-1:0] node5217;
	wire [14-1:0] node5220;
	wire [14-1:0] node5223;
	wire [14-1:0] node5224;
	wire [14-1:0] node5228;
	wire [14-1:0] node5229;
	wire [14-1:0] node5230;
	wire [14-1:0] node5233;
	wire [14-1:0] node5236;
	wire [14-1:0] node5237;
	wire [14-1:0] node5240;
	wire [14-1:0] node5243;
	wire [14-1:0] node5244;
	wire [14-1:0] node5245;
	wire [14-1:0] node5246;
	wire [14-1:0] node5249;
	wire [14-1:0] node5252;
	wire [14-1:0] node5253;
	wire [14-1:0] node5257;
	wire [14-1:0] node5258;
	wire [14-1:0] node5259;
	wire [14-1:0] node5262;
	wire [14-1:0] node5265;
	wire [14-1:0] node5266;
	wire [14-1:0] node5269;
	wire [14-1:0] node5272;
	wire [14-1:0] node5273;
	wire [14-1:0] node5274;
	wire [14-1:0] node5275;
	wire [14-1:0] node5277;
	wire [14-1:0] node5280;
	wire [14-1:0] node5281;
	wire [14-1:0] node5284;
	wire [14-1:0] node5287;
	wire [14-1:0] node5288;
	wire [14-1:0] node5289;
	wire [14-1:0] node5292;
	wire [14-1:0] node5295;
	wire [14-1:0] node5296;
	wire [14-1:0] node5299;
	wire [14-1:0] node5302;
	wire [14-1:0] node5303;
	wire [14-1:0] node5304;
	wire [14-1:0] node5305;
	wire [14-1:0] node5308;
	wire [14-1:0] node5311;
	wire [14-1:0] node5313;
	wire [14-1:0] node5316;
	wire [14-1:0] node5317;
	wire [14-1:0] node5319;
	wire [14-1:0] node5322;
	wire [14-1:0] node5323;
	wire [14-1:0] node5326;
	wire [14-1:0] node5329;
	wire [14-1:0] node5330;
	wire [14-1:0] node5331;
	wire [14-1:0] node5332;
	wire [14-1:0] node5333;
	wire [14-1:0] node5334;
	wire [14-1:0] node5335;
	wire [14-1:0] node5336;
	wire [14-1:0] node5339;
	wire [14-1:0] node5342;
	wire [14-1:0] node5343;
	wire [14-1:0] node5346;
	wire [14-1:0] node5349;
	wire [14-1:0] node5350;
	wire [14-1:0] node5351;
	wire [14-1:0] node5354;
	wire [14-1:0] node5357;
	wire [14-1:0] node5358;
	wire [14-1:0] node5361;
	wire [14-1:0] node5364;
	wire [14-1:0] node5365;
	wire [14-1:0] node5366;
	wire [14-1:0] node5367;
	wire [14-1:0] node5370;
	wire [14-1:0] node5373;
	wire [14-1:0] node5374;
	wire [14-1:0] node5377;
	wire [14-1:0] node5380;
	wire [14-1:0] node5381;
	wire [14-1:0] node5382;
	wire [14-1:0] node5385;
	wire [14-1:0] node5388;
	wire [14-1:0] node5389;
	wire [14-1:0] node5392;
	wire [14-1:0] node5395;
	wire [14-1:0] node5396;
	wire [14-1:0] node5397;
	wire [14-1:0] node5398;
	wire [14-1:0] node5399;
	wire [14-1:0] node5402;
	wire [14-1:0] node5405;
	wire [14-1:0] node5406;
	wire [14-1:0] node5409;
	wire [14-1:0] node5412;
	wire [14-1:0] node5413;
	wire [14-1:0] node5414;
	wire [14-1:0] node5417;
	wire [14-1:0] node5420;
	wire [14-1:0] node5421;
	wire [14-1:0] node5424;
	wire [14-1:0] node5427;
	wire [14-1:0] node5428;
	wire [14-1:0] node5429;
	wire [14-1:0] node5430;
	wire [14-1:0] node5433;
	wire [14-1:0] node5436;
	wire [14-1:0] node5437;
	wire [14-1:0] node5440;
	wire [14-1:0] node5443;
	wire [14-1:0] node5444;
	wire [14-1:0] node5445;
	wire [14-1:0] node5448;
	wire [14-1:0] node5451;
	wire [14-1:0] node5452;
	wire [14-1:0] node5455;
	wire [14-1:0] node5458;
	wire [14-1:0] node5459;
	wire [14-1:0] node5460;
	wire [14-1:0] node5461;
	wire [14-1:0] node5462;
	wire [14-1:0] node5463;
	wire [14-1:0] node5466;
	wire [14-1:0] node5469;
	wire [14-1:0] node5470;
	wire [14-1:0] node5473;
	wire [14-1:0] node5476;
	wire [14-1:0] node5477;
	wire [14-1:0] node5478;
	wire [14-1:0] node5481;
	wire [14-1:0] node5484;
	wire [14-1:0] node5485;
	wire [14-1:0] node5488;
	wire [14-1:0] node5491;
	wire [14-1:0] node5492;
	wire [14-1:0] node5493;
	wire [14-1:0] node5494;
	wire [14-1:0] node5497;
	wire [14-1:0] node5500;
	wire [14-1:0] node5501;
	wire [14-1:0] node5504;
	wire [14-1:0] node5507;
	wire [14-1:0] node5508;
	wire [14-1:0] node5509;
	wire [14-1:0] node5512;
	wire [14-1:0] node5515;
	wire [14-1:0] node5516;
	wire [14-1:0] node5519;
	wire [14-1:0] node5522;
	wire [14-1:0] node5523;
	wire [14-1:0] node5524;
	wire [14-1:0] node5525;
	wire [14-1:0] node5526;
	wire [14-1:0] node5529;
	wire [14-1:0] node5532;
	wire [14-1:0] node5533;
	wire [14-1:0] node5536;
	wire [14-1:0] node5539;
	wire [14-1:0] node5540;
	wire [14-1:0] node5541;
	wire [14-1:0] node5544;
	wire [14-1:0] node5547;
	wire [14-1:0] node5548;
	wire [14-1:0] node5551;
	wire [14-1:0] node5554;
	wire [14-1:0] node5555;
	wire [14-1:0] node5556;
	wire [14-1:0] node5557;
	wire [14-1:0] node5560;
	wire [14-1:0] node5563;
	wire [14-1:0] node5564;
	wire [14-1:0] node5567;
	wire [14-1:0] node5570;
	wire [14-1:0] node5571;
	wire [14-1:0] node5572;
	wire [14-1:0] node5575;
	wire [14-1:0] node5578;
	wire [14-1:0] node5579;
	wire [14-1:0] node5582;
	wire [14-1:0] node5585;
	wire [14-1:0] node5586;
	wire [14-1:0] node5587;
	wire [14-1:0] node5588;
	wire [14-1:0] node5589;
	wire [14-1:0] node5590;
	wire [14-1:0] node5591;
	wire [14-1:0] node5594;
	wire [14-1:0] node5597;
	wire [14-1:0] node5598;
	wire [14-1:0] node5601;
	wire [14-1:0] node5604;
	wire [14-1:0] node5605;
	wire [14-1:0] node5606;
	wire [14-1:0] node5609;
	wire [14-1:0] node5612;
	wire [14-1:0] node5613;
	wire [14-1:0] node5616;
	wire [14-1:0] node5619;
	wire [14-1:0] node5620;
	wire [14-1:0] node5621;
	wire [14-1:0] node5622;
	wire [14-1:0] node5625;
	wire [14-1:0] node5628;
	wire [14-1:0] node5629;
	wire [14-1:0] node5632;
	wire [14-1:0] node5635;
	wire [14-1:0] node5636;
	wire [14-1:0] node5637;
	wire [14-1:0] node5640;
	wire [14-1:0] node5643;
	wire [14-1:0] node5644;
	wire [14-1:0] node5647;
	wire [14-1:0] node5650;
	wire [14-1:0] node5651;
	wire [14-1:0] node5652;
	wire [14-1:0] node5653;
	wire [14-1:0] node5654;
	wire [14-1:0] node5658;
	wire [14-1:0] node5659;
	wire [14-1:0] node5662;
	wire [14-1:0] node5665;
	wire [14-1:0] node5666;
	wire [14-1:0] node5667;
	wire [14-1:0] node5670;
	wire [14-1:0] node5673;
	wire [14-1:0] node5674;
	wire [14-1:0] node5677;
	wire [14-1:0] node5680;
	wire [14-1:0] node5681;
	wire [14-1:0] node5682;
	wire [14-1:0] node5683;
	wire [14-1:0] node5686;
	wire [14-1:0] node5689;
	wire [14-1:0] node5690;
	wire [14-1:0] node5693;
	wire [14-1:0] node5696;
	wire [14-1:0] node5697;
	wire [14-1:0] node5698;
	wire [14-1:0] node5701;
	wire [14-1:0] node5704;
	wire [14-1:0] node5706;
	wire [14-1:0] node5709;
	wire [14-1:0] node5710;
	wire [14-1:0] node5711;
	wire [14-1:0] node5712;
	wire [14-1:0] node5713;
	wire [14-1:0] node5714;
	wire [14-1:0] node5717;
	wire [14-1:0] node5720;
	wire [14-1:0] node5721;
	wire [14-1:0] node5724;
	wire [14-1:0] node5727;
	wire [14-1:0] node5728;
	wire [14-1:0] node5729;
	wire [14-1:0] node5732;
	wire [14-1:0] node5735;
	wire [14-1:0] node5736;
	wire [14-1:0] node5739;
	wire [14-1:0] node5742;
	wire [14-1:0] node5743;
	wire [14-1:0] node5744;
	wire [14-1:0] node5745;
	wire [14-1:0] node5748;
	wire [14-1:0] node5751;
	wire [14-1:0] node5753;
	wire [14-1:0] node5756;
	wire [14-1:0] node5757;
	wire [14-1:0] node5758;
	wire [14-1:0] node5762;
	wire [14-1:0] node5763;
	wire [14-1:0] node5766;
	wire [14-1:0] node5769;
	wire [14-1:0] node5770;
	wire [14-1:0] node5771;
	wire [14-1:0] node5772;
	wire [14-1:0] node5773;
	wire [14-1:0] node5777;
	wire [14-1:0] node5778;
	wire [14-1:0] node5781;
	wire [14-1:0] node5784;
	wire [14-1:0] node5785;
	wire [14-1:0] node5786;
	wire [14-1:0] node5789;
	wire [14-1:0] node5792;
	wire [14-1:0] node5793;
	wire [14-1:0] node5796;
	wire [14-1:0] node5799;
	wire [14-1:0] node5800;
	wire [14-1:0] node5801;
	wire [14-1:0] node5802;
	wire [14-1:0] node5805;
	wire [14-1:0] node5808;
	wire [14-1:0] node5809;
	wire [14-1:0] node5812;
	wire [14-1:0] node5815;
	wire [14-1:0] node5816;
	wire [14-1:0] node5817;
	wire [14-1:0] node5820;
	wire [14-1:0] node5823;
	wire [14-1:0] node5824;
	wire [14-1:0] node5827;
	wire [14-1:0] node5830;
	wire [14-1:0] node5831;
	wire [14-1:0] node5832;
	wire [14-1:0] node5833;
	wire [14-1:0] node5834;
	wire [14-1:0] node5835;
	wire [14-1:0] node5836;
	wire [14-1:0] node5837;
	wire [14-1:0] node5838;
	wire [14-1:0] node5840;
	wire [14-1:0] node5843;
	wire [14-1:0] node5844;
	wire [14-1:0] node5847;
	wire [14-1:0] node5850;
	wire [14-1:0] node5851;
	wire [14-1:0] node5852;
	wire [14-1:0] node5855;
	wire [14-1:0] node5858;
	wire [14-1:0] node5859;
	wire [14-1:0] node5862;
	wire [14-1:0] node5865;
	wire [14-1:0] node5866;
	wire [14-1:0] node5867;
	wire [14-1:0] node5870;
	wire [14-1:0] node5871;
	wire [14-1:0] node5875;
	wire [14-1:0] node5876;
	wire [14-1:0] node5877;
	wire [14-1:0] node5880;
	wire [14-1:0] node5883;
	wire [14-1:0] node5884;
	wire [14-1:0] node5887;
	wire [14-1:0] node5890;
	wire [14-1:0] node5891;
	wire [14-1:0] node5892;
	wire [14-1:0] node5893;
	wire [14-1:0] node5895;
	wire [14-1:0] node5898;
	wire [14-1:0] node5899;
	wire [14-1:0] node5902;
	wire [14-1:0] node5905;
	wire [14-1:0] node5906;
	wire [14-1:0] node5907;
	wire [14-1:0] node5910;
	wire [14-1:0] node5913;
	wire [14-1:0] node5914;
	wire [14-1:0] node5917;
	wire [14-1:0] node5920;
	wire [14-1:0] node5921;
	wire [14-1:0] node5922;
	wire [14-1:0] node5923;
	wire [14-1:0] node5926;
	wire [14-1:0] node5929;
	wire [14-1:0] node5930;
	wire [14-1:0] node5933;
	wire [14-1:0] node5936;
	wire [14-1:0] node5937;
	wire [14-1:0] node5939;
	wire [14-1:0] node5942;
	wire [14-1:0] node5943;
	wire [14-1:0] node5946;
	wire [14-1:0] node5949;
	wire [14-1:0] node5950;
	wire [14-1:0] node5951;
	wire [14-1:0] node5952;
	wire [14-1:0] node5953;
	wire [14-1:0] node5954;
	wire [14-1:0] node5957;
	wire [14-1:0] node5960;
	wire [14-1:0] node5961;
	wire [14-1:0] node5964;
	wire [14-1:0] node5967;
	wire [14-1:0] node5968;
	wire [14-1:0] node5969;
	wire [14-1:0] node5972;
	wire [14-1:0] node5975;
	wire [14-1:0] node5976;
	wire [14-1:0] node5979;
	wire [14-1:0] node5982;
	wire [14-1:0] node5983;
	wire [14-1:0] node5984;
	wire [14-1:0] node5985;
	wire [14-1:0] node5988;
	wire [14-1:0] node5991;
	wire [14-1:0] node5992;
	wire [14-1:0] node5995;
	wire [14-1:0] node5998;
	wire [14-1:0] node5999;
	wire [14-1:0] node6001;
	wire [14-1:0] node6004;
	wire [14-1:0] node6005;
	wire [14-1:0] node6008;
	wire [14-1:0] node6011;
	wire [14-1:0] node6012;
	wire [14-1:0] node6013;
	wire [14-1:0] node6014;
	wire [14-1:0] node6015;
	wire [14-1:0] node6018;
	wire [14-1:0] node6021;
	wire [14-1:0] node6022;
	wire [14-1:0] node6025;
	wire [14-1:0] node6028;
	wire [14-1:0] node6029;
	wire [14-1:0] node6030;
	wire [14-1:0] node6033;
	wire [14-1:0] node6036;
	wire [14-1:0] node6037;
	wire [14-1:0] node6040;
	wire [14-1:0] node6043;
	wire [14-1:0] node6044;
	wire [14-1:0] node6045;
	wire [14-1:0] node6046;
	wire [14-1:0] node6049;
	wire [14-1:0] node6052;
	wire [14-1:0] node6053;
	wire [14-1:0] node6056;
	wire [14-1:0] node6059;
	wire [14-1:0] node6060;
	wire [14-1:0] node6061;
	wire [14-1:0] node6064;
	wire [14-1:0] node6067;
	wire [14-1:0] node6068;
	wire [14-1:0] node6071;
	wire [14-1:0] node6074;
	wire [14-1:0] node6075;
	wire [14-1:0] node6076;
	wire [14-1:0] node6077;
	wire [14-1:0] node6078;
	wire [14-1:0] node6079;
	wire [14-1:0] node6080;
	wire [14-1:0] node6083;
	wire [14-1:0] node6086;
	wire [14-1:0] node6087;
	wire [14-1:0] node6090;
	wire [14-1:0] node6093;
	wire [14-1:0] node6094;
	wire [14-1:0] node6095;
	wire [14-1:0] node6098;
	wire [14-1:0] node6101;
	wire [14-1:0] node6102;
	wire [14-1:0] node6105;
	wire [14-1:0] node6108;
	wire [14-1:0] node6109;
	wire [14-1:0] node6110;
	wire [14-1:0] node6111;
	wire [14-1:0] node6115;
	wire [14-1:0] node6116;
	wire [14-1:0] node6119;
	wire [14-1:0] node6122;
	wire [14-1:0] node6123;
	wire [14-1:0] node6124;
	wire [14-1:0] node6127;
	wire [14-1:0] node6130;
	wire [14-1:0] node6131;
	wire [14-1:0] node6134;
	wire [14-1:0] node6137;
	wire [14-1:0] node6138;
	wire [14-1:0] node6139;
	wire [14-1:0] node6140;
	wire [14-1:0] node6142;
	wire [14-1:0] node6145;
	wire [14-1:0] node6146;
	wire [14-1:0] node6149;
	wire [14-1:0] node6152;
	wire [14-1:0] node6153;
	wire [14-1:0] node6154;
	wire [14-1:0] node6157;
	wire [14-1:0] node6160;
	wire [14-1:0] node6161;
	wire [14-1:0] node6164;
	wire [14-1:0] node6167;
	wire [14-1:0] node6168;
	wire [14-1:0] node6169;
	wire [14-1:0] node6170;
	wire [14-1:0] node6173;
	wire [14-1:0] node6177;
	wire [14-1:0] node6178;
	wire [14-1:0] node6179;
	wire [14-1:0] node6183;
	wire [14-1:0] node6184;
	wire [14-1:0] node6187;
	wire [14-1:0] node6190;
	wire [14-1:0] node6191;
	wire [14-1:0] node6192;
	wire [14-1:0] node6193;
	wire [14-1:0] node6194;
	wire [14-1:0] node6195;
	wire [14-1:0] node6198;
	wire [14-1:0] node6201;
	wire [14-1:0] node6202;
	wire [14-1:0] node6205;
	wire [14-1:0] node6208;
	wire [14-1:0] node6209;
	wire [14-1:0] node6210;
	wire [14-1:0] node6213;
	wire [14-1:0] node6216;
	wire [14-1:0] node6217;
	wire [14-1:0] node6220;
	wire [14-1:0] node6223;
	wire [14-1:0] node6224;
	wire [14-1:0] node6225;
	wire [14-1:0] node6226;
	wire [14-1:0] node6229;
	wire [14-1:0] node6232;
	wire [14-1:0] node6233;
	wire [14-1:0] node6236;
	wire [14-1:0] node6239;
	wire [14-1:0] node6240;
	wire [14-1:0] node6241;
	wire [14-1:0] node6244;
	wire [14-1:0] node6247;
	wire [14-1:0] node6248;
	wire [14-1:0] node6251;
	wire [14-1:0] node6254;
	wire [14-1:0] node6255;
	wire [14-1:0] node6256;
	wire [14-1:0] node6257;
	wire [14-1:0] node6259;
	wire [14-1:0] node6262;
	wire [14-1:0] node6263;
	wire [14-1:0] node6266;
	wire [14-1:0] node6269;
	wire [14-1:0] node6270;
	wire [14-1:0] node6271;
	wire [14-1:0] node6274;
	wire [14-1:0] node6277;
	wire [14-1:0] node6278;
	wire [14-1:0] node6281;
	wire [14-1:0] node6284;
	wire [14-1:0] node6285;
	wire [14-1:0] node6286;
	wire [14-1:0] node6287;
	wire [14-1:0] node6290;
	wire [14-1:0] node6293;
	wire [14-1:0] node6294;
	wire [14-1:0] node6297;
	wire [14-1:0] node6300;
	wire [14-1:0] node6301;
	wire [14-1:0] node6302;
	wire [14-1:0] node6305;
	wire [14-1:0] node6308;
	wire [14-1:0] node6309;
	wire [14-1:0] node6312;
	wire [14-1:0] node6315;
	wire [14-1:0] node6316;
	wire [14-1:0] node6317;
	wire [14-1:0] node6318;
	wire [14-1:0] node6319;
	wire [14-1:0] node6320;
	wire [14-1:0] node6321;
	wire [14-1:0] node6322;
	wire [14-1:0] node6325;
	wire [14-1:0] node6328;
	wire [14-1:0] node6329;
	wire [14-1:0] node6332;
	wire [14-1:0] node6335;
	wire [14-1:0] node6336;
	wire [14-1:0] node6337;
	wire [14-1:0] node6340;
	wire [14-1:0] node6343;
	wire [14-1:0] node6344;
	wire [14-1:0] node6347;
	wire [14-1:0] node6350;
	wire [14-1:0] node6351;
	wire [14-1:0] node6352;
	wire [14-1:0] node6353;
	wire [14-1:0] node6356;
	wire [14-1:0] node6359;
	wire [14-1:0] node6360;
	wire [14-1:0] node6363;
	wire [14-1:0] node6366;
	wire [14-1:0] node6367;
	wire [14-1:0] node6368;
	wire [14-1:0] node6371;
	wire [14-1:0] node6374;
	wire [14-1:0] node6375;
	wire [14-1:0] node6378;
	wire [14-1:0] node6381;
	wire [14-1:0] node6382;
	wire [14-1:0] node6383;
	wire [14-1:0] node6384;
	wire [14-1:0] node6385;
	wire [14-1:0] node6388;
	wire [14-1:0] node6391;
	wire [14-1:0] node6392;
	wire [14-1:0] node6395;
	wire [14-1:0] node6398;
	wire [14-1:0] node6399;
	wire [14-1:0] node6401;
	wire [14-1:0] node6404;
	wire [14-1:0] node6405;
	wire [14-1:0] node6408;
	wire [14-1:0] node6411;
	wire [14-1:0] node6412;
	wire [14-1:0] node6413;
	wire [14-1:0] node6414;
	wire [14-1:0] node6417;
	wire [14-1:0] node6420;
	wire [14-1:0] node6421;
	wire [14-1:0] node6424;
	wire [14-1:0] node6427;
	wire [14-1:0] node6428;
	wire [14-1:0] node6429;
	wire [14-1:0] node6432;
	wire [14-1:0] node6435;
	wire [14-1:0] node6436;
	wire [14-1:0] node6439;
	wire [14-1:0] node6442;
	wire [14-1:0] node6443;
	wire [14-1:0] node6444;
	wire [14-1:0] node6445;
	wire [14-1:0] node6446;
	wire [14-1:0] node6447;
	wire [14-1:0] node6450;
	wire [14-1:0] node6453;
	wire [14-1:0] node6454;
	wire [14-1:0] node6457;
	wire [14-1:0] node6460;
	wire [14-1:0] node6461;
	wire [14-1:0] node6462;
	wire [14-1:0] node6465;
	wire [14-1:0] node6468;
	wire [14-1:0] node6471;
	wire [14-1:0] node6472;
	wire [14-1:0] node6473;
	wire [14-1:0] node6474;
	wire [14-1:0] node6477;
	wire [14-1:0] node6480;
	wire [14-1:0] node6481;
	wire [14-1:0] node6484;
	wire [14-1:0] node6487;
	wire [14-1:0] node6488;
	wire [14-1:0] node6490;
	wire [14-1:0] node6493;
	wire [14-1:0] node6494;
	wire [14-1:0] node6497;
	wire [14-1:0] node6500;
	wire [14-1:0] node6501;
	wire [14-1:0] node6502;
	wire [14-1:0] node6503;
	wire [14-1:0] node6504;
	wire [14-1:0] node6507;
	wire [14-1:0] node6510;
	wire [14-1:0] node6511;
	wire [14-1:0] node6514;
	wire [14-1:0] node6517;
	wire [14-1:0] node6518;
	wire [14-1:0] node6519;
	wire [14-1:0] node6522;
	wire [14-1:0] node6525;
	wire [14-1:0] node6526;
	wire [14-1:0] node6529;
	wire [14-1:0] node6532;
	wire [14-1:0] node6533;
	wire [14-1:0] node6534;
	wire [14-1:0] node6535;
	wire [14-1:0] node6538;
	wire [14-1:0] node6541;
	wire [14-1:0] node6542;
	wire [14-1:0] node6546;
	wire [14-1:0] node6547;
	wire [14-1:0] node6548;
	wire [14-1:0] node6551;
	wire [14-1:0] node6554;
	wire [14-1:0] node6555;
	wire [14-1:0] node6558;
	wire [14-1:0] node6561;
	wire [14-1:0] node6562;
	wire [14-1:0] node6563;
	wire [14-1:0] node6564;
	wire [14-1:0] node6565;
	wire [14-1:0] node6566;
	wire [14-1:0] node6567;
	wire [14-1:0] node6570;
	wire [14-1:0] node6573;
	wire [14-1:0] node6574;
	wire [14-1:0] node6577;
	wire [14-1:0] node6580;
	wire [14-1:0] node6581;
	wire [14-1:0] node6582;
	wire [14-1:0] node6585;
	wire [14-1:0] node6588;
	wire [14-1:0] node6589;
	wire [14-1:0] node6592;
	wire [14-1:0] node6595;
	wire [14-1:0] node6596;
	wire [14-1:0] node6597;
	wire [14-1:0] node6598;
	wire [14-1:0] node6602;
	wire [14-1:0] node6603;
	wire [14-1:0] node6606;
	wire [14-1:0] node6609;
	wire [14-1:0] node6610;
	wire [14-1:0] node6611;
	wire [14-1:0] node6614;
	wire [14-1:0] node6617;
	wire [14-1:0] node6618;
	wire [14-1:0] node6621;
	wire [14-1:0] node6624;
	wire [14-1:0] node6625;
	wire [14-1:0] node6626;
	wire [14-1:0] node6627;
	wire [14-1:0] node6629;
	wire [14-1:0] node6632;
	wire [14-1:0] node6633;
	wire [14-1:0] node6636;
	wire [14-1:0] node6639;
	wire [14-1:0] node6640;
	wire [14-1:0] node6641;
	wire [14-1:0] node6644;
	wire [14-1:0] node6647;
	wire [14-1:0] node6648;
	wire [14-1:0] node6651;
	wire [14-1:0] node6654;
	wire [14-1:0] node6655;
	wire [14-1:0] node6656;
	wire [14-1:0] node6657;
	wire [14-1:0] node6660;
	wire [14-1:0] node6663;
	wire [14-1:0] node6664;
	wire [14-1:0] node6667;
	wire [14-1:0] node6670;
	wire [14-1:0] node6671;
	wire [14-1:0] node6672;
	wire [14-1:0] node6675;
	wire [14-1:0] node6678;
	wire [14-1:0] node6679;
	wire [14-1:0] node6682;
	wire [14-1:0] node6685;
	wire [14-1:0] node6686;
	wire [14-1:0] node6687;
	wire [14-1:0] node6688;
	wire [14-1:0] node6689;
	wire [14-1:0] node6691;
	wire [14-1:0] node6694;
	wire [14-1:0] node6695;
	wire [14-1:0] node6698;
	wire [14-1:0] node6701;
	wire [14-1:0] node6702;
	wire [14-1:0] node6703;
	wire [14-1:0] node6706;
	wire [14-1:0] node6709;
	wire [14-1:0] node6710;
	wire [14-1:0] node6713;
	wire [14-1:0] node6716;
	wire [14-1:0] node6717;
	wire [14-1:0] node6718;
	wire [14-1:0] node6719;
	wire [14-1:0] node6722;
	wire [14-1:0] node6725;
	wire [14-1:0] node6726;
	wire [14-1:0] node6729;
	wire [14-1:0] node6732;
	wire [14-1:0] node6733;
	wire [14-1:0] node6734;
	wire [14-1:0] node6737;
	wire [14-1:0] node6740;
	wire [14-1:0] node6742;
	wire [14-1:0] node6745;
	wire [14-1:0] node6746;
	wire [14-1:0] node6747;
	wire [14-1:0] node6748;
	wire [14-1:0] node6749;
	wire [14-1:0] node6752;
	wire [14-1:0] node6755;
	wire [14-1:0] node6756;
	wire [14-1:0] node6759;
	wire [14-1:0] node6762;
	wire [14-1:0] node6763;
	wire [14-1:0] node6764;
	wire [14-1:0] node6767;
	wire [14-1:0] node6770;
	wire [14-1:0] node6771;
	wire [14-1:0] node6775;
	wire [14-1:0] node6776;
	wire [14-1:0] node6777;
	wire [14-1:0] node6779;
	wire [14-1:0] node6782;
	wire [14-1:0] node6783;
	wire [14-1:0] node6786;
	wire [14-1:0] node6789;
	wire [14-1:0] node6790;
	wire [14-1:0] node6791;
	wire [14-1:0] node6794;
	wire [14-1:0] node6797;
	wire [14-1:0] node6798;
	wire [14-1:0] node6801;
	wire [14-1:0] node6804;
	wire [14-1:0] node6805;
	wire [14-1:0] node6806;
	wire [14-1:0] node6807;
	wire [14-1:0] node6808;
	wire [14-1:0] node6809;
	wire [14-1:0] node6810;
	wire [14-1:0] node6811;
	wire [14-1:0] node6813;
	wire [14-1:0] node6816;
	wire [14-1:0] node6817;
	wire [14-1:0] node6820;
	wire [14-1:0] node6823;
	wire [14-1:0] node6824;
	wire [14-1:0] node6825;
	wire [14-1:0] node6828;
	wire [14-1:0] node6831;
	wire [14-1:0] node6832;
	wire [14-1:0] node6835;
	wire [14-1:0] node6838;
	wire [14-1:0] node6839;
	wire [14-1:0] node6840;
	wire [14-1:0] node6841;
	wire [14-1:0] node6844;
	wire [14-1:0] node6847;
	wire [14-1:0] node6848;
	wire [14-1:0] node6851;
	wire [14-1:0] node6854;
	wire [14-1:0] node6855;
	wire [14-1:0] node6856;
	wire [14-1:0] node6859;
	wire [14-1:0] node6862;
	wire [14-1:0] node6863;
	wire [14-1:0] node6866;
	wire [14-1:0] node6869;
	wire [14-1:0] node6870;
	wire [14-1:0] node6871;
	wire [14-1:0] node6872;
	wire [14-1:0] node6874;
	wire [14-1:0] node6877;
	wire [14-1:0] node6878;
	wire [14-1:0] node6882;
	wire [14-1:0] node6883;
	wire [14-1:0] node6884;
	wire [14-1:0] node6888;
	wire [14-1:0] node6889;
	wire [14-1:0] node6892;
	wire [14-1:0] node6895;
	wire [14-1:0] node6896;
	wire [14-1:0] node6897;
	wire [14-1:0] node6899;
	wire [14-1:0] node6902;
	wire [14-1:0] node6903;
	wire [14-1:0] node6906;
	wire [14-1:0] node6909;
	wire [14-1:0] node6910;
	wire [14-1:0] node6912;
	wire [14-1:0] node6915;
	wire [14-1:0] node6918;
	wire [14-1:0] node6919;
	wire [14-1:0] node6920;
	wire [14-1:0] node6921;
	wire [14-1:0] node6922;
	wire [14-1:0] node6923;
	wire [14-1:0] node6926;
	wire [14-1:0] node6929;
	wire [14-1:0] node6930;
	wire [14-1:0] node6933;
	wire [14-1:0] node6936;
	wire [14-1:0] node6937;
	wire [14-1:0] node6938;
	wire [14-1:0] node6941;
	wire [14-1:0] node6944;
	wire [14-1:0] node6945;
	wire [14-1:0] node6948;
	wire [14-1:0] node6951;
	wire [14-1:0] node6952;
	wire [14-1:0] node6953;
	wire [14-1:0] node6954;
	wire [14-1:0] node6957;
	wire [14-1:0] node6960;
	wire [14-1:0] node6961;
	wire [14-1:0] node6964;
	wire [14-1:0] node6967;
	wire [14-1:0] node6968;
	wire [14-1:0] node6969;
	wire [14-1:0] node6972;
	wire [14-1:0] node6975;
	wire [14-1:0] node6976;
	wire [14-1:0] node6979;
	wire [14-1:0] node6982;
	wire [14-1:0] node6983;
	wire [14-1:0] node6984;
	wire [14-1:0] node6985;
	wire [14-1:0] node6986;
	wire [14-1:0] node6989;
	wire [14-1:0] node6992;
	wire [14-1:0] node6993;
	wire [14-1:0] node6996;
	wire [14-1:0] node6999;
	wire [14-1:0] node7000;
	wire [14-1:0] node7001;
	wire [14-1:0] node7004;
	wire [14-1:0] node7007;
	wire [14-1:0] node7008;
	wire [14-1:0] node7011;
	wire [14-1:0] node7014;
	wire [14-1:0] node7015;
	wire [14-1:0] node7016;
	wire [14-1:0] node7017;
	wire [14-1:0] node7020;
	wire [14-1:0] node7023;
	wire [14-1:0] node7024;
	wire [14-1:0] node7027;
	wire [14-1:0] node7030;
	wire [14-1:0] node7031;
	wire [14-1:0] node7033;
	wire [14-1:0] node7036;
	wire [14-1:0] node7037;
	wire [14-1:0] node7040;
	wire [14-1:0] node7043;
	wire [14-1:0] node7044;
	wire [14-1:0] node7045;
	wire [14-1:0] node7046;
	wire [14-1:0] node7047;
	wire [14-1:0] node7048;
	wire [14-1:0] node7049;
	wire [14-1:0] node7053;
	wire [14-1:0] node7054;
	wire [14-1:0] node7057;
	wire [14-1:0] node7060;
	wire [14-1:0] node7061;
	wire [14-1:0] node7062;
	wire [14-1:0] node7065;
	wire [14-1:0] node7068;
	wire [14-1:0] node7069;
	wire [14-1:0] node7072;
	wire [14-1:0] node7075;
	wire [14-1:0] node7076;
	wire [14-1:0] node7077;
	wire [14-1:0] node7079;
	wire [14-1:0] node7082;
	wire [14-1:0] node7083;
	wire [14-1:0] node7086;
	wire [14-1:0] node7089;
	wire [14-1:0] node7090;
	wire [14-1:0] node7091;
	wire [14-1:0] node7094;
	wire [14-1:0] node7097;
	wire [14-1:0] node7098;
	wire [14-1:0] node7101;
	wire [14-1:0] node7104;
	wire [14-1:0] node7105;
	wire [14-1:0] node7106;
	wire [14-1:0] node7107;
	wire [14-1:0] node7108;
	wire [14-1:0] node7111;
	wire [14-1:0] node7114;
	wire [14-1:0] node7115;
	wire [14-1:0] node7118;
	wire [14-1:0] node7121;
	wire [14-1:0] node7122;
	wire [14-1:0] node7123;
	wire [14-1:0] node7126;
	wire [14-1:0] node7129;
	wire [14-1:0] node7130;
	wire [14-1:0] node7133;
	wire [14-1:0] node7136;
	wire [14-1:0] node7137;
	wire [14-1:0] node7139;
	wire [14-1:0] node7140;
	wire [14-1:0] node7144;
	wire [14-1:0] node7145;
	wire [14-1:0] node7146;
	wire [14-1:0] node7149;
	wire [14-1:0] node7152;
	wire [14-1:0] node7153;
	wire [14-1:0] node7156;
	wire [14-1:0] node7159;
	wire [14-1:0] node7160;
	wire [14-1:0] node7161;
	wire [14-1:0] node7162;
	wire [14-1:0] node7163;
	wire [14-1:0] node7164;
	wire [14-1:0] node7167;
	wire [14-1:0] node7170;
	wire [14-1:0] node7171;
	wire [14-1:0] node7174;
	wire [14-1:0] node7177;
	wire [14-1:0] node7178;
	wire [14-1:0] node7179;
	wire [14-1:0] node7182;
	wire [14-1:0] node7185;
	wire [14-1:0] node7186;
	wire [14-1:0] node7189;
	wire [14-1:0] node7192;
	wire [14-1:0] node7193;
	wire [14-1:0] node7194;
	wire [14-1:0] node7195;
	wire [14-1:0] node7198;
	wire [14-1:0] node7201;
	wire [14-1:0] node7203;
	wire [14-1:0] node7206;
	wire [14-1:0] node7207;
	wire [14-1:0] node7208;
	wire [14-1:0] node7211;
	wire [14-1:0] node7214;
	wire [14-1:0] node7215;
	wire [14-1:0] node7218;
	wire [14-1:0] node7221;
	wire [14-1:0] node7222;
	wire [14-1:0] node7223;
	wire [14-1:0] node7224;
	wire [14-1:0] node7225;
	wire [14-1:0] node7228;
	wire [14-1:0] node7231;
	wire [14-1:0] node7232;
	wire [14-1:0] node7235;
	wire [14-1:0] node7238;
	wire [14-1:0] node7239;
	wire [14-1:0] node7240;
	wire [14-1:0] node7243;
	wire [14-1:0] node7246;
	wire [14-1:0] node7248;
	wire [14-1:0] node7251;
	wire [14-1:0] node7252;
	wire [14-1:0] node7253;
	wire [14-1:0] node7254;
	wire [14-1:0] node7258;
	wire [14-1:0] node7259;
	wire [14-1:0] node7262;
	wire [14-1:0] node7265;
	wire [14-1:0] node7266;
	wire [14-1:0] node7267;
	wire [14-1:0] node7270;
	wire [14-1:0] node7273;
	wire [14-1:0] node7274;
	wire [14-1:0] node7277;
	wire [14-1:0] node7280;
	wire [14-1:0] node7281;
	wire [14-1:0] node7282;
	wire [14-1:0] node7283;
	wire [14-1:0] node7284;
	wire [14-1:0] node7285;
	wire [14-1:0] node7286;
	wire [14-1:0] node7287;
	wire [14-1:0] node7290;
	wire [14-1:0] node7293;
	wire [14-1:0] node7294;
	wire [14-1:0] node7297;
	wire [14-1:0] node7300;
	wire [14-1:0] node7301;
	wire [14-1:0] node7302;
	wire [14-1:0] node7305;
	wire [14-1:0] node7308;
	wire [14-1:0] node7310;
	wire [14-1:0] node7313;
	wire [14-1:0] node7314;
	wire [14-1:0] node7315;
	wire [14-1:0] node7316;
	wire [14-1:0] node7319;
	wire [14-1:0] node7322;
	wire [14-1:0] node7323;
	wire [14-1:0] node7326;
	wire [14-1:0] node7329;
	wire [14-1:0] node7330;
	wire [14-1:0] node7331;
	wire [14-1:0] node7334;
	wire [14-1:0] node7337;
	wire [14-1:0] node7338;
	wire [14-1:0] node7342;
	wire [14-1:0] node7343;
	wire [14-1:0] node7344;
	wire [14-1:0] node7345;
	wire [14-1:0] node7346;
	wire [14-1:0] node7349;
	wire [14-1:0] node7352;
	wire [14-1:0] node7353;
	wire [14-1:0] node7356;
	wire [14-1:0] node7359;
	wire [14-1:0] node7360;
	wire [14-1:0] node7361;
	wire [14-1:0] node7364;
	wire [14-1:0] node7367;
	wire [14-1:0] node7368;
	wire [14-1:0] node7372;
	wire [14-1:0] node7373;
	wire [14-1:0] node7374;
	wire [14-1:0] node7375;
	wire [14-1:0] node7378;
	wire [14-1:0] node7381;
	wire [14-1:0] node7382;
	wire [14-1:0] node7385;
	wire [14-1:0] node7388;
	wire [14-1:0] node7389;
	wire [14-1:0] node7390;
	wire [14-1:0] node7393;
	wire [14-1:0] node7396;
	wire [14-1:0] node7397;
	wire [14-1:0] node7400;
	wire [14-1:0] node7403;
	wire [14-1:0] node7404;
	wire [14-1:0] node7405;
	wire [14-1:0] node7406;
	wire [14-1:0] node7407;
	wire [14-1:0] node7408;
	wire [14-1:0] node7411;
	wire [14-1:0] node7414;
	wire [14-1:0] node7415;
	wire [14-1:0] node7418;
	wire [14-1:0] node7421;
	wire [14-1:0] node7422;
	wire [14-1:0] node7425;
	wire [14-1:0] node7426;
	wire [14-1:0] node7430;
	wire [14-1:0] node7431;
	wire [14-1:0] node7432;
	wire [14-1:0] node7433;
	wire [14-1:0] node7437;
	wire [14-1:0] node7438;
	wire [14-1:0] node7441;
	wire [14-1:0] node7444;
	wire [14-1:0] node7445;
	wire [14-1:0] node7446;
	wire [14-1:0] node7449;
	wire [14-1:0] node7452;
	wire [14-1:0] node7453;
	wire [14-1:0] node7456;
	wire [14-1:0] node7459;
	wire [14-1:0] node7460;
	wire [14-1:0] node7461;
	wire [14-1:0] node7462;
	wire [14-1:0] node7463;
	wire [14-1:0] node7466;
	wire [14-1:0] node7469;
	wire [14-1:0] node7470;
	wire [14-1:0] node7473;
	wire [14-1:0] node7476;
	wire [14-1:0] node7477;
	wire [14-1:0] node7478;
	wire [14-1:0] node7481;
	wire [14-1:0] node7484;
	wire [14-1:0] node7485;
	wire [14-1:0] node7488;
	wire [14-1:0] node7491;
	wire [14-1:0] node7492;
	wire [14-1:0] node7493;
	wire [14-1:0] node7494;
	wire [14-1:0] node7497;
	wire [14-1:0] node7500;
	wire [14-1:0] node7501;
	wire [14-1:0] node7504;
	wire [14-1:0] node7507;
	wire [14-1:0] node7508;
	wire [14-1:0] node7509;
	wire [14-1:0] node7512;
	wire [14-1:0] node7515;
	wire [14-1:0] node7516;
	wire [14-1:0] node7519;
	wire [14-1:0] node7522;
	wire [14-1:0] node7523;
	wire [14-1:0] node7524;
	wire [14-1:0] node7525;
	wire [14-1:0] node7526;
	wire [14-1:0] node7527;
	wire [14-1:0] node7528;
	wire [14-1:0] node7531;
	wire [14-1:0] node7534;
	wire [14-1:0] node7535;
	wire [14-1:0] node7538;
	wire [14-1:0] node7541;
	wire [14-1:0] node7542;
	wire [14-1:0] node7543;
	wire [14-1:0] node7546;
	wire [14-1:0] node7549;
	wire [14-1:0] node7550;
	wire [14-1:0] node7554;
	wire [14-1:0] node7555;
	wire [14-1:0] node7556;
	wire [14-1:0] node7557;
	wire [14-1:0] node7560;
	wire [14-1:0] node7563;
	wire [14-1:0] node7564;
	wire [14-1:0] node7567;
	wire [14-1:0] node7570;
	wire [14-1:0] node7571;
	wire [14-1:0] node7572;
	wire [14-1:0] node7575;
	wire [14-1:0] node7578;
	wire [14-1:0] node7579;
	wire [14-1:0] node7582;
	wire [14-1:0] node7585;
	wire [14-1:0] node7586;
	wire [14-1:0] node7587;
	wire [14-1:0] node7588;
	wire [14-1:0] node7589;
	wire [14-1:0] node7592;
	wire [14-1:0] node7595;
	wire [14-1:0] node7596;
	wire [14-1:0] node7599;
	wire [14-1:0] node7602;
	wire [14-1:0] node7603;
	wire [14-1:0] node7604;
	wire [14-1:0] node7607;
	wire [14-1:0] node7610;
	wire [14-1:0] node7611;
	wire [14-1:0] node7614;
	wire [14-1:0] node7617;
	wire [14-1:0] node7618;
	wire [14-1:0] node7619;
	wire [14-1:0] node7620;
	wire [14-1:0] node7623;
	wire [14-1:0] node7626;
	wire [14-1:0] node7627;
	wire [14-1:0] node7630;
	wire [14-1:0] node7633;
	wire [14-1:0] node7634;
	wire [14-1:0] node7635;
	wire [14-1:0] node7638;
	wire [14-1:0] node7641;
	wire [14-1:0] node7642;
	wire [14-1:0] node7645;
	wire [14-1:0] node7648;
	wire [14-1:0] node7649;
	wire [14-1:0] node7650;
	wire [14-1:0] node7651;
	wire [14-1:0] node7652;
	wire [14-1:0] node7653;
	wire [14-1:0] node7656;
	wire [14-1:0] node7659;
	wire [14-1:0] node7660;
	wire [14-1:0] node7663;
	wire [14-1:0] node7666;
	wire [14-1:0] node7667;
	wire [14-1:0] node7668;
	wire [14-1:0] node7671;
	wire [14-1:0] node7674;
	wire [14-1:0] node7675;
	wire [14-1:0] node7678;
	wire [14-1:0] node7681;
	wire [14-1:0] node7682;
	wire [14-1:0] node7683;
	wire [14-1:0] node7684;
	wire [14-1:0] node7687;
	wire [14-1:0] node7690;
	wire [14-1:0] node7691;
	wire [14-1:0] node7694;
	wire [14-1:0] node7697;
	wire [14-1:0] node7698;
	wire [14-1:0] node7699;
	wire [14-1:0] node7702;
	wire [14-1:0] node7705;
	wire [14-1:0] node7706;
	wire [14-1:0] node7709;
	wire [14-1:0] node7712;
	wire [14-1:0] node7713;
	wire [14-1:0] node7714;
	wire [14-1:0] node7715;
	wire [14-1:0] node7717;
	wire [14-1:0] node7720;
	wire [14-1:0] node7721;
	wire [14-1:0] node7724;
	wire [14-1:0] node7727;
	wire [14-1:0] node7728;
	wire [14-1:0] node7729;
	wire [14-1:0] node7732;
	wire [14-1:0] node7735;
	wire [14-1:0] node7736;
	wire [14-1:0] node7739;
	wire [14-1:0] node7742;
	wire [14-1:0] node7743;
	wire [14-1:0] node7744;
	wire [14-1:0] node7745;
	wire [14-1:0] node7748;
	wire [14-1:0] node7751;
	wire [14-1:0] node7752;
	wire [14-1:0] node7755;
	wire [14-1:0] node7758;
	wire [14-1:0] node7759;
	wire [14-1:0] node7760;
	wire [14-1:0] node7763;
	wire [14-1:0] node7766;
	wire [14-1:0] node7767;
	wire [14-1:0] node7770;

	assign outp = (inp[6]) ? node3882 : node1;
		assign node1 = (inp[12]) ? node1941 : node2;
			assign node2 = (inp[7]) ? node978 : node3;
				assign node3 = (inp[10]) ? node493 : node4;
					assign node4 = (inp[0]) ? node248 : node5;
						assign node5 = (inp[3]) ? node127 : node6;
							assign node6 = (inp[13]) ? node66 : node7;
								assign node7 = (inp[9]) ? node37 : node8;
									assign node8 = (inp[11]) ? node22 : node9;
										assign node9 = (inp[4]) ? node15 : node10;
											assign node10 = (inp[2]) ? 14'b00111111111111 : node11;
												assign node11 = (inp[8]) ? 14'b00111111111111 : 14'b01111111111111;
											assign node15 = (inp[1]) ? node19 : node16;
												assign node16 = (inp[2]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node19 = (inp[5]) ? 14'b00001111111111 : 14'b00011111111111;
										assign node22 = (inp[4]) ? node30 : node23;
											assign node23 = (inp[2]) ? node27 : node24;
												assign node24 = (inp[1]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node27 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node30 = (inp[5]) ? node34 : node31;
												assign node31 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node34 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node37 = (inp[4]) ? node53 : node38;
										assign node38 = (inp[11]) ? node46 : node39;
											assign node39 = (inp[2]) ? node43 : node40;
												assign node40 = (inp[8]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node43 = (inp[1]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node46 = (inp[2]) ? node50 : node47;
												assign node47 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node50 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node53 = (inp[2]) ? node61 : node54;
											assign node54 = (inp[8]) ? node58 : node55;
												assign node55 = (inp[5]) ? 14'b00001111111111 : 14'b00001111111111;
												assign node58 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node61 = (inp[5]) ? node63 : 14'b00001111111111;
												assign node63 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node66 = (inp[4]) ? node96 : node67;
									assign node67 = (inp[2]) ? node83 : node68;
										assign node68 = (inp[1]) ? node76 : node69;
											assign node69 = (inp[8]) ? node73 : node70;
												assign node70 = (inp[9]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node73 = (inp[9]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node76 = (inp[9]) ? node80 : node77;
												assign node77 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node80 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node83 = (inp[11]) ? node91 : node84;
											assign node84 = (inp[8]) ? node88 : node85;
												assign node85 = (inp[9]) ? 14'b00001111111111 : 14'b00001111111111;
												assign node88 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node91 = (inp[1]) ? node93 : 14'b00000111111111;
												assign node93 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node96 = (inp[9]) ? node112 : node97;
										assign node97 = (inp[11]) ? node105 : node98;
											assign node98 = (inp[1]) ? node102 : node99;
												assign node99 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node102 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node105 = (inp[5]) ? node109 : node106;
												assign node106 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node109 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node112 = (inp[2]) ? node120 : node113;
											assign node113 = (inp[5]) ? node117 : node114;
												assign node114 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node117 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node120 = (inp[1]) ? node124 : node121;
												assign node121 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node124 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node127 = (inp[9]) ? node189 : node128;
								assign node128 = (inp[4]) ? node158 : node129;
									assign node129 = (inp[8]) ? node145 : node130;
										assign node130 = (inp[2]) ? node138 : node131;
											assign node131 = (inp[1]) ? node135 : node132;
												assign node132 = (inp[13]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node135 = (inp[13]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node138 = (inp[5]) ? node142 : node139;
												assign node139 = (inp[13]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node142 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node145 = (inp[11]) ? node153 : node146;
											assign node146 = (inp[5]) ? node150 : node147;
												assign node147 = (inp[2]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node150 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node153 = (inp[5]) ? node155 : 14'b00000111111111;
												assign node155 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node158 = (inp[1]) ? node174 : node159;
										assign node159 = (inp[13]) ? node167 : node160;
											assign node160 = (inp[8]) ? node164 : node161;
												assign node161 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node164 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node167 = (inp[2]) ? node171 : node168;
												assign node168 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node171 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node174 = (inp[11]) ? node182 : node175;
											assign node175 = (inp[5]) ? node179 : node176;
												assign node176 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node179 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node182 = (inp[13]) ? node186 : node183;
												assign node183 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node186 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node189 = (inp[13]) ? node221 : node190;
									assign node190 = (inp[2]) ? node206 : node191;
										assign node191 = (inp[5]) ? node199 : node192;
											assign node192 = (inp[4]) ? node196 : node193;
												assign node193 = (inp[8]) ? 14'b00000111111111 : 14'b00011111111111;
												assign node196 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node199 = (inp[8]) ? node203 : node200;
												assign node200 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node203 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node206 = (inp[5]) ? node214 : node207;
											assign node207 = (inp[11]) ? node211 : node208;
												assign node208 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node211 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node214 = (inp[4]) ? node218 : node215;
												assign node215 = (inp[1]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node218 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node221 = (inp[1]) ? node235 : node222;
										assign node222 = (inp[5]) ? node228 : node223;
											assign node223 = (inp[11]) ? node225 : 14'b00001111111111;
												assign node225 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node228 = (inp[4]) ? node232 : node229;
												assign node229 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node232 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node235 = (inp[5]) ? node241 : node236;
											assign node236 = (inp[8]) ? node238 : 14'b00000011111111;
												assign node238 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node241 = (inp[2]) ? node245 : node242;
												assign node242 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node245 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node248 = (inp[5]) ? node368 : node249;
							assign node249 = (inp[11]) ? node307 : node250;
								assign node250 = (inp[1]) ? node278 : node251;
									assign node251 = (inp[3]) ? node265 : node252;
										assign node252 = (inp[9]) ? node258 : node253;
											assign node253 = (inp[4]) ? node255 : 14'b00111111111111;
												assign node255 = (inp[13]) ? 14'b00011111111111 : 14'b00011111111111;
											assign node258 = (inp[13]) ? node262 : node259;
												assign node259 = (inp[4]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node262 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node265 = (inp[2]) ? node273 : node266;
											assign node266 = (inp[9]) ? node270 : node267;
												assign node267 = (inp[13]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node270 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node273 = (inp[13]) ? 14'b00000111111111 : node274;
												assign node274 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node278 = (inp[8]) ? node294 : node279;
										assign node279 = (inp[4]) ? node287 : node280;
											assign node280 = (inp[2]) ? node284 : node281;
												assign node281 = (inp[3]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node284 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node287 = (inp[9]) ? node291 : node288;
												assign node288 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node291 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node294 = (inp[3]) ? node300 : node295;
											assign node295 = (inp[4]) ? 14'b00000011111111 : node296;
												assign node296 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node300 = (inp[9]) ? node304 : node301;
												assign node301 = (inp[2]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node304 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node307 = (inp[13]) ? node339 : node308;
									assign node308 = (inp[1]) ? node324 : node309;
										assign node309 = (inp[3]) ? node317 : node310;
											assign node310 = (inp[2]) ? node314 : node311;
												assign node311 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node314 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node317 = (inp[4]) ? node321 : node318;
												assign node318 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node321 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node324 = (inp[9]) ? node332 : node325;
											assign node325 = (inp[4]) ? node329 : node326;
												assign node326 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node329 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node332 = (inp[3]) ? node336 : node333;
												assign node333 = (inp[2]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node336 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node339 = (inp[8]) ? node355 : node340;
										assign node340 = (inp[3]) ? node348 : node341;
											assign node341 = (inp[4]) ? node345 : node342;
												assign node342 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node345 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node348 = (inp[9]) ? node352 : node349;
												assign node349 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node352 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node355 = (inp[4]) ? node363 : node356;
											assign node356 = (inp[9]) ? node360 : node357;
												assign node357 = (inp[1]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node360 = (inp[1]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node363 = (inp[9]) ? node365 : 14'b00000001111111;
												assign node365 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node368 = (inp[1]) ? node432 : node369;
								assign node369 = (inp[8]) ? node401 : node370;
									assign node370 = (inp[4]) ? node386 : node371;
										assign node371 = (inp[11]) ? node379 : node372;
											assign node372 = (inp[2]) ? node376 : node373;
												assign node373 = (inp[3]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node376 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node379 = (inp[3]) ? node383 : node380;
												assign node380 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node383 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node386 = (inp[11]) ? node394 : node387;
											assign node387 = (inp[2]) ? node391 : node388;
												assign node388 = (inp[9]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node391 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node394 = (inp[9]) ? node398 : node395;
												assign node395 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node398 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node401 = (inp[11]) ? node417 : node402;
										assign node402 = (inp[4]) ? node410 : node403;
											assign node403 = (inp[13]) ? node407 : node404;
												assign node404 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node407 = (inp[3]) ? 14'b00000011111111 : 14'b00001111111111;
											assign node410 = (inp[9]) ? node414 : node411;
												assign node411 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node414 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node417 = (inp[13]) ? node425 : node418;
											assign node418 = (inp[3]) ? node422 : node419;
												assign node419 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node422 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node425 = (inp[9]) ? node429 : node426;
												assign node426 = (inp[2]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node429 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node432 = (inp[13]) ? node464 : node433;
									assign node433 = (inp[2]) ? node449 : node434;
										assign node434 = (inp[3]) ? node442 : node435;
											assign node435 = (inp[11]) ? node439 : node436;
												assign node436 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node439 = (inp[9]) ? 14'b00000011111111 : 14'b00000011111111;
											assign node442 = (inp[9]) ? node446 : node443;
												assign node443 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node446 = (inp[4]) ? 14'b00000001111111 : 14'b00000001111111;
										assign node449 = (inp[4]) ? node457 : node450;
											assign node450 = (inp[11]) ? node454 : node451;
												assign node451 = (inp[3]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node454 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node457 = (inp[8]) ? node461 : node458;
												assign node458 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node461 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node464 = (inp[3]) ? node480 : node465;
										assign node465 = (inp[2]) ? node473 : node466;
											assign node466 = (inp[11]) ? node470 : node467;
												assign node467 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node470 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node473 = (inp[9]) ? node477 : node474;
												assign node474 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node477 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node480 = (inp[11]) ? node488 : node481;
											assign node481 = (inp[4]) ? node485 : node482;
												assign node482 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node485 = (inp[8]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node488 = (inp[8]) ? node490 : 14'b00000000111111;
												assign node490 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
					assign node493 = (inp[2]) ? node741 : node494;
						assign node494 = (inp[11]) ? node620 : node495;
							assign node495 = (inp[9]) ? node559 : node496;
								assign node496 = (inp[4]) ? node528 : node497;
									assign node497 = (inp[3]) ? node513 : node498;
										assign node498 = (inp[5]) ? node506 : node499;
											assign node499 = (inp[13]) ? node503 : node500;
												assign node500 = (inp[8]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node503 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node506 = (inp[0]) ? node510 : node507;
												assign node507 = (inp[1]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node510 = (inp[13]) ? 14'b00000011111111 : 14'b00001111111111;
										assign node513 = (inp[13]) ? node521 : node514;
											assign node514 = (inp[0]) ? node518 : node515;
												assign node515 = (inp[1]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node518 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node521 = (inp[0]) ? node525 : node522;
												assign node522 = (inp[1]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node525 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node528 = (inp[5]) ? node544 : node529;
										assign node529 = (inp[1]) ? node537 : node530;
											assign node530 = (inp[8]) ? node534 : node531;
												assign node531 = (inp[0]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node534 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node537 = (inp[13]) ? node541 : node538;
												assign node538 = (inp[8]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node541 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node544 = (inp[8]) ? node552 : node545;
											assign node545 = (inp[1]) ? node549 : node546;
												assign node546 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node549 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node552 = (inp[3]) ? node556 : node553;
												assign node553 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node556 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node559 = (inp[4]) ? node591 : node560;
									assign node560 = (inp[0]) ? node576 : node561;
										assign node561 = (inp[3]) ? node569 : node562;
											assign node562 = (inp[5]) ? node566 : node563;
												assign node563 = (inp[13]) ? 14'b00011111111111 : 14'b00011111111111;
												assign node566 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node569 = (inp[5]) ? node573 : node570;
												assign node570 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node573 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node576 = (inp[5]) ? node584 : node577;
											assign node577 = (inp[1]) ? node581 : node578;
												assign node578 = (inp[3]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node581 = (inp[13]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node584 = (inp[13]) ? node588 : node585;
												assign node585 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node588 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node591 = (inp[5]) ? node607 : node592;
										assign node592 = (inp[1]) ? node600 : node593;
											assign node593 = (inp[13]) ? node597 : node594;
												assign node594 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node597 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node600 = (inp[0]) ? node604 : node601;
												assign node601 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node604 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node607 = (inp[8]) ? node615 : node608;
											assign node608 = (inp[3]) ? node612 : node609;
												assign node609 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node612 = (inp[1]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node615 = (inp[0]) ? 14'b00000000111111 : node616;
												assign node616 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node620 = (inp[3]) ? node678 : node621;
								assign node621 = (inp[0]) ? node649 : node622;
									assign node622 = (inp[1]) ? node636 : node623;
										assign node623 = (inp[4]) ? node631 : node624;
											assign node624 = (inp[5]) ? node628 : node625;
												assign node625 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node628 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node631 = (inp[8]) ? node633 : 14'b00001111111111;
												assign node633 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node636 = (inp[4]) ? node644 : node637;
											assign node637 = (inp[9]) ? node641 : node638;
												assign node638 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node641 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node644 = (inp[13]) ? 14'b00000011111111 : node645;
												assign node645 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node649 = (inp[13]) ? node665 : node650;
										assign node650 = (inp[8]) ? node658 : node651;
											assign node651 = (inp[4]) ? node655 : node652;
												assign node652 = (inp[5]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node655 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node658 = (inp[1]) ? node662 : node659;
												assign node659 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node662 = (inp[5]) ? 14'b00000011111111 : 14'b00000001111111;
										assign node665 = (inp[4]) ? node673 : node666;
											assign node666 = (inp[9]) ? node670 : node667;
												assign node667 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node670 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node673 = (inp[5]) ? node675 : 14'b00000001111111;
												assign node675 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node678 = (inp[9]) ? node710 : node679;
									assign node679 = (inp[1]) ? node695 : node680;
										assign node680 = (inp[8]) ? node688 : node681;
											assign node681 = (inp[4]) ? node685 : node682;
												assign node682 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node685 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node688 = (inp[5]) ? node692 : node689;
												assign node689 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node692 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node695 = (inp[13]) ? node703 : node696;
											assign node696 = (inp[8]) ? node700 : node697;
												assign node697 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node700 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node703 = (inp[4]) ? node707 : node704;
												assign node704 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node707 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node710 = (inp[8]) ? node726 : node711;
										assign node711 = (inp[4]) ? node719 : node712;
											assign node712 = (inp[0]) ? node716 : node713;
												assign node713 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node716 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node719 = (inp[1]) ? node723 : node720;
												assign node720 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node723 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node726 = (inp[0]) ? node734 : node727;
											assign node727 = (inp[4]) ? node731 : node728;
												assign node728 = (inp[13]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node731 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node734 = (inp[13]) ? node738 : node735;
												assign node735 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node738 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node741 = (inp[1]) ? node857 : node742;
							assign node742 = (inp[3]) ? node796 : node743;
								assign node743 = (inp[0]) ? node771 : node744;
									assign node744 = (inp[5]) ? node758 : node745;
										assign node745 = (inp[9]) ? node751 : node746;
											assign node746 = (inp[4]) ? 14'b00001111111111 : node747;
												assign node747 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node751 = (inp[4]) ? node755 : node752;
												assign node752 = (inp[13]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node755 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node758 = (inp[11]) ? node764 : node759;
											assign node759 = (inp[4]) ? node761 : 14'b00000111111111;
												assign node761 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node764 = (inp[9]) ? node768 : node765;
												assign node765 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node768 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node771 = (inp[4]) ? node787 : node772;
										assign node772 = (inp[11]) ? node780 : node773;
											assign node773 = (inp[13]) ? node777 : node774;
												assign node774 = (inp[5]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node777 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node780 = (inp[8]) ? node784 : node781;
												assign node781 = (inp[5]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node784 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node787 = (inp[8]) ? 14'b00000001111111 : node788;
											assign node788 = (inp[5]) ? node792 : node789;
												assign node789 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node792 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node796 = (inp[13]) ? node828 : node797;
									assign node797 = (inp[8]) ? node813 : node798;
										assign node798 = (inp[11]) ? node806 : node799;
											assign node799 = (inp[9]) ? node803 : node800;
												assign node800 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node803 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node806 = (inp[4]) ? node810 : node807;
												assign node807 = (inp[5]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node810 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node813 = (inp[5]) ? node821 : node814;
											assign node814 = (inp[0]) ? node818 : node815;
												assign node815 = (inp[9]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node818 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node821 = (inp[4]) ? node825 : node822;
												assign node822 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node825 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node828 = (inp[9]) ? node842 : node829;
										assign node829 = (inp[4]) ? node837 : node830;
											assign node830 = (inp[8]) ? node834 : node831;
												assign node831 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node834 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node837 = (inp[11]) ? 14'b00000001111111 : node838;
												assign node838 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node842 = (inp[11]) ? node850 : node843;
											assign node843 = (inp[4]) ? node847 : node844;
												assign node844 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node847 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node850 = (inp[8]) ? node854 : node851;
												assign node851 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node854 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node857 = (inp[0]) ? node919 : node858;
								assign node858 = (inp[5]) ? node890 : node859;
									assign node859 = (inp[8]) ? node875 : node860;
										assign node860 = (inp[9]) ? node868 : node861;
											assign node861 = (inp[3]) ? node865 : node862;
												assign node862 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node865 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node868 = (inp[13]) ? node872 : node869;
												assign node869 = (inp[3]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node872 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node875 = (inp[4]) ? node883 : node876;
											assign node876 = (inp[3]) ? node880 : node877;
												assign node877 = (inp[13]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node880 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node883 = (inp[11]) ? node887 : node884;
												assign node884 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node887 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node890 = (inp[9]) ? node906 : node891;
										assign node891 = (inp[11]) ? node899 : node892;
											assign node892 = (inp[3]) ? node896 : node893;
												assign node893 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node896 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node899 = (inp[4]) ? node903 : node900;
												assign node900 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node903 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node906 = (inp[8]) ? node912 : node907;
											assign node907 = (inp[4]) ? node909 : 14'b00000001111111;
												assign node909 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node912 = (inp[3]) ? node916 : node913;
												assign node913 = (inp[11]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node916 = (inp[4]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node919 = (inp[8]) ? node951 : node920;
									assign node920 = (inp[9]) ? node936 : node921;
										assign node921 = (inp[13]) ? node929 : node922;
											assign node922 = (inp[5]) ? node926 : node923;
												assign node923 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node926 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node929 = (inp[4]) ? node933 : node930;
												assign node930 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node933 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node936 = (inp[11]) ? node944 : node937;
											assign node937 = (inp[13]) ? node941 : node938;
												assign node938 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node941 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node944 = (inp[4]) ? node948 : node945;
												assign node945 = (inp[5]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node948 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node951 = (inp[9]) ? node967 : node952;
										assign node952 = (inp[5]) ? node960 : node953;
											assign node953 = (inp[3]) ? node957 : node954;
												assign node954 = (inp[13]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node957 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node960 = (inp[11]) ? node964 : node961;
												assign node961 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node964 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node967 = (inp[4]) ? node973 : node968;
											assign node968 = (inp[11]) ? 14'b00000000011111 : node969;
												assign node969 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node973 = (inp[13]) ? node975 : 14'b00000000011111;
												assign node975 = (inp[5]) ? 14'b00000000000111 : 14'b00000000011111;
				assign node978 = (inp[8]) ? node1454 : node979;
					assign node979 = (inp[0]) ? node1219 : node980;
						assign node980 = (inp[1]) ? node1100 : node981;
							assign node981 = (inp[4]) ? node1041 : node982;
								assign node982 = (inp[13]) ? node1012 : node983;
									assign node983 = (inp[11]) ? node997 : node984;
										assign node984 = (inp[3]) ? node990 : node985;
											assign node985 = (inp[5]) ? 14'b00011111111111 : node986;
												assign node986 = (inp[2]) ? 14'b00011111111111 : 14'b00111111111111;
											assign node990 = (inp[9]) ? node994 : node991;
												assign node991 = (inp[5]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node994 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node997 = (inp[5]) ? node1005 : node998;
											assign node998 = (inp[2]) ? node1002 : node999;
												assign node999 = (inp[10]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node1002 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1005 = (inp[3]) ? node1009 : node1006;
												assign node1006 = (inp[2]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node1009 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node1012 = (inp[3]) ? node1026 : node1013;
										assign node1013 = (inp[11]) ? node1019 : node1014;
											assign node1014 = (inp[9]) ? 14'b00001111111111 : node1015;
												assign node1015 = (inp[5]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node1019 = (inp[2]) ? node1023 : node1020;
												assign node1020 = (inp[10]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node1023 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1026 = (inp[2]) ? node1034 : node1027;
											assign node1027 = (inp[10]) ? node1031 : node1028;
												assign node1028 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1031 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1034 = (inp[11]) ? node1038 : node1035;
												assign node1035 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1038 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1041 = (inp[3]) ? node1069 : node1042;
									assign node1042 = (inp[2]) ? node1056 : node1043;
										assign node1043 = (inp[9]) ? node1049 : node1044;
											assign node1044 = (inp[5]) ? 14'b00001111111111 : node1045;
												assign node1045 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node1049 = (inp[13]) ? node1053 : node1050;
												assign node1050 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1053 = (inp[5]) ? 14'b00000001111111 : 14'b00000111111111;
										assign node1056 = (inp[5]) ? node1062 : node1057;
											assign node1057 = (inp[9]) ? node1059 : 14'b00000111111111;
												assign node1059 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1062 = (inp[11]) ? node1066 : node1063;
												assign node1063 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1066 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1069 = (inp[9]) ? node1085 : node1070;
										assign node1070 = (inp[11]) ? node1078 : node1071;
											assign node1071 = (inp[2]) ? node1075 : node1072;
												assign node1072 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1075 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1078 = (inp[10]) ? node1082 : node1079;
												assign node1079 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1082 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1085 = (inp[5]) ? node1093 : node1086;
											assign node1086 = (inp[2]) ? node1090 : node1087;
												assign node1087 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1090 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1093 = (inp[10]) ? node1097 : node1094;
												assign node1094 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1097 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node1100 = (inp[11]) ? node1158 : node1101;
								assign node1101 = (inp[9]) ? node1131 : node1102;
									assign node1102 = (inp[4]) ? node1116 : node1103;
										assign node1103 = (inp[2]) ? node1111 : node1104;
											assign node1104 = (inp[13]) ? node1108 : node1105;
												assign node1105 = (inp[3]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node1108 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1111 = (inp[10]) ? 14'b00000011111111 : node1112;
												assign node1112 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node1116 = (inp[13]) ? node1124 : node1117;
											assign node1117 = (inp[10]) ? node1121 : node1118;
												assign node1118 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1121 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1124 = (inp[3]) ? node1128 : node1125;
												assign node1125 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1128 = (inp[2]) ? 14'b00000000111111 : 14'b00000011111111;
									assign node1131 = (inp[10]) ? node1143 : node1132;
										assign node1132 = (inp[2]) ? node1138 : node1133;
											assign node1133 = (inp[13]) ? node1135 : 14'b00000111111111;
												assign node1135 = (inp[3]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node1138 = (inp[4]) ? 14'b00000011111111 : node1139;
												assign node1139 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1143 = (inp[5]) ? node1151 : node1144;
											assign node1144 = (inp[4]) ? node1148 : node1145;
												assign node1145 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1148 = (inp[2]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node1151 = (inp[3]) ? node1155 : node1152;
												assign node1152 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1155 = (inp[2]) ? 14'b00000000011111 : 14'b00000001111111;
								assign node1158 = (inp[2]) ? node1190 : node1159;
									assign node1159 = (inp[4]) ? node1175 : node1160;
										assign node1160 = (inp[9]) ? node1168 : node1161;
											assign node1161 = (inp[10]) ? node1165 : node1162;
												assign node1162 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1165 = (inp[13]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node1168 = (inp[5]) ? node1172 : node1169;
												assign node1169 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1172 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1175 = (inp[3]) ? node1183 : node1176;
											assign node1176 = (inp[10]) ? node1180 : node1177;
												assign node1177 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1180 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1183 = (inp[13]) ? node1187 : node1184;
												assign node1184 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1187 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1190 = (inp[9]) ? node1206 : node1191;
										assign node1191 = (inp[4]) ? node1199 : node1192;
											assign node1192 = (inp[3]) ? node1196 : node1193;
												assign node1193 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1196 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1199 = (inp[10]) ? node1203 : node1200;
												assign node1200 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1203 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1206 = (inp[5]) ? node1214 : node1207;
											assign node1207 = (inp[13]) ? node1211 : node1208;
												assign node1208 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1211 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1214 = (inp[13]) ? 14'b00000000011111 : node1215;
												assign node1215 = (inp[4]) ? 14'b00000000011111 : 14'b00000001111111;
						assign node1219 = (inp[10]) ? node1341 : node1220;
							assign node1220 = (inp[5]) ? node1282 : node1221;
								assign node1221 = (inp[13]) ? node1251 : node1222;
									assign node1222 = (inp[4]) ? node1236 : node1223;
										assign node1223 = (inp[3]) ? node1231 : node1224;
											assign node1224 = (inp[9]) ? node1228 : node1225;
												assign node1225 = (inp[2]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node1228 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1231 = (inp[11]) ? 14'b00000111111111 : node1232;
												assign node1232 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node1236 = (inp[9]) ? node1244 : node1237;
											assign node1237 = (inp[3]) ? node1241 : node1238;
												assign node1238 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1241 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1244 = (inp[2]) ? node1248 : node1245;
												assign node1245 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1248 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1251 = (inp[1]) ? node1267 : node1252;
										assign node1252 = (inp[9]) ? node1260 : node1253;
											assign node1253 = (inp[3]) ? node1257 : node1254;
												assign node1254 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1257 = (inp[2]) ? 14'b00000011111111 : 14'b00000011111111;
											assign node1260 = (inp[2]) ? node1264 : node1261;
												assign node1261 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1264 = (inp[3]) ? 14'b00000000111111 : 14'b00000011111111;
										assign node1267 = (inp[4]) ? node1275 : node1268;
											assign node1268 = (inp[9]) ? node1272 : node1269;
												assign node1269 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1272 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1275 = (inp[11]) ? node1279 : node1276;
												assign node1276 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1279 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1282 = (inp[13]) ? node1312 : node1283;
									assign node1283 = (inp[1]) ? node1297 : node1284;
										assign node1284 = (inp[2]) ? node1292 : node1285;
											assign node1285 = (inp[11]) ? node1289 : node1286;
												assign node1286 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1289 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1292 = (inp[4]) ? 14'b00000011111111 : node1293;
												assign node1293 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1297 = (inp[4]) ? node1305 : node1298;
											assign node1298 = (inp[3]) ? node1302 : node1299;
												assign node1299 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1302 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1305 = (inp[9]) ? node1309 : node1306;
												assign node1306 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1309 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1312 = (inp[3]) ? node1326 : node1313;
										assign node1313 = (inp[2]) ? node1321 : node1314;
											assign node1314 = (inp[4]) ? node1318 : node1315;
												assign node1315 = (inp[9]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node1318 = (inp[9]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node1321 = (inp[4]) ? node1323 : 14'b00000001111111;
												assign node1323 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1326 = (inp[2]) ? node1334 : node1327;
											assign node1327 = (inp[4]) ? node1331 : node1328;
												assign node1328 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1331 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1334 = (inp[1]) ? node1338 : node1335;
												assign node1335 = (inp[9]) ? 14'b00000000011111 : 14'b00000001111111;
												assign node1338 = (inp[4]) ? 14'b00000000011111 : 14'b00000000011111;
							assign node1341 = (inp[3]) ? node1401 : node1342;
								assign node1342 = (inp[5]) ? node1370 : node1343;
									assign node1343 = (inp[11]) ? node1357 : node1344;
										assign node1344 = (inp[13]) ? node1350 : node1345;
											assign node1345 = (inp[9]) ? 14'b00000111111111 : node1346;
												assign node1346 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1350 = (inp[1]) ? node1354 : node1351;
												assign node1351 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1354 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1357 = (inp[9]) ? node1363 : node1358;
											assign node1358 = (inp[4]) ? node1360 : 14'b00000011111111;
												assign node1360 = (inp[1]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node1363 = (inp[2]) ? node1367 : node1364;
												assign node1364 = (inp[1]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node1367 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1370 = (inp[1]) ? node1386 : node1371;
										assign node1371 = (inp[13]) ? node1379 : node1372;
											assign node1372 = (inp[9]) ? node1376 : node1373;
												assign node1373 = (inp[11]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node1376 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1379 = (inp[4]) ? node1383 : node1380;
												assign node1380 = (inp[11]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node1383 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1386 = (inp[4]) ? node1394 : node1387;
											assign node1387 = (inp[2]) ? node1391 : node1388;
												assign node1388 = (inp[11]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node1391 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1394 = (inp[9]) ? node1398 : node1395;
												assign node1395 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1398 = (inp[13]) ? 14'b00000000001111 : 14'b00000000111111;
								assign node1401 = (inp[1]) ? node1425 : node1402;
									assign node1402 = (inp[2]) ? node1416 : node1403;
										assign node1403 = (inp[9]) ? node1409 : node1404;
											assign node1404 = (inp[4]) ? node1406 : 14'b00000011111111;
												assign node1406 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1409 = (inp[5]) ? node1413 : node1410;
												assign node1410 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1413 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1416 = (inp[11]) ? node1422 : node1417;
											assign node1417 = (inp[9]) ? 14'b00000000111111 : node1418;
												assign node1418 = (inp[4]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node1422 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node1425 = (inp[13]) ? node1439 : node1426;
										assign node1426 = (inp[9]) ? node1432 : node1427;
											assign node1427 = (inp[5]) ? node1429 : 14'b00000011111111;
												assign node1429 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1432 = (inp[4]) ? node1436 : node1433;
												assign node1433 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1436 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1439 = (inp[11]) ? node1447 : node1440;
											assign node1440 = (inp[9]) ? node1444 : node1441;
												assign node1441 = (inp[5]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node1444 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node1447 = (inp[4]) ? node1451 : node1448;
												assign node1448 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node1451 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
					assign node1454 = (inp[9]) ? node1698 : node1455;
						assign node1455 = (inp[1]) ? node1577 : node1456;
							assign node1456 = (inp[0]) ? node1518 : node1457;
								assign node1457 = (inp[5]) ? node1487 : node1458;
									assign node1458 = (inp[4]) ? node1472 : node1459;
										assign node1459 = (inp[13]) ? node1467 : node1460;
											assign node1460 = (inp[2]) ? node1464 : node1461;
												assign node1461 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node1464 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1467 = (inp[11]) ? 14'b00000111111111 : node1468;
												assign node1468 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node1472 = (inp[11]) ? node1480 : node1473;
											assign node1473 = (inp[13]) ? node1477 : node1474;
												assign node1474 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1477 = (inp[2]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node1480 = (inp[13]) ? node1484 : node1481;
												assign node1481 = (inp[3]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node1484 = (inp[10]) ? 14'b00000000111111 : 14'b00000011111111;
									assign node1487 = (inp[11]) ? node1503 : node1488;
										assign node1488 = (inp[13]) ? node1496 : node1489;
											assign node1489 = (inp[10]) ? node1493 : node1490;
												assign node1490 = (inp[4]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node1493 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1496 = (inp[10]) ? node1500 : node1497;
												assign node1497 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1500 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1503 = (inp[3]) ? node1511 : node1504;
											assign node1504 = (inp[2]) ? node1508 : node1505;
												assign node1505 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1508 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1511 = (inp[4]) ? node1515 : node1512;
												assign node1512 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1515 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1518 = (inp[11]) ? node1548 : node1519;
									assign node1519 = (inp[5]) ? node1533 : node1520;
										assign node1520 = (inp[13]) ? node1526 : node1521;
											assign node1521 = (inp[2]) ? 14'b00000111111111 : node1522;
												assign node1522 = (inp[3]) ? 14'b00000011111111 : 14'b00001111111111;
											assign node1526 = (inp[10]) ? node1530 : node1527;
												assign node1527 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1530 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1533 = (inp[3]) ? node1541 : node1534;
											assign node1534 = (inp[13]) ? node1538 : node1535;
												assign node1535 = (inp[10]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node1538 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1541 = (inp[10]) ? node1545 : node1542;
												assign node1542 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1545 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1548 = (inp[13]) ? node1564 : node1549;
										assign node1549 = (inp[4]) ? node1557 : node1550;
											assign node1550 = (inp[3]) ? node1554 : node1551;
												assign node1551 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1554 = (inp[5]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node1557 = (inp[2]) ? node1561 : node1558;
												assign node1558 = (inp[5]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node1561 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1564 = (inp[10]) ? node1570 : node1565;
											assign node1565 = (inp[2]) ? node1567 : 14'b00000001111111;
												assign node1567 = (inp[5]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node1570 = (inp[3]) ? node1574 : node1571;
												assign node1571 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1574 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node1577 = (inp[3]) ? node1637 : node1578;
								assign node1578 = (inp[13]) ? node1606 : node1579;
									assign node1579 = (inp[2]) ? node1595 : node1580;
										assign node1580 = (inp[0]) ? node1588 : node1581;
											assign node1581 = (inp[11]) ? node1585 : node1582;
												assign node1582 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1585 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1588 = (inp[5]) ? node1592 : node1589;
												assign node1589 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1592 = (inp[11]) ? 14'b00000001111111 : 14'b00000001111111;
										assign node1595 = (inp[10]) ? node1599 : node1596;
											assign node1596 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1599 = (inp[5]) ? node1603 : node1600;
												assign node1600 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1603 = (inp[0]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node1606 = (inp[5]) ? node1622 : node1607;
										assign node1607 = (inp[10]) ? node1615 : node1608;
											assign node1608 = (inp[0]) ? node1612 : node1609;
												assign node1609 = (inp[2]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node1612 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1615 = (inp[4]) ? node1619 : node1616;
												assign node1616 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1619 = (inp[11]) ? 14'b00000000111111 : 14'b00000011111111;
										assign node1622 = (inp[0]) ? node1630 : node1623;
											assign node1623 = (inp[4]) ? node1627 : node1624;
												assign node1624 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1627 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1630 = (inp[11]) ? node1634 : node1631;
												assign node1631 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1634 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node1637 = (inp[5]) ? node1667 : node1638;
									assign node1638 = (inp[10]) ? node1654 : node1639;
										assign node1639 = (inp[0]) ? node1647 : node1640;
											assign node1640 = (inp[4]) ? node1644 : node1641;
												assign node1641 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1644 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1647 = (inp[11]) ? node1651 : node1648;
												assign node1648 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1651 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1654 = (inp[4]) ? node1660 : node1655;
											assign node1655 = (inp[11]) ? node1657 : 14'b00000011111111;
												assign node1657 = (inp[0]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node1660 = (inp[2]) ? node1664 : node1661;
												assign node1661 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1664 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node1667 = (inp[13]) ? node1683 : node1668;
										assign node1668 = (inp[2]) ? node1676 : node1669;
											assign node1669 = (inp[11]) ? node1673 : node1670;
												assign node1670 = (inp[10]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node1673 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1676 = (inp[10]) ? node1680 : node1677;
												assign node1677 = (inp[11]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node1680 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1683 = (inp[0]) ? node1691 : node1684;
											assign node1684 = (inp[4]) ? node1688 : node1685;
												assign node1685 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1688 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node1691 = (inp[2]) ? node1695 : node1692;
												assign node1692 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node1695 = (inp[4]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node1698 = (inp[11]) ? node1818 : node1699;
							assign node1699 = (inp[4]) ? node1761 : node1700;
								assign node1700 = (inp[1]) ? node1730 : node1701;
									assign node1701 = (inp[10]) ? node1715 : node1702;
										assign node1702 = (inp[3]) ? node1708 : node1703;
											assign node1703 = (inp[13]) ? 14'b00000111111111 : node1704;
												assign node1704 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1708 = (inp[13]) ? node1712 : node1709;
												assign node1709 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1712 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node1715 = (inp[2]) ? node1723 : node1716;
											assign node1716 = (inp[3]) ? node1720 : node1717;
												assign node1717 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1720 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1723 = (inp[13]) ? node1727 : node1724;
												assign node1724 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1727 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node1730 = (inp[3]) ? node1746 : node1731;
										assign node1731 = (inp[10]) ? node1739 : node1732;
											assign node1732 = (inp[2]) ? node1736 : node1733;
												assign node1733 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1736 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1739 = (inp[13]) ? node1743 : node1740;
												assign node1740 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1743 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1746 = (inp[10]) ? node1754 : node1747;
											assign node1747 = (inp[5]) ? node1751 : node1748;
												assign node1748 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1751 = (inp[13]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node1754 = (inp[0]) ? node1758 : node1755;
												assign node1755 = (inp[2]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node1758 = (inp[2]) ? 14'b00000000001111 : 14'b00000000111111;
								assign node1761 = (inp[3]) ? node1789 : node1762;
									assign node1762 = (inp[13]) ? node1778 : node1763;
										assign node1763 = (inp[10]) ? node1771 : node1764;
											assign node1764 = (inp[0]) ? node1768 : node1765;
												assign node1765 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1768 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1771 = (inp[2]) ? node1775 : node1772;
												assign node1772 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1775 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1778 = (inp[1]) ? node1784 : node1779;
											assign node1779 = (inp[2]) ? node1781 : 14'b00000001111111;
												assign node1781 = (inp[10]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node1784 = (inp[0]) ? 14'b00000000111111 : node1785;
												assign node1785 = (inp[5]) ? 14'b00000000111111 : 14'b00000000111111;
									assign node1789 = (inp[2]) ? node1805 : node1790;
										assign node1790 = (inp[0]) ? node1798 : node1791;
											assign node1791 = (inp[10]) ? node1795 : node1792;
												assign node1792 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1795 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1798 = (inp[1]) ? node1802 : node1799;
												assign node1799 = (inp[13]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node1802 = (inp[5]) ? 14'b00000000001111 : 14'b00000000111111;
										assign node1805 = (inp[10]) ? node1813 : node1806;
											assign node1806 = (inp[1]) ? node1810 : node1807;
												assign node1807 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1810 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node1813 = (inp[13]) ? 14'b00000000011111 : node1814;
												assign node1814 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node1818 = (inp[13]) ? node1880 : node1819;
								assign node1819 = (inp[2]) ? node1851 : node1820;
									assign node1820 = (inp[4]) ? node1836 : node1821;
										assign node1821 = (inp[5]) ? node1829 : node1822;
											assign node1822 = (inp[3]) ? node1826 : node1823;
												assign node1823 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node1826 = (inp[0]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node1829 = (inp[0]) ? node1833 : node1830;
												assign node1830 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1833 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1836 = (inp[1]) ? node1844 : node1837;
											assign node1837 = (inp[5]) ? node1841 : node1838;
												assign node1838 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1841 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1844 = (inp[10]) ? node1848 : node1845;
												assign node1845 = (inp[3]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node1848 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node1851 = (inp[10]) ? node1865 : node1852;
										assign node1852 = (inp[4]) ? node1858 : node1853;
											assign node1853 = (inp[1]) ? 14'b00000000111111 : node1854;
												assign node1854 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node1858 = (inp[5]) ? node1862 : node1859;
												assign node1859 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1862 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node1865 = (inp[5]) ? node1873 : node1866;
											assign node1866 = (inp[4]) ? node1870 : node1867;
												assign node1867 = (inp[3]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node1870 = (inp[3]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node1873 = (inp[4]) ? node1877 : node1874;
												assign node1874 = (inp[1]) ? 14'b00000000001111 : 14'b00000000111111;
												assign node1877 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node1880 = (inp[5]) ? node1910 : node1881;
									assign node1881 = (inp[2]) ? node1895 : node1882;
										assign node1882 = (inp[0]) ? node1890 : node1883;
											assign node1883 = (inp[10]) ? node1887 : node1884;
												assign node1884 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node1887 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node1890 = (inp[4]) ? 14'b00000000111111 : node1891;
												assign node1891 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1895 = (inp[10]) ? node1903 : node1896;
											assign node1896 = (inp[1]) ? node1900 : node1897;
												assign node1897 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1900 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node1903 = (inp[3]) ? node1907 : node1904;
												assign node1904 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node1907 = (inp[1]) ? 14'b00000000001111 : 14'b00000000001111;
									assign node1910 = (inp[0]) ? node1926 : node1911;
										assign node1911 = (inp[3]) ? node1919 : node1912;
											assign node1912 = (inp[1]) ? node1916 : node1913;
												assign node1913 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node1916 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node1919 = (inp[10]) ? node1923 : node1920;
												assign node1920 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node1923 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node1926 = (inp[1]) ? node1934 : node1927;
											assign node1927 = (inp[3]) ? node1931 : node1928;
												assign node1928 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node1931 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node1934 = (inp[4]) ? node1938 : node1935;
												assign node1935 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node1938 = (inp[10]) ? 14'b00000000000011 : 14'b00000000001111;
			assign node1941 = (inp[3]) ? node2915 : node1942;
				assign node1942 = (inp[4]) ? node2430 : node1943;
					assign node1943 = (inp[2]) ? node2191 : node1944;
						assign node1944 = (inp[8]) ? node2068 : node1945;
							assign node1945 = (inp[9]) ? node2005 : node1946;
								assign node1946 = (inp[11]) ? node1976 : node1947;
									assign node1947 = (inp[1]) ? node1961 : node1948;
										assign node1948 = (inp[13]) ? node1956 : node1949;
											assign node1949 = (inp[5]) ? node1953 : node1950;
												assign node1950 = (inp[0]) ? 14'b00001111111111 : 14'b00111111111111;
												assign node1953 = (inp[7]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node1956 = (inp[0]) ? 14'b00001111111111 : node1957;
												assign node1957 = (inp[10]) ? 14'b00001111111111 : 14'b00111111111111;
										assign node1961 = (inp[0]) ? node1969 : node1962;
											assign node1962 = (inp[13]) ? node1966 : node1963;
												assign node1963 = (inp[5]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node1966 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1969 = (inp[7]) ? node1973 : node1970;
												assign node1970 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1973 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1976 = (inp[7]) ? node1992 : node1977;
										assign node1977 = (inp[0]) ? node1985 : node1978;
											assign node1978 = (inp[10]) ? node1982 : node1979;
												assign node1979 = (inp[1]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node1982 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node1985 = (inp[5]) ? node1989 : node1986;
												assign node1986 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node1989 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node1992 = (inp[10]) ? node1998 : node1993;
											assign node1993 = (inp[5]) ? node1995 : 14'b00000111111111;
												assign node1995 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node1998 = (inp[0]) ? node2002 : node1999;
												assign node1999 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2002 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node2005 = (inp[10]) ? node2037 : node2006;
									assign node2006 = (inp[13]) ? node2022 : node2007;
										assign node2007 = (inp[7]) ? node2015 : node2008;
											assign node2008 = (inp[0]) ? node2012 : node2009;
												assign node2009 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node2012 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node2015 = (inp[5]) ? node2019 : node2016;
												assign node2016 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2019 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2022 = (inp[7]) ? node2030 : node2023;
											assign node2023 = (inp[1]) ? node2027 : node2024;
												assign node2024 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2027 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2030 = (inp[0]) ? node2034 : node2031;
												assign node2031 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2034 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2037 = (inp[1]) ? node2053 : node2038;
										assign node2038 = (inp[5]) ? node2046 : node2039;
											assign node2039 = (inp[13]) ? node2043 : node2040;
												assign node2040 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2043 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2046 = (inp[13]) ? node2050 : node2047;
												assign node2047 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2050 = (inp[11]) ? 14'b00000000111111 : 14'b00000011111111;
										assign node2053 = (inp[0]) ? node2061 : node2054;
											assign node2054 = (inp[13]) ? node2058 : node2055;
												assign node2055 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2058 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2061 = (inp[7]) ? node2065 : node2062;
												assign node2062 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2065 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node2068 = (inp[11]) ? node2132 : node2069;
								assign node2069 = (inp[0]) ? node2101 : node2070;
									assign node2070 = (inp[7]) ? node2086 : node2071;
										assign node2071 = (inp[13]) ? node2079 : node2072;
											assign node2072 = (inp[10]) ? node2076 : node2073;
												assign node2073 = (inp[5]) ? 14'b00001111111111 : 14'b00001111111111;
												assign node2076 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node2079 = (inp[9]) ? node2083 : node2080;
												assign node2080 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2083 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2086 = (inp[9]) ? node2094 : node2087;
											assign node2087 = (inp[1]) ? node2091 : node2088;
												assign node2088 = (inp[10]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node2091 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2094 = (inp[10]) ? node2098 : node2095;
												assign node2095 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2098 = (inp[13]) ? 14'b00000000111111 : 14'b00000011111111;
									assign node2101 = (inp[13]) ? node2117 : node2102;
										assign node2102 = (inp[10]) ? node2110 : node2103;
											assign node2103 = (inp[1]) ? node2107 : node2104;
												assign node2104 = (inp[7]) ? 14'b00000111111111 : 14'b00011111111111;
												assign node2107 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2110 = (inp[1]) ? node2114 : node2111;
												assign node2111 = (inp[5]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node2114 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2117 = (inp[7]) ? node2125 : node2118;
											assign node2118 = (inp[9]) ? node2122 : node2119;
												assign node2119 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2122 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2125 = (inp[10]) ? node2129 : node2126;
												assign node2126 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2129 = (inp[9]) ? 14'b00000000011111 : 14'b00000001111111;
								assign node2132 = (inp[5]) ? node2162 : node2133;
									assign node2133 = (inp[9]) ? node2149 : node2134;
										assign node2134 = (inp[10]) ? node2142 : node2135;
											assign node2135 = (inp[7]) ? node2139 : node2136;
												assign node2136 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2139 = (inp[1]) ? 14'b00000111111111 : 14'b00000011111111;
											assign node2142 = (inp[0]) ? node2146 : node2143;
												assign node2143 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2146 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2149 = (inp[1]) ? node2157 : node2150;
											assign node2150 = (inp[7]) ? node2154 : node2151;
												assign node2151 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2154 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2157 = (inp[10]) ? 14'b00000000111111 : node2158;
												assign node2158 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2162 = (inp[10]) ? node2176 : node2163;
										assign node2163 = (inp[9]) ? node2171 : node2164;
											assign node2164 = (inp[1]) ? node2168 : node2165;
												assign node2165 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2168 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2171 = (inp[13]) ? 14'b00000001111111 : node2172;
												assign node2172 = (inp[0]) ? 14'b00000001111111 : 14'b00000001111111;
										assign node2176 = (inp[7]) ? node2184 : node2177;
											assign node2177 = (inp[13]) ? node2181 : node2178;
												assign node2178 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2181 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2184 = (inp[1]) ? node2188 : node2185;
												assign node2185 = (inp[0]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node2188 = (inp[13]) ? 14'b00000000011111 : 14'b00000000011111;
						assign node2191 = (inp[5]) ? node2309 : node2192;
							assign node2192 = (inp[10]) ? node2254 : node2193;
								assign node2193 = (inp[11]) ? node2225 : node2194;
									assign node2194 = (inp[13]) ? node2210 : node2195;
										assign node2195 = (inp[1]) ? node2203 : node2196;
											assign node2196 = (inp[8]) ? node2200 : node2197;
												assign node2197 = (inp[0]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node2200 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node2203 = (inp[8]) ? node2207 : node2204;
												assign node2204 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2207 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2210 = (inp[9]) ? node2218 : node2211;
											assign node2211 = (inp[8]) ? node2215 : node2212;
												assign node2212 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2215 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2218 = (inp[7]) ? node2222 : node2219;
												assign node2219 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2222 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2225 = (inp[0]) ? node2239 : node2226;
										assign node2226 = (inp[9]) ? node2232 : node2227;
											assign node2227 = (inp[1]) ? 14'b00000111111111 : node2228;
												assign node2228 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node2232 = (inp[8]) ? node2236 : node2233;
												assign node2233 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2236 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2239 = (inp[8]) ? node2247 : node2240;
											assign node2240 = (inp[1]) ? node2244 : node2241;
												assign node2241 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2244 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2247 = (inp[1]) ? node2251 : node2248;
												assign node2248 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2251 = (inp[13]) ? 14'b00000000111111 : 14'b00000000111111;
								assign node2254 = (inp[0]) ? node2286 : node2255;
									assign node2255 = (inp[8]) ? node2271 : node2256;
										assign node2256 = (inp[1]) ? node2264 : node2257;
											assign node2257 = (inp[9]) ? node2261 : node2258;
												assign node2258 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2261 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2264 = (inp[9]) ? node2268 : node2265;
												assign node2265 = (inp[7]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node2268 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2271 = (inp[7]) ? node2279 : node2272;
											assign node2272 = (inp[13]) ? node2276 : node2273;
												assign node2273 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2276 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2279 = (inp[1]) ? node2283 : node2280;
												assign node2280 = (inp[11]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node2283 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2286 = (inp[7]) ? node2296 : node2287;
										assign node2287 = (inp[9]) ? 14'b00000001111111 : node2288;
											assign node2288 = (inp[11]) ? node2292 : node2289;
												assign node2289 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2292 = (inp[13]) ? 14'b00000001111111 : 14'b00000001111111;
										assign node2296 = (inp[8]) ? node2302 : node2297;
											assign node2297 = (inp[11]) ? 14'b00000000011111 : node2298;
												assign node2298 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2302 = (inp[9]) ? node2306 : node2303;
												assign node2303 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2306 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node2309 = (inp[13]) ? node2371 : node2310;
								assign node2310 = (inp[9]) ? node2340 : node2311;
									assign node2311 = (inp[8]) ? node2327 : node2312;
										assign node2312 = (inp[11]) ? node2320 : node2313;
											assign node2313 = (inp[7]) ? node2317 : node2314;
												assign node2314 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2317 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2320 = (inp[0]) ? node2324 : node2321;
												assign node2321 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2324 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2327 = (inp[10]) ? node2333 : node2328;
											assign node2328 = (inp[1]) ? node2330 : 14'b00000011111111;
												assign node2330 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2333 = (inp[7]) ? node2337 : node2334;
												assign node2334 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2337 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2340 = (inp[10]) ? node2356 : node2341;
										assign node2341 = (inp[7]) ? node2349 : node2342;
											assign node2342 = (inp[0]) ? node2346 : node2343;
												assign node2343 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2346 = (inp[8]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node2349 = (inp[1]) ? node2353 : node2350;
												assign node2350 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2353 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2356 = (inp[1]) ? node2364 : node2357;
											assign node2357 = (inp[0]) ? node2361 : node2358;
												assign node2358 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2361 = (inp[7]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node2364 = (inp[8]) ? node2368 : node2365;
												assign node2365 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2368 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node2371 = (inp[11]) ? node2401 : node2372;
									assign node2372 = (inp[10]) ? node2388 : node2373;
										assign node2373 = (inp[8]) ? node2381 : node2374;
											assign node2374 = (inp[9]) ? node2378 : node2375;
												assign node2375 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2378 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2381 = (inp[7]) ? node2385 : node2382;
												assign node2382 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2385 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2388 = (inp[0]) ? node2394 : node2389;
											assign node2389 = (inp[8]) ? node2391 : 14'b00000001111111;
												assign node2391 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2394 = (inp[7]) ? node2398 : node2395;
												assign node2395 = (inp[1]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node2398 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2401 = (inp[9]) ? node2415 : node2402;
										assign node2402 = (inp[0]) ? node2408 : node2403;
											assign node2403 = (inp[10]) ? node2405 : 14'b00000001111111;
												assign node2405 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2408 = (inp[7]) ? node2412 : node2409;
												assign node2409 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2412 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2415 = (inp[0]) ? node2423 : node2416;
											assign node2416 = (inp[8]) ? node2420 : node2417;
												assign node2417 = (inp[10]) ? 14'b00000000011111 : 14'b00000001111111;
												assign node2420 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2423 = (inp[8]) ? node2427 : node2424;
												assign node2424 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node2427 = (inp[1]) ? 14'b00000000001111 : 14'b00000000001111;
					assign node2430 = (inp[1]) ? node2670 : node2431;
						assign node2431 = (inp[0]) ? node2547 : node2432;
							assign node2432 = (inp[13]) ? node2490 : node2433;
								assign node2433 = (inp[8]) ? node2461 : node2434;
									assign node2434 = (inp[2]) ? node2450 : node2435;
										assign node2435 = (inp[7]) ? node2443 : node2436;
											assign node2436 = (inp[11]) ? node2440 : node2437;
												assign node2437 = (inp[5]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node2440 = (inp[9]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node2443 = (inp[10]) ? node2447 : node2444;
												assign node2444 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2447 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2450 = (inp[9]) ? node2456 : node2451;
											assign node2451 = (inp[11]) ? 14'b00000111111111 : node2452;
												assign node2452 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node2456 = (inp[5]) ? 14'b00000011111111 : node2457;
												assign node2457 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node2461 = (inp[2]) ? node2477 : node2462;
										assign node2462 = (inp[7]) ? node2470 : node2463;
											assign node2463 = (inp[11]) ? node2467 : node2464;
												assign node2464 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2467 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2470 = (inp[10]) ? node2474 : node2471;
												assign node2471 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2474 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2477 = (inp[9]) ? node2485 : node2478;
											assign node2478 = (inp[5]) ? node2482 : node2479;
												assign node2479 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2482 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2485 = (inp[10]) ? node2487 : 14'b00000001111111;
												assign node2487 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node2490 = (inp[10]) ? node2516 : node2491;
									assign node2491 = (inp[2]) ? node2507 : node2492;
										assign node2492 = (inp[8]) ? node2500 : node2493;
											assign node2493 = (inp[7]) ? node2497 : node2494;
												assign node2494 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2497 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2500 = (inp[11]) ? node2504 : node2501;
												assign node2501 = (inp[5]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node2504 = (inp[7]) ? 14'b00000000111111 : 14'b00000011111111;
										assign node2507 = (inp[5]) ? node2509 : 14'b00000011111111;
											assign node2509 = (inp[11]) ? node2513 : node2510;
												assign node2510 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2513 = (inp[9]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node2516 = (inp[7]) ? node2532 : node2517;
										assign node2517 = (inp[9]) ? node2525 : node2518;
											assign node2518 = (inp[8]) ? node2522 : node2519;
												assign node2519 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2522 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2525 = (inp[11]) ? node2529 : node2526;
												assign node2526 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2529 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2532 = (inp[8]) ? node2540 : node2533;
											assign node2533 = (inp[11]) ? node2537 : node2534;
												assign node2534 = (inp[5]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node2537 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2540 = (inp[11]) ? node2544 : node2541;
												assign node2541 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2544 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node2547 = (inp[2]) ? node2607 : node2548;
								assign node2548 = (inp[9]) ? node2578 : node2549;
									assign node2549 = (inp[10]) ? node2565 : node2550;
										assign node2550 = (inp[7]) ? node2558 : node2551;
											assign node2551 = (inp[8]) ? node2555 : node2552;
												assign node2552 = (inp[5]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2555 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2558 = (inp[13]) ? node2562 : node2559;
												assign node2559 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2562 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2565 = (inp[5]) ? node2571 : node2566;
											assign node2566 = (inp[7]) ? node2568 : 14'b00000011111111;
												assign node2568 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2571 = (inp[8]) ? node2575 : node2572;
												assign node2572 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2575 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2578 = (inp[7]) ? node2594 : node2579;
										assign node2579 = (inp[10]) ? node2587 : node2580;
											assign node2580 = (inp[11]) ? node2584 : node2581;
												assign node2581 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2584 = (inp[13]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node2587 = (inp[13]) ? node2591 : node2588;
												assign node2588 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2591 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2594 = (inp[5]) ? node2600 : node2595;
											assign node2595 = (inp[8]) ? node2597 : 14'b00000011111111;
												assign node2597 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2600 = (inp[13]) ? node2604 : node2601;
												assign node2601 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2604 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node2607 = (inp[8]) ? node2639 : node2608;
									assign node2608 = (inp[10]) ? node2624 : node2609;
										assign node2609 = (inp[11]) ? node2617 : node2610;
											assign node2610 = (inp[13]) ? node2614 : node2611;
												assign node2611 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2614 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2617 = (inp[9]) ? node2621 : node2618;
												assign node2618 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2621 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2624 = (inp[5]) ? node2632 : node2625;
											assign node2625 = (inp[13]) ? node2629 : node2626;
												assign node2626 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2629 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2632 = (inp[7]) ? node2636 : node2633;
												assign node2633 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2636 = (inp[9]) ? 14'b00000000111111 : 14'b00000000111111;
									assign node2639 = (inp[7]) ? node2655 : node2640;
										assign node2640 = (inp[5]) ? node2648 : node2641;
											assign node2641 = (inp[11]) ? node2645 : node2642;
												assign node2642 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2645 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2648 = (inp[9]) ? node2652 : node2649;
												assign node2649 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2652 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2655 = (inp[10]) ? node2663 : node2656;
											assign node2656 = (inp[13]) ? node2660 : node2657;
												assign node2657 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2660 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2663 = (inp[9]) ? node2667 : node2664;
												assign node2664 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node2667 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node2670 = (inp[11]) ? node2792 : node2671;
							assign node2671 = (inp[10]) ? node2735 : node2672;
								assign node2672 = (inp[7]) ? node2704 : node2673;
									assign node2673 = (inp[0]) ? node2689 : node2674;
										assign node2674 = (inp[5]) ? node2682 : node2675;
											assign node2675 = (inp[8]) ? node2679 : node2676;
												assign node2676 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2679 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2682 = (inp[8]) ? node2686 : node2683;
												assign node2683 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2686 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2689 = (inp[13]) ? node2697 : node2690;
											assign node2690 = (inp[8]) ? node2694 : node2691;
												assign node2691 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2694 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2697 = (inp[5]) ? node2701 : node2698;
												assign node2698 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2701 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2704 = (inp[8]) ? node2720 : node2705;
										assign node2705 = (inp[9]) ? node2713 : node2706;
											assign node2706 = (inp[5]) ? node2710 : node2707;
												assign node2707 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2710 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2713 = (inp[2]) ? node2717 : node2714;
												assign node2714 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2717 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node2720 = (inp[2]) ? node2728 : node2721;
											assign node2721 = (inp[5]) ? node2725 : node2722;
												assign node2722 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2725 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2728 = (inp[0]) ? node2732 : node2729;
												assign node2729 = (inp[9]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node2732 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node2735 = (inp[0]) ? node2761 : node2736;
									assign node2736 = (inp[7]) ? node2748 : node2737;
										assign node2737 = (inp[5]) ? node2743 : node2738;
											assign node2738 = (inp[9]) ? node2740 : 14'b00000111111111;
												assign node2740 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2743 = (inp[9]) ? 14'b00000001111111 : node2744;
												assign node2744 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node2748 = (inp[8]) ? node2756 : node2749;
											assign node2749 = (inp[2]) ? node2753 : node2750;
												assign node2750 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2753 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2756 = (inp[9]) ? 14'b00000000011111 : node2757;
												assign node2757 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node2761 = (inp[5]) ? node2777 : node2762;
										assign node2762 = (inp[2]) ? node2770 : node2763;
											assign node2763 = (inp[8]) ? node2767 : node2764;
												assign node2764 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2767 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2770 = (inp[9]) ? node2774 : node2771;
												assign node2771 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2774 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node2777 = (inp[9]) ? node2785 : node2778;
											assign node2778 = (inp[2]) ? node2782 : node2779;
												assign node2779 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2782 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2785 = (inp[7]) ? node2789 : node2786;
												assign node2786 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node2789 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node2792 = (inp[7]) ? node2854 : node2793;
								assign node2793 = (inp[8]) ? node2825 : node2794;
									assign node2794 = (inp[9]) ? node2810 : node2795;
										assign node2795 = (inp[13]) ? node2803 : node2796;
											assign node2796 = (inp[10]) ? node2800 : node2797;
												assign node2797 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2800 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2803 = (inp[5]) ? node2807 : node2804;
												assign node2804 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2807 = (inp[0]) ? 14'b00000000011111 : 14'b00000001111111;
										assign node2810 = (inp[2]) ? node2818 : node2811;
											assign node2811 = (inp[10]) ? node2815 : node2812;
												assign node2812 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2815 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2818 = (inp[10]) ? node2822 : node2819;
												assign node2819 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2822 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node2825 = (inp[10]) ? node2841 : node2826;
										assign node2826 = (inp[9]) ? node2834 : node2827;
											assign node2827 = (inp[2]) ? node2831 : node2828;
												assign node2828 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2831 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node2834 = (inp[13]) ? node2838 : node2835;
												assign node2835 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2838 = (inp[2]) ? 14'b00000000011111 : 14'b00000000011111;
										assign node2841 = (inp[5]) ? node2849 : node2842;
											assign node2842 = (inp[2]) ? node2846 : node2843;
												assign node2843 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2846 = (inp[13]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node2849 = (inp[13]) ? node2851 : 14'b00000000011111;
												assign node2851 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node2854 = (inp[0]) ? node2886 : node2855;
									assign node2855 = (inp[2]) ? node2871 : node2856;
										assign node2856 = (inp[9]) ? node2864 : node2857;
											assign node2857 = (inp[5]) ? node2861 : node2858;
												assign node2858 = (inp[8]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node2861 = (inp[8]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node2864 = (inp[10]) ? node2868 : node2865;
												assign node2865 = (inp[13]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node2868 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node2871 = (inp[13]) ? node2879 : node2872;
											assign node2872 = (inp[9]) ? node2876 : node2873;
												assign node2873 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node2876 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node2879 = (inp[5]) ? node2883 : node2880;
												assign node2880 = (inp[10]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node2883 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node2886 = (inp[5]) ? node2900 : node2887;
										assign node2887 = (inp[13]) ? node2893 : node2888;
											assign node2888 = (inp[9]) ? node2890 : 14'b00000000111111;
												assign node2890 = (inp[8]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node2893 = (inp[10]) ? node2897 : node2894;
												assign node2894 = (inp[2]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node2897 = (inp[2]) ? 14'b00000000000111 : 14'b00000000011111;
										assign node2900 = (inp[9]) ? node2908 : node2901;
											assign node2901 = (inp[2]) ? node2905 : node2902;
												assign node2902 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node2905 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node2908 = (inp[2]) ? node2912 : node2909;
												assign node2909 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node2912 = (inp[10]) ? 14'b00000000000111 : 14'b00000000001111;
				assign node2915 = (inp[11]) ? node3397 : node2916;
					assign node2916 = (inp[9]) ? node3158 : node2917;
						assign node2917 = (inp[0]) ? node3041 : node2918;
							assign node2918 = (inp[13]) ? node2982 : node2919;
								assign node2919 = (inp[2]) ? node2951 : node2920;
									assign node2920 = (inp[1]) ? node2936 : node2921;
										assign node2921 = (inp[4]) ? node2929 : node2922;
											assign node2922 = (inp[7]) ? node2926 : node2923;
												assign node2923 = (inp[5]) ? 14'b00001111111111 : 14'b00001111111111;
												assign node2926 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node2929 = (inp[10]) ? node2933 : node2930;
												assign node2930 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2933 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2936 = (inp[4]) ? node2944 : node2937;
											assign node2937 = (inp[10]) ? node2941 : node2938;
												assign node2938 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node2941 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2944 = (inp[7]) ? node2948 : node2945;
												assign node2945 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2948 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node2951 = (inp[8]) ? node2967 : node2952;
										assign node2952 = (inp[5]) ? node2960 : node2953;
											assign node2953 = (inp[7]) ? node2957 : node2954;
												assign node2954 = (inp[1]) ? 14'b00001111111111 : 14'b00001111111111;
												assign node2957 = (inp[1]) ? 14'b00000011111111 : 14'b00001111111111;
											assign node2960 = (inp[1]) ? node2964 : node2961;
												assign node2961 = (inp[10]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node2964 = (inp[7]) ? 14'b00000000111111 : 14'b00000011111111;
										assign node2967 = (inp[7]) ? node2975 : node2968;
											assign node2968 = (inp[1]) ? node2972 : node2969;
												assign node2969 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node2972 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node2975 = (inp[10]) ? node2979 : node2976;
												assign node2976 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node2979 = (inp[5]) ? 14'b00000000111111 : 14'b00000000111111;
								assign node2982 = (inp[10]) ? node3012 : node2983;
									assign node2983 = (inp[8]) ? node2997 : node2984;
										assign node2984 = (inp[7]) ? node2992 : node2985;
											assign node2985 = (inp[1]) ? node2989 : node2986;
												assign node2986 = (inp[4]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node2989 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node2992 = (inp[1]) ? node2994 : 14'b00000001111111;
												assign node2994 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node2997 = (inp[5]) ? node3005 : node2998;
											assign node2998 = (inp[2]) ? node3002 : node2999;
												assign node2999 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3002 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3005 = (inp[2]) ? node3009 : node3006;
												assign node3006 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3009 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node3012 = (inp[2]) ? node3026 : node3013;
										assign node3013 = (inp[5]) ? node3019 : node3014;
											assign node3014 = (inp[7]) ? node3016 : 14'b00000011111111;
												assign node3016 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3019 = (inp[1]) ? node3023 : node3020;
												assign node3020 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3023 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3026 = (inp[4]) ? node3034 : node3027;
											assign node3027 = (inp[5]) ? node3031 : node3028;
												assign node3028 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3031 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3034 = (inp[1]) ? node3038 : node3035;
												assign node3035 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3038 = (inp[8]) ? 14'b00000000001111 : 14'b00000000111111;
							assign node3041 = (inp[8]) ? node3099 : node3042;
								assign node3042 = (inp[7]) ? node3068 : node3043;
									assign node3043 = (inp[2]) ? node3055 : node3044;
										assign node3044 = (inp[4]) ? node3050 : node3045;
											assign node3045 = (inp[13]) ? 14'b00000111111111 : node3046;
												assign node3046 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3050 = (inp[13]) ? 14'b00000011111111 : node3051;
												assign node3051 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node3055 = (inp[13]) ? node3063 : node3056;
											assign node3056 = (inp[4]) ? node3060 : node3057;
												assign node3057 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3060 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3063 = (inp[10]) ? 14'b00000000111111 : node3064;
												assign node3064 = (inp[5]) ? 14'b00000001111111 : 14'b00000001111111;
									assign node3068 = (inp[1]) ? node3084 : node3069;
										assign node3069 = (inp[5]) ? node3077 : node3070;
											assign node3070 = (inp[4]) ? node3074 : node3071;
												assign node3071 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3074 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3077 = (inp[10]) ? node3081 : node3078;
												assign node3078 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3081 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3084 = (inp[13]) ? node3092 : node3085;
											assign node3085 = (inp[5]) ? node3089 : node3086;
												assign node3086 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3089 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3092 = (inp[4]) ? node3096 : node3093;
												assign node3093 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3096 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node3099 = (inp[1]) ? node3127 : node3100;
									assign node3100 = (inp[10]) ? node3114 : node3101;
										assign node3101 = (inp[7]) ? node3107 : node3102;
											assign node3102 = (inp[13]) ? 14'b00000001111111 : node3103;
												assign node3103 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3107 = (inp[2]) ? node3111 : node3108;
												assign node3108 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3111 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3114 = (inp[5]) ? node3120 : node3115;
											assign node3115 = (inp[7]) ? 14'b00000001111111 : node3116;
												assign node3116 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3120 = (inp[13]) ? node3124 : node3121;
												assign node3121 = (inp[2]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node3124 = (inp[7]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node3127 = (inp[2]) ? node3143 : node3128;
										assign node3128 = (inp[5]) ? node3136 : node3129;
											assign node3129 = (inp[7]) ? node3133 : node3130;
												assign node3130 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3133 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3136 = (inp[4]) ? node3140 : node3137;
												assign node3137 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3140 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3143 = (inp[5]) ? node3151 : node3144;
											assign node3144 = (inp[10]) ? node3148 : node3145;
												assign node3145 = (inp[13]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node3148 = (inp[7]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node3151 = (inp[4]) ? node3155 : node3152;
												assign node3152 = (inp[10]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node3155 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node3158 = (inp[1]) ? node3276 : node3159;
							assign node3159 = (inp[2]) ? node3219 : node3160;
								assign node3160 = (inp[10]) ? node3188 : node3161;
									assign node3161 = (inp[8]) ? node3173 : node3162;
										assign node3162 = (inp[7]) ? node3168 : node3163;
											assign node3163 = (inp[4]) ? node3165 : 14'b00001111111111;
												assign node3165 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3168 = (inp[13]) ? 14'b00000011111111 : node3169;
												assign node3169 = (inp[0]) ? 14'b00000001111111 : 14'b00000111111111;
										assign node3173 = (inp[0]) ? node3181 : node3174;
											assign node3174 = (inp[4]) ? node3178 : node3175;
												assign node3175 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3178 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3181 = (inp[13]) ? node3185 : node3182;
												assign node3182 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3185 = (inp[4]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node3188 = (inp[7]) ? node3204 : node3189;
										assign node3189 = (inp[5]) ? node3197 : node3190;
											assign node3190 = (inp[4]) ? node3194 : node3191;
												assign node3191 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3194 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3197 = (inp[0]) ? node3201 : node3198;
												assign node3198 = (inp[8]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node3201 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3204 = (inp[13]) ? node3212 : node3205;
											assign node3205 = (inp[8]) ? node3209 : node3206;
												assign node3206 = (inp[4]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node3209 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3212 = (inp[5]) ? node3216 : node3213;
												assign node3213 = (inp[4]) ? 14'b00000001111111 : 14'b00000000111111;
												assign node3216 = (inp[4]) ? 14'b00000000011111 : 14'b00000001111111;
								assign node3219 = (inp[0]) ? node3249 : node3220;
									assign node3220 = (inp[4]) ? node3234 : node3221;
										assign node3221 = (inp[7]) ? node3227 : node3222;
											assign node3222 = (inp[5]) ? 14'b00000011111111 : node3223;
												assign node3223 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3227 = (inp[10]) ? node3231 : node3228;
												assign node3228 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3231 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3234 = (inp[13]) ? node3242 : node3235;
											assign node3235 = (inp[10]) ? node3239 : node3236;
												assign node3236 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3239 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3242 = (inp[7]) ? node3246 : node3243;
												assign node3243 = (inp[5]) ? 14'b00000000011111 : 14'b00000001111111;
												assign node3246 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node3249 = (inp[8]) ? node3263 : node3250;
										assign node3250 = (inp[5]) ? node3258 : node3251;
											assign node3251 = (inp[7]) ? node3255 : node3252;
												assign node3252 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3255 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3258 = (inp[7]) ? node3260 : 14'b00000000111111;
												assign node3260 = (inp[4]) ? 14'b00000000001111 : 14'b00000001111111;
										assign node3263 = (inp[10]) ? node3269 : node3264;
											assign node3264 = (inp[4]) ? node3266 : 14'b00000000111111;
												assign node3266 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3269 = (inp[4]) ? node3273 : node3270;
												assign node3270 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3273 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node3276 = (inp[4]) ? node3336 : node3277;
								assign node3277 = (inp[7]) ? node3307 : node3278;
									assign node3278 = (inp[8]) ? node3294 : node3279;
										assign node3279 = (inp[0]) ? node3287 : node3280;
											assign node3280 = (inp[2]) ? node3284 : node3281;
												assign node3281 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3284 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3287 = (inp[2]) ? node3291 : node3288;
												assign node3288 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3291 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3294 = (inp[2]) ? node3302 : node3295;
											assign node3295 = (inp[13]) ? node3299 : node3296;
												assign node3296 = (inp[10]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node3299 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3302 = (inp[5]) ? node3304 : 14'b00000000111111;
												assign node3304 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node3307 = (inp[10]) ? node3321 : node3308;
										assign node3308 = (inp[13]) ? node3316 : node3309;
											assign node3309 = (inp[5]) ? node3313 : node3310;
												assign node3310 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3313 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3316 = (inp[2]) ? 14'b00000000111111 : node3317;
												assign node3317 = (inp[8]) ? 14'b00000000111111 : 14'b00000000111111;
										assign node3321 = (inp[13]) ? node3329 : node3322;
											assign node3322 = (inp[5]) ? node3326 : node3323;
												assign node3323 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3326 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3329 = (inp[5]) ? node3333 : node3330;
												assign node3330 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3333 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node3336 = (inp[13]) ? node3368 : node3337;
									assign node3337 = (inp[5]) ? node3353 : node3338;
										assign node3338 = (inp[2]) ? node3346 : node3339;
											assign node3339 = (inp[0]) ? node3343 : node3340;
												assign node3340 = (inp[8]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node3343 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3346 = (inp[0]) ? node3350 : node3347;
												assign node3347 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3350 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3353 = (inp[0]) ? node3361 : node3354;
											assign node3354 = (inp[8]) ? node3358 : node3355;
												assign node3355 = (inp[2]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node3358 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3361 = (inp[2]) ? node3365 : node3362;
												assign node3362 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3365 = (inp[8]) ? 14'b00000000000111 : 14'b00000000011111;
									assign node3368 = (inp[0]) ? node3384 : node3369;
										assign node3369 = (inp[10]) ? node3377 : node3370;
											assign node3370 = (inp[8]) ? node3374 : node3371;
												assign node3371 = (inp[5]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node3374 = (inp[2]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node3377 = (inp[7]) ? node3381 : node3378;
												assign node3378 = (inp[2]) ? 14'b00000000001111 : 14'b00000000111111;
												assign node3381 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node3384 = (inp[5]) ? node3392 : node3385;
											assign node3385 = (inp[2]) ? node3389 : node3386;
												assign node3386 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3389 = (inp[10]) ? 14'b00000000001111 : 14'b00000000001111;
											assign node3392 = (inp[2]) ? node3394 : 14'b00000000001111;
												assign node3394 = (inp[8]) ? 14'b00000000000111 : 14'b00000000000111;
					assign node3397 = (inp[2]) ? node3639 : node3398;
						assign node3398 = (inp[9]) ? node3520 : node3399;
							assign node3399 = (inp[5]) ? node3459 : node3400;
								assign node3400 = (inp[13]) ? node3428 : node3401;
									assign node3401 = (inp[10]) ? node3413 : node3402;
										assign node3402 = (inp[4]) ? node3408 : node3403;
											assign node3403 = (inp[7]) ? node3405 : 14'b00000111111111;
												assign node3405 = (inp[8]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node3408 = (inp[7]) ? 14'b00000011111111 : node3409;
												assign node3409 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node3413 = (inp[0]) ? node3421 : node3414;
											assign node3414 = (inp[7]) ? node3418 : node3415;
												assign node3415 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3418 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3421 = (inp[8]) ? node3425 : node3422;
												assign node3422 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3425 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node3428 = (inp[8]) ? node3444 : node3429;
										assign node3429 = (inp[4]) ? node3437 : node3430;
											assign node3430 = (inp[10]) ? node3434 : node3431;
												assign node3431 = (inp[0]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node3434 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3437 = (inp[0]) ? node3441 : node3438;
												assign node3438 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3441 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3444 = (inp[10]) ? node3452 : node3445;
											assign node3445 = (inp[1]) ? node3449 : node3446;
												assign node3446 = (inp[7]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node3449 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3452 = (inp[0]) ? node3456 : node3453;
												assign node3453 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3456 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node3459 = (inp[0]) ? node3491 : node3460;
									assign node3460 = (inp[13]) ? node3476 : node3461;
										assign node3461 = (inp[1]) ? node3469 : node3462;
											assign node3462 = (inp[10]) ? node3466 : node3463;
												assign node3463 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3466 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3469 = (inp[7]) ? node3473 : node3470;
												assign node3470 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3473 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3476 = (inp[8]) ? node3484 : node3477;
											assign node3477 = (inp[7]) ? node3481 : node3478;
												assign node3478 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3481 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3484 = (inp[4]) ? node3488 : node3485;
												assign node3485 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3488 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node3491 = (inp[8]) ? node3505 : node3492;
										assign node3492 = (inp[10]) ? node3498 : node3493;
											assign node3493 = (inp[1]) ? node3495 : 14'b00000011111111;
												assign node3495 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3498 = (inp[7]) ? node3502 : node3499;
												assign node3499 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3502 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3505 = (inp[4]) ? node3513 : node3506;
											assign node3506 = (inp[1]) ? node3510 : node3507;
												assign node3507 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3510 = (inp[13]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node3513 = (inp[7]) ? node3517 : node3514;
												assign node3514 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3517 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node3520 = (inp[4]) ? node3580 : node3521;
								assign node3521 = (inp[7]) ? node3551 : node3522;
									assign node3522 = (inp[1]) ? node3536 : node3523;
										assign node3523 = (inp[10]) ? node3531 : node3524;
											assign node3524 = (inp[0]) ? node3528 : node3525;
												assign node3525 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3528 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3531 = (inp[5]) ? 14'b00000001111111 : node3532;
												assign node3532 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3536 = (inp[0]) ? node3544 : node3537;
											assign node3537 = (inp[13]) ? node3541 : node3538;
												assign node3538 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3541 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3544 = (inp[13]) ? node3548 : node3545;
												assign node3545 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3548 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node3551 = (inp[5]) ? node3565 : node3552;
										assign node3552 = (inp[10]) ? node3558 : node3553;
											assign node3553 = (inp[1]) ? node3555 : 14'b00000001111111;
												assign node3555 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3558 = (inp[0]) ? node3562 : node3559;
												assign node3559 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3562 = (inp[1]) ? 14'b00000000011111 : 14'b00000000011111;
										assign node3565 = (inp[8]) ? node3573 : node3566;
											assign node3566 = (inp[10]) ? node3570 : node3567;
												assign node3567 = (inp[1]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node3570 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3573 = (inp[13]) ? node3577 : node3574;
												assign node3574 = (inp[0]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node3577 = (inp[0]) ? 14'b00000000000111 : 14'b00000000001111;
								assign node3580 = (inp[1]) ? node3608 : node3581;
									assign node3581 = (inp[10]) ? node3593 : node3582;
										assign node3582 = (inp[5]) ? node3588 : node3583;
											assign node3583 = (inp[7]) ? 14'b00000001111111 : node3584;
												assign node3584 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node3588 = (inp[8]) ? node3590 : 14'b00000001111111;
												assign node3590 = (inp[0]) ? 14'b00000000111111 : 14'b00000000111111;
										assign node3593 = (inp[7]) ? node3601 : node3594;
											assign node3594 = (inp[8]) ? node3598 : node3595;
												assign node3595 = (inp[5]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node3598 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3601 = (inp[5]) ? node3605 : node3602;
												assign node3602 = (inp[8]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node3605 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node3608 = (inp[5]) ? node3624 : node3609;
										assign node3609 = (inp[10]) ? node3617 : node3610;
											assign node3610 = (inp[0]) ? node3614 : node3611;
												assign node3611 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3614 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3617 = (inp[7]) ? node3621 : node3618;
												assign node3618 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3621 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node3624 = (inp[10]) ? node3632 : node3625;
											assign node3625 = (inp[13]) ? node3629 : node3626;
												assign node3626 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3629 = (inp[7]) ? 14'b00000000000111 : 14'b00000000011111;
											assign node3632 = (inp[8]) ? node3636 : node3633;
												assign node3633 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node3636 = (inp[0]) ? 14'b00000000000111 : 14'b00000000001111;
						assign node3639 = (inp[13]) ? node3759 : node3640;
							assign node3640 = (inp[7]) ? node3702 : node3641;
								assign node3641 = (inp[4]) ? node3673 : node3642;
									assign node3642 = (inp[1]) ? node3658 : node3643;
										assign node3643 = (inp[10]) ? node3651 : node3644;
											assign node3644 = (inp[5]) ? node3648 : node3645;
												assign node3645 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3648 = (inp[9]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node3651 = (inp[8]) ? node3655 : node3652;
												assign node3652 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3655 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node3658 = (inp[0]) ? node3666 : node3659;
											assign node3659 = (inp[8]) ? node3663 : node3660;
												assign node3660 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3663 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3666 = (inp[10]) ? node3670 : node3667;
												assign node3667 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3670 = (inp[9]) ? 14'b00000000011111 : 14'b00000000011111;
									assign node3673 = (inp[5]) ? node3689 : node3674;
										assign node3674 = (inp[9]) ? node3682 : node3675;
											assign node3675 = (inp[0]) ? node3679 : node3676;
												assign node3676 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3679 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3682 = (inp[10]) ? node3686 : node3683;
												assign node3683 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3686 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3689 = (inp[8]) ? node3695 : node3690;
											assign node3690 = (inp[0]) ? node3692 : 14'b00000001111111;
												assign node3692 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3695 = (inp[1]) ? node3699 : node3696;
												assign node3696 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3699 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node3702 = (inp[5]) ? node3732 : node3703;
									assign node3703 = (inp[1]) ? node3719 : node3704;
										assign node3704 = (inp[9]) ? node3712 : node3705;
											assign node3705 = (inp[8]) ? node3709 : node3706;
												assign node3706 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node3709 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3712 = (inp[10]) ? node3716 : node3713;
												assign node3713 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3716 = (inp[0]) ? 14'b00000000001111 : 14'b00000000111111;
										assign node3719 = (inp[0]) ? node3725 : node3720;
											assign node3720 = (inp[10]) ? node3722 : 14'b00000001111111;
												assign node3722 = (inp[9]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node3725 = (inp[10]) ? node3729 : node3726;
												assign node3726 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3729 = (inp[4]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node3732 = (inp[8]) ? node3744 : node3733;
										assign node3733 = (inp[1]) ? node3739 : node3734;
											assign node3734 = (inp[9]) ? node3736 : 14'b00000000111111;
												assign node3736 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3739 = (inp[4]) ? node3741 : 14'b00000000011111;
												assign node3741 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node3744 = (inp[9]) ? node3752 : node3745;
											assign node3745 = (inp[10]) ? node3749 : node3746;
												assign node3746 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3749 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node3752 = (inp[4]) ? node3756 : node3753;
												assign node3753 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node3756 = (inp[0]) ? 14'b00000000000111 : 14'b00000000001111;
							assign node3759 = (inp[8]) ? node3821 : node3760;
								assign node3760 = (inp[7]) ? node3792 : node3761;
									assign node3761 = (inp[4]) ? node3777 : node3762;
										assign node3762 = (inp[10]) ? node3770 : node3763;
											assign node3763 = (inp[0]) ? node3767 : node3764;
												assign node3764 = (inp[1]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node3767 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node3770 = (inp[5]) ? node3774 : node3771;
												assign node3771 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3774 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node3777 = (inp[10]) ? node3785 : node3778;
											assign node3778 = (inp[1]) ? node3782 : node3779;
												assign node3779 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3782 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3785 = (inp[9]) ? node3789 : node3786;
												assign node3786 = (inp[5]) ? 14'b00000000001111 : 14'b00000000111111;
												assign node3789 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node3792 = (inp[0]) ? node3806 : node3793;
										assign node3793 = (inp[4]) ? node3799 : node3794;
											assign node3794 = (inp[9]) ? node3796 : 14'b00000000111111;
												assign node3796 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3799 = (inp[9]) ? node3803 : node3800;
												assign node3800 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3803 = (inp[5]) ? 14'b00000000000111 : 14'b00000000011111;
										assign node3806 = (inp[10]) ? node3814 : node3807;
											assign node3807 = (inp[5]) ? node3811 : node3808;
												assign node3808 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3811 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node3814 = (inp[5]) ? node3818 : node3815;
												assign node3815 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node3818 = (inp[4]) ? 14'b00000000000011 : 14'b00000000001111;
								assign node3821 = (inp[9]) ? node3853 : node3822;
									assign node3822 = (inp[4]) ? node3838 : node3823;
										assign node3823 = (inp[7]) ? node3831 : node3824;
											assign node3824 = (inp[1]) ? node3828 : node3825;
												assign node3825 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node3828 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node3831 = (inp[10]) ? node3835 : node3832;
												assign node3832 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3835 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node3838 = (inp[0]) ? node3846 : node3839;
											assign node3839 = (inp[7]) ? node3843 : node3840;
												assign node3840 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3843 = (inp[5]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node3846 = (inp[7]) ? node3850 : node3847;
												assign node3847 = (inp[1]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node3850 = (inp[5]) ? 14'b00000000000111 : 14'b00000000000111;
									assign node3853 = (inp[5]) ? node3867 : node3854;
										assign node3854 = (inp[10]) ? node3862 : node3855;
											assign node3855 = (inp[4]) ? node3859 : node3856;
												assign node3856 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node3859 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node3862 = (inp[7]) ? node3864 : 14'b00000000001111;
												assign node3864 = (inp[4]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node3867 = (inp[4]) ? node3875 : node3868;
											assign node3868 = (inp[10]) ? node3872 : node3869;
												assign node3869 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node3872 = (inp[0]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node3875 = (inp[1]) ? node3879 : node3876;
												assign node3876 = (inp[0]) ? 14'b00000000000111 : 14'b00000000001111;
												assign node3879 = (inp[0]) ? 14'b00000000000011 : 14'b00000000000111;
		assign node3882 = (inp[5]) ? node5830 : node3883;
			assign node3883 = (inp[11]) ? node4849 : node3884;
				assign node3884 = (inp[9]) ? node4366 : node3885;
					assign node3885 = (inp[4]) ? node4123 : node3886;
						assign node3886 = (inp[7]) ? node4010 : node3887;
							assign node3887 = (inp[0]) ? node3947 : node3888;
								assign node3888 = (inp[1]) ? node3920 : node3889;
									assign node3889 = (inp[3]) ? node3905 : node3890;
										assign node3890 = (inp[10]) ? node3898 : node3891;
											assign node3891 = (inp[12]) ? node3895 : node3892;
												assign node3892 = (inp[8]) ? 14'b00011111111111 : 14'b00111111111111;
												assign node3895 = (inp[2]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node3898 = (inp[13]) ? node3902 : node3899;
												assign node3899 = (inp[12]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node3902 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node3905 = (inp[12]) ? node3913 : node3906;
											assign node3906 = (inp[13]) ? node3910 : node3907;
												assign node3907 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node3910 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3913 = (inp[10]) ? node3917 : node3914;
												assign node3914 = (inp[8]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node3917 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node3920 = (inp[2]) ? node3932 : node3921;
										assign node3921 = (inp[10]) ? node3927 : node3922;
											assign node3922 = (inp[12]) ? 14'b00001111111111 : node3923;
												assign node3923 = (inp[3]) ? 14'b00001111111111 : 14'b00011111111111;
											assign node3927 = (inp[8]) ? 14'b00000111111111 : node3928;
												assign node3928 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node3932 = (inp[12]) ? node3940 : node3933;
											assign node3933 = (inp[13]) ? node3937 : node3934;
												assign node3934 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3937 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3940 = (inp[8]) ? node3944 : node3941;
												assign node3941 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3944 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node3947 = (inp[2]) ? node3979 : node3948;
									assign node3948 = (inp[8]) ? node3964 : node3949;
										assign node3949 = (inp[13]) ? node3957 : node3950;
											assign node3950 = (inp[1]) ? node3954 : node3951;
												assign node3951 = (inp[12]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node3954 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node3957 = (inp[12]) ? node3961 : node3958;
												assign node3958 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3961 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node3964 = (inp[12]) ? node3972 : node3965;
											assign node3965 = (inp[3]) ? node3969 : node3966;
												assign node3966 = (inp[13]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node3969 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3972 = (inp[10]) ? node3976 : node3973;
												assign node3973 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node3976 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node3979 = (inp[3]) ? node3995 : node3980;
										assign node3980 = (inp[10]) ? node3988 : node3981;
											assign node3981 = (inp[8]) ? node3985 : node3982;
												assign node3982 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node3985 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node3988 = (inp[1]) ? node3992 : node3989;
												assign node3989 = (inp[12]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node3992 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node3995 = (inp[1]) ? node4003 : node3996;
											assign node3996 = (inp[10]) ? node4000 : node3997;
												assign node3997 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4000 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4003 = (inp[12]) ? node4007 : node4004;
												assign node4004 = (inp[8]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node4007 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node4010 = (inp[0]) ? node4064 : node4011;
								assign node4011 = (inp[13]) ? node4033 : node4012;
									assign node4012 = (inp[8]) ? node4024 : node4013;
										assign node4013 = (inp[12]) ? node4021 : node4014;
											assign node4014 = (inp[10]) ? node4018 : node4015;
												assign node4015 = (inp[3]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node4018 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node4021 = (inp[2]) ? 14'b00000111111111 : 14'b00000011111111;
										assign node4024 = (inp[2]) ? node4026 : 14'b00000111111111;
											assign node4026 = (inp[12]) ? node4030 : node4027;
												assign node4027 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4030 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node4033 = (inp[10]) ? node4049 : node4034;
										assign node4034 = (inp[12]) ? node4042 : node4035;
											assign node4035 = (inp[2]) ? node4039 : node4036;
												assign node4036 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4039 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4042 = (inp[1]) ? node4046 : node4043;
												assign node4043 = (inp[2]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node4046 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4049 = (inp[12]) ? node4057 : node4050;
											assign node4050 = (inp[3]) ? node4054 : node4051;
												assign node4051 = (inp[2]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node4054 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4057 = (inp[2]) ? node4061 : node4058;
												assign node4058 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4061 = (inp[1]) ? 14'b00000000111111 : 14'b00000000111111;
								assign node4064 = (inp[8]) ? node4094 : node4065;
									assign node4065 = (inp[1]) ? node4081 : node4066;
										assign node4066 = (inp[10]) ? node4074 : node4067;
											assign node4067 = (inp[2]) ? node4071 : node4068;
												assign node4068 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4071 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4074 = (inp[12]) ? node4078 : node4075;
												assign node4075 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4078 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4081 = (inp[10]) ? node4089 : node4082;
											assign node4082 = (inp[13]) ? node4086 : node4083;
												assign node4083 = (inp[2]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node4086 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4089 = (inp[2]) ? node4091 : 14'b00000001111111;
												assign node4091 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node4094 = (inp[12]) ? node4110 : node4095;
										assign node4095 = (inp[13]) ? node4103 : node4096;
											assign node4096 = (inp[1]) ? node4100 : node4097;
												assign node4097 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4100 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4103 = (inp[3]) ? node4107 : node4104;
												assign node4104 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4107 = (inp[1]) ? 14'b00000000011111 : 14'b00000001111111;
										assign node4110 = (inp[2]) ? node4118 : node4111;
											assign node4111 = (inp[10]) ? node4115 : node4112;
												assign node4112 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4115 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4118 = (inp[3]) ? 14'b00000000111111 : node4119;
												assign node4119 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node4123 = (inp[8]) ? node4245 : node4124;
							assign node4124 = (inp[0]) ? node4186 : node4125;
								assign node4125 = (inp[12]) ? node4157 : node4126;
									assign node4126 = (inp[7]) ? node4142 : node4127;
										assign node4127 = (inp[13]) ? node4135 : node4128;
											assign node4128 = (inp[1]) ? node4132 : node4129;
												assign node4129 = (inp[3]) ? 14'b00011111111111 : 14'b00011111111111;
												assign node4132 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node4135 = (inp[10]) ? node4139 : node4136;
												assign node4136 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4139 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node4142 = (inp[1]) ? node4150 : node4143;
											assign node4143 = (inp[3]) ? node4147 : node4144;
												assign node4144 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4147 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4150 = (inp[13]) ? node4154 : node4151;
												assign node4151 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4154 = (inp[10]) ? 14'b00000001111111 : 14'b00000001111111;
									assign node4157 = (inp[1]) ? node4173 : node4158;
										assign node4158 = (inp[10]) ? node4166 : node4159;
											assign node4159 = (inp[13]) ? node4163 : node4160;
												assign node4160 = (inp[3]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node4163 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4166 = (inp[2]) ? node4170 : node4167;
												assign node4167 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4170 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4173 = (inp[7]) ? node4181 : node4174;
											assign node4174 = (inp[3]) ? node4178 : node4175;
												assign node4175 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4178 = (inp[2]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node4181 = (inp[13]) ? node4183 : 14'b00000001111111;
												assign node4183 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node4186 = (inp[10]) ? node4216 : node4187;
									assign node4187 = (inp[1]) ? node4201 : node4188;
										assign node4188 = (inp[3]) ? node4196 : node4189;
											assign node4189 = (inp[13]) ? node4193 : node4190;
												assign node4190 = (inp[7]) ? 14'b00001111111111 : 14'b00001111111111;
												assign node4193 = (inp[12]) ? 14'b00000011111111 : 14'b00001111111111;
											assign node4196 = (inp[13]) ? 14'b00000011111111 : node4197;
												assign node4197 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node4201 = (inp[7]) ? node4209 : node4202;
											assign node4202 = (inp[13]) ? node4206 : node4203;
												assign node4203 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4206 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4209 = (inp[2]) ? node4213 : node4210;
												assign node4210 = (inp[12]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node4213 = (inp[12]) ? 14'b00000000111111 : 14'b00000000111111;
									assign node4216 = (inp[3]) ? node4232 : node4217;
										assign node4217 = (inp[7]) ? node4225 : node4218;
											assign node4218 = (inp[13]) ? node4222 : node4219;
												assign node4219 = (inp[1]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node4222 = (inp[12]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node4225 = (inp[12]) ? node4229 : node4226;
												assign node4226 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4229 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4232 = (inp[12]) ? node4238 : node4233;
											assign node4233 = (inp[7]) ? node4235 : 14'b00000001111111;
												assign node4235 = (inp[13]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node4238 = (inp[2]) ? node4242 : node4239;
												assign node4239 = (inp[13]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node4242 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node4245 = (inp[3]) ? node4307 : node4246;
								assign node4246 = (inp[13]) ? node4278 : node4247;
									assign node4247 = (inp[7]) ? node4263 : node4248;
										assign node4248 = (inp[12]) ? node4256 : node4249;
											assign node4249 = (inp[2]) ? node4253 : node4250;
												assign node4250 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4253 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4256 = (inp[1]) ? node4260 : node4257;
												assign node4257 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4260 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4263 = (inp[2]) ? node4271 : node4264;
											assign node4264 = (inp[0]) ? node4268 : node4265;
												assign node4265 = (inp[10]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node4268 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4271 = (inp[0]) ? node4275 : node4272;
												assign node4272 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4275 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node4278 = (inp[10]) ? node4294 : node4279;
										assign node4279 = (inp[2]) ? node4287 : node4280;
											assign node4280 = (inp[7]) ? node4284 : node4281;
												assign node4281 = (inp[1]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node4284 = (inp[0]) ? 14'b00000001111111 : 14'b00000001111111;
											assign node4287 = (inp[1]) ? node4291 : node4288;
												assign node4288 = (inp[7]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node4291 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4294 = (inp[12]) ? node4300 : node4295;
											assign node4295 = (inp[1]) ? node4297 : 14'b00000001111111;
												assign node4297 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4300 = (inp[1]) ? node4304 : node4301;
												assign node4301 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4304 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node4307 = (inp[1]) ? node4335 : node4308;
									assign node4308 = (inp[13]) ? node4322 : node4309;
										assign node4309 = (inp[0]) ? node4315 : node4310;
											assign node4310 = (inp[7]) ? 14'b00000001111111 : node4311;
												assign node4311 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4315 = (inp[7]) ? node4319 : node4316;
												assign node4316 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4319 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4322 = (inp[0]) ? node4330 : node4323;
											assign node4323 = (inp[2]) ? node4327 : node4324;
												assign node4324 = (inp[7]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node4327 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4330 = (inp[12]) ? node4332 : 14'b00000000111111;
												assign node4332 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node4335 = (inp[12]) ? node4351 : node4336;
										assign node4336 = (inp[13]) ? node4344 : node4337;
											assign node4337 = (inp[0]) ? node4341 : node4338;
												assign node4338 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4341 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4344 = (inp[10]) ? node4348 : node4345;
												assign node4345 = (inp[0]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node4348 = (inp[0]) ? 14'b00000000001111 : 14'b00000000111111;
										assign node4351 = (inp[10]) ? node4359 : node4352;
											assign node4352 = (inp[2]) ? node4356 : node4353;
												assign node4353 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4356 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4359 = (inp[2]) ? node4363 : node4360;
												assign node4360 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4363 = (inp[7]) ? 14'b00000000001111 : 14'b00000000001111;
					assign node4366 = (inp[1]) ? node4602 : node4367;
						assign node4367 = (inp[10]) ? node4479 : node4368;
							assign node4368 = (inp[13]) ? node4424 : node4369;
								assign node4369 = (inp[7]) ? node4401 : node4370;
									assign node4370 = (inp[3]) ? node4386 : node4371;
										assign node4371 = (inp[0]) ? node4379 : node4372;
											assign node4372 = (inp[2]) ? node4376 : node4373;
												assign node4373 = (inp[12]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node4376 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node4379 = (inp[12]) ? node4383 : node4380;
												assign node4380 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4383 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node4386 = (inp[4]) ? node4394 : node4387;
											assign node4387 = (inp[8]) ? node4391 : node4388;
												assign node4388 = (inp[0]) ? 14'b00000111111111 : 14'b00011111111111;
												assign node4391 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4394 = (inp[0]) ? node4398 : node4395;
												assign node4395 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4398 = (inp[12]) ? 14'b00000000111111 : 14'b00000011111111;
									assign node4401 = (inp[2]) ? node4413 : node4402;
										assign node4402 = (inp[4]) ? node4408 : node4403;
											assign node4403 = (inp[3]) ? node4405 : 14'b00011111111111;
												assign node4405 = (inp[8]) ? 14'b00000111111111 : 14'b00000111111111;
											assign node4408 = (inp[12]) ? 14'b00000001111111 : node4409;
												assign node4409 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node4413 = (inp[12]) ? node4419 : node4414;
											assign node4414 = (inp[4]) ? node4416 : 14'b00000011111111;
												assign node4416 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4419 = (inp[3]) ? node4421 : 14'b00000011111111;
												assign node4421 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node4424 = (inp[12]) ? node4454 : node4425;
									assign node4425 = (inp[0]) ? node4439 : node4426;
										assign node4426 = (inp[3]) ? node4434 : node4427;
											assign node4427 = (inp[7]) ? node4431 : node4428;
												assign node4428 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4431 = (inp[4]) ? 14'b00000011111111 : 14'b00000011111111;
											assign node4434 = (inp[4]) ? 14'b00000011111111 : node4435;
												assign node4435 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node4439 = (inp[3]) ? node4447 : node4440;
											assign node4440 = (inp[2]) ? node4444 : node4441;
												assign node4441 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4444 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4447 = (inp[7]) ? node4451 : node4448;
												assign node4448 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4451 = (inp[8]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node4454 = (inp[8]) ? node4464 : node4455;
										assign node4455 = (inp[0]) ? 14'b00000001111111 : node4456;
											assign node4456 = (inp[7]) ? node4460 : node4457;
												assign node4457 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4460 = (inp[4]) ? 14'b00000001111111 : 14'b00000001111111;
										assign node4464 = (inp[2]) ? node4472 : node4465;
											assign node4465 = (inp[3]) ? node4469 : node4466;
												assign node4466 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4469 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4472 = (inp[3]) ? node4476 : node4473;
												assign node4473 = (inp[0]) ? 14'b00000000011111 : 14'b00000001111111;
												assign node4476 = (inp[7]) ? 14'b00000000011111 : 14'b00000000011111;
							assign node4479 = (inp[3]) ? node4541 : node4480;
								assign node4480 = (inp[12]) ? node4510 : node4481;
									assign node4481 = (inp[7]) ? node4497 : node4482;
										assign node4482 = (inp[8]) ? node4490 : node4483;
											assign node4483 = (inp[0]) ? node4487 : node4484;
												assign node4484 = (inp[4]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4487 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4490 = (inp[4]) ? node4494 : node4491;
												assign node4491 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4494 = (inp[13]) ? 14'b00000011111111 : 14'b00000001111111;
										assign node4497 = (inp[13]) ? node4505 : node4498;
											assign node4498 = (inp[2]) ? node4502 : node4499;
												assign node4499 = (inp[4]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node4502 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4505 = (inp[0]) ? 14'b00000000111111 : node4506;
												assign node4506 = (inp[4]) ? 14'b00000001111111 : 14'b00000001111111;
									assign node4510 = (inp[13]) ? node4526 : node4511;
										assign node4511 = (inp[4]) ? node4519 : node4512;
											assign node4512 = (inp[2]) ? node4516 : node4513;
												assign node4513 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4516 = (inp[7]) ? 14'b00000011111111 : 14'b00000001111111;
											assign node4519 = (inp[2]) ? node4523 : node4520;
												assign node4520 = (inp[7]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node4523 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4526 = (inp[8]) ? node4534 : node4527;
											assign node4527 = (inp[7]) ? node4531 : node4528;
												assign node4528 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4531 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4534 = (inp[7]) ? node4538 : node4535;
												assign node4535 = (inp[0]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node4538 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node4541 = (inp[0]) ? node4573 : node4542;
									assign node4542 = (inp[7]) ? node4558 : node4543;
										assign node4543 = (inp[2]) ? node4551 : node4544;
											assign node4544 = (inp[8]) ? node4548 : node4545;
												assign node4545 = (inp[12]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node4548 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4551 = (inp[8]) ? node4555 : node4552;
												assign node4552 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4555 = (inp[4]) ? 14'b00000000011111 : 14'b00000001111111;
										assign node4558 = (inp[13]) ? node4566 : node4559;
											assign node4559 = (inp[8]) ? node4563 : node4560;
												assign node4560 = (inp[12]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node4563 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4566 = (inp[4]) ? node4570 : node4567;
												assign node4567 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4570 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node4573 = (inp[13]) ? node4589 : node4574;
										assign node4574 = (inp[7]) ? node4582 : node4575;
											assign node4575 = (inp[2]) ? node4579 : node4576;
												assign node4576 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4579 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4582 = (inp[12]) ? node4586 : node4583;
												assign node4583 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4586 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4589 = (inp[2]) ? node4595 : node4590;
											assign node4590 = (inp[12]) ? 14'b00000000111111 : node4591;
												assign node4591 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4595 = (inp[12]) ? node4599 : node4596;
												assign node4596 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4599 = (inp[4]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node4602 = (inp[13]) ? node4730 : node4603;
							assign node4603 = (inp[8]) ? node4667 : node4604;
								assign node4604 = (inp[4]) ? node4636 : node4605;
									assign node4605 = (inp[2]) ? node4621 : node4606;
										assign node4606 = (inp[12]) ? node4614 : node4607;
											assign node4607 = (inp[0]) ? node4611 : node4608;
												assign node4608 = (inp[7]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4611 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4614 = (inp[10]) ? node4618 : node4615;
												assign node4615 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4618 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4621 = (inp[7]) ? node4629 : node4622;
											assign node4622 = (inp[12]) ? node4626 : node4623;
												assign node4623 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4626 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4629 = (inp[12]) ? node4633 : node4630;
												assign node4630 = (inp[0]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node4633 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node4636 = (inp[3]) ? node4652 : node4637;
										assign node4637 = (inp[12]) ? node4645 : node4638;
											assign node4638 = (inp[10]) ? node4642 : node4639;
												assign node4639 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4642 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4645 = (inp[2]) ? node4649 : node4646;
												assign node4646 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4649 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4652 = (inp[0]) ? node4660 : node4653;
											assign node4653 = (inp[12]) ? node4657 : node4654;
												assign node4654 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4657 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4660 = (inp[2]) ? node4664 : node4661;
												assign node4661 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4664 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node4667 = (inp[3]) ? node4699 : node4668;
									assign node4668 = (inp[7]) ? node4684 : node4669;
										assign node4669 = (inp[12]) ? node4677 : node4670;
											assign node4670 = (inp[0]) ? node4674 : node4671;
												assign node4671 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4674 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4677 = (inp[0]) ? node4681 : node4678;
												assign node4678 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4681 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4684 = (inp[10]) ? node4692 : node4685;
											assign node4685 = (inp[0]) ? node4689 : node4686;
												assign node4686 = (inp[2]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node4689 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4692 = (inp[4]) ? node4696 : node4693;
												assign node4693 = (inp[12]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node4696 = (inp[12]) ? 14'b00000000011111 : 14'b00000000011111;
									assign node4699 = (inp[2]) ? node4715 : node4700;
										assign node4700 = (inp[7]) ? node4708 : node4701;
											assign node4701 = (inp[10]) ? node4705 : node4702;
												assign node4702 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4705 = (inp[0]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node4708 = (inp[4]) ? node4712 : node4709;
												assign node4709 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4712 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4715 = (inp[4]) ? node4723 : node4716;
											assign node4716 = (inp[10]) ? node4720 : node4717;
												assign node4717 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4720 = (inp[12]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node4723 = (inp[0]) ? node4727 : node4724;
												assign node4724 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4727 = (inp[7]) ? 14'b00000000001111 : 14'b00000000001111;
							assign node4730 = (inp[10]) ? node4792 : node4731;
								assign node4731 = (inp[7]) ? node4761 : node4732;
									assign node4732 = (inp[2]) ? node4746 : node4733;
										assign node4733 = (inp[12]) ? node4741 : node4734;
											assign node4734 = (inp[0]) ? node4738 : node4735;
												assign node4735 = (inp[3]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node4738 = (inp[3]) ? 14'b00000011111111 : 14'b00000001111111;
											assign node4741 = (inp[4]) ? 14'b00000001111111 : node4742;
												assign node4742 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4746 = (inp[8]) ? node4754 : node4747;
											assign node4747 = (inp[4]) ? node4751 : node4748;
												assign node4748 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4751 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4754 = (inp[4]) ? node4758 : node4755;
												assign node4755 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4758 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node4761 = (inp[3]) ? node4777 : node4762;
										assign node4762 = (inp[0]) ? node4770 : node4763;
											assign node4763 = (inp[2]) ? node4767 : node4764;
												assign node4764 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4767 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4770 = (inp[12]) ? node4774 : node4771;
												assign node4771 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4774 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4777 = (inp[12]) ? node4785 : node4778;
											assign node4778 = (inp[8]) ? node4782 : node4779;
												assign node4779 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4782 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4785 = (inp[4]) ? node4789 : node4786;
												assign node4786 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4789 = (inp[2]) ? 14'b00000000001111 : 14'b00000000001111;
								assign node4792 = (inp[4]) ? node4818 : node4793;
									assign node4793 = (inp[7]) ? node4809 : node4794;
										assign node4794 = (inp[8]) ? node4802 : node4795;
											assign node4795 = (inp[2]) ? node4799 : node4796;
												assign node4796 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4799 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4802 = (inp[0]) ? node4806 : node4803;
												assign node4803 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4806 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node4809 = (inp[0]) ? node4811 : 14'b00000000111111;
											assign node4811 = (inp[8]) ? node4815 : node4812;
												assign node4812 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4815 = (inp[2]) ? 14'b00000000000111 : 14'b00000000011111;
									assign node4818 = (inp[3]) ? node4834 : node4819;
										assign node4819 = (inp[2]) ? node4827 : node4820;
											assign node4820 = (inp[12]) ? node4824 : node4821;
												assign node4821 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4824 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node4827 = (inp[7]) ? node4831 : node4828;
												assign node4828 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4831 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node4834 = (inp[8]) ? node4842 : node4835;
											assign node4835 = (inp[12]) ? node4839 : node4836;
												assign node4836 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node4839 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node4842 = (inp[7]) ? node4846 : node4843;
												assign node4843 = (inp[12]) ? 14'b00000000000111 : 14'b00000000011111;
												assign node4846 = (inp[2]) ? 14'b00000000000111 : 14'b00000000001111;
				assign node4849 = (inp[7]) ? node5329 : node4850;
					assign node4850 = (inp[8]) ? node5090 : node4851;
						assign node4851 = (inp[13]) ? node4973 : node4852;
							assign node4852 = (inp[4]) ? node4914 : node4853;
								assign node4853 = (inp[1]) ? node4885 : node4854;
									assign node4854 = (inp[9]) ? node4870 : node4855;
										assign node4855 = (inp[12]) ? node4863 : node4856;
											assign node4856 = (inp[10]) ? node4860 : node4857;
												assign node4857 = (inp[3]) ? 14'b00001111111111 : 14'b00011111111111;
												assign node4860 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node4863 = (inp[0]) ? node4867 : node4864;
												assign node4864 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4867 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node4870 = (inp[0]) ? node4878 : node4871;
											assign node4871 = (inp[12]) ? node4875 : node4872;
												assign node4872 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4875 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4878 = (inp[10]) ? node4882 : node4879;
												assign node4879 = (inp[3]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4882 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node4885 = (inp[0]) ? node4899 : node4886;
										assign node4886 = (inp[3]) ? node4894 : node4887;
											assign node4887 = (inp[10]) ? node4891 : node4888;
												assign node4888 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4891 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4894 = (inp[12]) ? node4896 : 14'b00000011111111;
												assign node4896 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4899 = (inp[12]) ? node4907 : node4900;
											assign node4900 = (inp[2]) ? node4904 : node4901;
												assign node4901 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4904 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4907 = (inp[3]) ? node4911 : node4908;
												assign node4908 = (inp[2]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node4911 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node4914 = (inp[2]) ? node4942 : node4915;
									assign node4915 = (inp[9]) ? node4929 : node4916;
										assign node4916 = (inp[10]) ? node4922 : node4917;
											assign node4917 = (inp[3]) ? node4919 : 14'b00001111111111;
												assign node4919 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4922 = (inp[12]) ? node4926 : node4923;
												assign node4923 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4926 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4929 = (inp[3]) ? node4937 : node4930;
											assign node4930 = (inp[1]) ? node4934 : node4931;
												assign node4931 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4934 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4937 = (inp[0]) ? 14'b00000001111111 : node4938;
												assign node4938 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node4942 = (inp[1]) ? node4958 : node4943;
										assign node4943 = (inp[10]) ? node4951 : node4944;
											assign node4944 = (inp[3]) ? node4948 : node4945;
												assign node4945 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4948 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4951 = (inp[3]) ? node4955 : node4952;
												assign node4952 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4955 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node4958 = (inp[0]) ? node4966 : node4959;
											assign node4959 = (inp[3]) ? node4963 : node4960;
												assign node4960 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node4963 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node4966 = (inp[9]) ? node4970 : node4967;
												assign node4967 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node4970 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node4973 = (inp[0]) ? node5035 : node4974;
								assign node4974 = (inp[3]) ? node5006 : node4975;
									assign node4975 = (inp[12]) ? node4991 : node4976;
										assign node4976 = (inp[1]) ? node4984 : node4977;
											assign node4977 = (inp[4]) ? node4981 : node4978;
												assign node4978 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node4981 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node4984 = (inp[9]) ? node4988 : node4985;
												assign node4985 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node4988 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node4991 = (inp[9]) ? node4999 : node4992;
											assign node4992 = (inp[2]) ? node4996 : node4993;
												assign node4993 = (inp[1]) ? 14'b00000111111111 : 14'b00000111111111;
												assign node4996 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node4999 = (inp[2]) ? node5003 : node5000;
												assign node5000 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5003 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node5006 = (inp[10]) ? node5022 : node5007;
										assign node5007 = (inp[1]) ? node5015 : node5008;
											assign node5008 = (inp[4]) ? node5012 : node5009;
												assign node5009 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5012 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5015 = (inp[4]) ? node5019 : node5016;
												assign node5016 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5019 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5022 = (inp[9]) ? node5030 : node5023;
											assign node5023 = (inp[12]) ? node5027 : node5024;
												assign node5024 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5027 = (inp[4]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node5030 = (inp[12]) ? node5032 : 14'b00000000111111;
												assign node5032 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node5035 = (inp[1]) ? node5061 : node5036;
									assign node5036 = (inp[12]) ? node5050 : node5037;
										assign node5037 = (inp[9]) ? node5045 : node5038;
											assign node5038 = (inp[2]) ? node5042 : node5039;
												assign node5039 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5042 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5045 = (inp[2]) ? node5047 : 14'b00000011111111;
												assign node5047 = (inp[4]) ? 14'b00000000111111 : 14'b00000000111111;
										assign node5050 = (inp[10]) ? node5056 : node5051;
											assign node5051 = (inp[4]) ? node5053 : 14'b00000001111111;
												assign node5053 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5056 = (inp[3]) ? 14'b00000000111111 : node5057;
												assign node5057 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node5061 = (inp[2]) ? node5075 : node5062;
										assign node5062 = (inp[10]) ? node5070 : node5063;
											assign node5063 = (inp[12]) ? node5067 : node5064;
												assign node5064 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5067 = (inp[3]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node5070 = (inp[3]) ? node5072 : 14'b00000000111111;
												assign node5072 = (inp[9]) ? 14'b00000000001111 : 14'b00000000111111;
										assign node5075 = (inp[4]) ? node5083 : node5076;
											assign node5076 = (inp[9]) ? node5080 : node5077;
												assign node5077 = (inp[3]) ? 14'b00000001111111 : 14'b00000000111111;
												assign node5080 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5083 = (inp[12]) ? node5087 : node5084;
												assign node5084 = (inp[9]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node5087 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node5090 = (inp[2]) ? node5212 : node5091;
							assign node5091 = (inp[12]) ? node5149 : node5092;
								assign node5092 = (inp[1]) ? node5122 : node5093;
									assign node5093 = (inp[4]) ? node5107 : node5094;
										assign node5094 = (inp[10]) ? node5102 : node5095;
											assign node5095 = (inp[9]) ? node5099 : node5096;
												assign node5096 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node5099 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5102 = (inp[13]) ? 14'b00000011111111 : node5103;
												assign node5103 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node5107 = (inp[3]) ? node5115 : node5108;
											assign node5108 = (inp[9]) ? node5112 : node5109;
												assign node5109 = (inp[10]) ? 14'b00000011111111 : 14'b00001111111111;
												assign node5112 = (inp[10]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node5115 = (inp[0]) ? node5119 : node5116;
												assign node5116 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5119 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node5122 = (inp[9]) ? node5136 : node5123;
										assign node5123 = (inp[0]) ? node5131 : node5124;
											assign node5124 = (inp[4]) ? node5128 : node5125;
												assign node5125 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5128 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5131 = (inp[13]) ? 14'b00000000111111 : node5132;
												assign node5132 = (inp[4]) ? 14'b00000001111111 : 14'b00000001111111;
										assign node5136 = (inp[3]) ? node5144 : node5137;
											assign node5137 = (inp[13]) ? node5141 : node5138;
												assign node5138 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5141 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5144 = (inp[10]) ? node5146 : 14'b00000001111111;
												assign node5146 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node5149 = (inp[4]) ? node5181 : node5150;
									assign node5150 = (inp[0]) ? node5166 : node5151;
										assign node5151 = (inp[10]) ? node5159 : node5152;
											assign node5152 = (inp[3]) ? node5156 : node5153;
												assign node5153 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5156 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5159 = (inp[9]) ? node5163 : node5160;
												assign node5160 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5163 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5166 = (inp[13]) ? node5174 : node5167;
											assign node5167 = (inp[1]) ? node5171 : node5168;
												assign node5168 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5171 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5174 = (inp[10]) ? node5178 : node5175;
												assign node5175 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5178 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5181 = (inp[1]) ? node5197 : node5182;
										assign node5182 = (inp[9]) ? node5190 : node5183;
											assign node5183 = (inp[10]) ? node5187 : node5184;
												assign node5184 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5187 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5190 = (inp[3]) ? node5194 : node5191;
												assign node5191 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5194 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5197 = (inp[0]) ? node5205 : node5198;
											assign node5198 = (inp[3]) ? node5202 : node5199;
												assign node5199 = (inp[9]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node5202 = (inp[13]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node5205 = (inp[9]) ? node5209 : node5206;
												assign node5206 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5209 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node5212 = (inp[4]) ? node5272 : node5213;
								assign node5213 = (inp[9]) ? node5243 : node5214;
									assign node5214 = (inp[13]) ? node5228 : node5215;
										assign node5215 = (inp[3]) ? node5223 : node5216;
											assign node5216 = (inp[12]) ? node5220 : node5217;
												assign node5217 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5220 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5223 = (inp[0]) ? 14'b00000001111111 : node5224;
												assign node5224 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node5228 = (inp[10]) ? node5236 : node5229;
											assign node5229 = (inp[0]) ? node5233 : node5230;
												assign node5230 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5233 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5236 = (inp[12]) ? node5240 : node5237;
												assign node5237 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5240 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5243 = (inp[10]) ? node5257 : node5244;
										assign node5244 = (inp[13]) ? node5252 : node5245;
											assign node5245 = (inp[0]) ? node5249 : node5246;
												assign node5246 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5249 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5252 = (inp[1]) ? 14'b00000000011111 : node5253;
												assign node5253 = (inp[12]) ? 14'b00000000011111 : 14'b00000001111111;
										assign node5257 = (inp[0]) ? node5265 : node5258;
											assign node5258 = (inp[12]) ? node5262 : node5259;
												assign node5259 = (inp[1]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node5262 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5265 = (inp[12]) ? node5269 : node5266;
												assign node5266 = (inp[3]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node5269 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node5272 = (inp[12]) ? node5302 : node5273;
									assign node5273 = (inp[1]) ? node5287 : node5274;
										assign node5274 = (inp[0]) ? node5280 : node5275;
											assign node5275 = (inp[3]) ? node5277 : 14'b00000001111111;
												assign node5277 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5280 = (inp[10]) ? node5284 : node5281;
												assign node5281 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5284 = (inp[3]) ? 14'b00000000001111 : 14'b00000000111111;
										assign node5287 = (inp[10]) ? node5295 : node5288;
											assign node5288 = (inp[3]) ? node5292 : node5289;
												assign node5289 = (inp[13]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node5292 = (inp[9]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node5295 = (inp[0]) ? node5299 : node5296;
												assign node5296 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node5299 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node5302 = (inp[0]) ? node5316 : node5303;
										assign node5303 = (inp[9]) ? node5311 : node5304;
											assign node5304 = (inp[13]) ? node5308 : node5305;
												assign node5305 = (inp[10]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node5308 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5311 = (inp[1]) ? node5313 : 14'b00000000011111;
												assign node5313 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5316 = (inp[13]) ? node5322 : node5317;
											assign node5317 = (inp[1]) ? node5319 : 14'b00000000011111;
												assign node5319 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5322 = (inp[1]) ? node5326 : node5323;
												assign node5323 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node5326 = (inp[3]) ? 14'b00000000000111 : 14'b00000000000111;
					assign node5329 = (inp[1]) ? node5585 : node5330;
						assign node5330 = (inp[13]) ? node5458 : node5331;
							assign node5331 = (inp[10]) ? node5395 : node5332;
								assign node5332 = (inp[12]) ? node5364 : node5333;
									assign node5333 = (inp[3]) ? node5349 : node5334;
										assign node5334 = (inp[8]) ? node5342 : node5335;
											assign node5335 = (inp[4]) ? node5339 : node5336;
												assign node5336 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node5339 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5342 = (inp[4]) ? node5346 : node5343;
												assign node5343 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5346 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node5349 = (inp[8]) ? node5357 : node5350;
											assign node5350 = (inp[2]) ? node5354 : node5351;
												assign node5351 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5354 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5357 = (inp[4]) ? node5361 : node5358;
												assign node5358 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5361 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5364 = (inp[9]) ? node5380 : node5365;
										assign node5365 = (inp[3]) ? node5373 : node5366;
											assign node5366 = (inp[0]) ? node5370 : node5367;
												assign node5367 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5370 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5373 = (inp[2]) ? node5377 : node5374;
												assign node5374 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5377 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5380 = (inp[3]) ? node5388 : node5381;
											assign node5381 = (inp[4]) ? node5385 : node5382;
												assign node5382 = (inp[8]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node5385 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5388 = (inp[4]) ? node5392 : node5389;
												assign node5389 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5392 = (inp[0]) ? 14'b00000000011111 : 14'b00000000011111;
								assign node5395 = (inp[4]) ? node5427 : node5396;
									assign node5396 = (inp[8]) ? node5412 : node5397;
										assign node5397 = (inp[9]) ? node5405 : node5398;
											assign node5398 = (inp[3]) ? node5402 : node5399;
												assign node5399 = (inp[2]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node5402 = (inp[0]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node5405 = (inp[12]) ? node5409 : node5406;
												assign node5406 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5409 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5412 = (inp[0]) ? node5420 : node5413;
											assign node5413 = (inp[2]) ? node5417 : node5414;
												assign node5414 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5417 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5420 = (inp[9]) ? node5424 : node5421;
												assign node5421 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5424 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5427 = (inp[9]) ? node5443 : node5428;
										assign node5428 = (inp[12]) ? node5436 : node5429;
											assign node5429 = (inp[8]) ? node5433 : node5430;
												assign node5430 = (inp[2]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node5433 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5436 = (inp[2]) ? node5440 : node5437;
												assign node5437 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5440 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5443 = (inp[3]) ? node5451 : node5444;
											assign node5444 = (inp[2]) ? node5448 : node5445;
												assign node5445 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5448 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5451 = (inp[8]) ? node5455 : node5452;
												assign node5452 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5455 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node5458 = (inp[12]) ? node5522 : node5459;
								assign node5459 = (inp[9]) ? node5491 : node5460;
									assign node5460 = (inp[10]) ? node5476 : node5461;
										assign node5461 = (inp[8]) ? node5469 : node5462;
											assign node5462 = (inp[0]) ? node5466 : node5463;
												assign node5463 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5466 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5469 = (inp[2]) ? node5473 : node5470;
												assign node5470 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5473 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5476 = (inp[3]) ? node5484 : node5477;
											assign node5477 = (inp[8]) ? node5481 : node5478;
												assign node5478 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5481 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5484 = (inp[0]) ? node5488 : node5485;
												assign node5485 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5488 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5491 = (inp[2]) ? node5507 : node5492;
										assign node5492 = (inp[0]) ? node5500 : node5493;
											assign node5493 = (inp[10]) ? node5497 : node5494;
												assign node5494 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5497 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5500 = (inp[8]) ? node5504 : node5501;
												assign node5501 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5504 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5507 = (inp[3]) ? node5515 : node5508;
											assign node5508 = (inp[8]) ? node5512 : node5509;
												assign node5509 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5512 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5515 = (inp[10]) ? node5519 : node5516;
												assign node5516 = (inp[0]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node5519 = (inp[8]) ? 14'b00000000001111 : 14'b00000000001111;
								assign node5522 = (inp[4]) ? node5554 : node5523;
									assign node5523 = (inp[10]) ? node5539 : node5524;
										assign node5524 = (inp[9]) ? node5532 : node5525;
											assign node5525 = (inp[2]) ? node5529 : node5526;
												assign node5526 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5529 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5532 = (inp[2]) ? node5536 : node5533;
												assign node5533 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5536 = (inp[3]) ? 14'b00000000011111 : 14'b00000000011111;
										assign node5539 = (inp[9]) ? node5547 : node5540;
											assign node5540 = (inp[3]) ? node5544 : node5541;
												assign node5541 = (inp[0]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node5544 = (inp[0]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node5547 = (inp[8]) ? node5551 : node5548;
												assign node5548 = (inp[3]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node5551 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node5554 = (inp[0]) ? node5570 : node5555;
										assign node5555 = (inp[9]) ? node5563 : node5556;
											assign node5556 = (inp[2]) ? node5560 : node5557;
												assign node5557 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5560 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5563 = (inp[3]) ? node5567 : node5564;
												assign node5564 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5567 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5570 = (inp[2]) ? node5578 : node5571;
											assign node5571 = (inp[8]) ? node5575 : node5572;
												assign node5572 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5575 = (inp[3]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5578 = (inp[9]) ? node5582 : node5579;
												assign node5579 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node5582 = (inp[8]) ? 14'b00000000000111 : 14'b00000000001111;
						assign node5585 = (inp[3]) ? node5709 : node5586;
							assign node5586 = (inp[0]) ? node5650 : node5587;
								assign node5587 = (inp[10]) ? node5619 : node5588;
									assign node5588 = (inp[8]) ? node5604 : node5589;
										assign node5589 = (inp[12]) ? node5597 : node5590;
											assign node5590 = (inp[9]) ? node5594 : node5591;
												assign node5591 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5594 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5597 = (inp[4]) ? node5601 : node5598;
												assign node5598 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5601 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5604 = (inp[4]) ? node5612 : node5605;
											assign node5605 = (inp[12]) ? node5609 : node5606;
												assign node5606 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5609 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5612 = (inp[2]) ? node5616 : node5613;
												assign node5613 = (inp[9]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node5616 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node5619 = (inp[2]) ? node5635 : node5620;
										assign node5620 = (inp[12]) ? node5628 : node5621;
											assign node5621 = (inp[4]) ? node5625 : node5622;
												assign node5622 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5625 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5628 = (inp[9]) ? node5632 : node5629;
												assign node5629 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5632 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5635 = (inp[9]) ? node5643 : node5636;
											assign node5636 = (inp[4]) ? node5640 : node5637;
												assign node5637 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5640 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5643 = (inp[8]) ? node5647 : node5644;
												assign node5644 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5647 = (inp[4]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node5650 = (inp[13]) ? node5680 : node5651;
									assign node5651 = (inp[4]) ? node5665 : node5652;
										assign node5652 = (inp[8]) ? node5658 : node5653;
											assign node5653 = (inp[2]) ? 14'b00000001111111 : node5654;
												assign node5654 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5658 = (inp[9]) ? node5662 : node5659;
												assign node5659 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5662 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5665 = (inp[12]) ? node5673 : node5666;
											assign node5666 = (inp[10]) ? node5670 : node5667;
												assign node5667 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5670 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5673 = (inp[2]) ? node5677 : node5674;
												assign node5674 = (inp[9]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node5677 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node5680 = (inp[4]) ? node5696 : node5681;
										assign node5681 = (inp[2]) ? node5689 : node5682;
											assign node5682 = (inp[9]) ? node5686 : node5683;
												assign node5683 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5686 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5689 = (inp[9]) ? node5693 : node5690;
												assign node5690 = (inp[8]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node5693 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5696 = (inp[9]) ? node5704 : node5697;
											assign node5697 = (inp[12]) ? node5701 : node5698;
												assign node5698 = (inp[8]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node5701 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5704 = (inp[8]) ? node5706 : 14'b00000000001111;
												assign node5706 = (inp[2]) ? 14'b00000000000011 : 14'b00000000001111;
							assign node5709 = (inp[4]) ? node5769 : node5710;
								assign node5710 = (inp[13]) ? node5742 : node5711;
									assign node5711 = (inp[2]) ? node5727 : node5712;
										assign node5712 = (inp[8]) ? node5720 : node5713;
											assign node5713 = (inp[0]) ? node5717 : node5714;
												assign node5714 = (inp[12]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node5717 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5720 = (inp[10]) ? node5724 : node5721;
												assign node5721 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5724 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node5727 = (inp[8]) ? node5735 : node5728;
											assign node5728 = (inp[12]) ? node5732 : node5729;
												assign node5729 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5732 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5735 = (inp[0]) ? node5739 : node5736;
												assign node5736 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5739 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node5742 = (inp[12]) ? node5756 : node5743;
										assign node5743 = (inp[9]) ? node5751 : node5744;
											assign node5744 = (inp[2]) ? node5748 : node5745;
												assign node5745 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5748 = (inp[8]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node5751 = (inp[0]) ? node5753 : 14'b00000000011111;
												assign node5753 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5756 = (inp[10]) ? node5762 : node5757;
											assign node5757 = (inp[8]) ? 14'b00000000001111 : node5758;
												assign node5758 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node5762 = (inp[0]) ? node5766 : node5763;
												assign node5763 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node5766 = (inp[8]) ? 14'b00000000000011 : 14'b00000000000111;
								assign node5769 = (inp[8]) ? node5799 : node5770;
									assign node5770 = (inp[9]) ? node5784 : node5771;
										assign node5771 = (inp[13]) ? node5777 : node5772;
											assign node5772 = (inp[10]) ? 14'b00000000111111 : node5773;
												assign node5773 = (inp[12]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node5777 = (inp[2]) ? node5781 : node5778;
												assign node5778 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5781 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node5784 = (inp[13]) ? node5792 : node5785;
											assign node5785 = (inp[10]) ? node5789 : node5786;
												assign node5786 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node5789 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5792 = (inp[2]) ? node5796 : node5793;
												assign node5793 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node5796 = (inp[12]) ? 14'b00000000000011 : 14'b00000000001111;
									assign node5799 = (inp[10]) ? node5815 : node5800;
										assign node5800 = (inp[13]) ? node5808 : node5801;
											assign node5801 = (inp[0]) ? node5805 : node5802;
												assign node5802 = (inp[12]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node5805 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node5808 = (inp[9]) ? node5812 : node5809;
												assign node5809 = (inp[0]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node5812 = (inp[12]) ? 14'b00000000000011 : 14'b00000000001111;
										assign node5815 = (inp[12]) ? node5823 : node5816;
											assign node5816 = (inp[2]) ? node5820 : node5817;
												assign node5817 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node5820 = (inp[9]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node5823 = (inp[0]) ? node5827 : node5824;
												assign node5824 = (inp[2]) ? 14'b00000000000111 : 14'b00000000001111;
												assign node5827 = (inp[2]) ? 14'b00000000000011 : 14'b00000000000111;
			assign node5830 = (inp[3]) ? node6804 : node5831;
				assign node5831 = (inp[10]) ? node6315 : node5832;
					assign node5832 = (inp[4]) ? node6074 : node5833;
						assign node5833 = (inp[1]) ? node5949 : node5834;
							assign node5834 = (inp[13]) ? node5890 : node5835;
								assign node5835 = (inp[12]) ? node5865 : node5836;
									assign node5836 = (inp[9]) ? node5850 : node5837;
										assign node5837 = (inp[7]) ? node5843 : node5838;
											assign node5838 = (inp[2]) ? node5840 : 14'b00011111111111;
												assign node5840 = (inp[0]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node5843 = (inp[11]) ? node5847 : node5844;
												assign node5844 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node5847 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node5850 = (inp[8]) ? node5858 : node5851;
											assign node5851 = (inp[0]) ? node5855 : node5852;
												assign node5852 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node5855 = (inp[2]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node5858 = (inp[2]) ? node5862 : node5859;
												assign node5859 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5862 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node5865 = (inp[7]) ? node5875 : node5866;
										assign node5866 = (inp[0]) ? node5870 : node5867;
											assign node5867 = (inp[2]) ? 14'b00000111111111 : 14'b00001111111111;
											assign node5870 = (inp[2]) ? 14'b00000001111111 : node5871;
												assign node5871 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node5875 = (inp[11]) ? node5883 : node5876;
											assign node5876 = (inp[2]) ? node5880 : node5877;
												assign node5877 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5880 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5883 = (inp[0]) ? node5887 : node5884;
												assign node5884 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5887 = (inp[9]) ? 14'b00000000011111 : 14'b00000001111111;
								assign node5890 = (inp[9]) ? node5920 : node5891;
									assign node5891 = (inp[12]) ? node5905 : node5892;
										assign node5892 = (inp[2]) ? node5898 : node5893;
											assign node5893 = (inp[7]) ? node5895 : 14'b00001111111111;
												assign node5895 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5898 = (inp[0]) ? node5902 : node5899;
												assign node5899 = (inp[11]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node5902 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node5905 = (inp[0]) ? node5913 : node5906;
											assign node5906 = (inp[7]) ? node5910 : node5907;
												assign node5907 = (inp[11]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node5910 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5913 = (inp[11]) ? node5917 : node5914;
												assign node5914 = (inp[7]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node5917 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node5920 = (inp[7]) ? node5936 : node5921;
										assign node5921 = (inp[2]) ? node5929 : node5922;
											assign node5922 = (inp[0]) ? node5926 : node5923;
												assign node5923 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5926 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5929 = (inp[0]) ? node5933 : node5930;
												assign node5930 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node5933 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5936 = (inp[8]) ? node5942 : node5937;
											assign node5937 = (inp[11]) ? node5939 : 14'b00000001111111;
												assign node5939 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node5942 = (inp[0]) ? node5946 : node5943;
												assign node5943 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node5946 = (inp[2]) ? 14'b00000000011111 : 14'b00000000011111;
							assign node5949 = (inp[11]) ? node6011 : node5950;
								assign node5950 = (inp[7]) ? node5982 : node5951;
									assign node5951 = (inp[12]) ? node5967 : node5952;
										assign node5952 = (inp[8]) ? node5960 : node5953;
											assign node5953 = (inp[0]) ? node5957 : node5954;
												assign node5954 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node5957 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node5960 = (inp[0]) ? node5964 : node5961;
												assign node5961 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5964 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node5967 = (inp[13]) ? node5975 : node5968;
											assign node5968 = (inp[9]) ? node5972 : node5969;
												assign node5969 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5972 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5975 = (inp[2]) ? node5979 : node5976;
												assign node5976 = (inp[8]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node5979 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node5982 = (inp[9]) ? node5998 : node5983;
										assign node5983 = (inp[2]) ? node5991 : node5984;
											assign node5984 = (inp[12]) ? node5988 : node5985;
												assign node5985 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node5988 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node5991 = (inp[8]) ? node5995 : node5992;
												assign node5992 = (inp[12]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node5995 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node5998 = (inp[13]) ? node6004 : node5999;
											assign node5999 = (inp[0]) ? node6001 : 14'b00000001111111;
												assign node6001 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node6004 = (inp[0]) ? node6008 : node6005;
												assign node6005 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6008 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node6011 = (inp[2]) ? node6043 : node6012;
									assign node6012 = (inp[13]) ? node6028 : node6013;
										assign node6013 = (inp[8]) ? node6021 : node6014;
											assign node6014 = (inp[7]) ? node6018 : node6015;
												assign node6015 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node6018 = (inp[12]) ? 14'b00000001111111 : 14'b00000111111111;
											assign node6021 = (inp[0]) ? node6025 : node6022;
												assign node6022 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6025 = (inp[9]) ? 14'b00000000011111 : 14'b00000001111111;
										assign node6028 = (inp[0]) ? node6036 : node6029;
											assign node6029 = (inp[8]) ? node6033 : node6030;
												assign node6030 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6033 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6036 = (inp[7]) ? node6040 : node6037;
												assign node6037 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6040 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node6043 = (inp[12]) ? node6059 : node6044;
										assign node6044 = (inp[0]) ? node6052 : node6045;
											assign node6045 = (inp[7]) ? node6049 : node6046;
												assign node6046 = (inp[13]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node6049 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6052 = (inp[8]) ? node6056 : node6053;
												assign node6053 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6056 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6059 = (inp[7]) ? node6067 : node6060;
											assign node6060 = (inp[9]) ? node6064 : node6061;
												assign node6061 = (inp[8]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node6064 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6067 = (inp[0]) ? node6071 : node6068;
												assign node6068 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node6071 = (inp[9]) ? 14'b00000000000111 : 14'b00000000001111;
						assign node6074 = (inp[7]) ? node6190 : node6075;
							assign node6075 = (inp[8]) ? node6137 : node6076;
								assign node6076 = (inp[11]) ? node6108 : node6077;
									assign node6077 = (inp[0]) ? node6093 : node6078;
										assign node6078 = (inp[13]) ? node6086 : node6079;
											assign node6079 = (inp[12]) ? node6083 : node6080;
												assign node6080 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node6083 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node6086 = (inp[9]) ? node6090 : node6087;
												assign node6087 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node6090 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node6093 = (inp[2]) ? node6101 : node6094;
											assign node6094 = (inp[1]) ? node6098 : node6095;
												assign node6095 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node6098 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node6101 = (inp[13]) ? node6105 : node6102;
												assign node6102 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6105 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node6108 = (inp[0]) ? node6122 : node6109;
										assign node6109 = (inp[13]) ? node6115 : node6110;
											assign node6110 = (inp[12]) ? 14'b00000011111111 : node6111;
												assign node6111 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node6115 = (inp[1]) ? node6119 : node6116;
												assign node6116 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6119 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node6122 = (inp[2]) ? node6130 : node6123;
											assign node6123 = (inp[12]) ? node6127 : node6124;
												assign node6124 = (inp[9]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node6127 = (inp[9]) ? 14'b00000000111111 : 14'b00000000111111;
											assign node6130 = (inp[13]) ? node6134 : node6131;
												assign node6131 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6134 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node6137 = (inp[12]) ? node6167 : node6138;
									assign node6138 = (inp[0]) ? node6152 : node6139;
										assign node6139 = (inp[11]) ? node6145 : node6140;
											assign node6140 = (inp[13]) ? node6142 : 14'b00000011111111;
												assign node6142 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node6145 = (inp[13]) ? node6149 : node6146;
												assign node6146 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6149 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node6152 = (inp[9]) ? node6160 : node6153;
											assign node6153 = (inp[1]) ? node6157 : node6154;
												assign node6154 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6157 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6160 = (inp[13]) ? node6164 : node6161;
												assign node6161 = (inp[2]) ? 14'b00000000011111 : 14'b00000001111111;
												assign node6164 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node6167 = (inp[9]) ? node6177 : node6168;
										assign node6168 = (inp[1]) ? 14'b00000000111111 : node6169;
											assign node6169 = (inp[0]) ? node6173 : node6170;
												assign node6170 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6173 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6177 = (inp[13]) ? node6183 : node6178;
											assign node6178 = (inp[11]) ? 14'b00000000111111 : node6179;
												assign node6179 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6183 = (inp[1]) ? node6187 : node6184;
												assign node6184 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6187 = (inp[11]) ? 14'b00000000001111 : 14'b00000000111111;
							assign node6190 = (inp[8]) ? node6254 : node6191;
								assign node6191 = (inp[13]) ? node6223 : node6192;
									assign node6192 = (inp[0]) ? node6208 : node6193;
										assign node6193 = (inp[12]) ? node6201 : node6194;
											assign node6194 = (inp[1]) ? node6198 : node6195;
												assign node6195 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node6198 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node6201 = (inp[1]) ? node6205 : node6202;
												assign node6202 = (inp[11]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node6205 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node6208 = (inp[11]) ? node6216 : node6209;
											assign node6209 = (inp[2]) ? node6213 : node6210;
												assign node6210 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6213 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6216 = (inp[1]) ? node6220 : node6217;
												assign node6217 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6220 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node6223 = (inp[9]) ? node6239 : node6224;
										assign node6224 = (inp[0]) ? node6232 : node6225;
											assign node6225 = (inp[2]) ? node6229 : node6226;
												assign node6226 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6229 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6232 = (inp[2]) ? node6236 : node6233;
												assign node6233 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6236 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6239 = (inp[12]) ? node6247 : node6240;
											assign node6240 = (inp[2]) ? node6244 : node6241;
												assign node6241 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6244 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6247 = (inp[11]) ? node6251 : node6248;
												assign node6248 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6251 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node6254 = (inp[11]) ? node6284 : node6255;
									assign node6255 = (inp[1]) ? node6269 : node6256;
										assign node6256 = (inp[9]) ? node6262 : node6257;
											assign node6257 = (inp[12]) ? node6259 : 14'b00000001111111;
												assign node6259 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6262 = (inp[0]) ? node6266 : node6263;
												assign node6263 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6266 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6269 = (inp[9]) ? node6277 : node6270;
											assign node6270 = (inp[13]) ? node6274 : node6271;
												assign node6271 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6274 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6277 = (inp[0]) ? node6281 : node6278;
												assign node6278 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6281 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node6284 = (inp[0]) ? node6300 : node6285;
										assign node6285 = (inp[2]) ? node6293 : node6286;
											assign node6286 = (inp[12]) ? node6290 : node6287;
												assign node6287 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6290 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6293 = (inp[13]) ? node6297 : node6294;
												assign node6294 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6297 = (inp[9]) ? 14'b00000000000111 : 14'b00000000011111;
										assign node6300 = (inp[12]) ? node6308 : node6301;
											assign node6301 = (inp[2]) ? node6305 : node6302;
												assign node6302 = (inp[1]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node6305 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node6308 = (inp[9]) ? node6312 : node6309;
												assign node6309 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node6312 = (inp[13]) ? 14'b00000000000111 : 14'b00000000001111;
					assign node6315 = (inp[9]) ? node6561 : node6316;
						assign node6316 = (inp[12]) ? node6442 : node6317;
							assign node6317 = (inp[0]) ? node6381 : node6318;
								assign node6318 = (inp[1]) ? node6350 : node6319;
									assign node6319 = (inp[8]) ? node6335 : node6320;
										assign node6320 = (inp[7]) ? node6328 : node6321;
											assign node6321 = (inp[4]) ? node6325 : node6322;
												assign node6322 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
												assign node6325 = (inp[2]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node6328 = (inp[11]) ? node6332 : node6329;
												assign node6329 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node6332 = (inp[13]) ? 14'b00000001111111 : 14'b00000001111111;
										assign node6335 = (inp[4]) ? node6343 : node6336;
											assign node6336 = (inp[2]) ? node6340 : node6337;
												assign node6337 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node6340 = (inp[11]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node6343 = (inp[11]) ? node6347 : node6344;
												assign node6344 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6347 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node6350 = (inp[11]) ? node6366 : node6351;
										assign node6351 = (inp[4]) ? node6359 : node6352;
											assign node6352 = (inp[7]) ? node6356 : node6353;
												assign node6353 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node6356 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node6359 = (inp[7]) ? node6363 : node6360;
												assign node6360 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6363 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node6366 = (inp[2]) ? node6374 : node6367;
											assign node6367 = (inp[8]) ? node6371 : node6368;
												assign node6368 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6371 = (inp[4]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node6374 = (inp[4]) ? node6378 : node6375;
												assign node6375 = (inp[8]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node6378 = (inp[7]) ? 14'b00000000001111 : 14'b00000000111111;
								assign node6381 = (inp[13]) ? node6411 : node6382;
									assign node6382 = (inp[7]) ? node6398 : node6383;
										assign node6383 = (inp[11]) ? node6391 : node6384;
											assign node6384 = (inp[4]) ? node6388 : node6385;
												assign node6385 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node6388 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node6391 = (inp[2]) ? node6395 : node6392;
												assign node6392 = (inp[4]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node6395 = (inp[4]) ? 14'b00000000111111 : 14'b00000000111111;
										assign node6398 = (inp[11]) ? node6404 : node6399;
											assign node6399 = (inp[4]) ? node6401 : 14'b00000001111111;
												assign node6401 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6404 = (inp[4]) ? node6408 : node6405;
												assign node6405 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6408 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node6411 = (inp[2]) ? node6427 : node6412;
										assign node6412 = (inp[1]) ? node6420 : node6413;
											assign node6413 = (inp[4]) ? node6417 : node6414;
												assign node6414 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6417 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6420 = (inp[4]) ? node6424 : node6421;
												assign node6421 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6424 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6427 = (inp[8]) ? node6435 : node6428;
											assign node6428 = (inp[4]) ? node6432 : node6429;
												assign node6429 = (inp[7]) ? 14'b00000000011111 : 14'b00000001111111;
												assign node6432 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6435 = (inp[7]) ? node6439 : node6436;
												assign node6436 = (inp[1]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node6439 = (inp[11]) ? 14'b00000000000111 : 14'b00000000011111;
							assign node6442 = (inp[4]) ? node6500 : node6443;
								assign node6443 = (inp[11]) ? node6471 : node6444;
									assign node6444 = (inp[8]) ? node6460 : node6445;
										assign node6445 = (inp[13]) ? node6453 : node6446;
											assign node6446 = (inp[2]) ? node6450 : node6447;
												assign node6447 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node6450 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node6453 = (inp[1]) ? node6457 : node6454;
												assign node6454 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6457 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node6460 = (inp[1]) ? node6468 : node6461;
											assign node6461 = (inp[13]) ? node6465 : node6462;
												assign node6462 = (inp[7]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node6465 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6468 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node6471 = (inp[0]) ? node6487 : node6472;
										assign node6472 = (inp[1]) ? node6480 : node6473;
											assign node6473 = (inp[2]) ? node6477 : node6474;
												assign node6474 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6477 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6480 = (inp[13]) ? node6484 : node6481;
												assign node6481 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6484 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6487 = (inp[7]) ? node6493 : node6488;
											assign node6488 = (inp[8]) ? node6490 : 14'b00000000111111;
												assign node6490 = (inp[1]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node6493 = (inp[13]) ? node6497 : node6494;
												assign node6494 = (inp[2]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node6497 = (inp[8]) ? 14'b00000000000111 : 14'b00000000001111;
								assign node6500 = (inp[13]) ? node6532 : node6501;
									assign node6501 = (inp[0]) ? node6517 : node6502;
										assign node6502 = (inp[1]) ? node6510 : node6503;
											assign node6503 = (inp[11]) ? node6507 : node6504;
												assign node6504 = (inp[8]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node6507 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6510 = (inp[8]) ? node6514 : node6511;
												assign node6511 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6514 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6517 = (inp[7]) ? node6525 : node6518;
											assign node6518 = (inp[1]) ? node6522 : node6519;
												assign node6519 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6522 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6525 = (inp[8]) ? node6529 : node6526;
												assign node6526 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6529 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node6532 = (inp[11]) ? node6546 : node6533;
										assign node6533 = (inp[2]) ? node6541 : node6534;
											assign node6534 = (inp[1]) ? node6538 : node6535;
												assign node6535 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6538 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6541 = (inp[0]) ? 14'b00000000001111 : node6542;
												assign node6542 = (inp[8]) ? 14'b00000000011111 : 14'b00000000011111;
										assign node6546 = (inp[8]) ? node6554 : node6547;
											assign node6547 = (inp[0]) ? node6551 : node6548;
												assign node6548 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6551 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node6554 = (inp[2]) ? node6558 : node6555;
												assign node6555 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node6558 = (inp[0]) ? 14'b00000000000111 : 14'b00000000001111;
						assign node6561 = (inp[2]) ? node6685 : node6562;
							assign node6562 = (inp[12]) ? node6624 : node6563;
								assign node6563 = (inp[11]) ? node6595 : node6564;
									assign node6564 = (inp[0]) ? node6580 : node6565;
										assign node6565 = (inp[8]) ? node6573 : node6566;
											assign node6566 = (inp[13]) ? node6570 : node6567;
												assign node6567 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node6570 = (inp[4]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node6573 = (inp[13]) ? node6577 : node6574;
												assign node6574 = (inp[4]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node6577 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node6580 = (inp[13]) ? node6588 : node6581;
											assign node6581 = (inp[8]) ? node6585 : node6582;
												assign node6582 = (inp[7]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node6585 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6588 = (inp[1]) ? node6592 : node6589;
												assign node6589 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6592 = (inp[4]) ? 14'b00000000001111 : 14'b00000000111111;
									assign node6595 = (inp[1]) ? node6609 : node6596;
										assign node6596 = (inp[4]) ? node6602 : node6597;
											assign node6597 = (inp[8]) ? 14'b00000001111111 : node6598;
												assign node6598 = (inp[13]) ? 14'b00000000111111 : 14'b00000011111111;
											assign node6602 = (inp[7]) ? node6606 : node6603;
												assign node6603 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6606 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6609 = (inp[4]) ? node6617 : node6610;
											assign node6610 = (inp[13]) ? node6614 : node6611;
												assign node6611 = (inp[7]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node6614 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6617 = (inp[0]) ? node6621 : node6618;
												assign node6618 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6621 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node6624 = (inp[7]) ? node6654 : node6625;
									assign node6625 = (inp[11]) ? node6639 : node6626;
										assign node6626 = (inp[13]) ? node6632 : node6627;
											assign node6627 = (inp[8]) ? node6629 : 14'b00000011111111;
												assign node6629 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6632 = (inp[4]) ? node6636 : node6633;
												assign node6633 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6636 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6639 = (inp[1]) ? node6647 : node6640;
											assign node6640 = (inp[0]) ? node6644 : node6641;
												assign node6641 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6644 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6647 = (inp[8]) ? node6651 : node6648;
												assign node6648 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6651 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node6654 = (inp[13]) ? node6670 : node6655;
										assign node6655 = (inp[1]) ? node6663 : node6656;
											assign node6656 = (inp[4]) ? node6660 : node6657;
												assign node6657 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6660 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6663 = (inp[8]) ? node6667 : node6664;
												assign node6664 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6667 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node6670 = (inp[4]) ? node6678 : node6671;
											assign node6671 = (inp[0]) ? node6675 : node6672;
												assign node6672 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6675 = (inp[11]) ? 14'b00000000001111 : 14'b00000000001111;
											assign node6678 = (inp[11]) ? node6682 : node6679;
												assign node6679 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node6682 = (inp[8]) ? 14'b00000000000111 : 14'b00000000001111;
							assign node6685 = (inp[13]) ? node6745 : node6686;
								assign node6686 = (inp[8]) ? node6716 : node6687;
									assign node6687 = (inp[11]) ? node6701 : node6688;
										assign node6688 = (inp[7]) ? node6694 : node6689;
											assign node6689 = (inp[12]) ? node6691 : 14'b00000011111111;
												assign node6691 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6694 = (inp[4]) ? node6698 : node6695;
												assign node6695 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6698 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6701 = (inp[7]) ? node6709 : node6702;
											assign node6702 = (inp[1]) ? node6706 : node6703;
												assign node6703 = (inp[12]) ? 14'b00000000011111 : 14'b00000001111111;
												assign node6706 = (inp[0]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node6709 = (inp[4]) ? node6713 : node6710;
												assign node6710 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6713 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node6716 = (inp[7]) ? node6732 : node6717;
										assign node6717 = (inp[1]) ? node6725 : node6718;
											assign node6718 = (inp[11]) ? node6722 : node6719;
												assign node6719 = (inp[12]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node6722 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6725 = (inp[12]) ? node6729 : node6726;
												assign node6726 = (inp[11]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6729 = (inp[4]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node6732 = (inp[1]) ? node6740 : node6733;
											assign node6733 = (inp[11]) ? node6737 : node6734;
												assign node6734 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6737 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node6740 = (inp[12]) ? node6742 : 14'b00000000001111;
												assign node6742 = (inp[11]) ? 14'b00000000000011 : 14'b00000000001111;
								assign node6745 = (inp[4]) ? node6775 : node6746;
									assign node6746 = (inp[12]) ? node6762 : node6747;
										assign node6747 = (inp[1]) ? node6755 : node6748;
											assign node6748 = (inp[0]) ? node6752 : node6749;
												assign node6749 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6752 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6755 = (inp[0]) ? node6759 : node6756;
												assign node6756 = (inp[7]) ? 14'b00000000001111 : 14'b00000000111111;
												assign node6759 = (inp[8]) ? 14'b00000000001111 : 14'b00000000001111;
										assign node6762 = (inp[8]) ? node6770 : node6763;
											assign node6763 = (inp[0]) ? node6767 : node6764;
												assign node6764 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6767 = (inp[7]) ? 14'b00000000001111 : 14'b00000000001111;
											assign node6770 = (inp[0]) ? 14'b00000000000111 : node6771;
												assign node6771 = (inp[7]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node6775 = (inp[8]) ? node6789 : node6776;
										assign node6776 = (inp[7]) ? node6782 : node6777;
											assign node6777 = (inp[1]) ? node6779 : 14'b00000000011111;
												assign node6779 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node6782 = (inp[1]) ? node6786 : node6783;
												assign node6783 = (inp[12]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node6786 = (inp[11]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node6789 = (inp[11]) ? node6797 : node6790;
											assign node6790 = (inp[12]) ? node6794 : node6791;
												assign node6791 = (inp[1]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node6794 = (inp[0]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node6797 = (inp[12]) ? node6801 : node6798;
												assign node6798 = (inp[7]) ? 14'b00000000000011 : 14'b00000000001111;
												assign node6801 = (inp[0]) ? 14'b00000000000011 : 14'b00000000000011;
				assign node6804 = (inp[11]) ? node7280 : node6805;
					assign node6805 = (inp[1]) ? node7043 : node6806;
						assign node6806 = (inp[8]) ? node6918 : node6807;
							assign node6807 = (inp[2]) ? node6869 : node6808;
								assign node6808 = (inp[4]) ? node6838 : node6809;
									assign node6809 = (inp[10]) ? node6823 : node6810;
										assign node6810 = (inp[7]) ? node6816 : node6811;
											assign node6811 = (inp[0]) ? node6813 : 14'b00001111111111;
												assign node6813 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node6816 = (inp[0]) ? node6820 : node6817;
												assign node6817 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node6820 = (inp[9]) ? 14'b00000001111111 : 14'b00000001111111;
										assign node6823 = (inp[9]) ? node6831 : node6824;
											assign node6824 = (inp[12]) ? node6828 : node6825;
												assign node6825 = (inp[0]) ? 14'b00000011111111 : 14'b00000011111111;
												assign node6828 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node6831 = (inp[12]) ? node6835 : node6832;
												assign node6832 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6835 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node6838 = (inp[12]) ? node6854 : node6839;
										assign node6839 = (inp[10]) ? node6847 : node6840;
											assign node6840 = (inp[13]) ? node6844 : node6841;
												assign node6841 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node6844 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node6847 = (inp[7]) ? node6851 : node6848;
												assign node6848 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6851 = (inp[9]) ? 14'b00000000011111 : 14'b00000001111111;
										assign node6854 = (inp[0]) ? node6862 : node6855;
											assign node6855 = (inp[9]) ? node6859 : node6856;
												assign node6856 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6859 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6862 = (inp[13]) ? node6866 : node6863;
												assign node6863 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6866 = (inp[9]) ? 14'b00000000011111 : 14'b00000000011111;
								assign node6869 = (inp[13]) ? node6895 : node6870;
									assign node6870 = (inp[0]) ? node6882 : node6871;
										assign node6871 = (inp[9]) ? node6877 : node6872;
											assign node6872 = (inp[12]) ? node6874 : 14'b00000111111111;
												assign node6874 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node6877 = (inp[10]) ? 14'b00000001111111 : node6878;
												assign node6878 = (inp[12]) ? 14'b00000001111111 : 14'b00000001111111;
										assign node6882 = (inp[12]) ? node6888 : node6883;
											assign node6883 = (inp[7]) ? 14'b00000000111111 : node6884;
												assign node6884 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node6888 = (inp[9]) ? node6892 : node6889;
												assign node6889 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6892 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node6895 = (inp[4]) ? node6909 : node6896;
										assign node6896 = (inp[0]) ? node6902 : node6897;
											assign node6897 = (inp[9]) ? node6899 : 14'b00000011111111;
												assign node6899 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6902 = (inp[12]) ? node6906 : node6903;
												assign node6903 = (inp[7]) ? 14'b00000000011111 : 14'b00000001111111;
												assign node6906 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6909 = (inp[10]) ? node6915 : node6910;
											assign node6910 = (inp[0]) ? node6912 : 14'b00000000111111;
												assign node6912 = (inp[7]) ? 14'b00000000001111 : 14'b00000000111111;
											assign node6915 = (inp[9]) ? 14'b00000000001111 : 14'b00000000111111;
							assign node6918 = (inp[10]) ? node6982 : node6919;
								assign node6919 = (inp[0]) ? node6951 : node6920;
									assign node6920 = (inp[2]) ? node6936 : node6921;
										assign node6921 = (inp[13]) ? node6929 : node6922;
											assign node6922 = (inp[4]) ? node6926 : node6923;
												assign node6923 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node6926 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node6929 = (inp[7]) ? node6933 : node6930;
												assign node6930 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6933 = (inp[4]) ? 14'b00000000011111 : 14'b00000001111111;
										assign node6936 = (inp[12]) ? node6944 : node6937;
											assign node6937 = (inp[9]) ? node6941 : node6938;
												assign node6938 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6941 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6944 = (inp[9]) ? node6948 : node6945;
												assign node6945 = (inp[4]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node6948 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node6951 = (inp[13]) ? node6967 : node6952;
										assign node6952 = (inp[7]) ? node6960 : node6953;
											assign node6953 = (inp[12]) ? node6957 : node6954;
												assign node6954 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6957 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6960 = (inp[4]) ? node6964 : node6961;
												assign node6961 = (inp[12]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node6964 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6967 = (inp[12]) ? node6975 : node6968;
											assign node6968 = (inp[7]) ? node6972 : node6969;
												assign node6969 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6972 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node6975 = (inp[9]) ? node6979 : node6976;
												assign node6976 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node6979 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node6982 = (inp[12]) ? node7014 : node6983;
									assign node6983 = (inp[9]) ? node6999 : node6984;
										assign node6984 = (inp[4]) ? node6992 : node6985;
											assign node6985 = (inp[7]) ? node6989 : node6986;
												assign node6986 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node6989 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node6992 = (inp[2]) ? node6996 : node6993;
												assign node6993 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node6996 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node6999 = (inp[7]) ? node7007 : node7000;
											assign node7000 = (inp[13]) ? node7004 : node7001;
												assign node7001 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7004 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node7007 = (inp[13]) ? node7011 : node7008;
												assign node7008 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7011 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node7014 = (inp[13]) ? node7030 : node7015;
										assign node7015 = (inp[0]) ? node7023 : node7016;
											assign node7016 = (inp[9]) ? node7020 : node7017;
												assign node7017 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7020 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node7023 = (inp[2]) ? node7027 : node7024;
												assign node7024 = (inp[7]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node7027 = (inp[4]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node7030 = (inp[2]) ? node7036 : node7031;
											assign node7031 = (inp[0]) ? node7033 : 14'b00000001111111;
												assign node7033 = (inp[4]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node7036 = (inp[7]) ? node7040 : node7037;
												assign node7037 = (inp[0]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node7040 = (inp[4]) ? 14'b00000000000011 : 14'b00000000001111;
						assign node7043 = (inp[10]) ? node7159 : node7044;
							assign node7044 = (inp[7]) ? node7104 : node7045;
								assign node7045 = (inp[13]) ? node7075 : node7046;
									assign node7046 = (inp[9]) ? node7060 : node7047;
										assign node7047 = (inp[2]) ? node7053 : node7048;
											assign node7048 = (inp[8]) ? 14'b00000011111111 : node7049;
												assign node7049 = (inp[4]) ? 14'b00000011111111 : 14'b00000111111111;
											assign node7053 = (inp[4]) ? node7057 : node7054;
												assign node7054 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node7057 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node7060 = (inp[4]) ? node7068 : node7061;
											assign node7061 = (inp[12]) ? node7065 : node7062;
												assign node7062 = (inp[8]) ? 14'b00000001111111 : 14'b00000111111111;
												assign node7065 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node7068 = (inp[12]) ? node7072 : node7069;
												assign node7069 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7072 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node7075 = (inp[8]) ? node7089 : node7076;
										assign node7076 = (inp[4]) ? node7082 : node7077;
											assign node7077 = (inp[9]) ? node7079 : 14'b00000001111111;
												assign node7079 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node7082 = (inp[2]) ? node7086 : node7083;
												assign node7083 = (inp[9]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node7086 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node7089 = (inp[0]) ? node7097 : node7090;
											assign node7090 = (inp[12]) ? node7094 : node7091;
												assign node7091 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7094 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node7097 = (inp[9]) ? node7101 : node7098;
												assign node7098 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7101 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node7104 = (inp[4]) ? node7136 : node7105;
									assign node7105 = (inp[8]) ? node7121 : node7106;
										assign node7106 = (inp[9]) ? node7114 : node7107;
											assign node7107 = (inp[2]) ? node7111 : node7108;
												assign node7108 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node7111 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node7114 = (inp[2]) ? node7118 : node7115;
												assign node7115 = (inp[13]) ? 14'b00000000111111 : 14'b00000011111111;
												assign node7118 = (inp[12]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node7121 = (inp[12]) ? node7129 : node7122;
											assign node7122 = (inp[13]) ? node7126 : node7123;
												assign node7123 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7126 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node7129 = (inp[2]) ? node7133 : node7130;
												assign node7130 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7133 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node7136 = (inp[0]) ? node7144 : node7137;
										assign node7137 = (inp[9]) ? node7139 : 14'b00000000111111;
											assign node7139 = (inp[12]) ? 14'b00000000011111 : node7140;
												assign node7140 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node7144 = (inp[8]) ? node7152 : node7145;
											assign node7145 = (inp[9]) ? node7149 : node7146;
												assign node7146 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7149 = (inp[12]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node7152 = (inp[2]) ? node7156 : node7153;
												assign node7153 = (inp[13]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node7156 = (inp[9]) ? 14'b00000000000011 : 14'b00000000001111;
							assign node7159 = (inp[13]) ? node7221 : node7160;
								assign node7160 = (inp[12]) ? node7192 : node7161;
									assign node7161 = (inp[8]) ? node7177 : node7162;
										assign node7162 = (inp[2]) ? node7170 : node7163;
											assign node7163 = (inp[4]) ? node7167 : node7164;
												assign node7164 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node7167 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node7170 = (inp[7]) ? node7174 : node7171;
												assign node7171 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7174 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node7177 = (inp[9]) ? node7185 : node7178;
											assign node7178 = (inp[7]) ? node7182 : node7179;
												assign node7179 = (inp[2]) ? 14'b00000001111111 : 14'b00000001111111;
												assign node7182 = (inp[4]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node7185 = (inp[2]) ? node7189 : node7186;
												assign node7186 = (inp[7]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node7189 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node7192 = (inp[7]) ? node7206 : node7193;
										assign node7193 = (inp[2]) ? node7201 : node7194;
											assign node7194 = (inp[4]) ? node7198 : node7195;
												assign node7195 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7198 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node7201 = (inp[9]) ? node7203 : 14'b00000000011111;
												assign node7203 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node7206 = (inp[9]) ? node7214 : node7207;
											assign node7207 = (inp[4]) ? node7211 : node7208;
												assign node7208 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7211 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node7214 = (inp[0]) ? node7218 : node7215;
												assign node7215 = (inp[2]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node7218 = (inp[2]) ? 14'b00000000000111 : 14'b00000000001111;
								assign node7221 = (inp[2]) ? node7251 : node7222;
									assign node7222 = (inp[4]) ? node7238 : node7223;
										assign node7223 = (inp[12]) ? node7231 : node7224;
											assign node7224 = (inp[7]) ? node7228 : node7225;
												assign node7225 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7228 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node7231 = (inp[9]) ? node7235 : node7232;
												assign node7232 = (inp[8]) ? 14'b00000000001111 : 14'b00000000111111;
												assign node7235 = (inp[8]) ? 14'b00000000001111 : 14'b00000000001111;
										assign node7238 = (inp[7]) ? node7246 : node7239;
											assign node7239 = (inp[0]) ? node7243 : node7240;
												assign node7240 = (inp[9]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node7243 = (inp[9]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node7246 = (inp[9]) ? node7248 : 14'b00000000001111;
												assign node7248 = (inp[12]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node7251 = (inp[9]) ? node7265 : node7252;
										assign node7252 = (inp[4]) ? node7258 : node7253;
											assign node7253 = (inp[12]) ? 14'b00000000011111 : node7254;
												assign node7254 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node7258 = (inp[12]) ? node7262 : node7259;
												assign node7259 = (inp[7]) ? 14'b00000000000111 : 14'b00000000011111;
												assign node7262 = (inp[8]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node7265 = (inp[0]) ? node7273 : node7266;
											assign node7266 = (inp[12]) ? node7270 : node7267;
												assign node7267 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node7270 = (inp[4]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node7273 = (inp[8]) ? node7277 : node7274;
												assign node7274 = (inp[4]) ? 14'b00000000000111 : 14'b00000000001111;
												assign node7277 = (inp[4]) ? 14'b00000000000011 : 14'b00000000000011;
					assign node7280 = (inp[12]) ? node7522 : node7281;
						assign node7281 = (inp[7]) ? node7403 : node7282;
							assign node7282 = (inp[9]) ? node7342 : node7283;
								assign node7283 = (inp[0]) ? node7313 : node7284;
									assign node7284 = (inp[4]) ? node7300 : node7285;
										assign node7285 = (inp[8]) ? node7293 : node7286;
											assign node7286 = (inp[1]) ? node7290 : node7287;
												assign node7287 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
												assign node7290 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
											assign node7293 = (inp[2]) ? node7297 : node7294;
												assign node7294 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node7297 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node7300 = (inp[10]) ? node7308 : node7301;
											assign node7301 = (inp[2]) ? node7305 : node7302;
												assign node7302 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node7305 = (inp[1]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node7308 = (inp[2]) ? node7310 : 14'b00000000111111;
												assign node7310 = (inp[1]) ? 14'b00000000011111 : 14'b00000000011111;
									assign node7313 = (inp[8]) ? node7329 : node7314;
										assign node7314 = (inp[2]) ? node7322 : node7315;
											assign node7315 = (inp[1]) ? node7319 : node7316;
												assign node7316 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node7319 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node7322 = (inp[13]) ? node7326 : node7323;
												assign node7323 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7326 = (inp[4]) ? 14'b00000000011111 : 14'b00000000011111;
										assign node7329 = (inp[10]) ? node7337 : node7330;
											assign node7330 = (inp[4]) ? node7334 : node7331;
												assign node7331 = (inp[2]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node7334 = (inp[1]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node7337 = (inp[1]) ? 14'b00000000011111 : node7338;
												assign node7338 = (inp[2]) ? 14'b00000000011111 : 14'b00000000011111;
								assign node7342 = (inp[13]) ? node7372 : node7343;
									assign node7343 = (inp[0]) ? node7359 : node7344;
										assign node7344 = (inp[8]) ? node7352 : node7345;
											assign node7345 = (inp[1]) ? node7349 : node7346;
												assign node7346 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node7349 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node7352 = (inp[10]) ? node7356 : node7353;
												assign node7353 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7356 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node7359 = (inp[2]) ? node7367 : node7360;
											assign node7360 = (inp[1]) ? node7364 : node7361;
												assign node7361 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7364 = (inp[10]) ? 14'b00000000011111 : 14'b00000000011111;
											assign node7367 = (inp[4]) ? 14'b00000000001111 : node7368;
												assign node7368 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node7372 = (inp[2]) ? node7388 : node7373;
										assign node7373 = (inp[10]) ? node7381 : node7374;
											assign node7374 = (inp[0]) ? node7378 : node7375;
												assign node7375 = (inp[4]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7378 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node7381 = (inp[8]) ? node7385 : node7382;
												assign node7382 = (inp[1]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7385 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node7388 = (inp[8]) ? node7396 : node7389;
											assign node7389 = (inp[1]) ? node7393 : node7390;
												assign node7390 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7393 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node7396 = (inp[10]) ? node7400 : node7397;
												assign node7397 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node7400 = (inp[4]) ? 14'b00000000000111 : 14'b00000000001111;
							assign node7403 = (inp[1]) ? node7459 : node7404;
								assign node7404 = (inp[4]) ? node7430 : node7405;
									assign node7405 = (inp[2]) ? node7421 : node7406;
										assign node7406 = (inp[10]) ? node7414 : node7407;
											assign node7407 = (inp[9]) ? node7411 : node7408;
												assign node7408 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node7411 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node7414 = (inp[8]) ? node7418 : node7415;
												assign node7415 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7418 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
										assign node7421 = (inp[0]) ? node7425 : node7422;
											assign node7422 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node7425 = (inp[9]) ? 14'b00000000001111 : node7426;
												assign node7426 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node7430 = (inp[8]) ? node7444 : node7431;
										assign node7431 = (inp[13]) ? node7437 : node7432;
											assign node7432 = (inp[10]) ? 14'b00000000111111 : node7433;
												assign node7433 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node7437 = (inp[9]) ? node7441 : node7438;
												assign node7438 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7441 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node7444 = (inp[0]) ? node7452 : node7445;
											assign node7445 = (inp[13]) ? node7449 : node7446;
												assign node7446 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7449 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node7452 = (inp[13]) ? node7456 : node7453;
												assign node7453 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node7456 = (inp[2]) ? 14'b00000000000011 : 14'b00000000001111;
								assign node7459 = (inp[10]) ? node7491 : node7460;
									assign node7460 = (inp[4]) ? node7476 : node7461;
										assign node7461 = (inp[13]) ? node7469 : node7462;
											assign node7462 = (inp[2]) ? node7466 : node7463;
												assign node7463 = (inp[8]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node7466 = (inp[0]) ? 14'b00000000011111 : 14'b00000001111111;
											assign node7469 = (inp[9]) ? node7473 : node7470;
												assign node7470 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7473 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node7476 = (inp[0]) ? node7484 : node7477;
											assign node7477 = (inp[8]) ? node7481 : node7478;
												assign node7478 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7481 = (inp[13]) ? 14'b00000000001111 : 14'b00000000001111;
											assign node7484 = (inp[9]) ? node7488 : node7485;
												assign node7485 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node7488 = (inp[13]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node7491 = (inp[0]) ? node7507 : node7492;
										assign node7492 = (inp[2]) ? node7500 : node7493;
											assign node7493 = (inp[8]) ? node7497 : node7494;
												assign node7494 = (inp[9]) ? 14'b00000000001111 : 14'b00000000111111;
												assign node7497 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node7500 = (inp[4]) ? node7504 : node7501;
												assign node7501 = (inp[8]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node7504 = (inp[9]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node7507 = (inp[8]) ? node7515 : node7508;
											assign node7508 = (inp[4]) ? node7512 : node7509;
												assign node7509 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node7512 = (inp[9]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node7515 = (inp[4]) ? node7519 : node7516;
												assign node7516 = (inp[2]) ? 14'b00000000000011 : 14'b00000000001111;
												assign node7519 = (inp[9]) ? 14'b00000000000011 : 14'b00000000000011;
						assign node7522 = (inp[1]) ? node7648 : node7523;
							assign node7523 = (inp[9]) ? node7585 : node7524;
								assign node7524 = (inp[4]) ? node7554 : node7525;
									assign node7525 = (inp[2]) ? node7541 : node7526;
										assign node7526 = (inp[7]) ? node7534 : node7527;
											assign node7527 = (inp[8]) ? node7531 : node7528;
												assign node7528 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
												assign node7531 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
											assign node7534 = (inp[0]) ? node7538 : node7535;
												assign node7535 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7538 = (inp[8]) ? 14'b00000000011111 : 14'b00000000011111;
										assign node7541 = (inp[13]) ? node7549 : node7542;
											assign node7542 = (inp[10]) ? node7546 : node7543;
												assign node7543 = (inp[0]) ? 14'b00000000111111 : 14'b00000000111111;
												assign node7546 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node7549 = (inp[0]) ? 14'b00000000011111 : node7550;
												assign node7550 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node7554 = (inp[10]) ? node7570 : node7555;
										assign node7555 = (inp[8]) ? node7563 : node7556;
											assign node7556 = (inp[7]) ? node7560 : node7557;
												assign node7557 = (inp[13]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7560 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node7563 = (inp[7]) ? node7567 : node7564;
												assign node7564 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7567 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node7570 = (inp[7]) ? node7578 : node7571;
											assign node7571 = (inp[8]) ? node7575 : node7572;
												assign node7572 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7575 = (inp[13]) ? 14'b00000000000111 : 14'b00000000011111;
											assign node7578 = (inp[13]) ? node7582 : node7579;
												assign node7579 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node7582 = (inp[0]) ? 14'b00000000000111 : 14'b00000000001111;
								assign node7585 = (inp[2]) ? node7617 : node7586;
									assign node7586 = (inp[4]) ? node7602 : node7587;
										assign node7587 = (inp[7]) ? node7595 : node7588;
											assign node7588 = (inp[10]) ? node7592 : node7589;
												assign node7589 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7592 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node7595 = (inp[13]) ? node7599 : node7596;
												assign node7596 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7599 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node7602 = (inp[10]) ? node7610 : node7603;
											assign node7603 = (inp[0]) ? node7607 : node7604;
												assign node7604 = (inp[8]) ? 14'b00000000011111 : 14'b00000000011111;
												assign node7607 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node7610 = (inp[7]) ? node7614 : node7611;
												assign node7611 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node7614 = (inp[0]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node7617 = (inp[10]) ? node7633 : node7618;
										assign node7618 = (inp[7]) ? node7626 : node7619;
											assign node7619 = (inp[4]) ? node7623 : node7620;
												assign node7620 = (inp[13]) ? 14'b00000000001111 : 14'b00000000111111;
												assign node7623 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node7626 = (inp[13]) ? node7630 : node7627;
												assign node7627 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node7630 = (inp[8]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node7633 = (inp[4]) ? node7641 : node7634;
											assign node7634 = (inp[8]) ? node7638 : node7635;
												assign node7635 = (inp[7]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node7638 = (inp[7]) ? 14'b00000000001111 : 14'b00000000000111;
											assign node7641 = (inp[7]) ? node7645 : node7642;
												assign node7642 = (inp[0]) ? 14'b00000000000111 : 14'b00000000000111;
												assign node7645 = (inp[13]) ? 14'b00000000000001 : 14'b00000000000111;
							assign node7648 = (inp[0]) ? node7712 : node7649;
								assign node7649 = (inp[4]) ? node7681 : node7650;
									assign node7650 = (inp[9]) ? node7666 : node7651;
										assign node7651 = (inp[13]) ? node7659 : node7652;
											assign node7652 = (inp[2]) ? node7656 : node7653;
												assign node7653 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
												assign node7656 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
											assign node7659 = (inp[7]) ? node7663 : node7660;
												assign node7660 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7663 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
										assign node7666 = (inp[2]) ? node7674 : node7667;
											assign node7667 = (inp[8]) ? node7671 : node7668;
												assign node7668 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7671 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node7674 = (inp[13]) ? node7678 : node7675;
												assign node7675 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node7678 = (inp[7]) ? 14'b00000000000111 : 14'b00000000001111;
									assign node7681 = (inp[10]) ? node7697 : node7682;
										assign node7682 = (inp[7]) ? node7690 : node7683;
											assign node7683 = (inp[9]) ? node7687 : node7684;
												assign node7684 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
												assign node7687 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node7690 = (inp[8]) ? node7694 : node7691;
												assign node7691 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node7694 = (inp[2]) ? 14'b00000000000111 : 14'b00000000000111;
										assign node7697 = (inp[9]) ? node7705 : node7698;
											assign node7698 = (inp[13]) ? node7702 : node7699;
												assign node7699 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node7702 = (inp[2]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node7705 = (inp[2]) ? node7709 : node7706;
												assign node7706 = (inp[8]) ? 14'b00000000000111 : 14'b00000000001111;
												assign node7709 = (inp[8]) ? 14'b00000000000011 : 14'b00000000000011;
								assign node7712 = (inp[10]) ? node7742 : node7713;
									assign node7713 = (inp[7]) ? node7727 : node7714;
										assign node7714 = (inp[4]) ? node7720 : node7715;
											assign node7715 = (inp[2]) ? node7717 : 14'b00000000111111;
												assign node7717 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
											assign node7720 = (inp[13]) ? node7724 : node7721;
												assign node7721 = (inp[9]) ? 14'b00000000001111 : 14'b00000000001111;
												assign node7724 = (inp[2]) ? 14'b00000000000111 : 14'b00000000001111;
										assign node7727 = (inp[13]) ? node7735 : node7728;
											assign node7728 = (inp[9]) ? node7732 : node7729;
												assign node7729 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node7732 = (inp[8]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node7735 = (inp[2]) ? node7739 : node7736;
												assign node7736 = (inp[4]) ? 14'b00000000000111 : 14'b00000000000111;
												assign node7739 = (inp[9]) ? 14'b00000000000011 : 14'b00000000000111;
									assign node7742 = (inp[13]) ? node7758 : node7743;
										assign node7743 = (inp[4]) ? node7751 : node7744;
											assign node7744 = (inp[7]) ? node7748 : node7745;
												assign node7745 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
												assign node7748 = (inp[8]) ? 14'b00000000000111 : 14'b00000000001111;
											assign node7751 = (inp[7]) ? node7755 : node7752;
												assign node7752 = (inp[9]) ? 14'b00000000000011 : 14'b00000000001111;
												assign node7755 = (inp[2]) ? 14'b00000000000011 : 14'b00000000000011;
										assign node7758 = (inp[9]) ? node7766 : node7759;
											assign node7759 = (inp[8]) ? node7763 : node7760;
												assign node7760 = (inp[4]) ? 14'b00000000000111 : 14'b00000000000111;
												assign node7763 = (inp[7]) ? 14'b00000000000011 : 14'b00000000000111;
											assign node7766 = (inp[4]) ? node7770 : node7767;
												assign node7767 = (inp[2]) ? 14'b00000000000001 : 14'b00000000000011;
												assign node7770 = (inp[2]) ? 14'b00000000000000 : 14'b00000000000001;

endmodule