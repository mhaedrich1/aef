module dtc_split5_bm88 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node87;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node133;
	wire [3-1:0] node135;
	wire [3-1:0] node137;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node161;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node258;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node266;
	wire [3-1:0] node268;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node294;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node356;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node363;
	wire [3-1:0] node366;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node400;
	wire [3-1:0] node402;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node411;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node420;
	wire [3-1:0] node423;
	wire [3-1:0] node425;
	wire [3-1:0] node428;
	wire [3-1:0] node430;
	wire [3-1:0] node432;
	wire [3-1:0] node434;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node441;
	wire [3-1:0] node443;
	wire [3-1:0] node445;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node452;
	wire [3-1:0] node454;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node485;
	wire [3-1:0] node488;
	wire [3-1:0] node490;
	wire [3-1:0] node492;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node502;
	wire [3-1:0] node505;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node511;
	wire [3-1:0] node514;
	wire [3-1:0] node516;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node536;
	wire [3-1:0] node539;
	wire [3-1:0] node541;
	wire [3-1:0] node543;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node556;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node568;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node576;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node583;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node590;
	wire [3-1:0] node593;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node627;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node636;
	wire [3-1:0] node639;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node652;
	wire [3-1:0] node653;
	wire [3-1:0] node656;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node663;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node682;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node689;
	wire [3-1:0] node692;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node703;
	wire [3-1:0] node706;
	wire [3-1:0] node708;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node715;
	wire [3-1:0] node717;
	wire [3-1:0] node719;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node731;
	wire [3-1:0] node734;
	wire [3-1:0] node736;
	wire [3-1:0] node739;
	wire [3-1:0] node741;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node746;
	wire [3-1:0] node748;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node759;
	wire [3-1:0] node762;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node769;
	wire [3-1:0] node772;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node782;
	wire [3-1:0] node785;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node789;
	wire [3-1:0] node792;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node814;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node829;
	wire [3-1:0] node831;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node841;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node850;
	wire [3-1:0] node852;
	wire [3-1:0] node855;
	wire [3-1:0] node857;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node864;
	wire [3-1:0] node867;
	wire [3-1:0] node868;
	wire [3-1:0] node871;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node879;
	wire [3-1:0] node882;
	wire [3-1:0] node884;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node894;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node900;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node915;
	wire [3-1:0] node916;
	wire [3-1:0] node918;
	wire [3-1:0] node919;
	wire [3-1:0] node922;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node931;
	wire [3-1:0] node932;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node938;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node943;
	wire [3-1:0] node946;
	wire [3-1:0] node949;
	wire [3-1:0] node950;
	wire [3-1:0] node953;
	wire [3-1:0] node955;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node966;
	wire [3-1:0] node967;
	wire [3-1:0] node968;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node981;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node985;
	wire [3-1:0] node989;
	wire [3-1:0] node990;
	wire [3-1:0] node993;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node998;
	wire [3-1:0] node999;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1009;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1018;
	wire [3-1:0] node1019;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1034;
	wire [3-1:0] node1035;
	wire [3-1:0] node1037;
	wire [3-1:0] node1041;
	wire [3-1:0] node1043;
	wire [3-1:0] node1044;
	wire [3-1:0] node1046;
	wire [3-1:0] node1049;
	wire [3-1:0] node1051;
	wire [3-1:0] node1054;
	wire [3-1:0] node1055;
	wire [3-1:0] node1056;
	wire [3-1:0] node1057;
	wire [3-1:0] node1059;
	wire [3-1:0] node1060;
	wire [3-1:0] node1062;
	wire [3-1:0] node1066;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1070;
	wire [3-1:0] node1073;
	wire [3-1:0] node1076;
	wire [3-1:0] node1077;
	wire [3-1:0] node1081;
	wire [3-1:0] node1082;
	wire [3-1:0] node1083;
	wire [3-1:0] node1085;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1092;
	wire [3-1:0] node1093;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1100;
	wire [3-1:0] node1101;
	wire [3-1:0] node1103;
	wire [3-1:0] node1106;
	wire [3-1:0] node1107;
	wire [3-1:0] node1110;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1116;
	wire [3-1:0] node1118;
	wire [3-1:0] node1121;
	wire [3-1:0] node1122;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1128;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1134;
	wire [3-1:0] node1138;
	wire [3-1:0] node1139;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1142;
	wire [3-1:0] node1146;
	wire [3-1:0] node1148;
	wire [3-1:0] node1149;
	wire [3-1:0] node1152;
	wire [3-1:0] node1155;
	wire [3-1:0] node1157;
	wire [3-1:0] node1160;
	wire [3-1:0] node1161;
	wire [3-1:0] node1162;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1167;
	wire [3-1:0] node1170;
	wire [3-1:0] node1173;
	wire [3-1:0] node1175;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1181;
	wire [3-1:0] node1183;

	assign outp = (inp[6]) ? node394 : node1;
		assign node1 = (inp[3]) ? node249 : node2;
			assign node2 = (inp[0]) ? node64 : node3;
				assign node3 = (inp[9]) ? node39 : node4;
					assign node4 = (inp[7]) ? node26 : node5;
						assign node5 = (inp[5]) ? node11 : node6;
							assign node6 = (inp[8]) ? 3'b000 : node7;
								assign node7 = (inp[10]) ? 3'b010 : 3'b000;
							assign node11 = (inp[10]) ? node19 : node12;
								assign node12 = (inp[8]) ? 3'b000 : node13;
									assign node13 = (inp[4]) ? 3'b010 : node14;
										assign node14 = (inp[11]) ? 3'b000 : 3'b010;
								assign node19 = (inp[8]) ? 3'b010 : node20;
									assign node20 = (inp[11]) ? node22 : 3'b100;
										assign node22 = (inp[4]) ? 3'b100 : 3'b110;
						assign node26 = (inp[8]) ? 3'b000 : node27;
							assign node27 = (inp[5]) ? node29 : 3'b000;
								assign node29 = (inp[4]) ? node33 : node30;
									assign node30 = (inp[10]) ? 3'b010 : 3'b000;
									assign node33 = (inp[11]) ? 3'b000 : node34;
										assign node34 = (inp[2]) ? 3'b010 : 3'b000;
					assign node39 = (inp[8]) ? 3'b000 : node40;
						assign node40 = (inp[5]) ? node42 : 3'b000;
							assign node42 = (inp[7]) ? node52 : node43;
								assign node43 = (inp[2]) ? 3'b000 : node44;
									assign node44 = (inp[4]) ? 3'b000 : node45;
										assign node45 = (inp[11]) ? 3'b000 : node46;
											assign node46 = (inp[10]) ? 3'b000 : 3'b010;
								assign node52 = (inp[10]) ? node60 : node53;
									assign node53 = (inp[2]) ? node55 : 3'b000;
										assign node55 = (inp[11]) ? 3'b000 : node56;
											assign node56 = (inp[1]) ? 3'b010 : 3'b000;
									assign node60 = (inp[4]) ? 3'b000 : 3'b010;
				assign node64 = (inp[4]) ? node164 : node65;
					assign node65 = (inp[9]) ? node125 : node66;
						assign node66 = (inp[7]) ? node92 : node67;
							assign node67 = (inp[8]) ? node77 : node68;
								assign node68 = (inp[5]) ? node74 : node69;
									assign node69 = (inp[10]) ? 3'b100 : node70;
										assign node70 = (inp[11]) ? 3'b010 : 3'b110;
									assign node74 = (inp[1]) ? 3'b100 : 3'b000;
								assign node77 = (inp[10]) ? node85 : node78;
									assign node78 = (inp[5]) ? node82 : node79;
										assign node79 = (inp[1]) ? 3'b110 : 3'b100;
										assign node82 = (inp[11]) ? 3'b010 : 3'b110;
									assign node85 = (inp[1]) ? node87 : 3'b000;
										assign node87 = (inp[11]) ? node89 : 3'b010;
											assign node89 = (inp[2]) ? 3'b010 : 3'b100;
							assign node92 = (inp[5]) ? node110 : node93;
								assign node93 = (inp[10]) ? node105 : node94;
									assign node94 = (inp[8]) ? node100 : node95;
										assign node95 = (inp[1]) ? 3'b001 : node96;
											assign node96 = (inp[11]) ? 3'b000 : 3'b001;
										assign node100 = (inp[1]) ? node102 : 3'b010;
											assign node102 = (inp[11]) ? 3'b000 : 3'b100;
									assign node105 = (inp[1]) ? node107 : 3'b100;
										assign node107 = (inp[11]) ? 3'b110 : 3'b000;
								assign node110 = (inp[1]) ? node118 : node111;
									assign node111 = (inp[8]) ? node115 : node112;
										assign node112 = (inp[11]) ? 3'b100 : 3'b000;
										assign node115 = (inp[11]) ? 3'b000 : 3'b100;
									assign node118 = (inp[8]) ? node122 : node119;
										assign node119 = (inp[10]) ? 3'b010 : 3'b110;
										assign node122 = (inp[10]) ? 3'b110 : 3'b001;
						assign node125 = (inp[7]) ? node141 : node126;
							assign node126 = (inp[10]) ? 3'b000 : node127;
								assign node127 = (inp[5]) ? node133 : node128;
									assign node128 = (inp[8]) ? 3'b100 : node129;
										assign node129 = (inp[1]) ? 3'b100 : 3'b000;
									assign node133 = (inp[2]) ? node135 : 3'b000;
										assign node135 = (inp[8]) ? node137 : 3'b000;
											assign node137 = (inp[1]) ? 3'b100 : 3'b000;
							assign node141 = (inp[5]) ? node155 : node142;
								assign node142 = (inp[10]) ? node152 : node143;
									assign node143 = (inp[1]) ? node147 : node144;
										assign node144 = (inp[8]) ? 3'b000 : 3'b010;
										assign node147 = (inp[8]) ? node149 : 3'b010;
											assign node149 = (inp[11]) ? 3'b010 : 3'b110;
									assign node152 = (inp[1]) ? 3'b100 : 3'b110;
								assign node155 = (inp[8]) ? node159 : node156;
									assign node156 = (inp[10]) ? 3'b000 : 3'b100;
									assign node159 = (inp[10]) ? node161 : 3'b010;
										assign node161 = (inp[1]) ? 3'b100 : 3'b110;
					assign node164 = (inp[10]) ? node222 : node165;
						assign node165 = (inp[9]) ? node199 : node166;
							assign node166 = (inp[7]) ? node182 : node167;
								assign node167 = (inp[5]) ? node175 : node168;
									assign node168 = (inp[1]) ? node172 : node169;
										assign node169 = (inp[8]) ? 3'b100 : 3'b110;
										assign node172 = (inp[8]) ? 3'b010 : 3'b100;
									assign node175 = (inp[8]) ? 3'b110 : node176;
										assign node176 = (inp[11]) ? 3'b000 : node177;
											assign node177 = (inp[2]) ? 3'b100 : 3'b000;
								assign node182 = (inp[1]) ? node194 : node183;
									assign node183 = (inp[5]) ? node189 : node184;
										assign node184 = (inp[8]) ? node186 : 3'b010;
											assign node186 = (inp[2]) ? 3'b000 : 3'b100;
										assign node189 = (inp[8]) ? node191 : 3'b100;
											assign node191 = (inp[2]) ? 3'b111 : 3'b001;
									assign node194 = (inp[11]) ? 3'b010 : node195;
										assign node195 = (inp[8]) ? 3'b110 : 3'b010;
							assign node199 = (inp[8]) ? node207 : node200;
								assign node200 = (inp[2]) ? node202 : 3'b000;
									assign node202 = (inp[7]) ? node204 : 3'b000;
										assign node204 = (inp[1]) ? 3'b000 : 3'b100;
								assign node207 = (inp[11]) ? node217 : node208;
									assign node208 = (inp[7]) ? node210 : 3'b000;
										assign node210 = (inp[5]) ? node214 : node211;
											assign node211 = (inp[2]) ? 3'b010 : 3'b110;
											assign node214 = (inp[2]) ? 3'b100 : 3'b010;
									assign node217 = (inp[5]) ? 3'b000 : node218;
										assign node218 = (inp[2]) ? 3'b100 : 3'b000;
						assign node222 = (inp[7]) ? node230 : node223;
							assign node223 = (inp[11]) ? 3'b000 : node224;
								assign node224 = (inp[8]) ? node226 : 3'b000;
									assign node226 = (inp[2]) ? 3'b100 : 3'b000;
							assign node230 = (inp[9]) ? node242 : node231;
								assign node231 = (inp[8]) ? node237 : node232;
									assign node232 = (inp[5]) ? 3'b000 : node233;
										assign node233 = (inp[1]) ? 3'b000 : 3'b010;
									assign node237 = (inp[1]) ? 3'b010 : node238;
										assign node238 = (inp[11]) ? 3'b110 : 3'b000;
								assign node242 = (inp[5]) ? 3'b000 : node243;
									assign node243 = (inp[2]) ? 3'b000 : node244;
										assign node244 = (inp[1]) ? 3'b000 : 3'b010;
			assign node249 = (inp[7]) ? node283 : node250;
				assign node250 = (inp[4]) ? 3'b000 : node251;
					assign node251 = (inp[9]) ? 3'b000 : node252;
						assign node252 = (inp[5]) ? 3'b000 : node253;
							assign node253 = (inp[11]) ? node271 : node254;
								assign node254 = (inp[1]) ? node262 : node255;
									assign node255 = (inp[10]) ? 3'b000 : node256;
										assign node256 = (inp[0]) ? node258 : 3'b000;
											assign node258 = (inp[8]) ? 3'b100 : 3'b000;
									assign node262 = (inp[0]) ? node266 : node263;
										assign node263 = (inp[8]) ? 3'b000 : 3'b100;
										assign node266 = (inp[8]) ? node268 : 3'b000;
											assign node268 = (inp[10]) ? 3'b000 : 3'b100;
								assign node271 = (inp[0]) ? 3'b000 : node272;
									assign node272 = (inp[10]) ? 3'b000 : node273;
										assign node273 = (inp[8]) ? 3'b000 : node274;
											assign node274 = (inp[2]) ? 3'b000 : 3'b100;
				assign node283 = (inp[8]) ? node321 : node284;
					assign node284 = (inp[9]) ? 3'b000 : node285;
						assign node285 = (inp[4]) ? node307 : node286;
							assign node286 = (inp[1]) ? node298 : node287;
								assign node287 = (inp[10]) ? 3'b000 : node288;
									assign node288 = (inp[2]) ? node294 : node289;
										assign node289 = (inp[11]) ? 3'b000 : node290;
											assign node290 = (inp[5]) ? 3'b000 : 3'b100;
										assign node294 = (inp[11]) ? 3'b000 : 3'b010;
								assign node298 = (inp[0]) ? node304 : node299;
									assign node299 = (inp[5]) ? node301 : 3'b010;
										assign node301 = (inp[10]) ? 3'b100 : 3'b110;
									assign node304 = (inp[2]) ? 3'b000 : 3'b100;
							assign node307 = (inp[10]) ? 3'b000 : node308;
								assign node308 = (inp[0]) ? node312 : node309;
									assign node309 = (inp[11]) ? 3'b000 : 3'b010;
									assign node312 = (inp[1]) ? 3'b000 : node313;
										assign node313 = (inp[5]) ? 3'b000 : node314;
											assign node314 = (inp[11]) ? 3'b000 : 3'b100;
					assign node321 = (inp[9]) ? node373 : node322;
						assign node322 = (inp[0]) ? node348 : node323;
							assign node323 = (inp[5]) ? node325 : 3'b100;
								assign node325 = (inp[1]) ? node337 : node326;
									assign node326 = (inp[4]) ? node332 : node327;
										assign node327 = (inp[10]) ? 3'b000 : node328;
											assign node328 = (inp[11]) ? 3'b100 : 3'b000;
										assign node332 = (inp[11]) ? 3'b100 : node333;
											assign node333 = (inp[10]) ? 3'b100 : 3'b000;
									assign node337 = (inp[4]) ? node343 : node338;
										assign node338 = (inp[11]) ? 3'b010 : node339;
											assign node339 = (inp[10]) ? 3'b110 : 3'b010;
										assign node343 = (inp[11]) ? 3'b100 : node344;
											assign node344 = (inp[10]) ? 3'b100 : 3'b010;
							assign node348 = (inp[10]) ? node366 : node349;
								assign node349 = (inp[5]) ? node359 : node350;
									assign node350 = (inp[4]) ? node356 : node351;
										assign node351 = (inp[11]) ? 3'b100 : node352;
											assign node352 = (inp[1]) ? 3'b010 : 3'b110;
										assign node356 = (inp[1]) ? 3'b000 : 3'b100;
									assign node359 = (inp[1]) ? node363 : node360;
										assign node360 = (inp[11]) ? 3'b000 : 3'b100;
										assign node363 = (inp[4]) ? 3'b000 : 3'b100;
								assign node366 = (inp[1]) ? node368 : 3'b000;
									assign node368 = (inp[4]) ? 3'b000 : node369;
										assign node369 = (inp[5]) ? 3'b000 : 3'b100;
						assign node373 = (inp[0]) ? node385 : node374;
							assign node374 = (inp[5]) ? 3'b000 : node375;
								assign node375 = (inp[1]) ? node379 : node376;
									assign node376 = (inp[10]) ? 3'b000 : 3'b100;
									assign node379 = (inp[2]) ? node381 : 3'b100;
										assign node381 = (inp[10]) ? 3'b100 : 3'b000;
							assign node385 = (inp[4]) ? 3'b000 : node386;
								assign node386 = (inp[10]) ? 3'b000 : node387;
									assign node387 = (inp[5]) ? 3'b000 : node388;
										assign node388 = (inp[11]) ? 3'b000 : 3'b010;
		assign node394 = (inp[3]) ? node722 : node395;
			assign node395 = (inp[0]) ? node495 : node396;
				assign node396 = (inp[7]) ? node406 : node397;
					assign node397 = (inp[8]) ? 3'b001 : node398;
						assign node398 = (inp[5]) ? node400 : 3'b001;
							assign node400 = (inp[10]) ? node402 : 3'b000;
								assign node402 = (inp[9]) ? 3'b000 : 3'b001;
					assign node406 = (inp[8]) ? node438 : node407;
						assign node407 = (inp[5]) ? 3'b000 : node408;
							assign node408 = (inp[9]) ? node416 : node409;
								assign node409 = (inp[2]) ? node411 : 3'b111;
									assign node411 = (inp[10]) ? node413 : 3'b111;
										assign node413 = (inp[1]) ? 3'b011 : 3'b111;
								assign node416 = (inp[2]) ? node428 : node417;
									assign node417 = (inp[1]) ? node423 : node418;
										assign node418 = (inp[4]) ? node420 : 3'b011;
											assign node420 = (inp[11]) ? 3'b011 : 3'b111;
										assign node423 = (inp[4]) ? node425 : 3'b011;
											assign node425 = (inp[10]) ? 3'b001 : 3'b011;
									assign node428 = (inp[4]) ? node430 : 3'b111;
										assign node430 = (inp[1]) ? node432 : 3'b011;
											assign node432 = (inp[11]) ? node434 : 3'b111;
												assign node434 = (inp[10]) ? 3'b001 : 3'b101;
						assign node438 = (inp[9]) ? node448 : node439;
							assign node439 = (inp[5]) ? node441 : 3'b111;
								assign node441 = (inp[10]) ? node443 : 3'b111;
									assign node443 = (inp[1]) ? node445 : 3'b111;
										assign node445 = (inp[4]) ? 3'b011 : 3'b111;
							assign node448 = (inp[4]) ? node466 : node449;
								assign node449 = (inp[2]) ? node457 : node450;
									assign node450 = (inp[11]) ? node452 : 3'b111;
										assign node452 = (inp[10]) ? node454 : 3'b111;
											assign node454 = (inp[1]) ? 3'b011 : 3'b111;
									assign node457 = (inp[10]) ? node461 : node458;
										assign node458 = (inp[11]) ? 3'b111 : 3'b011;
										assign node461 = (inp[1]) ? 3'b011 : node462;
											assign node462 = (inp[5]) ? 3'b111 : 3'b011;
								assign node466 = (inp[11]) ? node480 : node467;
									assign node467 = (inp[2]) ? node469 : 3'b011;
										assign node469 = (inp[1]) ? node475 : node470;
											assign node470 = (inp[5]) ? 3'b011 : node471;
												assign node471 = (inp[10]) ? 3'b011 : 3'b111;
											assign node475 = (inp[10]) ? 3'b101 : node476;
												assign node476 = (inp[5]) ? 3'b111 : 3'b011;
									assign node480 = (inp[10]) ? node488 : node481;
										assign node481 = (inp[1]) ? node485 : node482;
											assign node482 = (inp[5]) ? 3'b011 : 3'b111;
											assign node485 = (inp[5]) ? 3'b101 : 3'b001;
										assign node488 = (inp[2]) ? node490 : 3'b101;
											assign node490 = (inp[1]) ? node492 : 3'b101;
												assign node492 = (inp[5]) ? 3'b001 : 3'b101;
				assign node495 = (inp[10]) ? node619 : node496;
					assign node496 = (inp[4]) ? node546 : node497;
						assign node497 = (inp[5]) ? node521 : node498;
							assign node498 = (inp[8]) ? node514 : node499;
								assign node499 = (inp[11]) ? node505 : node500;
									assign node500 = (inp[7]) ? node502 : 3'b011;
										assign node502 = (inp[1]) ? 3'b101 : 3'b011;
									assign node505 = (inp[7]) ? node507 : 3'b111;
										assign node507 = (inp[9]) ? node511 : node508;
											assign node508 = (inp[2]) ? 3'b011 : 3'b111;
											assign node511 = (inp[1]) ? 3'b110 : 3'b011;
								assign node514 = (inp[7]) ? node516 : 3'b111;
									assign node516 = (inp[1]) ? node518 : 3'b111;
										assign node518 = (inp[11]) ? 3'b111 : 3'b011;
							assign node521 = (inp[8]) ? node533 : node522;
								assign node522 = (inp[7]) ? node526 : node523;
									assign node523 = (inp[11]) ? 3'b001 : 3'b101;
									assign node526 = (inp[9]) ? 3'b111 : node527;
										assign node527 = (inp[1]) ? 3'b011 : node528;
											assign node528 = (inp[11]) ? 3'b111 : 3'b011;
								assign node533 = (inp[11]) ? node539 : node534;
									assign node534 = (inp[7]) ? node536 : 3'b011;
										assign node536 = (inp[1]) ? 3'b101 : 3'b011;
									assign node539 = (inp[7]) ? node541 : 3'b111;
										assign node541 = (inp[9]) ? node543 : 3'b011;
											assign node543 = (inp[1]) ? 3'b110 : 3'b011;
						assign node546 = (inp[11]) ? node586 : node547;
							assign node547 = (inp[7]) ? node559 : node548;
								assign node548 = (inp[8]) ? node556 : node549;
									assign node549 = (inp[5]) ? node551 : 3'b001;
										assign node551 = (inp[2]) ? 3'b110 : node552;
											assign node552 = (inp[1]) ? 3'b100 : 3'b000;
									assign node556 = (inp[5]) ? 3'b001 : 3'b101;
								assign node559 = (inp[1]) ? node571 : node560;
									assign node560 = (inp[8]) ? node568 : node561;
										assign node561 = (inp[5]) ? node563 : 3'b111;
											assign node563 = (inp[9]) ? 3'b111 : node564;
												assign node564 = (inp[2]) ? 3'b001 : 3'b011;
										assign node568 = (inp[9]) ? 3'b011 : 3'b111;
									assign node571 = (inp[8]) ? node579 : node572;
										assign node572 = (inp[5]) ? node576 : node573;
											assign node573 = (inp[9]) ? 3'b001 : 3'b101;
											assign node576 = (inp[2]) ? 3'b101 : 3'b111;
										assign node579 = (inp[5]) ? node583 : node580;
											assign node580 = (inp[9]) ? 3'b001 : 3'b011;
											assign node583 = (inp[9]) ? 3'b001 : 3'b101;
							assign node586 = (inp[7]) ? node596 : node587;
								assign node587 = (inp[8]) ? node593 : node588;
									assign node588 = (inp[5]) ? node590 : 3'b011;
										assign node590 = (inp[2]) ? 3'b110 : 3'b010;
									assign node593 = (inp[5]) ? 3'b011 : 3'b111;
								assign node596 = (inp[9]) ? node608 : node597;
									assign node597 = (inp[5]) ? node603 : node598;
										assign node598 = (inp[1]) ? 3'b011 : node599;
											assign node599 = (inp[8]) ? 3'b111 : 3'b011;
										assign node603 = (inp[1]) ? 3'b101 : node604;
											assign node604 = (inp[8]) ? 3'b011 : 3'b101;
									assign node608 = (inp[1]) ? node614 : node609;
										assign node609 = (inp[8]) ? node611 : 3'b001;
											assign node611 = (inp[5]) ? 3'b001 : 3'b101;
										assign node614 = (inp[2]) ? 3'b000 : node615;
											assign node615 = (inp[8]) ? 3'b001 : 3'b101;
					assign node619 = (inp[7]) ? node647 : node620;
						assign node620 = (inp[11]) ? node632 : node621;
							assign node621 = (inp[8]) ? 3'b110 : node622;
								assign node622 = (inp[5]) ? node624 : 3'b110;
									assign node624 = (inp[4]) ? 3'b110 : node625;
										assign node625 = (inp[2]) ? node627 : 3'b100;
											assign node627 = (inp[1]) ? 3'b000 : 3'b100;
							assign node632 = (inp[4]) ? node642 : node633;
								assign node633 = (inp[8]) ? node639 : node634;
									assign node634 = (inp[5]) ? node636 : 3'b010;
										assign node636 = (inp[1]) ? 3'b000 : 3'b100;
									assign node639 = (inp[5]) ? 3'b010 : 3'b110;
								assign node642 = (inp[8]) ? 3'b100 : node643;
									assign node643 = (inp[5]) ? 3'b110 : 3'b100;
						assign node647 = (inp[5]) ? node685 : node648;
							assign node648 = (inp[1]) ? node666 : node649;
								assign node649 = (inp[9]) ? node659 : node650;
									assign node650 = (inp[4]) ? node652 : 3'b111;
										assign node652 = (inp[11]) ? node656 : node653;
											assign node653 = (inp[8]) ? 3'b111 : 3'b011;
											assign node656 = (inp[8]) ? 3'b011 : 3'b101;
									assign node659 = (inp[8]) ? node663 : node660;
										assign node660 = (inp[4]) ? 3'b001 : 3'b101;
										assign node663 = (inp[4]) ? 3'b001 : 3'b011;
								assign node666 = (inp[9]) ? node672 : node667;
									assign node667 = (inp[8]) ? 3'b101 : node668;
										assign node668 = (inp[4]) ? 3'b001 : 3'b011;
									assign node672 = (inp[8]) ? node678 : node673;
										assign node673 = (inp[4]) ? node675 : 3'b110;
											assign node675 = (inp[11]) ? 3'b010 : 3'b110;
										assign node678 = (inp[4]) ? node682 : node679;
											assign node679 = (inp[11]) ? 3'b001 : 3'b101;
											assign node682 = (inp[11]) ? 3'b110 : 3'b100;
							assign node685 = (inp[8]) ? node697 : node686;
								assign node686 = (inp[4]) ? node692 : node687;
									assign node687 = (inp[1]) ? node689 : 3'b110;
										assign node689 = (inp[9]) ? 3'b110 : 3'b010;
									assign node692 = (inp[1]) ? node694 : 3'b100;
										assign node694 = (inp[9]) ? 3'b100 : 3'b000;
								assign node697 = (inp[9]) ? node711 : node698;
									assign node698 = (inp[11]) ? node706 : node699;
										assign node699 = (inp[2]) ? node703 : node700;
											assign node700 = (inp[1]) ? 3'b001 : 3'b011;
											assign node703 = (inp[1]) ? 3'b011 : 3'b111;
										assign node706 = (inp[1]) ? node708 : 3'b101;
											assign node708 = (inp[4]) ? 3'b001 : 3'b101;
									assign node711 = (inp[4]) ? node715 : node712;
										assign node712 = (inp[1]) ? 3'b110 : 3'b101;
										assign node715 = (inp[2]) ? node717 : 3'b110;
											assign node717 = (inp[11]) ? node719 : 3'b110;
												assign node719 = (inp[1]) ? 3'b010 : 3'b110;
			assign node722 = (inp[7]) ? node912 : node723;
				assign node723 = (inp[9]) ? node845 : node724;
					assign node724 = (inp[10]) ? node796 : node725;
						assign node725 = (inp[11]) ? node765 : node726;
							assign node726 = (inp[4]) ? node744 : node727;
								assign node727 = (inp[2]) ? node739 : node728;
									assign node728 = (inp[0]) ? node734 : node729;
										assign node729 = (inp[8]) ? node731 : 3'b110;
											assign node731 = (inp[5]) ? 3'b110 : 3'b000;
										assign node734 = (inp[1]) ? node736 : 3'b010;
											assign node736 = (inp[8]) ? 3'b110 : 3'b010;
									assign node739 = (inp[8]) ? node741 : 3'b110;
										assign node741 = (inp[5]) ? 3'b110 : 3'b100;
								assign node744 = (inp[0]) ? node756 : node745;
									assign node745 = (inp[2]) ? node751 : node746;
										assign node746 = (inp[5]) ? node748 : 3'b110;
											assign node748 = (inp[8]) ? 3'b110 : 3'b000;
										assign node751 = (inp[5]) ? 3'b110 : node752;
											assign node752 = (inp[8]) ? 3'b000 : 3'b110;
									assign node756 = (inp[1]) ? node762 : node757;
										assign node757 = (inp[2]) ? node759 : 3'b010;
											assign node759 = (inp[8]) ? 3'b010 : 3'b100;
										assign node762 = (inp[5]) ? 3'b000 : 3'b100;
							assign node765 = (inp[0]) ? node775 : node766;
								assign node766 = (inp[8]) ? node772 : node767;
									assign node767 = (inp[5]) ? node769 : 3'b010;
										assign node769 = (inp[4]) ? 3'b010 : 3'b000;
									assign node772 = (inp[5]) ? 3'b010 : 3'b000;
								assign node775 = (inp[4]) ? node785 : node776;
									assign node776 = (inp[1]) ? node778 : 3'b010;
										assign node778 = (inp[5]) ? node782 : node779;
											assign node779 = (inp[8]) ? 3'b110 : 3'b010;
											assign node782 = (inp[8]) ? 3'b010 : 3'b100;
									assign node785 = (inp[2]) ? 3'b100 : node786;
										assign node786 = (inp[1]) ? node792 : node787;
											assign node787 = (inp[8]) ? node789 : 3'b010;
												assign node789 = (inp[5]) ? 3'b010 : 3'b000;
											assign node792 = (inp[8]) ? 3'b000 : 3'b100;
						assign node796 = (inp[0]) ? node814 : node797;
							assign node797 = (inp[5]) ? node803 : node798;
								assign node798 = (inp[8]) ? 3'b000 : node799;
									assign node799 = (inp[2]) ? 3'b010 : 3'b100;
								assign node803 = (inp[11]) ? node809 : node804;
									assign node804 = (inp[8]) ? 3'b010 : node805;
										assign node805 = (inp[1]) ? 3'b100 : 3'b110;
									assign node809 = (inp[8]) ? 3'b100 : node810;
										assign node810 = (inp[1]) ? 3'b100 : 3'b110;
							assign node814 = (inp[1]) ? node826 : node815;
								assign node815 = (inp[8]) ? node819 : node816;
									assign node816 = (inp[5]) ? 3'b000 : 3'b100;
									assign node819 = (inp[5]) ? 3'b100 : node820;
										assign node820 = (inp[11]) ? 3'b000 : node821;
											assign node821 = (inp[2]) ? 3'b100 : 3'b000;
								assign node826 = (inp[4]) ? node834 : node827;
									assign node827 = (inp[8]) ? node829 : 3'b100;
										assign node829 = (inp[11]) ? node831 : 3'b010;
											assign node831 = (inp[5]) ? 3'b000 : 3'b010;
									assign node834 = (inp[11]) ? 3'b000 : node835;
										assign node835 = (inp[8]) ? node837 : 3'b000;
											assign node837 = (inp[2]) ? node841 : node838;
												assign node838 = (inp[5]) ? 3'b100 : 3'b000;
												assign node841 = (inp[5]) ? 3'b000 : 3'b100;
					assign node845 = (inp[0]) ? node887 : node846;
						assign node846 = (inp[10]) ? node874 : node847;
							assign node847 = (inp[11]) ? node867 : node848;
								assign node848 = (inp[2]) ? node860 : node849;
									assign node849 = (inp[4]) ? node855 : node850;
										assign node850 = (inp[8]) ? node852 : 3'b000;
											assign node852 = (inp[5]) ? 3'b110 : 3'b000;
										assign node855 = (inp[5]) ? node857 : 3'b110;
											assign node857 = (inp[8]) ? 3'b110 : 3'b000;
									assign node860 = (inp[8]) ? node864 : node861;
										assign node861 = (inp[5]) ? 3'b000 : 3'b110;
										assign node864 = (inp[5]) ? 3'b110 : 3'b000;
								assign node867 = (inp[5]) ? node871 : node868;
									assign node868 = (inp[8]) ? 3'b000 : 3'b010;
									assign node871 = (inp[8]) ? 3'b010 : 3'b000;
							assign node874 = (inp[11]) ? node882 : node875;
								assign node875 = (inp[5]) ? node879 : node876;
									assign node876 = (inp[8]) ? 3'b000 : 3'b010;
									assign node879 = (inp[8]) ? 3'b010 : 3'b100;
								assign node882 = (inp[8]) ? node884 : 3'b100;
									assign node884 = (inp[5]) ? 3'b100 : 3'b000;
						assign node887 = (inp[5]) ? node903 : node888;
							assign node888 = (inp[8]) ? node890 : 3'b000;
								assign node890 = (inp[4]) ? node894 : node891;
									assign node891 = (inp[10]) ? 3'b000 : 3'b100;
									assign node894 = (inp[2]) ? node896 : 3'b000;
										assign node896 = (inp[11]) ? node900 : node897;
											assign node897 = (inp[10]) ? 3'b100 : 3'b000;
											assign node900 = (inp[10]) ? 3'b000 : 3'b100;
							assign node903 = (inp[8]) ? 3'b000 : node904;
								assign node904 = (inp[4]) ? 3'b000 : node905;
									assign node905 = (inp[11]) ? 3'b000 : node906;
										assign node906 = (inp[10]) ? 3'b000 : 3'b010;
				assign node912 = (inp[9]) ? node1054 : node913;
					assign node913 = (inp[0]) ? node981 : node914;
						assign node914 = (inp[4]) ? node936 : node915;
							assign node915 = (inp[1]) ? node925 : node916;
								assign node916 = (inp[10]) ? node918 : 3'b111;
									assign node918 = (inp[8]) ? node922 : node919;
										assign node919 = (inp[5]) ? 3'b110 : 3'b011;
										assign node922 = (inp[11]) ? 3'b011 : 3'b111;
								assign node925 = (inp[10]) ? node931 : node926;
									assign node926 = (inp[8]) ? 3'b011 : node927;
										assign node927 = (inp[11]) ? 3'b111 : 3'b001;
									assign node931 = (inp[8]) ? 3'b101 : node932;
										assign node932 = (inp[5]) ? 3'b111 : 3'b101;
							assign node936 = (inp[5]) ? node958 : node937;
								assign node937 = (inp[10]) ? node949 : node938;
									assign node938 = (inp[11]) ? node940 : 3'b011;
										assign node940 = (inp[2]) ? node946 : node941;
											assign node941 = (inp[8]) ? node943 : 3'b001;
												assign node943 = (inp[1]) ? 3'b111 : 3'b001;
											assign node946 = (inp[1]) ? 3'b111 : 3'b101;
									assign node949 = (inp[11]) ? node953 : node950;
										assign node950 = (inp[1]) ? 3'b110 : 3'b101;
										assign node953 = (inp[8]) ? node955 : 3'b001;
											assign node955 = (inp[1]) ? 3'b001 : 3'b101;
								assign node958 = (inp[8]) ? node966 : node959;
									assign node959 = (inp[11]) ? 3'b110 : node960;
										assign node960 = (inp[10]) ? 3'b110 : node961;
											assign node961 = (inp[1]) ? 3'b001 : 3'b000;
									assign node966 = (inp[1]) ? node972 : node967;
										assign node967 = (inp[2]) ? 3'b101 : node968;
											assign node968 = (inp[11]) ? 3'b001 : 3'b101;
										assign node972 = (inp[10]) ? node976 : node973;
											assign node973 = (inp[11]) ? 3'b001 : 3'b101;
											assign node976 = (inp[11]) ? 3'b110 : node977;
												assign node977 = (inp[2]) ? 3'b110 : 3'b001;
						assign node981 = (inp[1]) ? node1023 : node982;
							assign node982 = (inp[4]) ? node996 : node983;
								assign node983 = (inp[10]) ? node989 : node984;
									assign node984 = (inp[5]) ? 3'b101 : node985;
										assign node985 = (inp[8]) ? 3'b011 : 3'b101;
									assign node989 = (inp[8]) ? node993 : node990;
										assign node990 = (inp[5]) ? 3'b010 : 3'b001;
										assign node993 = (inp[5]) ? 3'b001 : 3'b101;
								assign node996 = (inp[11]) ? node1012 : node997;
									assign node997 = (inp[8]) ? node1003 : node998;
										assign node998 = (inp[5]) ? 3'b110 : node999;
											assign node999 = (inp[10]) ? 3'b110 : 3'b001;
										assign node1003 = (inp[5]) ? node1009 : node1004;
											assign node1004 = (inp[2]) ? 3'b001 : node1005;
												assign node1005 = (inp[10]) ? 3'b001 : 3'b101;
											assign node1009 = (inp[2]) ? 3'b110 : 3'b001;
									assign node1012 = (inp[8]) ? node1018 : node1013;
										assign node1013 = (inp[10]) ? 3'b010 : node1014;
											assign node1014 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1018 = (inp[5]) ? 3'b110 : node1019;
											assign node1019 = (inp[10]) ? 3'b110 : 3'b001;
							assign node1023 = (inp[10]) ? node1041 : node1024;
								assign node1024 = (inp[4]) ? node1034 : node1025;
									assign node1025 = (inp[8]) ? node1029 : node1026;
										assign node1026 = (inp[5]) ? 3'b110 : 3'b001;
										assign node1029 = (inp[11]) ? 3'b001 : node1030;
											assign node1030 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1034 = (inp[8]) ? 3'b110 : node1035;
										assign node1035 = (inp[5]) ? node1037 : 3'b010;
											assign node1037 = (inp[2]) ? 3'b100 : 3'b010;
								assign node1041 = (inp[4]) ? node1043 : 3'b110;
									assign node1043 = (inp[8]) ? node1049 : node1044;
										assign node1044 = (inp[5]) ? node1046 : 3'b100;
											assign node1046 = (inp[2]) ? 3'b000 : 3'b100;
										assign node1049 = (inp[5]) ? node1051 : 3'b010;
											assign node1051 = (inp[11]) ? 3'b100 : 3'b110;
					assign node1054 = (inp[0]) ? node1126 : node1055;
						assign node1055 = (inp[4]) ? node1081 : node1056;
							assign node1056 = (inp[10]) ? node1066 : node1057;
								assign node1057 = (inp[1]) ? node1059 : 3'b101;
									assign node1059 = (inp[8]) ? 3'b001 : node1060;
										assign node1060 = (inp[5]) ? node1062 : 3'b001;
											assign node1062 = (inp[11]) ? 3'b110 : 3'b000;
								assign node1066 = (inp[5]) ? node1076 : node1067;
									assign node1067 = (inp[1]) ? node1073 : node1068;
										assign node1068 = (inp[8]) ? node1070 : 3'b001;
											assign node1070 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1073 = (inp[8]) ? 3'b001 : 3'b110;
									assign node1076 = (inp[11]) ? 3'b110 : node1077;
										assign node1077 = (inp[1]) ? 3'b110 : 3'b001;
							assign node1081 = (inp[10]) ? node1097 : node1082;
								assign node1082 = (inp[1]) ? node1088 : node1083;
									assign node1083 = (inp[8]) ? node1085 : 3'b110;
										assign node1085 = (inp[11]) ? 3'b000 : 3'b001;
									assign node1088 = (inp[8]) ? node1092 : node1089;
										assign node1089 = (inp[5]) ? 3'b000 : 3'b010;
										assign node1092 = (inp[2]) ? 3'b010 : node1093;
											assign node1093 = (inp[11]) ? 3'b010 : 3'b110;
								assign node1097 = (inp[1]) ? node1113 : node1098;
									assign node1098 = (inp[11]) ? node1100 : 3'b110;
										assign node1100 = (inp[2]) ? node1106 : node1101;
											assign node1101 = (inp[5]) ? node1103 : 3'b110;
												assign node1103 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1106 = (inp[5]) ? node1110 : node1107;
												assign node1107 = (inp[8]) ? 3'b110 : 3'b010;
												assign node1110 = (inp[8]) ? 3'b010 : 3'b110;
									assign node1113 = (inp[11]) ? node1121 : node1114;
										assign node1114 = (inp[8]) ? node1116 : 3'b110;
											assign node1116 = (inp[5]) ? node1118 : 3'b010;
												assign node1118 = (inp[2]) ? 3'b110 : 3'b010;
										assign node1121 = (inp[8]) ? 3'b100 : node1122;
											assign node1122 = (inp[5]) ? 3'b110 : 3'b100;
						assign node1126 = (inp[8]) ? node1138 : node1127;
							assign node1127 = (inp[5]) ? 3'b000 : node1128;
								assign node1128 = (inp[2]) ? node1130 : 3'b000;
									assign node1130 = (inp[1]) ? node1134 : node1131;
										assign node1131 = (inp[4]) ? 3'b100 : 3'b110;
										assign node1134 = (inp[4]) ? 3'b000 : 3'b100;
							assign node1138 = (inp[4]) ? node1160 : node1139;
								assign node1139 = (inp[11]) ? node1155 : node1140;
									assign node1140 = (inp[2]) ? node1146 : node1141;
										assign node1141 = (inp[10]) ? 3'b010 : node1142;
											assign node1142 = (inp[5]) ? 3'b110 : 3'b001;
										assign node1146 = (inp[10]) ? node1148 : 3'b110;
											assign node1148 = (inp[5]) ? node1152 : node1149;
												assign node1149 = (inp[1]) ? 3'b010 : 3'b110;
												assign node1152 = (inp[1]) ? 3'b100 : 3'b010;
									assign node1155 = (inp[1]) ? node1157 : 3'b110;
										assign node1157 = (inp[10]) ? 3'b100 : 3'b010;
								assign node1160 = (inp[1]) ? node1178 : node1161;
									assign node1161 = (inp[10]) ? node1173 : node1162;
										assign node1162 = (inp[5]) ? node1170 : node1163;
											assign node1163 = (inp[11]) ? node1167 : node1164;
												assign node1164 = (inp[2]) ? 3'b010 : 3'b110;
												assign node1167 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1170 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1173 = (inp[11]) ? node1175 : 3'b100;
											assign node1175 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1178 = (inp[10]) ? 3'b000 : node1179;
										assign node1179 = (inp[5]) ? node1181 : 3'b100;
											assign node1181 = (inp[2]) ? node1183 : 3'b000;
												assign node1183 = (inp[11]) ? 3'b000 : 3'b100;

endmodule