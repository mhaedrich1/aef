module dtc_split25_bm73 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node196;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node232;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node240;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node272;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node289;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node303;
	wire [3-1:0] node305;
	wire [3-1:0] node307;
	wire [3-1:0] node309;
	wire [3-1:0] node312;
	wire [3-1:0] node314;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node337;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node344;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node359;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node370;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node379;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node389;
	wire [3-1:0] node392;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node403;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node410;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node419;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node427;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node439;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node446;
	wire [3-1:0] node448;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node463;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node480;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node486;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node493;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node509;
	wire [3-1:0] node510;
	wire [3-1:0] node513;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node523;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node538;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node550;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node557;
	wire [3-1:0] node560;
	wire [3-1:0] node562;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node570;
	wire [3-1:0] node572;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node599;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node622;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node640;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node648;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node668;
	wire [3-1:0] node672;
	wire [3-1:0] node673;

	assign outp = (inp[9]) ? node250 : node1;
		assign node1 = (inp[3]) ? node183 : node2;
			assign node2 = (inp[6]) ? node110 : node3;
				assign node3 = (inp[10]) ? node61 : node4;
					assign node4 = (inp[4]) ? node32 : node5;
						assign node5 = (inp[7]) ? node19 : node6;
							assign node6 = (inp[11]) ? node12 : node7;
								assign node7 = (inp[5]) ? 3'b110 : node8;
									assign node8 = (inp[8]) ? 3'b001 : 3'b101;
								assign node12 = (inp[5]) ? node16 : node13;
									assign node13 = (inp[8]) ? 3'b101 : 3'b011;
									assign node16 = (inp[8]) ? 3'b001 : 3'b101;
							assign node19 = (inp[8]) ? node27 : node20;
								assign node20 = (inp[11]) ? node24 : node21;
									assign node21 = (inp[5]) ? 3'b010 : 3'b110;
									assign node24 = (inp[0]) ? 3'b001 : 3'b110;
								assign node27 = (inp[11]) ? node29 : 3'b010;
									assign node29 = (inp[1]) ? 3'b110 : 3'b010;
						assign node32 = (inp[7]) ? node48 : node33;
							assign node33 = (inp[8]) ? node41 : node34;
								assign node34 = (inp[0]) ? 3'b110 : node35;
									assign node35 = (inp[1]) ? 3'b110 : node36;
										assign node36 = (inp[11]) ? 3'b110 : 3'b010;
								assign node41 = (inp[5]) ? node45 : node42;
									assign node42 = (inp[11]) ? 3'b110 : 3'b010;
									assign node45 = (inp[11]) ? 3'b010 : 3'b100;
							assign node48 = (inp[8]) ? node56 : node49;
								assign node49 = (inp[11]) ? node53 : node50;
									assign node50 = (inp[1]) ? 3'b000 : 3'b100;
									assign node53 = (inp[5]) ? 3'b100 : 3'b010;
								assign node56 = (inp[11]) ? node58 : 3'b000;
									assign node58 = (inp[5]) ? 3'b000 : 3'b100;
					assign node61 = (inp[4]) ? node87 : node62;
						assign node62 = (inp[7]) ? node76 : node63;
							assign node63 = (inp[11]) ? node71 : node64;
								assign node64 = (inp[2]) ? node68 : node65;
									assign node65 = (inp[5]) ? 3'b101 : 3'b011;
									assign node68 = (inp[5]) ? 3'b011 : 3'b111;
								assign node71 = (inp[8]) ? node73 : 3'b111;
									assign node73 = (inp[5]) ? 3'b011 : 3'b111;
							assign node76 = (inp[5]) ? node82 : node77;
								assign node77 = (inp[11]) ? 3'b011 : node78;
									assign node78 = (inp[8]) ? 3'b001 : 3'b101;
								assign node82 = (inp[1]) ? 3'b001 : node83;
									assign node83 = (inp[8]) ? 3'b001 : 3'b101;
						assign node87 = (inp[7]) ? node101 : node88;
							assign node88 = (inp[8]) ? node94 : node89;
								assign node89 = (inp[5]) ? node91 : 3'b011;
									assign node91 = (inp[0]) ? 3'b001 : 3'b101;
								assign node94 = (inp[5]) ? node98 : node95;
									assign node95 = (inp[11]) ? 3'b101 : 3'b001;
									assign node98 = (inp[11]) ? 3'b001 : 3'b110;
							assign node101 = (inp[8]) ? node107 : node102;
								assign node102 = (inp[5]) ? node104 : 3'b001;
									assign node104 = (inp[11]) ? 3'b110 : 3'b010;
								assign node107 = (inp[11]) ? 3'b110 : 3'b100;
				assign node110 = (inp[10]) ? node130 : node111;
					assign node111 = (inp[4]) ? 3'b000 : node112;
						assign node112 = (inp[7]) ? 3'b000 : node113;
							assign node113 = (inp[11]) ? node121 : node114;
								assign node114 = (inp[2]) ? node116 : 3'b000;
									assign node116 = (inp[8]) ? 3'b000 : node117;
										assign node117 = (inp[5]) ? 3'b000 : 3'b100;
								assign node121 = (inp[8]) ? node125 : node122;
									assign node122 = (inp[5]) ? 3'b100 : 3'b010;
									assign node125 = (inp[5]) ? 3'b000 : 3'b100;
					assign node130 = (inp[7]) ? node160 : node131;
						assign node131 = (inp[4]) ? node147 : node132;
							assign node132 = (inp[8]) ? node140 : node133;
								assign node133 = (inp[5]) ? node137 : node134;
									assign node134 = (inp[11]) ? 3'b001 : 3'b110;
									assign node137 = (inp[11]) ? 3'b110 : 3'b010;
								assign node140 = (inp[5]) ? node144 : node141;
									assign node141 = (inp[11]) ? 3'b110 : 3'b010;
									assign node144 = (inp[11]) ? 3'b010 : 3'b100;
							assign node147 = (inp[8]) ? node155 : node148;
								assign node148 = (inp[11]) ? node152 : node149;
									assign node149 = (inp[5]) ? 3'b000 : 3'b100;
									assign node152 = (inp[5]) ? 3'b100 : 3'b010;
								assign node155 = (inp[5]) ? 3'b000 : node156;
									assign node156 = (inp[11]) ? 3'b100 : 3'b000;
						assign node160 = (inp[4]) ? 3'b000 : node161;
							assign node161 = (inp[5]) ? node175 : node162;
								assign node162 = (inp[1]) ? node168 : node163;
									assign node163 = (inp[2]) ? node165 : 3'b100;
										assign node165 = (inp[11]) ? 3'b000 : 3'b100;
									assign node168 = (inp[11]) ? node172 : node169;
										assign node169 = (inp[8]) ? 3'b000 : 3'b100;
										assign node172 = (inp[8]) ? 3'b100 : 3'b010;
								assign node175 = (inp[11]) ? node177 : 3'b000;
									assign node177 = (inp[1]) ? 3'b100 : node178;
										assign node178 = (inp[8]) ? 3'b000 : 3'b010;
			assign node183 = (inp[6]) ? 3'b000 : node184;
				assign node184 = (inp[7]) ? node232 : node185;
					assign node185 = (inp[10]) ? node201 : node186;
						assign node186 = (inp[4]) ? 3'b000 : node187;
							assign node187 = (inp[11]) ? node193 : node188;
								assign node188 = (inp[8]) ? 3'b000 : node189;
									assign node189 = (inp[5]) ? 3'b000 : 3'b100;
								assign node193 = (inp[0]) ? 3'b100 : node194;
									assign node194 = (inp[2]) ? node196 : 3'b100;
										assign node196 = (inp[5]) ? 3'b000 : 3'b010;
						assign node201 = (inp[4]) ? node219 : node202;
							assign node202 = (inp[11]) ? node212 : node203;
								assign node203 = (inp[2]) ? node209 : node204;
									assign node204 = (inp[8]) ? 3'b010 : node205;
										assign node205 = (inp[5]) ? 3'b010 : 3'b110;
									assign node209 = (inp[8]) ? 3'b100 : 3'b110;
								assign node212 = (inp[8]) ? node216 : node213;
									assign node213 = (inp[5]) ? 3'b110 : 3'b001;
									assign node216 = (inp[5]) ? 3'b010 : 3'b110;
							assign node219 = (inp[11]) ? node225 : node220;
								assign node220 = (inp[5]) ? 3'b000 : node221;
									assign node221 = (inp[2]) ? 3'b000 : 3'b100;
								assign node225 = (inp[0]) ? 3'b100 : node226;
									assign node226 = (inp[8]) ? 3'b100 : node227;
										assign node227 = (inp[5]) ? 3'b100 : 3'b010;
					assign node232 = (inp[10]) ? node234 : 3'b000;
						assign node234 = (inp[4]) ? 3'b000 : node235;
							assign node235 = (inp[5]) ? node243 : node236;
								assign node236 = (inp[11]) ? node240 : node237;
									assign node237 = (inp[8]) ? 3'b000 : 3'b100;
									assign node240 = (inp[8]) ? 3'b100 : 3'b010;
								assign node243 = (inp[11]) ? node245 : 3'b000;
									assign node245 = (inp[8]) ? 3'b000 : 3'b100;
		assign node250 = (inp[3]) ? node466 : node251;
			assign node251 = (inp[6]) ? node329 : node252;
				assign node252 = (inp[10]) ? node300 : node253;
					assign node253 = (inp[4]) ? node265 : node254;
						assign node254 = (inp[7]) ? node256 : 3'b111;
							assign node256 = (inp[8]) ? node262 : node257;
								assign node257 = (inp[5]) ? node259 : 3'b111;
									assign node259 = (inp[11]) ? 3'b111 : 3'b011;
								assign node262 = (inp[11]) ? 3'b011 : 3'b101;
						assign node265 = (inp[7]) ? node285 : node266;
							assign node266 = (inp[2]) ? node276 : node267;
								assign node267 = (inp[11]) ? 3'b011 : node268;
									assign node268 = (inp[8]) ? node272 : node269;
										assign node269 = (inp[5]) ? 3'b011 : 3'b111;
										assign node272 = (inp[5]) ? 3'b101 : 3'b011;
								assign node276 = (inp[11]) ? node280 : node277;
									assign node277 = (inp[5]) ? 3'b101 : 3'b011;
									assign node280 = (inp[8]) ? node282 : 3'b111;
										assign node282 = (inp[5]) ? 3'b011 : 3'b111;
							assign node285 = (inp[0]) ? node293 : node286;
								assign node286 = (inp[5]) ? 3'b110 : node287;
									assign node287 = (inp[2]) ? node289 : 3'b101;
										assign node289 = (inp[1]) ? 3'b001 : 3'b011;
								assign node293 = (inp[8]) ? node297 : node294;
									assign node294 = (inp[5]) ? 3'b101 : 3'b011;
									assign node297 = (inp[5]) ? 3'b001 : 3'b101;
					assign node300 = (inp[0]) ? node312 : node301;
						assign node301 = (inp[1]) ? node303 : 3'b111;
							assign node303 = (inp[7]) ? node305 : 3'b111;
								assign node305 = (inp[5]) ? node307 : 3'b111;
									assign node307 = (inp[8]) ? node309 : 3'b111;
										assign node309 = (inp[11]) ? 3'b111 : 3'b101;
						assign node312 = (inp[7]) ? node314 : 3'b111;
							assign node314 = (inp[4]) ? node316 : 3'b111;
								assign node316 = (inp[11]) ? node324 : node317;
									assign node317 = (inp[1]) ? node321 : node318;
										assign node318 = (inp[5]) ? 3'b011 : 3'b011;
										assign node321 = (inp[5]) ? 3'b101 : 3'b011;
									assign node324 = (inp[1]) ? node326 : 3'b111;
										assign node326 = (inp[8]) ? 3'b011 : 3'b111;
				assign node329 = (inp[10]) ? node397 : node330;
					assign node330 = (inp[7]) ? node362 : node331;
						assign node331 = (inp[4]) ? node349 : node332;
							assign node332 = (inp[11]) ? node342 : node333;
								assign node333 = (inp[0]) ? node337 : node334;
									assign node334 = (inp[8]) ? 3'b001 : 3'b101;
									assign node337 = (inp[8]) ? node339 : 3'b001;
										assign node339 = (inp[5]) ? 3'b110 : 3'b001;
								assign node342 = (inp[8]) ? node344 : 3'b011;
									assign node344 = (inp[5]) ? node346 : 3'b011;
										assign node346 = (inp[1]) ? 3'b001 : 3'b101;
							assign node349 = (inp[2]) ? node355 : node350;
								assign node350 = (inp[8]) ? 3'b010 : node351;
									assign node351 = (inp[1]) ? 3'b110 : 3'b001;
								assign node355 = (inp[8]) ? node359 : node356;
									assign node356 = (inp[5]) ? 3'b010 : 3'b110;
									assign node359 = (inp[0]) ? 3'b100 : 3'b110;
						assign node362 = (inp[4]) ? node382 : node363;
							assign node363 = (inp[0]) ? node373 : node364;
								assign node364 = (inp[5]) ? node370 : node365;
									assign node365 = (inp[11]) ? 3'b001 : node366;
										assign node366 = (inp[1]) ? 3'b010 : 3'b001;
									assign node370 = (inp[11]) ? 3'b110 : 3'b010;
								assign node373 = (inp[2]) ? node379 : node374;
									assign node374 = (inp[5]) ? 3'b010 : node375;
										assign node375 = (inp[11]) ? 3'b110 : 3'b010;
									assign node379 = (inp[11]) ? 3'b110 : 3'b100;
							assign node382 = (inp[11]) ? node392 : node383;
								assign node383 = (inp[1]) ? node387 : node384;
									assign node384 = (inp[8]) ? 3'b000 : 3'b010;
									assign node387 = (inp[0]) ? node389 : 3'b100;
										assign node389 = (inp[5]) ? 3'b000 : 3'b100;
								assign node392 = (inp[5]) ? node394 : 3'b010;
									assign node394 = (inp[0]) ? 3'b100 : 3'b010;
					assign node397 = (inp[4]) ? node431 : node398;
						assign node398 = (inp[8]) ? node414 : node399;
							assign node399 = (inp[7]) ? node407 : node400;
								assign node400 = (inp[11]) ? 3'b111 : node401;
									assign node401 = (inp[0]) ? node403 : 3'b111;
										assign node403 = (inp[2]) ? 3'b011 : 3'b111;
								assign node407 = (inp[2]) ? 3'b101 : node408;
									assign node408 = (inp[1]) ? node410 : 3'b011;
										assign node410 = (inp[11]) ? 3'b111 : 3'b011;
							assign node414 = (inp[7]) ? node424 : node415;
								assign node415 = (inp[11]) ? node419 : node416;
									assign node416 = (inp[5]) ? 3'b101 : 3'b011;
									assign node419 = (inp[0]) ? node421 : 3'b111;
										assign node421 = (inp[5]) ? 3'b011 : 3'b111;
								assign node424 = (inp[1]) ? 3'b110 : node425;
									assign node425 = (inp[2]) ? node427 : 3'b101;
										assign node427 = (inp[11]) ? 3'b101 : 3'b110;
						assign node431 = (inp[7]) ? node451 : node432;
							assign node432 = (inp[0]) ? node442 : node433;
								assign node433 = (inp[1]) ? node439 : node434;
									assign node434 = (inp[8]) ? 3'b101 : node435;
										assign node435 = (inp[11]) ? 3'b011 : 3'b001;
									assign node439 = (inp[5]) ? 3'b001 : 3'b011;
								assign node442 = (inp[8]) ? node446 : node443;
									assign node443 = (inp[11]) ? 3'b011 : 3'b101;
									assign node446 = (inp[11]) ? node448 : 3'b001;
										assign node448 = (inp[1]) ? 3'b001 : 3'b101;
							assign node451 = (inp[11]) ? node457 : node452;
								assign node452 = (inp[8]) ? 3'b010 : node453;
									assign node453 = (inp[0]) ? 3'b010 : 3'b110;
								assign node457 = (inp[0]) ? node463 : node458;
									assign node458 = (inp[8]) ? 3'b001 : node459;
										assign node459 = (inp[5]) ? 3'b001 : 3'b101;
									assign node463 = (inp[8]) ? 3'b110 : 3'b101;
			assign node466 = (inp[6]) ? node592 : node467;
				assign node467 = (inp[10]) ? node527 : node468;
					assign node468 = (inp[4]) ? node496 : node469;
						assign node469 = (inp[7]) ? node483 : node470;
							assign node470 = (inp[5]) ? node478 : node471;
								assign node471 = (inp[8]) ? node475 : node472;
									assign node472 = (inp[11]) ? 3'b011 : 3'b101;
									assign node475 = (inp[2]) ? 3'b001 : 3'b101;
								assign node478 = (inp[8]) ? node480 : 3'b001;
									assign node480 = (inp[11]) ? 3'b001 : 3'b110;
							assign node483 = (inp[0]) ? node489 : node484;
								assign node484 = (inp[8]) ? node486 : 3'b110;
									assign node486 = (inp[1]) ? 3'b110 : 3'b010;
								assign node489 = (inp[5]) ? node493 : node490;
									assign node490 = (inp[11]) ? 3'b001 : 3'b110;
									assign node493 = (inp[11]) ? 3'b110 : 3'b010;
						assign node496 = (inp[7]) ? node516 : node497;
							assign node497 = (inp[0]) ? node509 : node498;
								assign node498 = (inp[2]) ? node504 : node499;
									assign node499 = (inp[5]) ? 3'b010 : node500;
										assign node500 = (inp[8]) ? 3'b010 : 3'b110;
									assign node504 = (inp[11]) ? 3'b010 : node505;
										assign node505 = (inp[8]) ? 3'b100 : 3'b010;
								assign node509 = (inp[1]) ? node513 : node510;
									assign node510 = (inp[11]) ? 3'b001 : 3'b110;
									assign node513 = (inp[2]) ? 3'b110 : 3'b100;
							assign node516 = (inp[8]) ? node520 : node517;
								assign node517 = (inp[11]) ? 3'b010 : 3'b100;
								assign node520 = (inp[0]) ? 3'b000 : node521;
									assign node521 = (inp[5]) ? node523 : 3'b100;
										assign node523 = (inp[2]) ? 3'b000 : 3'b000;
					assign node527 = (inp[11]) ? node565 : node528;
						assign node528 = (inp[4]) ? node546 : node529;
							assign node529 = (inp[7]) ? node535 : node530;
								assign node530 = (inp[5]) ? node532 : 3'b011;
									assign node532 = (inp[2]) ? 3'b111 : 3'b101;
								assign node535 = (inp[8]) ? node541 : node536;
									assign node536 = (inp[2]) ? node538 : 3'b101;
										assign node538 = (inp[5]) ? 3'b001 : 3'b101;
									assign node541 = (inp[1]) ? 3'b001 : node542;
										assign node542 = (inp[5]) ? 3'b000 : 3'b001;
							assign node546 = (inp[7]) ? node560 : node547;
								assign node547 = (inp[2]) ? node553 : node548;
									assign node548 = (inp[5]) ? node550 : 3'b011;
										assign node550 = (inp[8]) ? 3'b001 : 3'b101;
									assign node553 = (inp[5]) ? node557 : node554;
										assign node554 = (inp[1]) ? 3'b001 : 3'b101;
										assign node557 = (inp[1]) ? 3'b110 : 3'b101;
								assign node560 = (inp[2]) ? node562 : 3'b100;
									assign node562 = (inp[0]) ? 3'b010 : 3'b110;
						assign node565 = (inp[5]) ? node575 : node566;
							assign node566 = (inp[2]) ? node570 : node567;
								assign node567 = (inp[4]) ? 3'b001 : 3'b011;
								assign node570 = (inp[4]) ? node572 : 3'b111;
									assign node572 = (inp[8]) ? 3'b101 : 3'b011;
							assign node575 = (inp[4]) ? node587 : node576;
								assign node576 = (inp[7]) ? node580 : node577;
									assign node577 = (inp[2]) ? 3'b011 : 3'b111;
									assign node580 = (inp[0]) ? node584 : node581;
										assign node581 = (inp[8]) ? 3'b101 : 3'b011;
										assign node584 = (inp[8]) ? 3'b001 : 3'b101;
								assign node587 = (inp[8]) ? 3'b110 : node588;
									assign node588 = (inp[0]) ? 3'b101 : 3'b001;
				assign node592 = (inp[10]) ? node616 : node593;
					assign node593 = (inp[7]) ? 3'b000 : node594;
						assign node594 = (inp[4]) ? node608 : node595;
							assign node595 = (inp[11]) ? node603 : node596;
								assign node596 = (inp[8]) ? 3'b000 : node597;
									assign node597 = (inp[5]) ? node599 : 3'b100;
										assign node599 = (inp[0]) ? 3'b000 : 3'b100;
								assign node603 = (inp[0]) ? 3'b010 : node604;
									assign node604 = (inp[1]) ? 3'b110 : 3'b010;
							assign node608 = (inp[8]) ? 3'b000 : node609;
								assign node609 = (inp[2]) ? 3'b000 : node610;
									assign node610 = (inp[1]) ? 3'b000 : 3'b100;
					assign node616 = (inp[11]) ? node644 : node617;
						assign node617 = (inp[4]) ? node637 : node618;
							assign node618 = (inp[7]) ? node626 : node619;
								assign node619 = (inp[2]) ? 3'b110 : node620;
									assign node620 = (inp[1]) ? node622 : 3'b001;
										assign node622 = (inp[0]) ? 3'b100 : 3'b010;
								assign node626 = (inp[0]) ? node632 : node627;
									assign node627 = (inp[1]) ? 3'b100 : node628;
										assign node628 = (inp[2]) ? 3'b000 : 3'b100;
									assign node632 = (inp[1]) ? 3'b000 : node633;
										assign node633 = (inp[5]) ? 3'b000 : 3'b010;
							assign node637 = (inp[5]) ? 3'b000 : node638;
								assign node638 = (inp[1]) ? node640 : 3'b100;
									assign node640 = (inp[7]) ? 3'b000 : 3'b010;
						assign node644 = (inp[4]) ? node664 : node645;
							assign node645 = (inp[7]) ? node653 : node646;
								assign node646 = (inp[8]) ? node648 : 3'b001;
									assign node648 = (inp[2]) ? node650 : 3'b110;
										assign node650 = (inp[0]) ? 3'b010 : 3'b110;
								assign node653 = (inp[8]) ? node659 : node654;
									assign node654 = (inp[5]) ? 3'b010 : node655;
										assign node655 = (inp[1]) ? 3'b010 : 3'b110;
									assign node659 = (inp[5]) ? 3'b100 : node660;
										assign node660 = (inp[0]) ? 3'b000 : 3'b010;
							assign node664 = (inp[7]) ? node672 : node665;
								assign node665 = (inp[8]) ? 3'b100 : node666;
									assign node666 = (inp[1]) ? node668 : 3'b010;
										assign node668 = (inp[5]) ? 3'b100 : 3'b110;
								assign node672 = (inp[8]) ? 3'b000 : node673;
									assign node673 = (inp[5]) ? 3'b000 : 3'b100;

endmodule