module dtc_split33_bm37 (
	input  wire [8-1:0] inp,
	output wire [63-1:0] outp
);

	wire [63-1:0] node1;
	wire [63-1:0] node2;
	wire [63-1:0] node3;
	wire [63-1:0] node4;
	wire [63-1:0] node5;
	wire [63-1:0] node7;
	wire [63-1:0] node11;
	wire [63-1:0] node13;
	wire [63-1:0] node16;
	wire [63-1:0] node17;
	wire [63-1:0] node20;
	wire [63-1:0] node21;
	wire [63-1:0] node24;
	wire [63-1:0] node26;
	wire [63-1:0] node27;
	wire [63-1:0] node31;
	wire [63-1:0] node32;
	wire [63-1:0] node33;
	wire [63-1:0] node34;
	wire [63-1:0] node36;
	wire [63-1:0] node40;
	wire [63-1:0] node43;
	wire [63-1:0] node44;
	wire [63-1:0] node45;
	wire [63-1:0] node46;
	wire [63-1:0] node49;
	wire [63-1:0] node52;
	wire [63-1:0] node55;
	wire [63-1:0] node57;
	wire [63-1:0] node60;
	wire [63-1:0] node61;
	wire [63-1:0] node62;
	wire [63-1:0] node63;
	wire [63-1:0] node66;
	wire [63-1:0] node69;
	wire [63-1:0] node70;
	wire [63-1:0] node71;
	wire [63-1:0] node75;
	wire [63-1:0] node76;
	wire [63-1:0] node78;
	wire [63-1:0] node82;
	wire [63-1:0] node83;
	wire [63-1:0] node84;
	wire [63-1:0] node85;
	wire [63-1:0] node87;
	wire [63-1:0] node90;
	wire [63-1:0] node92;
	wire [63-1:0] node95;
	wire [63-1:0] node96;
	wire [63-1:0] node97;
	wire [63-1:0] node101;
	wire [63-1:0] node104;
	wire [63-1:0] node105;
	wire [63-1:0] node106;
	wire [63-1:0] node110;
	wire [63-1:0] node111;
	wire [63-1:0] node114;
	wire [63-1:0] node115;

	assign outp = (inp[7]) ? node60 : node1;
		assign node1 = (inp[6]) ? node31 : node2;
			assign node2 = (inp[1]) ? node16 : node3;
				assign node3 = (inp[3]) ? node11 : node4;
					assign node4 = (inp[2]) ? 63'b100111101001100000110001101110110010010101011101001101001010101 : node5;
						assign node5 = (inp[0]) ? node7 : 63'b100111101001100000110001101110110010010101001100001101001010101;
							assign node7 = (inp[4]) ? 63'b100111101001100000110001101110110010010101001101001101001010101 : 63'b100111101001100000110001101110110010010101001100001101001010101;
					assign node11 = (inp[2]) ? node13 : 63'b100110101001100000110001101110110011010101001100000101001010101;
						assign node13 = (inp[5]) ? 63'b100111101001000000110001101110110011000110001100101001001010101 : 63'b100110101001100000110001101110110011010101011100000101001010101;
				assign node16 = (inp[2]) ? node20 : node17;
					assign node17 = (inp[3]) ? 63'b100001101001100000010001101110010010010101001100101101000010101 : 63'b100111101001100000010001101110010010010101001100101101000000101;
					assign node20 = (inp[0]) ? node24 : node21;
						assign node21 = (inp[4]) ? 63'b110111100001000000110001101100110011010101001100111101001010101 : 63'b101110100001100000110001101110110011010101001100101101001010100;
						assign node24 = (inp[4]) ? node26 : 63'b100111101001000000110001101110110011010100001100101101001110101;
							assign node26 = (inp[3]) ? 63'b100001101001100000110001101110010010010101011101101101000010101 : node27;
								assign node27 = (inp[5]) ? 63'b100111101001100000110001101110010010010101011101101101000000101 : 63'b100111101001100000110001101110010010010101011100101101000000101;
			assign node31 = (inp[2]) ? node43 : node32;
				assign node32 = (inp[3]) ? node40 : node33;
					assign node33 = (inp[1]) ? 63'b100110101001100000110001101110110011010101000100001101001010001 : node34;
						assign node34 = (inp[0]) ? node36 : 63'b100110101001100000110001101110110001010101000100101101001010000;
							assign node36 = (inp[5]) ? 63'b100110101001100000110001101110110001010101000101101101001010000 : 63'b100110101001100000110001101110110001010101000100101101001010000;
					assign node40 = (inp[1]) ? 63'b100110101001100000110001101110100011010101001100100101001010100 : 63'b100110101001100000110001101110110011010001001100001101001010101;
				assign node43 = (inp[5]) ? node55 : node44;
					assign node44 = (inp[4]) ? node52 : node45;
						assign node45 = (inp[3]) ? node49 : node46;
							assign node46 = (inp[0]) ? 63'b100111101001100000110001101110110011010101001100101101001010101 : 63'b100111101001100000111001101110110011010001001100100101001010100;
							assign node49 = (inp[1]) ? 63'b100111101001100000110011101110110011010101001100001101001010101 : 63'b100111101001100000110001101110110011010101001100101101011010100;
						assign node52 = (inp[3]) ? 63'b100111001001100000110001101110110011010001001100101101001000101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
					assign node55 = (inp[4]) ? node57 : 63'b100111101001100100110001101110110011010101001100101101001010101;
						assign node57 = (inp[3]) ? 63'b100111101001100000110101101110110011010101001100101101001010101 : 63'b100111101001100001110001101110110011010101001100101101001010101;
		assign node60 = (inp[2]) ? node82 : node61;
			assign node61 = (inp[6]) ? node69 : node62;
				assign node62 = (inp[3]) ? node66 : node63;
					assign node63 = (inp[1]) ? 63'b100111101001100000110001101110110011010101001100101101000010101 : 63'b100111101001100000110001101110110011010101001000101101001000101;
					assign node66 = (inp[4]) ? 63'b000111101001001000110001101010110011000101001100101101001010101 : 63'b100111101000000000110001100000110011010101001100101100001010101;
				assign node69 = (inp[3]) ? node75 : node70;
					assign node70 = (inp[1]) ? 63'b100111101001100000110001001110110011010101001100101101000010101 : node71;
						assign node71 = (inp[4]) ? 63'b100111101001000000110001101000110111010101001101101100001010101 : 63'b100111101000000000110001100000110011010101001100101100001010101;
					assign node75 = (inp[1]) ? 63'b100111101001000000110000100100110011010101101100101101001010101 : node76;
						assign node76 = (inp[4]) ? node78 : 63'b100111101011100000100001101110110010010101001100101101000010101;
							assign node78 = (inp[5]) ? 63'b100111101001100000100001101110110010010101001101101101000010101 : 63'b100111101001100000100001101110110010010101001100101101000010101;
			assign node82 = (inp[4]) ? node104 : node83;
				assign node83 = (inp[5]) ? node95 : node84;
					assign node84 = (inp[6]) ? node90 : node85;
						assign node85 = (inp[3]) ? node87 : 63'b100111101001100000110001101110110011010101001100101101001010101;
							assign node87 = (inp[1]) ? 63'b100111101001100000110001101110110011010101001100101101001010101 : 63'b100001101001100000110001101110110011010101001100101101001010101;
						assign node90 = (inp[1]) ? node92 : 63'b100111101011100000100001101110110011010101001100101101001010100;
							assign node92 = (inp[0]) ? 63'b100111101001100000110001101110110011010101001100101101001010101 : 63'b100111101001100000110001101110110011010001001100101101001010100;
					assign node95 = (inp[0]) ? node101 : node96;
						assign node96 = (inp[1]) ? 63'b100111101001100100110001101110110011010101001100101101001010101 : node97;
							assign node97 = (inp[3]) ? 63'b100111101011100100110001101110110011010101001100101101001010101 : 63'b100111101001100100110001101110110011010101001100101101001010101;
						assign node101 = (inp[3]) ? 63'b100111101011000000110001101110110011000110001100101001001010101 : 63'b100111101001000000110001101110110011010100001100101101001110101;
				assign node104 = (inp[0]) ? node110 : node105;
					assign node105 = (inp[1]) ? 63'b100111101001000000110001101000110011010101001100101100101010101 : node106;
						assign node106 = (inp[3]) ? 63'b100101101001110000110001101110110011010101001100101101001010101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
					assign node110 = (inp[1]) ? node114 : node111;
						assign node111 = (inp[5]) ? 63'b100111101001100000110001001110111010010101011101101101000010101 : 63'b100111101001100000110001001110111010010101011100101101000010101;
						assign node114 = (inp[3]) ? 63'b100111101001100000110001101110110011010101011101101101001010101 : node115;
							assign node115 = (inp[5]) ? 63'b100111101001100000110001001110110011010101011101101101000010101 : 63'b100111101001100000110001101110110011010101011100101101000010101;

endmodule