module dtc_split66_bm86 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node160;
	wire [3-1:0] node162;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node197;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node251;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node282;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node296;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node314;
	wire [3-1:0] node317;
	wire [3-1:0] node319;
	wire [3-1:0] node322;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node332;
	wire [3-1:0] node334;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node342;
	wire [3-1:0] node344;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node351;
	wire [3-1:0] node353;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node382;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node389;
	wire [3-1:0] node392;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node402;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node410;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node432;
	wire [3-1:0] node434;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node440;

	assign outp = (inp[3]) ? node332 : node1;
		assign node1 = (inp[0]) ? node135 : node2;
			assign node2 = (inp[6]) ? 3'b000 : node3;
				assign node3 = (inp[4]) ? node103 : node4;
					assign node4 = (inp[9]) ? node58 : node5;
						assign node5 = (inp[7]) ? node39 : node6;
							assign node6 = (inp[1]) ? node14 : node7;
								assign node7 = (inp[2]) ? node9 : 3'b000;
									assign node9 = (inp[10]) ? node11 : 3'b000;
										assign node11 = (inp[5]) ? 3'b000 : 3'b100;
								assign node14 = (inp[5]) ? node28 : node15;
									assign node15 = (inp[2]) ? node21 : node16;
										assign node16 = (inp[10]) ? node18 : 3'b100;
											assign node18 = (inp[8]) ? 3'b110 : 3'b010;
										assign node21 = (inp[8]) ? node25 : node22;
											assign node22 = (inp[10]) ? 3'b110 : 3'b010;
											assign node25 = (inp[11]) ? 3'b000 : 3'b010;
									assign node28 = (inp[11]) ? node34 : node29;
										assign node29 = (inp[8]) ? 3'b000 : node30;
											assign node30 = (inp[2]) ? 3'b100 : 3'b000;
										assign node34 = (inp[10]) ? 3'b010 : node35;
											assign node35 = (inp[8]) ? 3'b000 : 3'b100;
							assign node39 = (inp[1]) ? node47 : node40;
								assign node40 = (inp[2]) ? node42 : 3'b010;
									assign node42 = (inp[11]) ? node44 : 3'b010;
										assign node44 = (inp[5]) ? 3'b010 : 3'b000;
								assign node47 = (inp[5]) ? node53 : node48;
									assign node48 = (inp[11]) ? node50 : 3'b110;
										assign node50 = (inp[2]) ? 3'b100 : 3'b110;
									assign node53 = (inp[2]) ? node55 : 3'b010;
										assign node55 = (inp[11]) ? 3'b110 : 3'b010;
						assign node58 = (inp[7]) ? node98 : node59;
							assign node59 = (inp[1]) ? node65 : node60;
								assign node60 = (inp[8]) ? node62 : 3'b110;
									assign node62 = (inp[11]) ? 3'b001 : 3'b110;
								assign node65 = (inp[5]) ? node79 : node66;
									assign node66 = (inp[2]) ? node74 : node67;
										assign node67 = (inp[10]) ? node69 : 3'b110;
											assign node69 = (inp[8]) ? 3'b101 : node70;
												assign node70 = (inp[11]) ? 3'b101 : 3'b001;
										assign node74 = (inp[10]) ? 3'b011 : node75;
											assign node75 = (inp[11]) ? 3'b101 : 3'b001;
									assign node79 = (inp[10]) ? node89 : node80;
										assign node80 = (inp[2]) ? node84 : node81;
											assign node81 = (inp[11]) ? 3'b010 : 3'b100;
											assign node84 = (inp[8]) ? 3'b110 : node85;
												assign node85 = (inp[11]) ? 3'b110 : 3'b010;
										assign node89 = (inp[2]) ? node93 : node90;
											assign node90 = (inp[11]) ? 3'b110 : 3'b000;
											assign node93 = (inp[11]) ? node95 : 3'b110;
												assign node95 = (inp[8]) ? 3'b101 : 3'b001;
							assign node98 = (inp[11]) ? node100 : 3'b011;
								assign node100 = (inp[2]) ? 3'b111 : 3'b011;
					assign node103 = (inp[9]) ? node105 : 3'b000;
						assign node105 = (inp[7]) ? 3'b000 : node106;
							assign node106 = (inp[10]) ? node116 : node107;
								assign node107 = (inp[8]) ? 3'b000 : node108;
									assign node108 = (inp[2]) ? node110 : 3'b000;
										assign node110 = (inp[1]) ? node112 : 3'b000;
											assign node112 = (inp[5]) ? 3'b000 : 3'b100;
								assign node116 = (inp[1]) ? node122 : node117;
									assign node117 = (inp[5]) ? 3'b000 : node118;
										assign node118 = (inp[8]) ? 3'b000 : 3'b010;
									assign node122 = (inp[5]) ? node130 : node123;
										assign node123 = (inp[2]) ? node127 : node124;
											assign node124 = (inp[11]) ? 3'b100 : 3'b000;
											assign node127 = (inp[8]) ? 3'b010 : 3'b110;
										assign node130 = (inp[2]) ? 3'b100 : 3'b000;
			assign node135 = (inp[6]) ? node327 : node136;
				assign node136 = (inp[4]) ? node202 : node137;
					assign node137 = (inp[7]) ? 3'b111 : node138;
						assign node138 = (inp[1]) ? node186 : node139;
							assign node139 = (inp[9]) ? node165 : node140;
								assign node140 = (inp[5]) ? node154 : node141;
									assign node141 = (inp[2]) ? node147 : node142;
										assign node142 = (inp[11]) ? node144 : 3'b001;
											assign node144 = (inp[10]) ? 3'b101 : 3'b001;
										assign node147 = (inp[11]) ? node151 : node148;
											assign node148 = (inp[8]) ? 3'b001 : 3'b101;
											assign node151 = (inp[8]) ? 3'b011 : 3'b111;
									assign node154 = (inp[11]) ? node160 : node155;
										assign node155 = (inp[8]) ? 3'b010 : node156;
											assign node156 = (inp[2]) ? 3'b110 : 3'b010;
										assign node160 = (inp[2]) ? node162 : 3'b110;
											assign node162 = (inp[8]) ? 3'b001 : 3'b101;
								assign node165 = (inp[5]) ? node177 : node166;
									assign node166 = (inp[10]) ? node172 : node167;
										assign node167 = (inp[2]) ? node169 : 3'b011;
											assign node169 = (inp[8]) ? 3'b111 : 3'b011;
										assign node172 = (inp[8]) ? 3'b111 : node173;
											assign node173 = (inp[2]) ? 3'b111 : 3'b011;
									assign node177 = (inp[10]) ? node181 : node178;
										assign node178 = (inp[2]) ? 3'b101 : 3'b011;
										assign node181 = (inp[2]) ? 3'b011 : node182;
											assign node182 = (inp[8]) ? 3'b011 : 3'b101;
							assign node186 = (inp[9]) ? node194 : node187;
								assign node187 = (inp[5]) ? node189 : 3'b111;
									assign node189 = (inp[11]) ? node191 : 3'b101;
										assign node191 = (inp[2]) ? 3'b111 : 3'b101;
								assign node194 = (inp[10]) ? 3'b111 : node195;
									assign node195 = (inp[5]) ? node197 : 3'b111;
										assign node197 = (inp[2]) ? 3'b111 : 3'b011;
					assign node202 = (inp[9]) ? node268 : node203;
						assign node203 = (inp[1]) ? node227 : node204;
							assign node204 = (inp[5]) ? node212 : node205;
								assign node205 = (inp[2]) ? node207 : 3'b100;
									assign node207 = (inp[10]) ? node209 : 3'b100;
										assign node209 = (inp[11]) ? 3'b100 : 3'b110;
								assign node212 = (inp[2]) ? node218 : node213;
									assign node213 = (inp[7]) ? 3'b100 : node214;
										assign node214 = (inp[10]) ? 3'b000 : 3'b100;
									assign node218 = (inp[11]) ? node222 : node219;
										assign node219 = (inp[10]) ? 3'b000 : 3'b100;
										assign node222 = (inp[7]) ? 3'b000 : node223;
											assign node223 = (inp[10]) ? 3'b100 : 3'b000;
							assign node227 = (inp[5]) ? node243 : node228;
								assign node228 = (inp[7]) ? 3'b110 : node229;
									assign node229 = (inp[2]) ? node239 : node230;
										assign node230 = (inp[10]) ? node232 : 3'b110;
											assign node232 = (inp[11]) ? node236 : node233;
												assign node233 = (inp[8]) ? 3'b110 : 3'b100;
												assign node236 = (inp[8]) ? 3'b010 : 3'b000;
										assign node239 = (inp[8]) ? 3'b100 : 3'b000;
								assign node243 = (inp[2]) ? node255 : node244;
									assign node244 = (inp[7]) ? 3'b100 : node245;
										assign node245 = (inp[8]) ? node251 : node246;
											assign node246 = (inp[11]) ? 3'b010 : node247;
												assign node247 = (inp[10]) ? 3'b100 : 3'b000;
											assign node251 = (inp[10]) ? 3'b110 : 3'b100;
									assign node255 = (inp[11]) ? node259 : node256;
										assign node256 = (inp[7]) ? 3'b100 : 3'b000;
										assign node259 = (inp[7]) ? 3'b010 : node260;
											assign node260 = (inp[10]) ? node264 : node261;
												assign node261 = (inp[8]) ? 3'b000 : 3'b010;
												assign node264 = (inp[8]) ? 3'b000 : 3'b100;
						assign node268 = (inp[5]) ? node300 : node269;
							assign node269 = (inp[7]) ? 3'b111 : node270;
								assign node270 = (inp[1]) ? node276 : node271;
									assign node271 = (inp[11]) ? node273 : 3'b110;
										assign node273 = (inp[2]) ? 3'b101 : 3'b110;
									assign node276 = (inp[8]) ? node290 : node277;
										assign node277 = (inp[2]) ? node285 : node278;
											assign node278 = (inp[10]) ? node282 : node279;
												assign node279 = (inp[11]) ? 3'b101 : 3'b111;
												assign node282 = (inp[11]) ? 3'b011 : 3'b101;
											assign node285 = (inp[10]) ? 3'b011 : node286;
												assign node286 = (inp[11]) ? 3'b011 : 3'b001;
										assign node290 = (inp[10]) ? node294 : node291;
											assign node291 = (inp[2]) ? 3'b111 : 3'b101;
											assign node294 = (inp[11]) ? node296 : 3'b111;
												assign node296 = (inp[2]) ? 3'b111 : 3'b011;
							assign node300 = (inp[7]) ? node322 : node301;
								assign node301 = (inp[10]) ? node311 : node302;
									assign node302 = (inp[2]) ? node306 : node303;
										assign node303 = (inp[1]) ? 3'b110 : 3'b100;
										assign node306 = (inp[1]) ? 3'b001 : node307;
											assign node307 = (inp[8]) ? 3'b110 : 3'b100;
									assign node311 = (inp[1]) ? node317 : node312;
										assign node312 = (inp[11]) ? node314 : 3'b010;
											assign node314 = (inp[8]) ? 3'b110 : 3'b010;
										assign node317 = (inp[11]) ? node319 : 3'b110;
											assign node319 = (inp[2]) ? 3'b011 : 3'b101;
								assign node322 = (inp[2]) ? node324 : 3'b101;
									assign node324 = (inp[11]) ? 3'b011 : 3'b101;
				assign node327 = (inp[4]) ? 3'b000 : node328;
					assign node328 = (inp[9]) ? 3'b111 : 3'b000;
		assign node332 = (inp[9]) ? node334 : 3'b000;
			assign node334 = (inp[0]) ? node336 : 3'b000;
				assign node336 = (inp[6]) ? node410 : node337;
					assign node337 = (inp[4]) ? node397 : node338;
						assign node338 = (inp[7]) ? node378 : node339;
							assign node339 = (inp[1]) ? node347 : node340;
								assign node340 = (inp[10]) ? node342 : 3'b000;
									assign node342 = (inp[2]) ? node344 : 3'b000;
										assign node344 = (inp[5]) ? 3'b000 : 3'b100;
								assign node347 = (inp[5]) ? node365 : node348;
									assign node348 = (inp[11]) ? node356 : node349;
										assign node349 = (inp[10]) ? node351 : 3'b010;
											assign node351 = (inp[2]) ? node353 : 3'b010;
												assign node353 = (inp[8]) ? 3'b010 : 3'b110;
										assign node356 = (inp[2]) ? node360 : node357;
											assign node357 = (inp[10]) ? 3'b110 : 3'b100;
											assign node360 = (inp[8]) ? 3'b001 : node361;
												assign node361 = (inp[10]) ? 3'b110 : 3'b010;
									assign node365 = (inp[10]) ? node371 : node366;
										assign node366 = (inp[8]) ? 3'b000 : node367;
											assign node367 = (inp[2]) ? 3'b100 : 3'b000;
										assign node371 = (inp[8]) ? 3'b100 : node372;
											assign node372 = (inp[11]) ? 3'b010 : node373;
												assign node373 = (inp[2]) ? 3'b100 : 3'b000;
							assign node378 = (inp[1]) ? node386 : node379;
								assign node379 = (inp[5]) ? 3'b010 : node380;
									assign node380 = (inp[11]) ? node382 : 3'b010;
										assign node382 = (inp[2]) ? 3'b000 : 3'b010;
								assign node386 = (inp[5]) ? node392 : node387;
									assign node387 = (inp[2]) ? node389 : 3'b110;
										assign node389 = (inp[11]) ? 3'b101 : 3'b110;
									assign node392 = (inp[2]) ? node394 : 3'b010;
										assign node394 = (inp[11]) ? 3'b110 : 3'b010;
						assign node397 = (inp[1]) ? node399 : 3'b000;
							assign node399 = (inp[5]) ? 3'b000 : node400;
								assign node400 = (inp[11]) ? node402 : 3'b000;
									assign node402 = (inp[2]) ? node404 : 3'b000;
										assign node404 = (inp[8]) ? 3'b100 : node405;
											assign node405 = (inp[7]) ? 3'b100 : 3'b000;
					assign node410 = (inp[5]) ? node412 : 3'b000;
						assign node412 = (inp[4]) ? node432 : node413;
							assign node413 = (inp[1]) ? node415 : 3'b000;
								assign node415 = (inp[2]) ? node421 : node416;
									assign node416 = (inp[11]) ? node418 : 3'b000;
										assign node418 = (inp[7]) ? 3'b001 : 3'b000;
									assign node421 = (inp[8]) ? node427 : node422;
										assign node422 = (inp[11]) ? 3'b000 : node423;
											assign node423 = (inp[7]) ? 3'b001 : 3'b000;
										assign node427 = (inp[7]) ? 3'b000 : node428;
											assign node428 = (inp[10]) ? 3'b000 : 3'b001;
							assign node432 = (inp[2]) ? node434 : 3'b000;
								assign node434 = (inp[1]) ? node436 : 3'b000;
									assign node436 = (inp[11]) ? node440 : node437;
										assign node437 = (inp[7]) ? 3'b100 : 3'b000;
										assign node440 = (inp[7]) ? 3'b010 : 3'b100;

endmodule