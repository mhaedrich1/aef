module dtc_split125_bm27 (
	input  wire [16-1:0] inp,
	output wire [16-1:0] outp
);

	wire [16-1:0] node1;
	wire [16-1:0] node2;
	wire [16-1:0] node3;
	wire [16-1:0] node4;
	wire [16-1:0] node5;
	wire [16-1:0] node6;
	wire [16-1:0] node7;
	wire [16-1:0] node8;
	wire [16-1:0] node9;
	wire [16-1:0] node10;
	wire [16-1:0] node12;
	wire [16-1:0] node13;
	wire [16-1:0] node14;
	wire [16-1:0] node16;
	wire [16-1:0] node21;
	wire [16-1:0] node23;
	wire [16-1:0] node24;
	wire [16-1:0] node25;
	wire [16-1:0] node30;
	wire [16-1:0] node31;
	wire [16-1:0] node32;
	wire [16-1:0] node33;
	wire [16-1:0] node37;
	wire [16-1:0] node39;
	wire [16-1:0] node41;
	wire [16-1:0] node44;
	wire [16-1:0] node46;
	wire [16-1:0] node49;
	wire [16-1:0] node50;
	wire [16-1:0] node51;
	wire [16-1:0] node52;
	wire [16-1:0] node53;
	wire [16-1:0] node54;
	wire [16-1:0] node59;
	wire [16-1:0] node60;
	wire [16-1:0] node61;
	wire [16-1:0] node65;
	wire [16-1:0] node66;
	wire [16-1:0] node70;
	wire [16-1:0] node71;
	wire [16-1:0] node72;
	wire [16-1:0] node74;
	wire [16-1:0] node78;
	wire [16-1:0] node79;
	wire [16-1:0] node83;
	wire [16-1:0] node84;
	wire [16-1:0] node85;
	wire [16-1:0] node87;
	wire [16-1:0] node88;
	wire [16-1:0] node93;
	wire [16-1:0] node95;
	wire [16-1:0] node98;
	wire [16-1:0] node99;
	wire [16-1:0] node100;
	wire [16-1:0] node101;
	wire [16-1:0] node102;
	wire [16-1:0] node104;
	wire [16-1:0] node105;
	wire [16-1:0] node110;
	wire [16-1:0] node111;
	wire [16-1:0] node114;
	wire [16-1:0] node116;
	wire [16-1:0] node119;
	wire [16-1:0] node120;
	wire [16-1:0] node121;
	wire [16-1:0] node124;
	wire [16-1:0] node125;
	wire [16-1:0] node128;
	wire [16-1:0] node129;
	wire [16-1:0] node133;
	wire [16-1:0] node134;
	wire [16-1:0] node135;
	wire [16-1:0] node139;
	wire [16-1:0] node140;
	wire [16-1:0] node141;
	wire [16-1:0] node145;
	wire [16-1:0] node148;
	wire [16-1:0] node149;
	wire [16-1:0] node150;
	wire [16-1:0] node151;
	wire [16-1:0] node154;
	wire [16-1:0] node156;
	wire [16-1:0] node159;
	wire [16-1:0] node160;
	wire [16-1:0] node163;
	wire [16-1:0] node165;
	wire [16-1:0] node168;
	wire [16-1:0] node169;
	wire [16-1:0] node170;
	wire [16-1:0] node171;
	wire [16-1:0] node175;
	wire [16-1:0] node176;
	wire [16-1:0] node180;
	wire [16-1:0] node181;
	wire [16-1:0] node182;
	wire [16-1:0] node186;
	wire [16-1:0] node189;
	wire [16-1:0] node190;
	wire [16-1:0] node191;
	wire [16-1:0] node192;
	wire [16-1:0] node193;
	wire [16-1:0] node195;
	wire [16-1:0] node198;
	wire [16-1:0] node199;
	wire [16-1:0] node201;
	wire [16-1:0] node202;
	wire [16-1:0] node206;
	wire [16-1:0] node209;
	wire [16-1:0] node210;
	wire [16-1:0] node211;
	wire [16-1:0] node214;
	wire [16-1:0] node215;
	wire [16-1:0] node217;
	wire [16-1:0] node221;
	wire [16-1:0] node222;
	wire [16-1:0] node224;
	wire [16-1:0] node227;
	wire [16-1:0] node230;
	wire [16-1:0] node231;
	wire [16-1:0] node232;
	wire [16-1:0] node233;
	wire [16-1:0] node235;
	wire [16-1:0] node237;
	wire [16-1:0] node241;
	wire [16-1:0] node242;
	wire [16-1:0] node244;
	wire [16-1:0] node247;
	wire [16-1:0] node250;
	wire [16-1:0] node251;
	wire [16-1:0] node252;
	wire [16-1:0] node255;
	wire [16-1:0] node258;
	wire [16-1:0] node259;
	wire [16-1:0] node262;
	wire [16-1:0] node265;
	wire [16-1:0] node266;
	wire [16-1:0] node267;
	wire [16-1:0] node268;
	wire [16-1:0] node269;
	wire [16-1:0] node273;
	wire [16-1:0] node274;
	wire [16-1:0] node275;
	wire [16-1:0] node276;
	wire [16-1:0] node281;
	wire [16-1:0] node283;
	wire [16-1:0] node286;
	wire [16-1:0] node287;
	wire [16-1:0] node288;
	wire [16-1:0] node289;
	wire [16-1:0] node290;
	wire [16-1:0] node295;
	wire [16-1:0] node297;
	wire [16-1:0] node300;
	wire [16-1:0] node301;
	wire [16-1:0] node303;
	wire [16-1:0] node306;
	wire [16-1:0] node309;
	wire [16-1:0] node310;
	wire [16-1:0] node311;
	wire [16-1:0] node312;
	wire [16-1:0] node315;
	wire [16-1:0] node318;
	wire [16-1:0] node319;
	wire [16-1:0] node321;
	wire [16-1:0] node323;
	wire [16-1:0] node326;
	wire [16-1:0] node329;
	wire [16-1:0] node330;
	wire [16-1:0] node332;
	wire [16-1:0] node334;
	wire [16-1:0] node335;
	wire [16-1:0] node339;
	wire [16-1:0] node340;
	wire [16-1:0] node342;
	wire [16-1:0] node343;
	wire [16-1:0] node348;
	wire [16-1:0] node349;
	wire [16-1:0] node350;
	wire [16-1:0] node351;
	wire [16-1:0] node352;
	wire [16-1:0] node353;
	wire [16-1:0] node354;
	wire [16-1:0] node358;
	wire [16-1:0] node359;
	wire [16-1:0] node363;
	wire [16-1:0] node364;
	wire [16-1:0] node365;
	wire [16-1:0] node368;
	wire [16-1:0] node369;
	wire [16-1:0] node373;
	wire [16-1:0] node374;
	wire [16-1:0] node375;
	wire [16-1:0] node378;
	wire [16-1:0] node379;
	wire [16-1:0] node381;
	wire [16-1:0] node385;
	wire [16-1:0] node387;
	wire [16-1:0] node390;
	wire [16-1:0] node391;
	wire [16-1:0] node392;
	wire [16-1:0] node393;
	wire [16-1:0] node396;
	wire [16-1:0] node398;
	wire [16-1:0] node400;
	wire [16-1:0] node401;
	wire [16-1:0] node405;
	wire [16-1:0] node406;
	wire [16-1:0] node407;
	wire [16-1:0] node409;
	wire [16-1:0] node413;
	wire [16-1:0] node416;
	wire [16-1:0] node417;
	wire [16-1:0] node418;
	wire [16-1:0] node420;
	wire [16-1:0] node423;
	wire [16-1:0] node424;
	wire [16-1:0] node426;
	wire [16-1:0] node430;
	wire [16-1:0] node432;
	wire [16-1:0] node434;
	wire [16-1:0] node435;
	wire [16-1:0] node439;
	wire [16-1:0] node440;
	wire [16-1:0] node441;
	wire [16-1:0] node442;
	wire [16-1:0] node443;
	wire [16-1:0] node446;
	wire [16-1:0] node447;
	wire [16-1:0] node451;
	wire [16-1:0] node452;
	wire [16-1:0] node453;
	wire [16-1:0] node455;
	wire [16-1:0] node458;
	wire [16-1:0] node459;
	wire [16-1:0] node464;
	wire [16-1:0] node465;
	wire [16-1:0] node466;
	wire [16-1:0] node470;
	wire [16-1:0] node471;
	wire [16-1:0] node474;
	wire [16-1:0] node475;
	wire [16-1:0] node477;
	wire [16-1:0] node481;
	wire [16-1:0] node482;
	wire [16-1:0] node483;
	wire [16-1:0] node484;
	wire [16-1:0] node487;
	wire [16-1:0] node488;
	wire [16-1:0] node489;
	wire [16-1:0] node492;
	wire [16-1:0] node495;
	wire [16-1:0] node496;
	wire [16-1:0] node500;
	wire [16-1:0] node501;
	wire [16-1:0] node502;
	wire [16-1:0] node505;
	wire [16-1:0] node508;
	wire [16-1:0] node509;
	wire [16-1:0] node513;
	wire [16-1:0] node514;
	wire [16-1:0] node515;
	wire [16-1:0] node518;
	wire [16-1:0] node520;
	wire [16-1:0] node521;
	wire [16-1:0] node525;
	wire [16-1:0] node527;
	wire [16-1:0] node529;
	wire [16-1:0] node531;
	wire [16-1:0] node534;
	wire [16-1:0] node535;
	wire [16-1:0] node536;
	wire [16-1:0] node537;
	wire [16-1:0] node538;
	wire [16-1:0] node539;
	wire [16-1:0] node540;
	wire [16-1:0] node544;
	wire [16-1:0] node546;
	wire [16-1:0] node549;
	wire [16-1:0] node550;
	wire [16-1:0] node552;
	wire [16-1:0] node556;
	wire [16-1:0] node557;
	wire [16-1:0] node559;
	wire [16-1:0] node560;
	wire [16-1:0] node561;
	wire [16-1:0] node566;
	wire [16-1:0] node567;
	wire [16-1:0] node568;
	wire [16-1:0] node573;
	wire [16-1:0] node574;
	wire [16-1:0] node575;
	wire [16-1:0] node576;
	wire [16-1:0] node578;
	wire [16-1:0] node579;
	wire [16-1:0] node583;
	wire [16-1:0] node585;
	wire [16-1:0] node588;
	wire [16-1:0] node589;
	wire [16-1:0] node590;
	wire [16-1:0] node594;
	wire [16-1:0] node596;
	wire [16-1:0] node599;
	wire [16-1:0] node600;
	wire [16-1:0] node601;
	wire [16-1:0] node602;
	wire [16-1:0] node605;
	wire [16-1:0] node606;
	wire [16-1:0] node610;
	wire [16-1:0] node612;
	wire [16-1:0] node615;
	wire [16-1:0] node616;
	wire [16-1:0] node617;
	wire [16-1:0] node621;
	wire [16-1:0] node623;
	wire [16-1:0] node626;
	wire [16-1:0] node627;
	wire [16-1:0] node628;
	wire [16-1:0] node629;
	wire [16-1:0] node630;
	wire [16-1:0] node632;
	wire [16-1:0] node636;
	wire [16-1:0] node637;
	wire [16-1:0] node638;
	wire [16-1:0] node639;
	wire [16-1:0] node644;
	wire [16-1:0] node647;
	wire [16-1:0] node648;
	wire [16-1:0] node650;
	wire [16-1:0] node652;
	wire [16-1:0] node655;
	wire [16-1:0] node656;
	wire [16-1:0] node657;
	wire [16-1:0] node661;
	wire [16-1:0] node663;
	wire [16-1:0] node664;
	wire [16-1:0] node668;
	wire [16-1:0] node669;
	wire [16-1:0] node670;
	wire [16-1:0] node672;
	wire [16-1:0] node675;
	wire [16-1:0] node676;
	wire [16-1:0] node678;
	wire [16-1:0] node679;
	wire [16-1:0] node682;
	wire [16-1:0] node686;
	wire [16-1:0] node687;
	wire [16-1:0] node688;
	wire [16-1:0] node692;
	wire [16-1:0] node693;
	wire [16-1:0] node696;
	wire [16-1:0] node697;
	wire [16-1:0] node699;
	wire [16-1:0] node702;
	wire [16-1:0] node705;
	wire [16-1:0] node706;
	wire [16-1:0] node707;
	wire [16-1:0] node708;
	wire [16-1:0] node709;
	wire [16-1:0] node710;
	wire [16-1:0] node711;
	wire [16-1:0] node712;
	wire [16-1:0] node714;
	wire [16-1:0] node717;
	wire [16-1:0] node718;
	wire [16-1:0] node720;
	wire [16-1:0] node724;
	wire [16-1:0] node725;
	wire [16-1:0] node729;
	wire [16-1:0] node730;
	wire [16-1:0] node731;
	wire [16-1:0] node734;
	wire [16-1:0] node736;
	wire [16-1:0] node739;
	wire [16-1:0] node740;
	wire [16-1:0] node741;
	wire [16-1:0] node743;
	wire [16-1:0] node746;
	wire [16-1:0] node748;
	wire [16-1:0] node751;
	wire [16-1:0] node753;
	wire [16-1:0] node756;
	wire [16-1:0] node757;
	wire [16-1:0] node758;
	wire [16-1:0] node759;
	wire [16-1:0] node761;
	wire [16-1:0] node765;
	wire [16-1:0] node766;
	wire [16-1:0] node768;
	wire [16-1:0] node771;
	wire [16-1:0] node773;
	wire [16-1:0] node774;
	wire [16-1:0] node778;
	wire [16-1:0] node779;
	wire [16-1:0] node780;
	wire [16-1:0] node782;
	wire [16-1:0] node785;
	wire [16-1:0] node788;
	wire [16-1:0] node789;
	wire [16-1:0] node792;
	wire [16-1:0] node794;
	wire [16-1:0] node795;
	wire [16-1:0] node799;
	wire [16-1:0] node800;
	wire [16-1:0] node801;
	wire [16-1:0] node802;
	wire [16-1:0] node803;
	wire [16-1:0] node804;
	wire [16-1:0] node806;
	wire [16-1:0] node809;
	wire [16-1:0] node812;
	wire [16-1:0] node815;
	wire [16-1:0] node816;
	wire [16-1:0] node818;
	wire [16-1:0] node820;
	wire [16-1:0] node823;
	wire [16-1:0] node826;
	wire [16-1:0] node827;
	wire [16-1:0] node828;
	wire [16-1:0] node830;
	wire [16-1:0] node834;
	wire [16-1:0] node835;
	wire [16-1:0] node837;
	wire [16-1:0] node840;
	wire [16-1:0] node841;
	wire [16-1:0] node842;
	wire [16-1:0] node846;
	wire [16-1:0] node849;
	wire [16-1:0] node850;
	wire [16-1:0] node851;
	wire [16-1:0] node852;
	wire [16-1:0] node853;
	wire [16-1:0] node855;
	wire [16-1:0] node859;
	wire [16-1:0] node860;
	wire [16-1:0] node861;
	wire [16-1:0] node865;
	wire [16-1:0] node866;
	wire [16-1:0] node870;
	wire [16-1:0] node871;
	wire [16-1:0] node874;
	wire [16-1:0] node877;
	wire [16-1:0] node879;
	wire [16-1:0] node880;
	wire [16-1:0] node882;
	wire [16-1:0] node886;
	wire [16-1:0] node887;
	wire [16-1:0] node888;
	wire [16-1:0] node889;
	wire [16-1:0] node890;
	wire [16-1:0] node891;
	wire [16-1:0] node893;
	wire [16-1:0] node894;
	wire [16-1:0] node896;
	wire [16-1:0] node900;
	wire [16-1:0] node903;
	wire [16-1:0] node904;
	wire [16-1:0] node908;
	wire [16-1:0] node909;
	wire [16-1:0] node910;
	wire [16-1:0] node911;
	wire [16-1:0] node915;
	wire [16-1:0] node916;
	wire [16-1:0] node920;
	wire [16-1:0] node922;
	wire [16-1:0] node923;
	wire [16-1:0] node927;
	wire [16-1:0] node928;
	wire [16-1:0] node929;
	wire [16-1:0] node931;
	wire [16-1:0] node933;
	wire [16-1:0] node934;
	wire [16-1:0] node938;
	wire [16-1:0] node939;
	wire [16-1:0] node940;
	wire [16-1:0] node941;
	wire [16-1:0] node946;
	wire [16-1:0] node948;
	wire [16-1:0] node951;
	wire [16-1:0] node952;
	wire [16-1:0] node953;
	wire [16-1:0] node955;
	wire [16-1:0] node956;
	wire [16-1:0] node960;
	wire [16-1:0] node961;
	wire [16-1:0] node964;
	wire [16-1:0] node967;
	wire [16-1:0] node968;
	wire [16-1:0] node971;
	wire [16-1:0] node972;
	wire [16-1:0] node975;
	wire [16-1:0] node978;
	wire [16-1:0] node979;
	wire [16-1:0] node980;
	wire [16-1:0] node981;
	wire [16-1:0] node982;
	wire [16-1:0] node985;
	wire [16-1:0] node987;
	wire [16-1:0] node990;
	wire [16-1:0] node991;
	wire [16-1:0] node994;
	wire [16-1:0] node997;
	wire [16-1:0] node998;
	wire [16-1:0] node999;
	wire [16-1:0] node1003;
	wire [16-1:0] node1004;
	wire [16-1:0] node1006;
	wire [16-1:0] node1009;
	wire [16-1:0] node1010;
	wire [16-1:0] node1013;
	wire [16-1:0] node1016;
	wire [16-1:0] node1017;
	wire [16-1:0] node1018;
	wire [16-1:0] node1019;
	wire [16-1:0] node1020;
	wire [16-1:0] node1025;
	wire [16-1:0] node1026;
	wire [16-1:0] node1027;
	wire [16-1:0] node1029;
	wire [16-1:0] node1033;
	wire [16-1:0] node1034;
	wire [16-1:0] node1035;
	wire [16-1:0] node1037;
	wire [16-1:0] node1042;
	wire [16-1:0] node1043;
	wire [16-1:0] node1044;
	wire [16-1:0] node1047;
	wire [16-1:0] node1048;
	wire [16-1:0] node1052;
	wire [16-1:0] node1053;
	wire [16-1:0] node1054;
	wire [16-1:0] node1056;
	wire [16-1:0] node1060;
	wire [16-1:0] node1061;
	wire [16-1:0] node1062;
	wire [16-1:0] node1065;
	wire [16-1:0] node1068;
	wire [16-1:0] node1069;
	wire [16-1:0] node1072;
	wire [16-1:0] node1075;
	wire [16-1:0] node1076;
	wire [16-1:0] node1077;
	wire [16-1:0] node1078;
	wire [16-1:0] node1079;
	wire [16-1:0] node1080;
	wire [16-1:0] node1081;
	wire [16-1:0] node1082;
	wire [16-1:0] node1085;
	wire [16-1:0] node1088;
	wire [16-1:0] node1089;
	wire [16-1:0] node1090;
	wire [16-1:0] node1094;
	wire [16-1:0] node1097;
	wire [16-1:0] node1098;
	wire [16-1:0] node1101;
	wire [16-1:0] node1103;
	wire [16-1:0] node1106;
	wire [16-1:0] node1107;
	wire [16-1:0] node1108;
	wire [16-1:0] node1109;
	wire [16-1:0] node1110;
	wire [16-1:0] node1115;
	wire [16-1:0] node1117;
	wire [16-1:0] node1120;
	wire [16-1:0] node1121;
	wire [16-1:0] node1124;
	wire [16-1:0] node1127;
	wire [16-1:0] node1128;
	wire [16-1:0] node1129;
	wire [16-1:0] node1130;
	wire [16-1:0] node1132;
	wire [16-1:0] node1133;
	wire [16-1:0] node1136;
	wire [16-1:0] node1139;
	wire [16-1:0] node1140;
	wire [16-1:0] node1144;
	wire [16-1:0] node1146;
	wire [16-1:0] node1149;
	wire [16-1:0] node1150;
	wire [16-1:0] node1152;
	wire [16-1:0] node1155;
	wire [16-1:0] node1157;
	wire [16-1:0] node1158;
	wire [16-1:0] node1162;
	wire [16-1:0] node1163;
	wire [16-1:0] node1164;
	wire [16-1:0] node1165;
	wire [16-1:0] node1166;
	wire [16-1:0] node1167;
	wire [16-1:0] node1168;
	wire [16-1:0] node1173;
	wire [16-1:0] node1174;
	wire [16-1:0] node1177;
	wire [16-1:0] node1180;
	wire [16-1:0] node1181;
	wire [16-1:0] node1182;
	wire [16-1:0] node1185;
	wire [16-1:0] node1186;
	wire [16-1:0] node1187;
	wire [16-1:0] node1192;
	wire [16-1:0] node1195;
	wire [16-1:0] node1196;
	wire [16-1:0] node1197;
	wire [16-1:0] node1198;
	wire [16-1:0] node1200;
	wire [16-1:0] node1204;
	wire [16-1:0] node1207;
	wire [16-1:0] node1208;
	wire [16-1:0] node1210;
	wire [16-1:0] node1212;
	wire [16-1:0] node1213;
	wire [16-1:0] node1217;
	wire [16-1:0] node1218;
	wire [16-1:0] node1219;
	wire [16-1:0] node1223;
	wire [16-1:0] node1225;
	wire [16-1:0] node1227;
	wire [16-1:0] node1230;
	wire [16-1:0] node1231;
	wire [16-1:0] node1232;
	wire [16-1:0] node1233;
	wire [16-1:0] node1234;
	wire [16-1:0] node1235;
	wire [16-1:0] node1240;
	wire [16-1:0] node1241;
	wire [16-1:0] node1244;
	wire [16-1:0] node1247;
	wire [16-1:0] node1248;
	wire [16-1:0] node1250;
	wire [16-1:0] node1252;
	wire [16-1:0] node1255;
	wire [16-1:0] node1256;
	wire [16-1:0] node1257;
	wire [16-1:0] node1262;
	wire [16-1:0] node1263;
	wire [16-1:0] node1264;
	wire [16-1:0] node1266;
	wire [16-1:0] node1268;
	wire [16-1:0] node1271;
	wire [16-1:0] node1274;
	wire [16-1:0] node1275;
	wire [16-1:0] node1276;
	wire [16-1:0] node1280;
	wire [16-1:0] node1281;
	wire [16-1:0] node1283;
	wire [16-1:0] node1286;
	wire [16-1:0] node1289;
	wire [16-1:0] node1290;
	wire [16-1:0] node1291;
	wire [16-1:0] node1292;
	wire [16-1:0] node1293;
	wire [16-1:0] node1294;
	wire [16-1:0] node1296;
	wire [16-1:0] node1297;
	wire [16-1:0] node1301;
	wire [16-1:0] node1303;
	wire [16-1:0] node1306;
	wire [16-1:0] node1307;
	wire [16-1:0] node1310;
	wire [16-1:0] node1312;
	wire [16-1:0] node1313;
	wire [16-1:0] node1317;
	wire [16-1:0] node1318;
	wire [16-1:0] node1319;
	wire [16-1:0] node1322;
	wire [16-1:0] node1324;
	wire [16-1:0] node1327;
	wire [16-1:0] node1328;
	wire [16-1:0] node1331;
	wire [16-1:0] node1334;
	wire [16-1:0] node1335;
	wire [16-1:0] node1336;
	wire [16-1:0] node1337;
	wire [16-1:0] node1339;
	wire [16-1:0] node1342;
	wire [16-1:0] node1343;
	wire [16-1:0] node1347;
	wire [16-1:0] node1350;
	wire [16-1:0] node1351;
	wire [16-1:0] node1352;
	wire [16-1:0] node1353;
	wire [16-1:0] node1356;
	wire [16-1:0] node1357;
	wire [16-1:0] node1361;
	wire [16-1:0] node1363;
	wire [16-1:0] node1365;
	wire [16-1:0] node1368;
	wire [16-1:0] node1369;
	wire [16-1:0] node1370;
	wire [16-1:0] node1371;
	wire [16-1:0] node1372;
	wire [16-1:0] node1377;
	wire [16-1:0] node1378;
	wire [16-1:0] node1382;
	wire [16-1:0] node1383;
	wire [16-1:0] node1385;
	wire [16-1:0] node1386;
	wire [16-1:0] node1390;
	wire [16-1:0] node1391;
	wire [16-1:0] node1395;
	wire [16-1:0] node1396;
	wire [16-1:0] node1397;
	wire [16-1:0] node1398;
	wire [16-1:0] node1399;
	wire [16-1:0] node1401;
	wire [16-1:0] node1402;
	wire [16-1:0] node1406;
	wire [16-1:0] node1407;
	wire [16-1:0] node1410;
	wire [16-1:0] node1412;
	wire [16-1:0] node1413;
	wire [16-1:0] node1417;
	wire [16-1:0] node1419;
	wire [16-1:0] node1420;
	wire [16-1:0] node1422;
	wire [16-1:0] node1424;
	wire [16-1:0] node1428;
	wire [16-1:0] node1429;
	wire [16-1:0] node1431;
	wire [16-1:0] node1432;
	wire [16-1:0] node1434;
	wire [16-1:0] node1438;
	wire [16-1:0] node1439;
	wire [16-1:0] node1441;
	wire [16-1:0] node1444;
	wire [16-1:0] node1445;
	wire [16-1:0] node1447;
	wire [16-1:0] node1451;
	wire [16-1:0] node1452;
	wire [16-1:0] node1453;
	wire [16-1:0] node1456;
	wire [16-1:0] node1458;
	wire [16-1:0] node1459;
	wire [16-1:0] node1461;
	wire [16-1:0] node1465;
	wire [16-1:0] node1467;
	wire [16-1:0] node1468;
	wire [16-1:0] node1469;
	wire [16-1:0] node1472;
	wire [16-1:0] node1475;
	wire [16-1:0] node1476;
	wire [16-1:0] node1478;
	wire [16-1:0] node1482;
	wire [16-1:0] node1483;
	wire [16-1:0] node1484;
	wire [16-1:0] node1485;
	wire [16-1:0] node1486;
	wire [16-1:0] node1487;
	wire [16-1:0] node1488;
	wire [16-1:0] node1489;
	wire [16-1:0] node1490;
	wire [16-1:0] node1492;
	wire [16-1:0] node1495;
	wire [16-1:0] node1498;
	wire [16-1:0] node1500;
	wire [16-1:0] node1501;
	wire [16-1:0] node1505;
	wire [16-1:0] node1506;
	wire [16-1:0] node1508;
	wire [16-1:0] node1511;
	wire [16-1:0] node1512;
	wire [16-1:0] node1515;
	wire [16-1:0] node1516;
	wire [16-1:0] node1519;
	wire [16-1:0] node1522;
	wire [16-1:0] node1523;
	wire [16-1:0] node1524;
	wire [16-1:0] node1525;
	wire [16-1:0] node1526;
	wire [16-1:0] node1530;
	wire [16-1:0] node1533;
	wire [16-1:0] node1534;
	wire [16-1:0] node1535;
	wire [16-1:0] node1539;
	wire [16-1:0] node1542;
	wire [16-1:0] node1543;
	wire [16-1:0] node1544;
	wire [16-1:0] node1547;
	wire [16-1:0] node1549;
	wire [16-1:0] node1551;
	wire [16-1:0] node1554;
	wire [16-1:0] node1556;
	wire [16-1:0] node1558;
	wire [16-1:0] node1559;
	wire [16-1:0] node1561;
	wire [16-1:0] node1565;
	wire [16-1:0] node1566;
	wire [16-1:0] node1567;
	wire [16-1:0] node1568;
	wire [16-1:0] node1569;
	wire [16-1:0] node1570;
	wire [16-1:0] node1574;
	wire [16-1:0] node1575;
	wire [16-1:0] node1577;
	wire [16-1:0] node1581;
	wire [16-1:0] node1582;
	wire [16-1:0] node1583;
	wire [16-1:0] node1587;
	wire [16-1:0] node1588;
	wire [16-1:0] node1590;
	wire [16-1:0] node1594;
	wire [16-1:0] node1595;
	wire [16-1:0] node1596;
	wire [16-1:0] node1598;
	wire [16-1:0] node1601;
	wire [16-1:0] node1604;
	wire [16-1:0] node1605;
	wire [16-1:0] node1606;
	wire [16-1:0] node1608;
	wire [16-1:0] node1612;
	wire [16-1:0] node1615;
	wire [16-1:0] node1616;
	wire [16-1:0] node1617;
	wire [16-1:0] node1618;
	wire [16-1:0] node1619;
	wire [16-1:0] node1621;
	wire [16-1:0] node1624;
	wire [16-1:0] node1625;
	wire [16-1:0] node1628;
	wire [16-1:0] node1630;
	wire [16-1:0] node1634;
	wire [16-1:0] node1635;
	wire [16-1:0] node1637;
	wire [16-1:0] node1638;
	wire [16-1:0] node1639;
	wire [16-1:0] node1644;
	wire [16-1:0] node1646;
	wire [16-1:0] node1649;
	wire [16-1:0] node1650;
	wire [16-1:0] node1651;
	wire [16-1:0] node1654;
	wire [16-1:0] node1655;
	wire [16-1:0] node1658;
	wire [16-1:0] node1659;
	wire [16-1:0] node1661;
	wire [16-1:0] node1665;
	wire [16-1:0] node1666;
	wire [16-1:0] node1668;
	wire [16-1:0] node1672;
	wire [16-1:0] node1673;
	wire [16-1:0] node1674;
	wire [16-1:0] node1675;
	wire [16-1:0] node1676;
	wire [16-1:0] node1678;
	wire [16-1:0] node1681;
	wire [16-1:0] node1682;
	wire [16-1:0] node1683;
	wire [16-1:0] node1687;
	wire [16-1:0] node1690;
	wire [16-1:0] node1691;
	wire [16-1:0] node1692;
	wire [16-1:0] node1695;
	wire [16-1:0] node1696;
	wire [16-1:0] node1699;
	wire [16-1:0] node1700;
	wire [16-1:0] node1704;
	wire [16-1:0] node1705;
	wire [16-1:0] node1707;
	wire [16-1:0] node1709;
	wire [16-1:0] node1712;
	wire [16-1:0] node1714;
	wire [16-1:0] node1716;
	wire [16-1:0] node1719;
	wire [16-1:0] node1720;
	wire [16-1:0] node1721;
	wire [16-1:0] node1723;
	wire [16-1:0] node1725;
	wire [16-1:0] node1728;
	wire [16-1:0] node1729;
	wire [16-1:0] node1733;
	wire [16-1:0] node1734;
	wire [16-1:0] node1735;
	wire [16-1:0] node1738;
	wire [16-1:0] node1740;
	wire [16-1:0] node1741;
	wire [16-1:0] node1745;
	wire [16-1:0] node1746;
	wire [16-1:0] node1747;
	wire [16-1:0] node1751;
	wire [16-1:0] node1754;
	wire [16-1:0] node1755;
	wire [16-1:0] node1756;
	wire [16-1:0] node1757;
	wire [16-1:0] node1758;
	wire [16-1:0] node1759;
	wire [16-1:0] node1761;
	wire [16-1:0] node1766;
	wire [16-1:0] node1767;
	wire [16-1:0] node1768;
	wire [16-1:0] node1769;
	wire [16-1:0] node1773;
	wire [16-1:0] node1775;
	wire [16-1:0] node1778;
	wire [16-1:0] node1779;
	wire [16-1:0] node1782;
	wire [16-1:0] node1783;
	wire [16-1:0] node1787;
	wire [16-1:0] node1788;
	wire [16-1:0] node1789;
	wire [16-1:0] node1792;
	wire [16-1:0] node1795;
	wire [16-1:0] node1797;
	wire [16-1:0] node1799;
	wire [16-1:0] node1802;
	wire [16-1:0] node1803;
	wire [16-1:0] node1804;
	wire [16-1:0] node1805;
	wire [16-1:0] node1807;
	wire [16-1:0] node1808;
	wire [16-1:0] node1810;
	wire [16-1:0] node1814;
	wire [16-1:0] node1816;
	wire [16-1:0] node1819;
	wire [16-1:0] node1821;
	wire [16-1:0] node1822;
	wire [16-1:0] node1826;
	wire [16-1:0] node1827;
	wire [16-1:0] node1829;
	wire [16-1:0] node1830;
	wire [16-1:0] node1831;
	wire [16-1:0] node1836;
	wire [16-1:0] node1837;
	wire [16-1:0] node1840;
	wire [16-1:0] node1843;
	wire [16-1:0] node1844;
	wire [16-1:0] node1845;
	wire [16-1:0] node1846;
	wire [16-1:0] node1847;
	wire [16-1:0] node1848;
	wire [16-1:0] node1849;
	wire [16-1:0] node1850;
	wire [16-1:0] node1854;
	wire [16-1:0] node1857;
	wire [16-1:0] node1858;
	wire [16-1:0] node1859;
	wire [16-1:0] node1862;
	wire [16-1:0] node1865;
	wire [16-1:0] node1866;
	wire [16-1:0] node1870;
	wire [16-1:0] node1871;
	wire [16-1:0] node1872;
	wire [16-1:0] node1874;
	wire [16-1:0] node1876;
	wire [16-1:0] node1879;
	wire [16-1:0] node1882;
	wire [16-1:0] node1883;
	wire [16-1:0] node1884;
	wire [16-1:0] node1885;
	wire [16-1:0] node1889;
	wire [16-1:0] node1890;
	wire [16-1:0] node1894;
	wire [16-1:0] node1895;
	wire [16-1:0] node1898;
	wire [16-1:0] node1900;
	wire [16-1:0] node1903;
	wire [16-1:0] node1904;
	wire [16-1:0] node1905;
	wire [16-1:0] node1906;
	wire [16-1:0] node1907;
	wire [16-1:0] node1910;
	wire [16-1:0] node1912;
	wire [16-1:0] node1915;
	wire [16-1:0] node1918;
	wire [16-1:0] node1919;
	wire [16-1:0] node1920;
	wire [16-1:0] node1922;
	wire [16-1:0] node1925;
	wire [16-1:0] node1928;
	wire [16-1:0] node1930;
	wire [16-1:0] node1933;
	wire [16-1:0] node1934;
	wire [16-1:0] node1935;
	wire [16-1:0] node1937;
	wire [16-1:0] node1939;
	wire [16-1:0] node1942;
	wire [16-1:0] node1943;
	wire [16-1:0] node1947;
	wire [16-1:0] node1948;
	wire [16-1:0] node1951;
	wire [16-1:0] node1954;
	wire [16-1:0] node1955;
	wire [16-1:0] node1956;
	wire [16-1:0] node1957;
	wire [16-1:0] node1958;
	wire [16-1:0] node1960;
	wire [16-1:0] node1963;
	wire [16-1:0] node1964;
	wire [16-1:0] node1968;
	wire [16-1:0] node1969;
	wire [16-1:0] node1973;
	wire [16-1:0] node1974;
	wire [16-1:0] node1975;
	wire [16-1:0] node1976;
	wire [16-1:0] node1979;
	wire [16-1:0] node1982;
	wire [16-1:0] node1984;
	wire [16-1:0] node1986;
	wire [16-1:0] node1989;
	wire [16-1:0] node1990;
	wire [16-1:0] node1992;
	wire [16-1:0] node1993;
	wire [16-1:0] node1996;
	wire [16-1:0] node1999;
	wire [16-1:0] node2000;
	wire [16-1:0] node2001;
	wire [16-1:0] node2004;
	wire [16-1:0] node2008;
	wire [16-1:0] node2009;
	wire [16-1:0] node2010;
	wire [16-1:0] node2011;
	wire [16-1:0] node2013;
	wire [16-1:0] node2016;
	wire [16-1:0] node2018;
	wire [16-1:0] node2021;
	wire [16-1:0] node2022;
	wire [16-1:0] node2023;
	wire [16-1:0] node2025;
	wire [16-1:0] node2028;
	wire [16-1:0] node2031;
	wire [16-1:0] node2033;
	wire [16-1:0] node2036;
	wire [16-1:0] node2037;
	wire [16-1:0] node2039;
	wire [16-1:0] node2040;
	wire [16-1:0] node2044;
	wire [16-1:0] node2045;
	wire [16-1:0] node2047;
	wire [16-1:0] node2048;
	wire [16-1:0] node2052;
	wire [16-1:0] node2053;
	wire [16-1:0] node2056;
	wire [16-1:0] node2058;
	wire [16-1:0] node2059;
	wire [16-1:0] node2063;
	wire [16-1:0] node2064;
	wire [16-1:0] node2065;
	wire [16-1:0] node2066;
	wire [16-1:0] node2067;
	wire [16-1:0] node2068;
	wire [16-1:0] node2071;
	wire [16-1:0] node2072;
	wire [16-1:0] node2076;
	wire [16-1:0] node2078;
	wire [16-1:0] node2079;
	wire [16-1:0] node2082;
	wire [16-1:0] node2084;
	wire [16-1:0] node2086;
	wire [16-1:0] node2089;
	wire [16-1:0] node2090;
	wire [16-1:0] node2091;
	wire [16-1:0] node2095;
	wire [16-1:0] node2096;
	wire [16-1:0] node2098;
	wire [16-1:0] node2099;
	wire [16-1:0] node2103;
	wire [16-1:0] node2106;
	wire [16-1:0] node2107;
	wire [16-1:0] node2108;
	wire [16-1:0] node2109;
	wire [16-1:0] node2110;
	wire [16-1:0] node2114;
	wire [16-1:0] node2115;
	wire [16-1:0] node2116;
	wire [16-1:0] node2121;
	wire [16-1:0] node2122;
	wire [16-1:0] node2124;
	wire [16-1:0] node2125;
	wire [16-1:0] node2127;
	wire [16-1:0] node2130;
	wire [16-1:0] node2133;
	wire [16-1:0] node2136;
	wire [16-1:0] node2137;
	wire [16-1:0] node2138;
	wire [16-1:0] node2140;
	wire [16-1:0] node2143;
	wire [16-1:0] node2145;
	wire [16-1:0] node2148;
	wire [16-1:0] node2149;
	wire [16-1:0] node2150;
	wire [16-1:0] node2154;
	wire [16-1:0] node2157;
	wire [16-1:0] node2158;
	wire [16-1:0] node2159;
	wire [16-1:0] node2160;
	wire [16-1:0] node2161;
	wire [16-1:0] node2162;
	wire [16-1:0] node2165;
	wire [16-1:0] node2169;
	wire [16-1:0] node2170;
	wire [16-1:0] node2171;
	wire [16-1:0] node2175;
	wire [16-1:0] node2178;
	wire [16-1:0] node2179;
	wire [16-1:0] node2180;
	wire [16-1:0] node2183;
	wire [16-1:0] node2185;
	wire [16-1:0] node2186;
	wire [16-1:0] node2190;
	wire [16-1:0] node2192;
	wire [16-1:0] node2194;
	wire [16-1:0] node2195;
	wire [16-1:0] node2199;
	wire [16-1:0] node2200;
	wire [16-1:0] node2201;
	wire [16-1:0] node2202;
	wire [16-1:0] node2203;
	wire [16-1:0] node2204;
	wire [16-1:0] node2206;
	wire [16-1:0] node2210;
	wire [16-1:0] node2214;
	wire [16-1:0] node2215;
	wire [16-1:0] node2216;
	wire [16-1:0] node2219;
	wire [16-1:0] node2221;
	wire [16-1:0] node2224;
	wire [16-1:0] node2225;
	wire [16-1:0] node2227;
	wire [16-1:0] node2231;
	wire [16-1:0] node2232;
	wire [16-1:0] node2233;
	wire [16-1:0] node2235;
	wire [16-1:0] node2236;
	wire [16-1:0] node2240;
	wire [16-1:0] node2243;
	wire [16-1:0] node2244;
	wire [16-1:0] node2246;
	wire [16-1:0] node2249;
	wire [16-1:0] node2251;
	wire [16-1:0] node2253;
	wire [16-1:0] node2256;
	wire [16-1:0] node2257;
	wire [16-1:0] node2258;
	wire [16-1:0] node2259;
	wire [16-1:0] node2260;
	wire [16-1:0] node2261;
	wire [16-1:0] node2262;
	wire [16-1:0] node2263;
	wire [16-1:0] node2265;
	wire [16-1:0] node2266;
	wire [16-1:0] node2270;
	wire [16-1:0] node2273;
	wire [16-1:0] node2274;
	wire [16-1:0] node2275;
	wire [16-1:0] node2277;
	wire [16-1:0] node2278;
	wire [16-1:0] node2282;
	wire [16-1:0] node2286;
	wire [16-1:0] node2287;
	wire [16-1:0] node2288;
	wire [16-1:0] node2289;
	wire [16-1:0] node2293;
	wire [16-1:0] node2295;
	wire [16-1:0] node2298;
	wire [16-1:0] node2299;
	wire [16-1:0] node2300;
	wire [16-1:0] node2304;
	wire [16-1:0] node2307;
	wire [16-1:0] node2308;
	wire [16-1:0] node2309;
	wire [16-1:0] node2310;
	wire [16-1:0] node2311;
	wire [16-1:0] node2313;
	wire [16-1:0] node2314;
	wire [16-1:0] node2319;
	wire [16-1:0] node2322;
	wire [16-1:0] node2323;
	wire [16-1:0] node2324;
	wire [16-1:0] node2327;
	wire [16-1:0] node2330;
	wire [16-1:0] node2331;
	wire [16-1:0] node2335;
	wire [16-1:0] node2336;
	wire [16-1:0] node2337;
	wire [16-1:0] node2338;
	wire [16-1:0] node2341;
	wire [16-1:0] node2344;
	wire [16-1:0] node2347;
	wire [16-1:0] node2349;
	wire [16-1:0] node2351;
	wire [16-1:0] node2354;
	wire [16-1:0] node2355;
	wire [16-1:0] node2356;
	wire [16-1:0] node2357;
	wire [16-1:0] node2358;
	wire [16-1:0] node2359;
	wire [16-1:0] node2360;
	wire [16-1:0] node2365;
	wire [16-1:0] node2368;
	wire [16-1:0] node2369;
	wire [16-1:0] node2371;
	wire [16-1:0] node2372;
	wire [16-1:0] node2374;
	wire [16-1:0] node2379;
	wire [16-1:0] node2380;
	wire [16-1:0] node2382;
	wire [16-1:0] node2385;
	wire [16-1:0] node2386;
	wire [16-1:0] node2388;
	wire [16-1:0] node2389;
	wire [16-1:0] node2391;
	wire [16-1:0] node2395;
	wire [16-1:0] node2396;
	wire [16-1:0] node2399;
	wire [16-1:0] node2401;
	wire [16-1:0] node2404;
	wire [16-1:0] node2405;
	wire [16-1:0] node2406;
	wire [16-1:0] node2407;
	wire [16-1:0] node2409;
	wire [16-1:0] node2412;
	wire [16-1:0] node2413;
	wire [16-1:0] node2414;
	wire [16-1:0] node2418;
	wire [16-1:0] node2421;
	wire [16-1:0] node2422;
	wire [16-1:0] node2425;
	wire [16-1:0] node2426;
	wire [16-1:0] node2429;
	wire [16-1:0] node2431;
	wire [16-1:0] node2434;
	wire [16-1:0] node2435;
	wire [16-1:0] node2436;
	wire [16-1:0] node2438;
	wire [16-1:0] node2441;
	wire [16-1:0] node2442;
	wire [16-1:0] node2444;
	wire [16-1:0] node2447;
	wire [16-1:0] node2450;
	wire [16-1:0] node2451;
	wire [16-1:0] node2454;
	wire [16-1:0] node2456;
	wire [16-1:0] node2459;
	wire [16-1:0] node2460;
	wire [16-1:0] node2461;
	wire [16-1:0] node2462;
	wire [16-1:0] node2463;
	wire [16-1:0] node2464;
	wire [16-1:0] node2467;
	wire [16-1:0] node2470;
	wire [16-1:0] node2471;
	wire [16-1:0] node2472;
	wire [16-1:0] node2476;
	wire [16-1:0] node2477;
	wire [16-1:0] node2479;
	wire [16-1:0] node2483;
	wire [16-1:0] node2484;
	wire [16-1:0] node2485;
	wire [16-1:0] node2489;
	wire [16-1:0] node2491;
	wire [16-1:0] node2492;
	wire [16-1:0] node2493;
	wire [16-1:0] node2497;
	wire [16-1:0] node2498;
	wire [16-1:0] node2502;
	wire [16-1:0] node2503;
	wire [16-1:0] node2504;
	wire [16-1:0] node2505;
	wire [16-1:0] node2507;
	wire [16-1:0] node2508;
	wire [16-1:0] node2512;
	wire [16-1:0] node2515;
	wire [16-1:0] node2516;
	wire [16-1:0] node2519;
	wire [16-1:0] node2521;
	wire [16-1:0] node2522;
	wire [16-1:0] node2526;
	wire [16-1:0] node2527;
	wire [16-1:0] node2528;
	wire [16-1:0] node2531;
	wire [16-1:0] node2532;
	wire [16-1:0] node2534;
	wire [16-1:0] node2538;
	wire [16-1:0] node2539;
	wire [16-1:0] node2541;
	wire [16-1:0] node2542;
	wire [16-1:0] node2546;
	wire [16-1:0] node2548;
	wire [16-1:0] node2551;
	wire [16-1:0] node2552;
	wire [16-1:0] node2553;
	wire [16-1:0] node2554;
	wire [16-1:0] node2555;
	wire [16-1:0] node2558;
	wire [16-1:0] node2559;
	wire [16-1:0] node2562;
	wire [16-1:0] node2564;
	wire [16-1:0] node2567;
	wire [16-1:0] node2569;
	wire [16-1:0] node2571;
	wire [16-1:0] node2574;
	wire [16-1:0] node2575;
	wire [16-1:0] node2576;
	wire [16-1:0] node2579;
	wire [16-1:0] node2582;
	wire [16-1:0] node2583;
	wire [16-1:0] node2585;
	wire [16-1:0] node2588;
	wire [16-1:0] node2590;
	wire [16-1:0] node2593;
	wire [16-1:0] node2594;
	wire [16-1:0] node2595;
	wire [16-1:0] node2596;
	wire [16-1:0] node2598;
	wire [16-1:0] node2601;
	wire [16-1:0] node2603;
	wire [16-1:0] node2604;
	wire [16-1:0] node2607;
	wire [16-1:0] node2610;
	wire [16-1:0] node2611;
	wire [16-1:0] node2614;
	wire [16-1:0] node2615;
	wire [16-1:0] node2616;
	wire [16-1:0] node2621;
	wire [16-1:0] node2622;
	wire [16-1:0] node2623;
	wire [16-1:0] node2626;
	wire [16-1:0] node2628;
	wire [16-1:0] node2631;
	wire [16-1:0] node2632;
	wire [16-1:0] node2636;
	wire [16-1:0] node2637;
	wire [16-1:0] node2638;
	wire [16-1:0] node2639;
	wire [16-1:0] node2640;
	wire [16-1:0] node2641;
	wire [16-1:0] node2642;
	wire [16-1:0] node2643;
	wire [16-1:0] node2644;
	wire [16-1:0] node2646;
	wire [16-1:0] node2651;
	wire [16-1:0] node2654;
	wire [16-1:0] node2655;
	wire [16-1:0] node2658;
	wire [16-1:0] node2661;
	wire [16-1:0] node2662;
	wire [16-1:0] node2663;
	wire [16-1:0] node2664;
	wire [16-1:0] node2666;
	wire [16-1:0] node2670;
	wire [16-1:0] node2673;
	wire [16-1:0] node2674;
	wire [16-1:0] node2675;
	wire [16-1:0] node2677;
	wire [16-1:0] node2681;
	wire [16-1:0] node2682;
	wire [16-1:0] node2684;
	wire [16-1:0] node2688;
	wire [16-1:0] node2689;
	wire [16-1:0] node2690;
	wire [16-1:0] node2691;
	wire [16-1:0] node2694;
	wire [16-1:0] node2696;
	wire [16-1:0] node2699;
	wire [16-1:0] node2700;
	wire [16-1:0] node2701;
	wire [16-1:0] node2705;
	wire [16-1:0] node2708;
	wire [16-1:0] node2710;
	wire [16-1:0] node2711;
	wire [16-1:0] node2714;
	wire [16-1:0] node2716;
	wire [16-1:0] node2719;
	wire [16-1:0] node2720;
	wire [16-1:0] node2721;
	wire [16-1:0] node2722;
	wire [16-1:0] node2723;
	wire [16-1:0] node2724;
	wire [16-1:0] node2729;
	wire [16-1:0] node2730;
	wire [16-1:0] node2733;
	wire [16-1:0] node2735;
	wire [16-1:0] node2736;
	wire [16-1:0] node2740;
	wire [16-1:0] node2741;
	wire [16-1:0] node2742;
	wire [16-1:0] node2743;
	wire [16-1:0] node2747;
	wire [16-1:0] node2748;
	wire [16-1:0] node2752;
	wire [16-1:0] node2753;
	wire [16-1:0] node2756;
	wire [16-1:0] node2759;
	wire [16-1:0] node2760;
	wire [16-1:0] node2761;
	wire [16-1:0] node2762;
	wire [16-1:0] node2763;
	wire [16-1:0] node2764;
	wire [16-1:0] node2769;
	wire [16-1:0] node2771;
	wire [16-1:0] node2774;
	wire [16-1:0] node2775;
	wire [16-1:0] node2778;
	wire [16-1:0] node2781;
	wire [16-1:0] node2782;
	wire [16-1:0] node2784;
	wire [16-1:0] node2785;
	wire [16-1:0] node2788;
	wire [16-1:0] node2791;
	wire [16-1:0] node2792;
	wire [16-1:0] node2793;
	wire [16-1:0] node2795;
	wire [16-1:0] node2796;
	wire [16-1:0] node2801;
	wire [16-1:0] node2803;
	wire [16-1:0] node2804;
	wire [16-1:0] node2806;
	wire [16-1:0] node2810;
	wire [16-1:0] node2811;
	wire [16-1:0] node2812;
	wire [16-1:0] node2813;
	wire [16-1:0] node2814;
	wire [16-1:0] node2815;
	wire [16-1:0] node2817;
	wire [16-1:0] node2821;
	wire [16-1:0] node2822;
	wire [16-1:0] node2824;
	wire [16-1:0] node2827;
	wire [16-1:0] node2830;
	wire [16-1:0] node2831;
	wire [16-1:0] node2832;
	wire [16-1:0] node2833;
	wire [16-1:0] node2837;
	wire [16-1:0] node2838;
	wire [16-1:0] node2842;
	wire [16-1:0] node2843;
	wire [16-1:0] node2846;
	wire [16-1:0] node2848;
	wire [16-1:0] node2850;
	wire [16-1:0] node2853;
	wire [16-1:0] node2854;
	wire [16-1:0] node2855;
	wire [16-1:0] node2856;
	wire [16-1:0] node2857;
	wire [16-1:0] node2860;
	wire [16-1:0] node2862;
	wire [16-1:0] node2864;
	wire [16-1:0] node2867;
	wire [16-1:0] node2868;
	wire [16-1:0] node2872;
	wire [16-1:0] node2874;
	wire [16-1:0] node2875;
	wire [16-1:0] node2879;
	wire [16-1:0] node2880;
	wire [16-1:0] node2881;
	wire [16-1:0] node2882;
	wire [16-1:0] node2886;
	wire [16-1:0] node2889;
	wire [16-1:0] node2890;
	wire [16-1:0] node2891;
	wire [16-1:0] node2893;
	wire [16-1:0] node2897;
	wire [16-1:0] node2899;
	wire [16-1:0] node2901;
	wire [16-1:0] node2904;
	wire [16-1:0] node2905;
	wire [16-1:0] node2906;
	wire [16-1:0] node2907;
	wire [16-1:0] node2909;
	wire [16-1:0] node2910;
	wire [16-1:0] node2911;
	wire [16-1:0] node2916;
	wire [16-1:0] node2917;
	wire [16-1:0] node2918;
	wire [16-1:0] node2921;
	wire [16-1:0] node2923;
	wire [16-1:0] node2927;
	wire [16-1:0] node2928;
	wire [16-1:0] node2931;
	wire [16-1:0] node2932;
	wire [16-1:0] node2934;
	wire [16-1:0] node2937;
	wire [16-1:0] node2938;
	wire [16-1:0] node2942;
	wire [16-1:0] node2943;
	wire [16-1:0] node2944;
	wire [16-1:0] node2945;
	wire [16-1:0] node2946;
	wire [16-1:0] node2950;
	wire [16-1:0] node2953;
	wire [16-1:0] node2954;
	wire [16-1:0] node2955;
	wire [16-1:0] node2959;
	wire [16-1:0] node2960;
	wire [16-1:0] node2964;
	wire [16-1:0] node2965;
	wire [16-1:0] node2966;
	wire [16-1:0] node2967;
	wire [16-1:0] node2971;
	wire [16-1:0] node2973;
	wire [16-1:0] node2976;
	wire [16-1:0] node2977;
	wire [16-1:0] node2979;
	wire [16-1:0] node2981;
	wire [16-1:0] node2984;
	wire [16-1:0] node2986;
	wire [16-1:0] node2989;
	wire [16-1:0] node2990;
	wire [16-1:0] node2991;
	wire [16-1:0] node2992;
	wire [16-1:0] node2993;
	wire [16-1:0] node2994;
	wire [16-1:0] node2995;
	wire [16-1:0] node2996;
	wire [16-1:0] node2997;
	wire [16-1:0] node2998;
	wire [16-1:0] node2999;
	wire [16-1:0] node3000;
	wire [16-1:0] node3002;
	wire [16-1:0] node3006;
	wire [16-1:0] node3010;
	wire [16-1:0] node3011;
	wire [16-1:0] node3013;
	wire [16-1:0] node3014;
	wire [16-1:0] node3019;
	wire [16-1:0] node3020;
	wire [16-1:0] node3021;
	wire [16-1:0] node3022;
	wire [16-1:0] node3023;
	wire [16-1:0] node3027;
	wire [16-1:0] node3030;
	wire [16-1:0] node3032;
	wire [16-1:0] node3033;
	wire [16-1:0] node3037;
	wire [16-1:0] node3040;
	wire [16-1:0] node3041;
	wire [16-1:0] node3042;
	wire [16-1:0] node3043;
	wire [16-1:0] node3046;
	wire [16-1:0] node3047;
	wire [16-1:0] node3048;
	wire [16-1:0] node3053;
	wire [16-1:0] node3054;
	wire [16-1:0] node3055;
	wire [16-1:0] node3058;
	wire [16-1:0] node3061;
	wire [16-1:0] node3063;
	wire [16-1:0] node3066;
	wire [16-1:0] node3067;
	wire [16-1:0] node3068;
	wire [16-1:0] node3069;
	wire [16-1:0] node3071;
	wire [16-1:0] node3074;
	wire [16-1:0] node3076;
	wire [16-1:0] node3079;
	wire [16-1:0] node3082;
	wire [16-1:0] node3083;
	wire [16-1:0] node3084;
	wire [16-1:0] node3087;
	wire [16-1:0] node3088;
	wire [16-1:0] node3092;
	wire [16-1:0] node3095;
	wire [16-1:0] node3096;
	wire [16-1:0] node3097;
	wire [16-1:0] node3098;
	wire [16-1:0] node3099;
	wire [16-1:0] node3102;
	wire [16-1:0] node3103;
	wire [16-1:0] node3107;
	wire [16-1:0] node3108;
	wire [16-1:0] node3110;
	wire [16-1:0] node3113;
	wire [16-1:0] node3116;
	wire [16-1:0] node3117;
	wire [16-1:0] node3118;
	wire [16-1:0] node3119;
	wire [16-1:0] node3122;
	wire [16-1:0] node3123;
	wire [16-1:0] node3127;
	wire [16-1:0] node3130;
	wire [16-1:0] node3131;
	wire [16-1:0] node3134;
	wire [16-1:0] node3137;
	wire [16-1:0] node3138;
	wire [16-1:0] node3139;
	wire [16-1:0] node3140;
	wire [16-1:0] node3142;
	wire [16-1:0] node3143;
	wire [16-1:0] node3147;
	wire [16-1:0] node3150;
	wire [16-1:0] node3151;
	wire [16-1:0] node3152;
	wire [16-1:0] node3154;
	wire [16-1:0] node3158;
	wire [16-1:0] node3160;
	wire [16-1:0] node3163;
	wire [16-1:0] node3164;
	wire [16-1:0] node3165;
	wire [16-1:0] node3167;
	wire [16-1:0] node3170;
	wire [16-1:0] node3171;
	wire [16-1:0] node3174;
	wire [16-1:0] node3175;
	wire [16-1:0] node3179;
	wire [16-1:0] node3180;
	wire [16-1:0] node3181;
	wire [16-1:0] node3185;
	wire [16-1:0] node3187;
	wire [16-1:0] node3190;
	wire [16-1:0] node3191;
	wire [16-1:0] node3192;
	wire [16-1:0] node3193;
	wire [16-1:0] node3194;
	wire [16-1:0] node3195;
	wire [16-1:0] node3197;
	wire [16-1:0] node3201;
	wire [16-1:0] node3203;
	wire [16-1:0] node3204;
	wire [16-1:0] node3205;
	wire [16-1:0] node3206;
	wire [16-1:0] node3211;
	wire [16-1:0] node3214;
	wire [16-1:0] node3215;
	wire [16-1:0] node3216;
	wire [16-1:0] node3217;
	wire [16-1:0] node3220;
	wire [16-1:0] node3221;
	wire [16-1:0] node3225;
	wire [16-1:0] node3227;
	wire [16-1:0] node3228;
	wire [16-1:0] node3232;
	wire [16-1:0] node3233;
	wire [16-1:0] node3236;
	wire [16-1:0] node3237;
	wire [16-1:0] node3241;
	wire [16-1:0] node3242;
	wire [16-1:0] node3243;
	wire [16-1:0] node3246;
	wire [16-1:0] node3247;
	wire [16-1:0] node3248;
	wire [16-1:0] node3250;
	wire [16-1:0] node3254;
	wire [16-1:0] node3255;
	wire [16-1:0] node3259;
	wire [16-1:0] node3260;
	wire [16-1:0] node3261;
	wire [16-1:0] node3264;
	wire [16-1:0] node3267;
	wire [16-1:0] node3268;
	wire [16-1:0] node3269;
	wire [16-1:0] node3274;
	wire [16-1:0] node3275;
	wire [16-1:0] node3276;
	wire [16-1:0] node3277;
	wire [16-1:0] node3279;
	wire [16-1:0] node3280;
	wire [16-1:0] node3284;
	wire [16-1:0] node3285;
	wire [16-1:0] node3286;
	wire [16-1:0] node3287;
	wire [16-1:0] node3291;
	wire [16-1:0] node3294;
	wire [16-1:0] node3297;
	wire [16-1:0] node3298;
	wire [16-1:0] node3299;
	wire [16-1:0] node3302;
	wire [16-1:0] node3304;
	wire [16-1:0] node3307;
	wire [16-1:0] node3308;
	wire [16-1:0] node3311;
	wire [16-1:0] node3312;
	wire [16-1:0] node3316;
	wire [16-1:0] node3317;
	wire [16-1:0] node3318;
	wire [16-1:0] node3320;
	wire [16-1:0] node3322;
	wire [16-1:0] node3325;
	wire [16-1:0] node3328;
	wire [16-1:0] node3329;
	wire [16-1:0] node3330;
	wire [16-1:0] node3333;
	wire [16-1:0] node3335;
	wire [16-1:0] node3338;
	wire [16-1:0] node3339;
	wire [16-1:0] node3340;
	wire [16-1:0] node3343;
	wire [16-1:0] node3344;
	wire [16-1:0] node3349;
	wire [16-1:0] node3350;
	wire [16-1:0] node3351;
	wire [16-1:0] node3352;
	wire [16-1:0] node3353;
	wire [16-1:0] node3354;
	wire [16-1:0] node3355;
	wire [16-1:0] node3358;
	wire [16-1:0] node3361;
	wire [16-1:0] node3363;
	wire [16-1:0] node3366;
	wire [16-1:0] node3367;
	wire [16-1:0] node3368;
	wire [16-1:0] node3371;
	wire [16-1:0] node3374;
	wire [16-1:0] node3375;
	wire [16-1:0] node3379;
	wire [16-1:0] node3380;
	wire [16-1:0] node3381;
	wire [16-1:0] node3382;
	wire [16-1:0] node3384;
	wire [16-1:0] node3387;
	wire [16-1:0] node3388;
	wire [16-1:0] node3391;
	wire [16-1:0] node3392;
	wire [16-1:0] node3396;
	wire [16-1:0] node3397;
	wire [16-1:0] node3400;
	wire [16-1:0] node3401;
	wire [16-1:0] node3402;
	wire [16-1:0] node3407;
	wire [16-1:0] node3408;
	wire [16-1:0] node3411;
	wire [16-1:0] node3412;
	wire [16-1:0] node3413;
	wire [16-1:0] node3415;
	wire [16-1:0] node3417;
	wire [16-1:0] node3420;
	wire [16-1:0] node3421;
	wire [16-1:0] node3422;
	wire [16-1:0] node3425;
	wire [16-1:0] node3430;
	wire [16-1:0] node3431;
	wire [16-1:0] node3432;
	wire [16-1:0] node3433;
	wire [16-1:0] node3434;
	wire [16-1:0] node3435;
	wire [16-1:0] node3437;
	wire [16-1:0] node3440;
	wire [16-1:0] node3442;
	wire [16-1:0] node3444;
	wire [16-1:0] node3447;
	wire [16-1:0] node3450;
	wire [16-1:0] node3451;
	wire [16-1:0] node3453;
	wire [16-1:0] node3454;
	wire [16-1:0] node3459;
	wire [16-1:0] node3460;
	wire [16-1:0] node3461;
	wire [16-1:0] node3464;
	wire [16-1:0] node3465;
	wire [16-1:0] node3467;
	wire [16-1:0] node3471;
	wire [16-1:0] node3472;
	wire [16-1:0] node3473;
	wire [16-1:0] node3474;
	wire [16-1:0] node3479;
	wire [16-1:0] node3481;
	wire [16-1:0] node3483;
	wire [16-1:0] node3486;
	wire [16-1:0] node3487;
	wire [16-1:0] node3488;
	wire [16-1:0] node3489;
	wire [16-1:0] node3492;
	wire [16-1:0] node3493;
	wire [16-1:0] node3494;
	wire [16-1:0] node3498;
	wire [16-1:0] node3501;
	wire [16-1:0] node3502;
	wire [16-1:0] node3503;
	wire [16-1:0] node3505;
	wire [16-1:0] node3506;
	wire [16-1:0] node3511;
	wire [16-1:0] node3513;
	wire [16-1:0] node3514;
	wire [16-1:0] node3518;
	wire [16-1:0] node3519;
	wire [16-1:0] node3520;
	wire [16-1:0] node3521;
	wire [16-1:0] node3522;
	wire [16-1:0] node3526;
	wire [16-1:0] node3528;
	wire [16-1:0] node3531;
	wire [16-1:0] node3534;
	wire [16-1:0] node3536;
	wire [16-1:0] node3538;
	wire [16-1:0] node3541;
	wire [16-1:0] node3542;
	wire [16-1:0] node3543;
	wire [16-1:0] node3544;
	wire [16-1:0] node3545;
	wire [16-1:0] node3548;
	wire [16-1:0] node3549;
	wire [16-1:0] node3552;
	wire [16-1:0] node3554;
	wire [16-1:0] node3557;
	wire [16-1:0] node3558;
	wire [16-1:0] node3559;
	wire [16-1:0] node3560;
	wire [16-1:0] node3561;
	wire [16-1:0] node3566;
	wire [16-1:0] node3568;
	wire [16-1:0] node3571;
	wire [16-1:0] node3572;
	wire [16-1:0] node3573;
	wire [16-1:0] node3576;
	wire [16-1:0] node3580;
	wire [16-1:0] node3581;
	wire [16-1:0] node3582;
	wire [16-1:0] node3583;
	wire [16-1:0] node3586;
	wire [16-1:0] node3589;
	wire [16-1:0] node3590;
	wire [16-1:0] node3594;
	wire [16-1:0] node3595;
	wire [16-1:0] node3597;
	wire [16-1:0] node3598;
	wire [16-1:0] node3601;
	wire [16-1:0] node3604;
	wire [16-1:0] node3605;
	wire [16-1:0] node3606;
	wire [16-1:0] node3608;
	wire [16-1:0] node3610;
	wire [16-1:0] node3613;
	wire [16-1:0] node3616;
	wire [16-1:0] node3617;
	wire [16-1:0] node3620;
	wire [16-1:0] node3623;
	wire [16-1:0] node3624;
	wire [16-1:0] node3625;
	wire [16-1:0] node3626;
	wire [16-1:0] node3627;
	wire [16-1:0] node3631;
	wire [16-1:0] node3632;
	wire [16-1:0] node3633;
	wire [16-1:0] node3637;
	wire [16-1:0] node3639;
	wire [16-1:0] node3642;
	wire [16-1:0] node3643;
	wire [16-1:0] node3644;
	wire [16-1:0] node3647;
	wire [16-1:0] node3648;
	wire [16-1:0] node3651;
	wire [16-1:0] node3654;
	wire [16-1:0] node3655;
	wire [16-1:0] node3657;
	wire [16-1:0] node3661;
	wire [16-1:0] node3662;
	wire [16-1:0] node3663;
	wire [16-1:0] node3664;
	wire [16-1:0] node3665;
	wire [16-1:0] node3669;
	wire [16-1:0] node3670;
	wire [16-1:0] node3674;
	wire [16-1:0] node3675;
	wire [16-1:0] node3677;
	wire [16-1:0] node3678;
	wire [16-1:0] node3680;
	wire [16-1:0] node3684;
	wire [16-1:0] node3685;
	wire [16-1:0] node3689;
	wire [16-1:0] node3690;
	wire [16-1:0] node3692;
	wire [16-1:0] node3695;
	wire [16-1:0] node3696;
	wire [16-1:0] node3697;
	wire [16-1:0] node3699;
	wire [16-1:0] node3701;
	wire [16-1:0] node3705;
	wire [16-1:0] node3708;
	wire [16-1:0] node3709;
	wire [16-1:0] node3710;
	wire [16-1:0] node3711;
	wire [16-1:0] node3712;
	wire [16-1:0] node3713;
	wire [16-1:0] node3714;
	wire [16-1:0] node3715;
	wire [16-1:0] node3716;
	wire [16-1:0] node3721;
	wire [16-1:0] node3722;
	wire [16-1:0] node3723;
	wire [16-1:0] node3727;
	wire [16-1:0] node3730;
	wire [16-1:0] node3732;
	wire [16-1:0] node3733;
	wire [16-1:0] node3734;
	wire [16-1:0] node3736;
	wire [16-1:0] node3740;
	wire [16-1:0] node3743;
	wire [16-1:0] node3744;
	wire [16-1:0] node3745;
	wire [16-1:0] node3746;
	wire [16-1:0] node3747;
	wire [16-1:0] node3751;
	wire [16-1:0] node3754;
	wire [16-1:0] node3755;
	wire [16-1:0] node3756;
	wire [16-1:0] node3757;
	wire [16-1:0] node3762;
	wire [16-1:0] node3763;
	wire [16-1:0] node3764;
	wire [16-1:0] node3765;
	wire [16-1:0] node3770;
	wire [16-1:0] node3771;
	wire [16-1:0] node3773;
	wire [16-1:0] node3777;
	wire [16-1:0] node3778;
	wire [16-1:0] node3779;
	wire [16-1:0] node3781;
	wire [16-1:0] node3782;
	wire [16-1:0] node3784;
	wire [16-1:0] node3788;
	wire [16-1:0] node3791;
	wire [16-1:0] node3792;
	wire [16-1:0] node3794;
	wire [16-1:0] node3795;
	wire [16-1:0] node3799;
	wire [16-1:0] node3801;
	wire [16-1:0] node3803;
	wire [16-1:0] node3804;
	wire [16-1:0] node3808;
	wire [16-1:0] node3809;
	wire [16-1:0] node3810;
	wire [16-1:0] node3811;
	wire [16-1:0] node3812;
	wire [16-1:0] node3814;
	wire [16-1:0] node3815;
	wire [16-1:0] node3817;
	wire [16-1:0] node3821;
	wire [16-1:0] node3823;
	wire [16-1:0] node3826;
	wire [16-1:0] node3827;
	wire [16-1:0] node3828;
	wire [16-1:0] node3833;
	wire [16-1:0] node3834;
	wire [16-1:0] node3835;
	wire [16-1:0] node3836;
	wire [16-1:0] node3839;
	wire [16-1:0] node3840;
	wire [16-1:0] node3844;
	wire [16-1:0] node3845;
	wire [16-1:0] node3849;
	wire [16-1:0] node3851;
	wire [16-1:0] node3852;
	wire [16-1:0] node3855;
	wire [16-1:0] node3858;
	wire [16-1:0] node3859;
	wire [16-1:0] node3860;
	wire [16-1:0] node3861;
	wire [16-1:0] node3862;
	wire [16-1:0] node3866;
	wire [16-1:0] node3867;
	wire [16-1:0] node3869;
	wire [16-1:0] node3870;
	wire [16-1:0] node3875;
	wire [16-1:0] node3877;
	wire [16-1:0] node3880;
	wire [16-1:0] node3882;
	wire [16-1:0] node3883;
	wire [16-1:0] node3886;
	wire [16-1:0] node3887;
	wire [16-1:0] node3889;
	wire [16-1:0] node3893;
	wire [16-1:0] node3894;
	wire [16-1:0] node3895;
	wire [16-1:0] node3896;
	wire [16-1:0] node3897;
	wire [16-1:0] node3898;
	wire [16-1:0] node3899;
	wire [16-1:0] node3901;
	wire [16-1:0] node3904;
	wire [16-1:0] node3908;
	wire [16-1:0] node3909;
	wire [16-1:0] node3911;
	wire [16-1:0] node3914;
	wire [16-1:0] node3917;
	wire [16-1:0] node3918;
	wire [16-1:0] node3919;
	wire [16-1:0] node3922;
	wire [16-1:0] node3924;
	wire [16-1:0] node3927;
	wire [16-1:0] node3928;
	wire [16-1:0] node3930;
	wire [16-1:0] node3931;
	wire [16-1:0] node3933;
	wire [16-1:0] node3937;
	wire [16-1:0] node3939;
	wire [16-1:0] node3940;
	wire [16-1:0] node3944;
	wire [16-1:0] node3945;
	wire [16-1:0] node3946;
	wire [16-1:0] node3948;
	wire [16-1:0] node3950;
	wire [16-1:0] node3951;
	wire [16-1:0] node3955;
	wire [16-1:0] node3956;
	wire [16-1:0] node3957;
	wire [16-1:0] node3958;
	wire [16-1:0] node3963;
	wire [16-1:0] node3966;
	wire [16-1:0] node3967;
	wire [16-1:0] node3968;
	wire [16-1:0] node3971;
	wire [16-1:0] node3974;
	wire [16-1:0] node3975;
	wire [16-1:0] node3976;
	wire [16-1:0] node3980;
	wire [16-1:0] node3983;
	wire [16-1:0] node3984;
	wire [16-1:0] node3985;
	wire [16-1:0] node3986;
	wire [16-1:0] node3987;
	wire [16-1:0] node3988;
	wire [16-1:0] node3991;
	wire [16-1:0] node3993;
	wire [16-1:0] node3996;
	wire [16-1:0] node3998;
	wire [16-1:0] node3999;
	wire [16-1:0] node4001;
	wire [16-1:0] node4005;
	wire [16-1:0] node4006;
	wire [16-1:0] node4008;
	wire [16-1:0] node4009;
	wire [16-1:0] node4014;
	wire [16-1:0] node4015;
	wire [16-1:0] node4018;
	wire [16-1:0] node4019;
	wire [16-1:0] node4021;
	wire [16-1:0] node4024;
	wire [16-1:0] node4025;
	wire [16-1:0] node4028;
	wire [16-1:0] node4029;
	wire [16-1:0] node4033;
	wire [16-1:0] node4034;
	wire [16-1:0] node4035;
	wire [16-1:0] node4036;
	wire [16-1:0] node4037;
	wire [16-1:0] node4039;
	wire [16-1:0] node4043;
	wire [16-1:0] node4046;
	wire [16-1:0] node4047;
	wire [16-1:0] node4050;
	wire [16-1:0] node4051;
	wire [16-1:0] node4054;
	wire [16-1:0] node4055;
	wire [16-1:0] node4059;
	wire [16-1:0] node4060;
	wire [16-1:0] node4061;
	wire [16-1:0] node4064;
	wire [16-1:0] node4066;
	wire [16-1:0] node4067;
	wire [16-1:0] node4071;
	wire [16-1:0] node4072;
	wire [16-1:0] node4074;
	wire [16-1:0] node4075;
	wire [16-1:0] node4076;
	wire [16-1:0] node4081;
	wire [16-1:0] node4083;
	wire [16-1:0] node4084;
	wire [16-1:0] node4085;
	wire [16-1:0] node4090;
	wire [16-1:0] node4091;
	wire [16-1:0] node4092;
	wire [16-1:0] node4093;
	wire [16-1:0] node4094;
	wire [16-1:0] node4095;
	wire [16-1:0] node4096;
	wire [16-1:0] node4098;
	wire [16-1:0] node4099;
	wire [16-1:0] node4101;
	wire [16-1:0] node4105;
	wire [16-1:0] node4106;
	wire [16-1:0] node4108;
	wire [16-1:0] node4112;
	wire [16-1:0] node4113;
	wire [16-1:0] node4114;
	wire [16-1:0] node4116;
	wire [16-1:0] node4120;
	wire [16-1:0] node4121;
	wire [16-1:0] node4123;
	wire [16-1:0] node4126;
	wire [16-1:0] node4129;
	wire [16-1:0] node4130;
	wire [16-1:0] node4131;
	wire [16-1:0] node4134;
	wire [16-1:0] node4135;
	wire [16-1:0] node4136;
	wire [16-1:0] node4140;
	wire [16-1:0] node4142;
	wire [16-1:0] node4145;
	wire [16-1:0] node4146;
	wire [16-1:0] node4147;
	wire [16-1:0] node4151;
	wire [16-1:0] node4154;
	wire [16-1:0] node4155;
	wire [16-1:0] node4156;
	wire [16-1:0] node4158;
	wire [16-1:0] node4161;
	wire [16-1:0] node4162;
	wire [16-1:0] node4164;
	wire [16-1:0] node4167;
	wire [16-1:0] node4169;
	wire [16-1:0] node4170;
	wire [16-1:0] node4174;
	wire [16-1:0] node4175;
	wire [16-1:0] node4177;
	wire [16-1:0] node4178;
	wire [16-1:0] node4182;
	wire [16-1:0] node4183;
	wire [16-1:0] node4186;
	wire [16-1:0] node4188;
	wire [16-1:0] node4189;
	wire [16-1:0] node4193;
	wire [16-1:0] node4194;
	wire [16-1:0] node4195;
	wire [16-1:0] node4196;
	wire [16-1:0] node4198;
	wire [16-1:0] node4199;
	wire [16-1:0] node4203;
	wire [16-1:0] node4204;
	wire [16-1:0] node4208;
	wire [16-1:0] node4209;
	wire [16-1:0] node4211;
	wire [16-1:0] node4212;
	wire [16-1:0] node4215;
	wire [16-1:0] node4216;
	wire [16-1:0] node4220;
	wire [16-1:0] node4221;
	wire [16-1:0] node4222;
	wire [16-1:0] node4226;
	wire [16-1:0] node4229;
	wire [16-1:0] node4230;
	wire [16-1:0] node4231;
	wire [16-1:0] node4233;
	wire [16-1:0] node4236;
	wire [16-1:0] node4237;
	wire [16-1:0] node4241;
	wire [16-1:0] node4242;
	wire [16-1:0] node4243;
	wire [16-1:0] node4244;
	wire [16-1:0] node4249;
	wire [16-1:0] node4250;
	wire [16-1:0] node4251;
	wire [16-1:0] node4255;
	wire [16-1:0] node4256;
	wire [16-1:0] node4257;
	wire [16-1:0] node4262;
	wire [16-1:0] node4263;
	wire [16-1:0] node4264;
	wire [16-1:0] node4265;
	wire [16-1:0] node4266;
	wire [16-1:0] node4267;
	wire [16-1:0] node4270;
	wire [16-1:0] node4271;
	wire [16-1:0] node4273;
	wire [16-1:0] node4276;
	wire [16-1:0] node4279;
	wire [16-1:0] node4280;
	wire [16-1:0] node4282;
	wire [16-1:0] node4283;
	wire [16-1:0] node4287;
	wire [16-1:0] node4288;
	wire [16-1:0] node4291;
	wire [16-1:0] node4294;
	wire [16-1:0] node4295;
	wire [16-1:0] node4296;
	wire [16-1:0] node4298;
	wire [16-1:0] node4301;
	wire [16-1:0] node4303;
	wire [16-1:0] node4306;
	wire [16-1:0] node4307;
	wire [16-1:0] node4309;
	wire [16-1:0] node4312;
	wire [16-1:0] node4314;
	wire [16-1:0] node4317;
	wire [16-1:0] node4318;
	wire [16-1:0] node4319;
	wire [16-1:0] node4320;
	wire [16-1:0] node4321;
	wire [16-1:0] node4325;
	wire [16-1:0] node4328;
	wire [16-1:0] node4329;
	wire [16-1:0] node4333;
	wire [16-1:0] node4334;
	wire [16-1:0] node4335;
	wire [16-1:0] node4338;
	wire [16-1:0] node4340;
	wire [16-1:0] node4343;
	wire [16-1:0] node4344;
	wire [16-1:0] node4347;
	wire [16-1:0] node4348;
	wire [16-1:0] node4350;
	wire [16-1:0] node4354;
	wire [16-1:0] node4355;
	wire [16-1:0] node4356;
	wire [16-1:0] node4357;
	wire [16-1:0] node4358;
	wire [16-1:0] node4360;
	wire [16-1:0] node4363;
	wire [16-1:0] node4366;
	wire [16-1:0] node4367;
	wire [16-1:0] node4370;
	wire [16-1:0] node4372;
	wire [16-1:0] node4375;
	wire [16-1:0] node4376;
	wire [16-1:0] node4377;
	wire [16-1:0] node4378;
	wire [16-1:0] node4380;
	wire [16-1:0] node4385;
	wire [16-1:0] node4386;
	wire [16-1:0] node4387;
	wire [16-1:0] node4389;
	wire [16-1:0] node4393;
	wire [16-1:0] node4394;
	wire [16-1:0] node4398;
	wire [16-1:0] node4399;
	wire [16-1:0] node4400;
	wire [16-1:0] node4401;
	wire [16-1:0] node4405;
	wire [16-1:0] node4407;
	wire [16-1:0] node4408;
	wire [16-1:0] node4409;
	wire [16-1:0] node4410;
	wire [16-1:0] node4414;
	wire [16-1:0] node4418;
	wire [16-1:0] node4419;
	wire [16-1:0] node4420;
	wire [16-1:0] node4423;
	wire [16-1:0] node4424;
	wire [16-1:0] node4426;
	wire [16-1:0] node4429;
	wire [16-1:0] node4432;
	wire [16-1:0] node4433;
	wire [16-1:0] node4434;
	wire [16-1:0] node4437;
	wire [16-1:0] node4439;
	wire [16-1:0] node4442;
	wire [16-1:0] node4443;
	wire [16-1:0] node4446;
	wire [16-1:0] node4448;
	wire [16-1:0] node4451;
	wire [16-1:0] node4452;
	wire [16-1:0] node4453;
	wire [16-1:0] node4454;
	wire [16-1:0] node4455;
	wire [16-1:0] node4456;
	wire [16-1:0] node4457;
	wire [16-1:0] node4458;
	wire [16-1:0] node4459;
	wire [16-1:0] node4460;
	wire [16-1:0] node4462;
	wire [16-1:0] node4467;
	wire [16-1:0] node4468;
	wire [16-1:0] node4469;
	wire [16-1:0] node4470;
	wire [16-1:0] node4474;
	wire [16-1:0] node4477;
	wire [16-1:0] node4478;
	wire [16-1:0] node4482;
	wire [16-1:0] node4483;
	wire [16-1:0] node4484;
	wire [16-1:0] node4486;
	wire [16-1:0] node4487;
	wire [16-1:0] node4489;
	wire [16-1:0] node4493;
	wire [16-1:0] node4496;
	wire [16-1:0] node4497;
	wire [16-1:0] node4498;
	wire [16-1:0] node4499;
	wire [16-1:0] node4503;
	wire [16-1:0] node4505;
	wire [16-1:0] node4509;
	wire [16-1:0] node4510;
	wire [16-1:0] node4511;
	wire [16-1:0] node4512;
	wire [16-1:0] node4515;
	wire [16-1:0] node4518;
	wire [16-1:0] node4519;
	wire [16-1:0] node4520;
	wire [16-1:0] node4524;
	wire [16-1:0] node4525;
	wire [16-1:0] node4529;
	wire [16-1:0] node4530;
	wire [16-1:0] node4531;
	wire [16-1:0] node4533;
	wire [16-1:0] node4535;
	wire [16-1:0] node4538;
	wire [16-1:0] node4539;
	wire [16-1:0] node4543;
	wire [16-1:0] node4544;
	wire [16-1:0] node4546;
	wire [16-1:0] node4548;
	wire [16-1:0] node4549;
	wire [16-1:0] node4554;
	wire [16-1:0] node4555;
	wire [16-1:0] node4556;
	wire [16-1:0] node4557;
	wire [16-1:0] node4558;
	wire [16-1:0] node4560;
	wire [16-1:0] node4562;
	wire [16-1:0] node4565;
	wire [16-1:0] node4568;
	wire [16-1:0] node4569;
	wire [16-1:0] node4572;
	wire [16-1:0] node4573;
	wire [16-1:0] node4576;
	wire [16-1:0] node4578;
	wire [16-1:0] node4581;
	wire [16-1:0] node4582;
	wire [16-1:0] node4583;
	wire [16-1:0] node4584;
	wire [16-1:0] node4588;
	wire [16-1:0] node4590;
	wire [16-1:0] node4593;
	wire [16-1:0] node4594;
	wire [16-1:0] node4596;
	wire [16-1:0] node4597;
	wire [16-1:0] node4601;
	wire [16-1:0] node4603;
	wire [16-1:0] node4606;
	wire [16-1:0] node4607;
	wire [16-1:0] node4608;
	wire [16-1:0] node4609;
	wire [16-1:0] node4611;
	wire [16-1:0] node4614;
	wire [16-1:0] node4616;
	wire [16-1:0] node4619;
	wire [16-1:0] node4621;
	wire [16-1:0] node4622;
	wire [16-1:0] node4623;
	wire [16-1:0] node4628;
	wire [16-1:0] node4629;
	wire [16-1:0] node4630;
	wire [16-1:0] node4631;
	wire [16-1:0] node4635;
	wire [16-1:0] node4636;
	wire [16-1:0] node4640;
	wire [16-1:0] node4641;
	wire [16-1:0] node4644;
	wire [16-1:0] node4645;
	wire [16-1:0] node4649;
	wire [16-1:0] node4650;
	wire [16-1:0] node4651;
	wire [16-1:0] node4652;
	wire [16-1:0] node4653;
	wire [16-1:0] node4654;
	wire [16-1:0] node4657;
	wire [16-1:0] node4660;
	wire [16-1:0] node4661;
	wire [16-1:0] node4664;
	wire [16-1:0] node4665;
	wire [16-1:0] node4667;
	wire [16-1:0] node4671;
	wire [16-1:0] node4672;
	wire [16-1:0] node4673;
	wire [16-1:0] node4677;
	wire [16-1:0] node4678;
	wire [16-1:0] node4682;
	wire [16-1:0] node4683;
	wire [16-1:0] node4684;
	wire [16-1:0] node4685;
	wire [16-1:0] node4687;
	wire [16-1:0] node4688;
	wire [16-1:0] node4693;
	wire [16-1:0] node4694;
	wire [16-1:0] node4697;
	wire [16-1:0] node4700;
	wire [16-1:0] node4701;
	wire [16-1:0] node4702;
	wire [16-1:0] node4704;
	wire [16-1:0] node4705;
	wire [16-1:0] node4709;
	wire [16-1:0] node4710;
	wire [16-1:0] node4712;
	wire [16-1:0] node4716;
	wire [16-1:0] node4717;
	wire [16-1:0] node4719;
	wire [16-1:0] node4722;
	wire [16-1:0] node4723;
	wire [16-1:0] node4724;
	wire [16-1:0] node4728;
	wire [16-1:0] node4731;
	wire [16-1:0] node4732;
	wire [16-1:0] node4733;
	wire [16-1:0] node4734;
	wire [16-1:0] node4735;
	wire [16-1:0] node4738;
	wire [16-1:0] node4739;
	wire [16-1:0] node4743;
	wire [16-1:0] node4744;
	wire [16-1:0] node4748;
	wire [16-1:0] node4749;
	wire [16-1:0] node4750;
	wire [16-1:0] node4751;
	wire [16-1:0] node4752;
	wire [16-1:0] node4756;
	wire [16-1:0] node4759;
	wire [16-1:0] node4760;
	wire [16-1:0] node4763;
	wire [16-1:0] node4766;
	wire [16-1:0] node4768;
	wire [16-1:0] node4771;
	wire [16-1:0] node4772;
	wire [16-1:0] node4773;
	wire [16-1:0] node4774;
	wire [16-1:0] node4776;
	wire [16-1:0] node4779;
	wire [16-1:0] node4782;
	wire [16-1:0] node4783;
	wire [16-1:0] node4784;
	wire [16-1:0] node4786;
	wire [16-1:0] node4789;
	wire [16-1:0] node4791;
	wire [16-1:0] node4794;
	wire [16-1:0] node4795;
	wire [16-1:0] node4799;
	wire [16-1:0] node4800;
	wire [16-1:0] node4801;
	wire [16-1:0] node4804;
	wire [16-1:0] node4805;
	wire [16-1:0] node4807;
	wire [16-1:0] node4808;
	wire [16-1:0] node4812;
	wire [16-1:0] node4815;
	wire [16-1:0] node4816;
	wire [16-1:0] node4819;
	wire [16-1:0] node4820;
	wire [16-1:0] node4821;
	wire [16-1:0] node4825;
	wire [16-1:0] node4827;
	wire [16-1:0] node4830;
	wire [16-1:0] node4831;
	wire [16-1:0] node4832;
	wire [16-1:0] node4833;
	wire [16-1:0] node4834;
	wire [16-1:0] node4835;
	wire [16-1:0] node4837;
	wire [16-1:0] node4839;
	wire [16-1:0] node4842;
	wire [16-1:0] node4843;
	wire [16-1:0] node4844;
	wire [16-1:0] node4848;
	wire [16-1:0] node4851;
	wire [16-1:0] node4852;
	wire [16-1:0] node4853;
	wire [16-1:0] node4854;
	wire [16-1:0] node4858;
	wire [16-1:0] node4859;
	wire [16-1:0] node4863;
	wire [16-1:0] node4864;
	wire [16-1:0] node4868;
	wire [16-1:0] node4869;
	wire [16-1:0] node4870;
	wire [16-1:0] node4871;
	wire [16-1:0] node4875;
	wire [16-1:0] node4876;
	wire [16-1:0] node4878;
	wire [16-1:0] node4879;
	wire [16-1:0] node4883;
	wire [16-1:0] node4886;
	wire [16-1:0] node4887;
	wire [16-1:0] node4888;
	wire [16-1:0] node4889;
	wire [16-1:0] node4891;
	wire [16-1:0] node4895;
	wire [16-1:0] node4897;
	wire [16-1:0] node4898;
	wire [16-1:0] node4902;
	wire [16-1:0] node4903;
	wire [16-1:0] node4904;
	wire [16-1:0] node4906;
	wire [16-1:0] node4909;
	wire [16-1:0] node4910;
	wire [16-1:0] node4913;
	wire [16-1:0] node4916;
	wire [16-1:0] node4917;
	wire [16-1:0] node4921;
	wire [16-1:0] node4922;
	wire [16-1:0] node4923;
	wire [16-1:0] node4924;
	wire [16-1:0] node4925;
	wire [16-1:0] node4926;
	wire [16-1:0] node4930;
	wire [16-1:0] node4933;
	wire [16-1:0] node4934;
	wire [16-1:0] node4935;
	wire [16-1:0] node4939;
	wire [16-1:0] node4940;
	wire [16-1:0] node4943;
	wire [16-1:0] node4946;
	wire [16-1:0] node4947;
	wire [16-1:0] node4948;
	wire [16-1:0] node4951;
	wire [16-1:0] node4954;
	wire [16-1:0] node4955;
	wire [16-1:0] node4959;
	wire [16-1:0] node4960;
	wire [16-1:0] node4961;
	wire [16-1:0] node4962;
	wire [16-1:0] node4964;
	wire [16-1:0] node4968;
	wire [16-1:0] node4969;
	wire [16-1:0] node4970;
	wire [16-1:0] node4971;
	wire [16-1:0] node4976;
	wire [16-1:0] node4977;
	wire [16-1:0] node4980;
	wire [16-1:0] node4982;
	wire [16-1:0] node4985;
	wire [16-1:0] node4986;
	wire [16-1:0] node4987;
	wire [16-1:0] node4989;
	wire [16-1:0] node4992;
	wire [16-1:0] node4993;
	wire [16-1:0] node4995;
	wire [16-1:0] node4999;
	wire [16-1:0] node5001;
	wire [16-1:0] node5003;
	wire [16-1:0] node5004;
	wire [16-1:0] node5008;
	wire [16-1:0] node5009;
	wire [16-1:0] node5010;
	wire [16-1:0] node5011;
	wire [16-1:0] node5012;
	wire [16-1:0] node5013;
	wire [16-1:0] node5017;
	wire [16-1:0] node5018;
	wire [16-1:0] node5022;
	wire [16-1:0] node5023;
	wire [16-1:0] node5024;
	wire [16-1:0] node5026;
	wire [16-1:0] node5030;
	wire [16-1:0] node5031;
	wire [16-1:0] node5034;
	wire [16-1:0] node5036;
	wire [16-1:0] node5038;
	wire [16-1:0] node5041;
	wire [16-1:0] node5042;
	wire [16-1:0] node5043;
	wire [16-1:0] node5044;
	wire [16-1:0] node5046;
	wire [16-1:0] node5047;
	wire [16-1:0] node5051;
	wire [16-1:0] node5053;
	wire [16-1:0] node5056;
	wire [16-1:0] node5057;
	wire [16-1:0] node5058;
	wire [16-1:0] node5062;
	wire [16-1:0] node5065;
	wire [16-1:0] node5066;
	wire [16-1:0] node5068;
	wire [16-1:0] node5069;
	wire [16-1:0] node5071;
	wire [16-1:0] node5075;
	wire [16-1:0] node5077;
	wire [16-1:0] node5078;
	wire [16-1:0] node5080;
	wire [16-1:0] node5083;
	wire [16-1:0] node5086;
	wire [16-1:0] node5087;
	wire [16-1:0] node5088;
	wire [16-1:0] node5089;
	wire [16-1:0] node5091;
	wire [16-1:0] node5094;
	wire [16-1:0] node5095;
	wire [16-1:0] node5096;
	wire [16-1:0] node5099;
	wire [16-1:0] node5102;
	wire [16-1:0] node5103;
	wire [16-1:0] node5107;
	wire [16-1:0] node5108;
	wire [16-1:0] node5109;
	wire [16-1:0] node5112;
	wire [16-1:0] node5114;
	wire [16-1:0] node5115;
	wire [16-1:0] node5118;
	wire [16-1:0] node5121;
	wire [16-1:0] node5122;
	wire [16-1:0] node5125;
	wire [16-1:0] node5126;
	wire [16-1:0] node5130;
	wire [16-1:0] node5131;
	wire [16-1:0] node5132;
	wire [16-1:0] node5133;
	wire [16-1:0] node5137;
	wire [16-1:0] node5138;
	wire [16-1:0] node5139;
	wire [16-1:0] node5141;
	wire [16-1:0] node5145;
	wire [16-1:0] node5147;
	wire [16-1:0] node5150;
	wire [16-1:0] node5151;
	wire [16-1:0] node5153;
	wire [16-1:0] node5154;
	wire [16-1:0] node5155;
	wire [16-1:0] node5160;
	wire [16-1:0] node5161;
	wire [16-1:0] node5163;
	wire [16-1:0] node5165;
	wire [16-1:0] node5168;
	wire [16-1:0] node5171;
	wire [16-1:0] node5172;
	wire [16-1:0] node5173;
	wire [16-1:0] node5174;
	wire [16-1:0] node5175;
	wire [16-1:0] node5176;
	wire [16-1:0] node5177;
	wire [16-1:0] node5178;
	wire [16-1:0] node5181;
	wire [16-1:0] node5183;
	wire [16-1:0] node5186;
	wire [16-1:0] node5187;
	wire [16-1:0] node5190;
	wire [16-1:0] node5192;
	wire [16-1:0] node5195;
	wire [16-1:0] node5196;
	wire [16-1:0] node5197;
	wire [16-1:0] node5198;
	wire [16-1:0] node5199;
	wire [16-1:0] node5204;
	wire [16-1:0] node5206;
	wire [16-1:0] node5209;
	wire [16-1:0] node5210;
	wire [16-1:0] node5213;
	wire [16-1:0] node5216;
	wire [16-1:0] node5217;
	wire [16-1:0] node5218;
	wire [16-1:0] node5220;
	wire [16-1:0] node5223;
	wire [16-1:0] node5225;
	wire [16-1:0] node5226;
	wire [16-1:0] node5228;
	wire [16-1:0] node5232;
	wire [16-1:0] node5233;
	wire [16-1:0] node5234;
	wire [16-1:0] node5237;
	wire [16-1:0] node5239;
	wire [16-1:0] node5240;
	wire [16-1:0] node5244;
	wire [16-1:0] node5245;
	wire [16-1:0] node5246;
	wire [16-1:0] node5248;
	wire [16-1:0] node5251;
	wire [16-1:0] node5253;
	wire [16-1:0] node5256;
	wire [16-1:0] node5259;
	wire [16-1:0] node5260;
	wire [16-1:0] node5261;
	wire [16-1:0] node5262;
	wire [16-1:0] node5264;
	wire [16-1:0] node5265;
	wire [16-1:0] node5269;
	wire [16-1:0] node5270;
	wire [16-1:0] node5273;
	wire [16-1:0] node5276;
	wire [16-1:0] node5277;
	wire [16-1:0] node5278;
	wire [16-1:0] node5283;
	wire [16-1:0] node5284;
	wire [16-1:0] node5285;
	wire [16-1:0] node5287;
	wire [16-1:0] node5288;
	wire [16-1:0] node5290;
	wire [16-1:0] node5293;
	wire [16-1:0] node5296;
	wire [16-1:0] node5297;
	wire [16-1:0] node5298;
	wire [16-1:0] node5300;
	wire [16-1:0] node5304;
	wire [16-1:0] node5306;
	wire [16-1:0] node5307;
	wire [16-1:0] node5310;
	wire [16-1:0] node5313;
	wire [16-1:0] node5314;
	wire [16-1:0] node5315;
	wire [16-1:0] node5316;
	wire [16-1:0] node5318;
	wire [16-1:0] node5319;
	wire [16-1:0] node5324;
	wire [16-1:0] node5327;
	wire [16-1:0] node5328;
	wire [16-1:0] node5329;
	wire [16-1:0] node5332;
	wire [16-1:0] node5335;
	wire [16-1:0] node5336;
	wire [16-1:0] node5337;
	wire [16-1:0] node5340;
	wire [16-1:0] node5343;
	wire [16-1:0] node5346;
	wire [16-1:0] node5347;
	wire [16-1:0] node5348;
	wire [16-1:0] node5349;
	wire [16-1:0] node5350;
	wire [16-1:0] node5351;
	wire [16-1:0] node5352;
	wire [16-1:0] node5353;
	wire [16-1:0] node5358;
	wire [16-1:0] node5359;
	wire [16-1:0] node5363;
	wire [16-1:0] node5366;
	wire [16-1:0] node5367;
	wire [16-1:0] node5368;
	wire [16-1:0] node5369;
	wire [16-1:0] node5372;
	wire [16-1:0] node5373;
	wire [16-1:0] node5375;
	wire [16-1:0] node5378;
	wire [16-1:0] node5381;
	wire [16-1:0] node5382;
	wire [16-1:0] node5386;
	wire [16-1:0] node5387;
	wire [16-1:0] node5390;
	wire [16-1:0] node5392;
	wire [16-1:0] node5395;
	wire [16-1:0] node5396;
	wire [16-1:0] node5397;
	wire [16-1:0] node5398;
	wire [16-1:0] node5402;
	wire [16-1:0] node5403;
	wire [16-1:0] node5404;
	wire [16-1:0] node5406;
	wire [16-1:0] node5410;
	wire [16-1:0] node5411;
	wire [16-1:0] node5413;
	wire [16-1:0] node5416;
	wire [16-1:0] node5419;
	wire [16-1:0] node5420;
	wire [16-1:0] node5421;
	wire [16-1:0] node5424;
	wire [16-1:0] node5425;
	wire [16-1:0] node5427;
	wire [16-1:0] node5429;
	wire [16-1:0] node5433;
	wire [16-1:0] node5434;
	wire [16-1:0] node5438;
	wire [16-1:0] node5439;
	wire [16-1:0] node5440;
	wire [16-1:0] node5441;
	wire [16-1:0] node5442;
	wire [16-1:0] node5443;
	wire [16-1:0] node5444;
	wire [16-1:0] node5449;
	wire [16-1:0] node5452;
	wire [16-1:0] node5453;
	wire [16-1:0] node5456;
	wire [16-1:0] node5459;
	wire [16-1:0] node5460;
	wire [16-1:0] node5461;
	wire [16-1:0] node5464;
	wire [16-1:0] node5466;
	wire [16-1:0] node5467;
	wire [16-1:0] node5471;
	wire [16-1:0] node5472;
	wire [16-1:0] node5473;
	wire [16-1:0] node5474;
	wire [16-1:0] node5476;
	wire [16-1:0] node5479;
	wire [16-1:0] node5483;
	wire [16-1:0] node5484;
	wire [16-1:0] node5487;
	wire [16-1:0] node5488;
	wire [16-1:0] node5490;
	wire [16-1:0] node5493;
	wire [16-1:0] node5496;
	wire [16-1:0] node5497;
	wire [16-1:0] node5498;
	wire [16-1:0] node5499;
	wire [16-1:0] node5500;
	wire [16-1:0] node5504;
	wire [16-1:0] node5505;
	wire [16-1:0] node5509;
	wire [16-1:0] node5510;
	wire [16-1:0] node5511;
	wire [16-1:0] node5515;
	wire [16-1:0] node5518;
	wire [16-1:0] node5519;
	wire [16-1:0] node5520;
	wire [16-1:0] node5522;
	wire [16-1:0] node5524;
	wire [16-1:0] node5527;
	wire [16-1:0] node5530;
	wire [16-1:0] node5532;
	wire [16-1:0] node5535;
	wire [16-1:0] node5536;
	wire [16-1:0] node5537;
	wire [16-1:0] node5538;
	wire [16-1:0] node5539;
	wire [16-1:0] node5540;
	wire [16-1:0] node5541;
	wire [16-1:0] node5542;
	wire [16-1:0] node5543;
	wire [16-1:0] node5544;
	wire [16-1:0] node5549;
	wire [16-1:0] node5552;
	wire [16-1:0] node5553;
	wire [16-1:0] node5556;
	wire [16-1:0] node5559;
	wire [16-1:0] node5560;
	wire [16-1:0] node5562;
	wire [16-1:0] node5565;
	wire [16-1:0] node5568;
	wire [16-1:0] node5569;
	wire [16-1:0] node5571;
	wire [16-1:0] node5574;
	wire [16-1:0] node5575;
	wire [16-1:0] node5578;
	wire [16-1:0] node5581;
	wire [16-1:0] node5582;
	wire [16-1:0] node5583;
	wire [16-1:0] node5584;
	wire [16-1:0] node5586;
	wire [16-1:0] node5587;
	wire [16-1:0] node5591;
	wire [16-1:0] node5593;
	wire [16-1:0] node5596;
	wire [16-1:0] node5597;
	wire [16-1:0] node5598;
	wire [16-1:0] node5599;
	wire [16-1:0] node5600;
	wire [16-1:0] node5604;
	wire [16-1:0] node5608;
	wire [16-1:0] node5610;
	wire [16-1:0] node5613;
	wire [16-1:0] node5614;
	wire [16-1:0] node5616;
	wire [16-1:0] node5618;
	wire [16-1:0] node5621;
	wire [16-1:0] node5622;
	wire [16-1:0] node5625;
	wire [16-1:0] node5626;
	wire [16-1:0] node5629;
	wire [16-1:0] node5631;
	wire [16-1:0] node5634;
	wire [16-1:0] node5635;
	wire [16-1:0] node5636;
	wire [16-1:0] node5637;
	wire [16-1:0] node5638;
	wire [16-1:0] node5641;
	wire [16-1:0] node5644;
	wire [16-1:0] node5645;
	wire [16-1:0] node5646;
	wire [16-1:0] node5647;
	wire [16-1:0] node5652;
	wire [16-1:0] node5653;
	wire [16-1:0] node5657;
	wire [16-1:0] node5658;
	wire [16-1:0] node5659;
	wire [16-1:0] node5662;
	wire [16-1:0] node5664;
	wire [16-1:0] node5665;
	wire [16-1:0] node5668;
	wire [16-1:0] node5670;
	wire [16-1:0] node5673;
	wire [16-1:0] node5676;
	wire [16-1:0] node5677;
	wire [16-1:0] node5678;
	wire [16-1:0] node5680;
	wire [16-1:0] node5682;
	wire [16-1:0] node5685;
	wire [16-1:0] node5686;
	wire [16-1:0] node5688;
	wire [16-1:0] node5689;
	wire [16-1:0] node5692;
	wire [16-1:0] node5696;
	wire [16-1:0] node5697;
	wire [16-1:0] node5698;
	wire [16-1:0] node5699;
	wire [16-1:0] node5703;
	wire [16-1:0] node5705;
	wire [16-1:0] node5708;
	wire [16-1:0] node5709;
	wire [16-1:0] node5710;
	wire [16-1:0] node5712;
	wire [16-1:0] node5716;
	wire [16-1:0] node5717;
	wire [16-1:0] node5719;
	wire [16-1:0] node5723;
	wire [16-1:0] node5724;
	wire [16-1:0] node5725;
	wire [16-1:0] node5726;
	wire [16-1:0] node5727;
	wire [16-1:0] node5728;
	wire [16-1:0] node5729;
	wire [16-1:0] node5733;
	wire [16-1:0] node5736;
	wire [16-1:0] node5737;
	wire [16-1:0] node5738;
	wire [16-1:0] node5741;
	wire [16-1:0] node5744;
	wire [16-1:0] node5745;
	wire [16-1:0] node5746;
	wire [16-1:0] node5750;
	wire [16-1:0] node5751;
	wire [16-1:0] node5754;
	wire [16-1:0] node5757;
	wire [16-1:0] node5758;
	wire [16-1:0] node5759;
	wire [16-1:0] node5760;
	wire [16-1:0] node5762;
	wire [16-1:0] node5764;
	wire [16-1:0] node5767;
	wire [16-1:0] node5769;
	wire [16-1:0] node5772;
	wire [16-1:0] node5774;
	wire [16-1:0] node5777;
	wire [16-1:0] node5778;
	wire [16-1:0] node5779;
	wire [16-1:0] node5783;
	wire [16-1:0] node5786;
	wire [16-1:0] node5787;
	wire [16-1:0] node5788;
	wire [16-1:0] node5789;
	wire [16-1:0] node5790;
	wire [16-1:0] node5793;
	wire [16-1:0] node5795;
	wire [16-1:0] node5798;
	wire [16-1:0] node5799;
	wire [16-1:0] node5801;
	wire [16-1:0] node5802;
	wire [16-1:0] node5807;
	wire [16-1:0] node5808;
	wire [16-1:0] node5810;
	wire [16-1:0] node5813;
	wire [16-1:0] node5815;
	wire [16-1:0] node5817;
	wire [16-1:0] node5820;
	wire [16-1:0] node5821;
	wire [16-1:0] node5822;
	wire [16-1:0] node5824;
	wire [16-1:0] node5826;
	wire [16-1:0] node5829;
	wire [16-1:0] node5830;
	wire [16-1:0] node5834;
	wire [16-1:0] node5835;
	wire [16-1:0] node5837;
	wire [16-1:0] node5839;
	wire [16-1:0] node5842;
	wire [16-1:0] node5845;
	wire [16-1:0] node5846;
	wire [16-1:0] node5847;
	wire [16-1:0] node5848;
	wire [16-1:0] node5849;
	wire [16-1:0] node5850;
	wire [16-1:0] node5851;
	wire [16-1:0] node5856;
	wire [16-1:0] node5857;
	wire [16-1:0] node5861;
	wire [16-1:0] node5862;
	wire [16-1:0] node5865;
	wire [16-1:0] node5867;
	wire [16-1:0] node5869;
	wire [16-1:0] node5872;
	wire [16-1:0] node5873;
	wire [16-1:0] node5874;
	wire [16-1:0] node5875;
	wire [16-1:0] node5879;
	wire [16-1:0] node5882;
	wire [16-1:0] node5883;
	wire [16-1:0] node5884;
	wire [16-1:0] node5887;
	wire [16-1:0] node5890;
	wire [16-1:0] node5891;
	wire [16-1:0] node5894;
	wire [16-1:0] node5897;
	wire [16-1:0] node5898;
	wire [16-1:0] node5899;
	wire [16-1:0] node5900;
	wire [16-1:0] node5901;
	wire [16-1:0] node5905;
	wire [16-1:0] node5907;
	wire [16-1:0] node5908;
	wire [16-1:0] node5912;
	wire [16-1:0] node5913;
	wire [16-1:0] node5914;
	wire [16-1:0] node5916;
	wire [16-1:0] node5919;
	wire [16-1:0] node5921;
	wire [16-1:0] node5925;
	wire [16-1:0] node5926;
	wire [16-1:0] node5927;
	wire [16-1:0] node5930;
	wire [16-1:0] node5931;
	wire [16-1:0] node5932;
	wire [16-1:0] node5935;
	wire [16-1:0] node5938;
	wire [16-1:0] node5941;
	wire [16-1:0] node5942;
	wire [16-1:0] node5943;
	wire [16-1:0] node5944;
	wire [16-1:0] node5946;
	wire [16-1:0] node5951;
	wire [16-1:0] node5952;
	wire [16-1:0] node5954;
	wire [16-1:0] node5957;
	wire [16-1:0] node5960;
	wire [16-1:0] node5961;
	wire [16-1:0] node5962;
	wire [16-1:0] node5963;
	wire [16-1:0] node5964;
	wire [16-1:0] node5965;
	wire [16-1:0] node5966;
	wire [16-1:0] node5967;
	wire [16-1:0] node5968;
	wire [16-1:0] node5969;
	wire [16-1:0] node5972;
	wire [16-1:0] node5973;
	wire [16-1:0] node5975;
	wire [16-1:0] node5976;
	wire [16-1:0] node5979;
	wire [16-1:0] node5982;
	wire [16-1:0] node5984;
	wire [16-1:0] node5987;
	wire [16-1:0] node5988;
	wire [16-1:0] node5989;
	wire [16-1:0] node5992;
	wire [16-1:0] node5994;
	wire [16-1:0] node5997;
	wire [16-1:0] node5998;
	wire [16-1:0] node6002;
	wire [16-1:0] node6003;
	wire [16-1:0] node6004;
	wire [16-1:0] node6005;
	wire [16-1:0] node6007;
	wire [16-1:0] node6008;
	wire [16-1:0] node6013;
	wire [16-1:0] node6014;
	wire [16-1:0] node6018;
	wire [16-1:0] node6019;
	wire [16-1:0] node6020;
	wire [16-1:0] node6024;
	wire [16-1:0] node6025;
	wire [16-1:0] node6026;
	wire [16-1:0] node6030;
	wire [16-1:0] node6032;
	wire [16-1:0] node6033;
	wire [16-1:0] node6037;
	wire [16-1:0] node6038;
	wire [16-1:0] node6039;
	wire [16-1:0] node6040;
	wire [16-1:0] node6041;
	wire [16-1:0] node6043;
	wire [16-1:0] node6045;
	wire [16-1:0] node6048;
	wire [16-1:0] node6050;
	wire [16-1:0] node6051;
	wire [16-1:0] node6056;
	wire [16-1:0] node6057;
	wire [16-1:0] node6058;
	wire [16-1:0] node6061;
	wire [16-1:0] node6063;
	wire [16-1:0] node6064;
	wire [16-1:0] node6068;
	wire [16-1:0] node6069;
	wire [16-1:0] node6072;
	wire [16-1:0] node6074;
	wire [16-1:0] node6077;
	wire [16-1:0] node6078;
	wire [16-1:0] node6079;
	wire [16-1:0] node6081;
	wire [16-1:0] node6084;
	wire [16-1:0] node6085;
	wire [16-1:0] node6087;
	wire [16-1:0] node6088;
	wire [16-1:0] node6090;
	wire [16-1:0] node6094;
	wire [16-1:0] node6097;
	wire [16-1:0] node6098;
	wire [16-1:0] node6099;
	wire [16-1:0] node6101;
	wire [16-1:0] node6104;
	wire [16-1:0] node6106;
	wire [16-1:0] node6107;
	wire [16-1:0] node6111;
	wire [16-1:0] node6112;
	wire [16-1:0] node6115;
	wire [16-1:0] node6118;
	wire [16-1:0] node6119;
	wire [16-1:0] node6120;
	wire [16-1:0] node6121;
	wire [16-1:0] node6122;
	wire [16-1:0] node6123;
	wire [16-1:0] node6125;
	wire [16-1:0] node6128;
	wire [16-1:0] node6129;
	wire [16-1:0] node6133;
	wire [16-1:0] node6134;
	wire [16-1:0] node6135;
	wire [16-1:0] node6137;
	wire [16-1:0] node6141;
	wire [16-1:0] node6144;
	wire [16-1:0] node6145;
	wire [16-1:0] node6146;
	wire [16-1:0] node6148;
	wire [16-1:0] node6149;
	wire [16-1:0] node6150;
	wire [16-1:0] node6155;
	wire [16-1:0] node6157;
	wire [16-1:0] node6160;
	wire [16-1:0] node6161;
	wire [16-1:0] node6162;
	wire [16-1:0] node6164;
	wire [16-1:0] node6167;
	wire [16-1:0] node6168;
	wire [16-1:0] node6171;
	wire [16-1:0] node6174;
	wire [16-1:0] node6176;
	wire [16-1:0] node6179;
	wire [16-1:0] node6180;
	wire [16-1:0] node6181;
	wire [16-1:0] node6182;
	wire [16-1:0] node6184;
	wire [16-1:0] node6188;
	wire [16-1:0] node6189;
	wire [16-1:0] node6190;
	wire [16-1:0] node6191;
	wire [16-1:0] node6196;
	wire [16-1:0] node6197;
	wire [16-1:0] node6199;
	wire [16-1:0] node6202;
	wire [16-1:0] node6205;
	wire [16-1:0] node6206;
	wire [16-1:0] node6207;
	wire [16-1:0] node6208;
	wire [16-1:0] node6212;
	wire [16-1:0] node6214;
	wire [16-1:0] node6217;
	wire [16-1:0] node6218;
	wire [16-1:0] node6220;
	wire [16-1:0] node6224;
	wire [16-1:0] node6225;
	wire [16-1:0] node6226;
	wire [16-1:0] node6227;
	wire [16-1:0] node6228;
	wire [16-1:0] node6229;
	wire [16-1:0] node6233;
	wire [16-1:0] node6234;
	wire [16-1:0] node6237;
	wire [16-1:0] node6238;
	wire [16-1:0] node6243;
	wire [16-1:0] node6244;
	wire [16-1:0] node6245;
	wire [16-1:0] node6246;
	wire [16-1:0] node6248;
	wire [16-1:0] node6251;
	wire [16-1:0] node6252;
	wire [16-1:0] node6256;
	wire [16-1:0] node6258;
	wire [16-1:0] node6261;
	wire [16-1:0] node6262;
	wire [16-1:0] node6265;
	wire [16-1:0] node6267;
	wire [16-1:0] node6270;
	wire [16-1:0] node6271;
	wire [16-1:0] node6272;
	wire [16-1:0] node6273;
	wire [16-1:0] node6276;
	wire [16-1:0] node6278;
	wire [16-1:0] node6281;
	wire [16-1:0] node6282;
	wire [16-1:0] node6283;
	wire [16-1:0] node6285;
	wire [16-1:0] node6289;
	wire [16-1:0] node6291;
	wire [16-1:0] node6294;
	wire [16-1:0] node6295;
	wire [16-1:0] node6296;
	wire [16-1:0] node6297;
	wire [16-1:0] node6301;
	wire [16-1:0] node6303;
	wire [16-1:0] node6304;
	wire [16-1:0] node6308;
	wire [16-1:0] node6309;
	wire [16-1:0] node6312;
	wire [16-1:0] node6314;
	wire [16-1:0] node6317;
	wire [16-1:0] node6318;
	wire [16-1:0] node6319;
	wire [16-1:0] node6320;
	wire [16-1:0] node6321;
	wire [16-1:0] node6322;
	wire [16-1:0] node6323;
	wire [16-1:0] node6324;
	wire [16-1:0] node6328;
	wire [16-1:0] node6329;
	wire [16-1:0] node6333;
	wire [16-1:0] node6334;
	wire [16-1:0] node6337;
	wire [16-1:0] node6340;
	wire [16-1:0] node6341;
	wire [16-1:0] node6344;
	wire [16-1:0] node6345;
	wire [16-1:0] node6347;
	wire [16-1:0] node6351;
	wire [16-1:0] node6352;
	wire [16-1:0] node6353;
	wire [16-1:0] node6354;
	wire [16-1:0] node6357;
	wire [16-1:0] node6359;
	wire [16-1:0] node6362;
	wire [16-1:0] node6363;
	wire [16-1:0] node6367;
	wire [16-1:0] node6368;
	wire [16-1:0] node6369;
	wire [16-1:0] node6371;
	wire [16-1:0] node6374;
	wire [16-1:0] node6376;
	wire [16-1:0] node6379;
	wire [16-1:0] node6380;
	wire [16-1:0] node6384;
	wire [16-1:0] node6385;
	wire [16-1:0] node6386;
	wire [16-1:0] node6387;
	wire [16-1:0] node6388;
	wire [16-1:0] node6392;
	wire [16-1:0] node6393;
	wire [16-1:0] node6396;
	wire [16-1:0] node6398;
	wire [16-1:0] node6400;
	wire [16-1:0] node6403;
	wire [16-1:0] node6404;
	wire [16-1:0] node6405;
	wire [16-1:0] node6407;
	wire [16-1:0] node6408;
	wire [16-1:0] node6412;
	wire [16-1:0] node6414;
	wire [16-1:0] node6415;
	wire [16-1:0] node6419;
	wire [16-1:0] node6420;
	wire [16-1:0] node6423;
	wire [16-1:0] node6426;
	wire [16-1:0] node6427;
	wire [16-1:0] node6428;
	wire [16-1:0] node6429;
	wire [16-1:0] node6430;
	wire [16-1:0] node6434;
	wire [16-1:0] node6437;
	wire [16-1:0] node6440;
	wire [16-1:0] node6441;
	wire [16-1:0] node6442;
	wire [16-1:0] node6443;
	wire [16-1:0] node6444;
	wire [16-1:0] node6446;
	wire [16-1:0] node6450;
	wire [16-1:0] node6453;
	wire [16-1:0] node6455;
	wire [16-1:0] node6458;
	wire [16-1:0] node6459;
	wire [16-1:0] node6462;
	wire [16-1:0] node6465;
	wire [16-1:0] node6466;
	wire [16-1:0] node6467;
	wire [16-1:0] node6468;
	wire [16-1:0] node6469;
	wire [16-1:0] node6470;
	wire [16-1:0] node6471;
	wire [16-1:0] node6474;
	wire [16-1:0] node6476;
	wire [16-1:0] node6479;
	wire [16-1:0] node6480;
	wire [16-1:0] node6481;
	wire [16-1:0] node6485;
	wire [16-1:0] node6486;
	wire [16-1:0] node6490;
	wire [16-1:0] node6492;
	wire [16-1:0] node6495;
	wire [16-1:0] node6496;
	wire [16-1:0] node6497;
	wire [16-1:0] node6498;
	wire [16-1:0] node6502;
	wire [16-1:0] node6503;
	wire [16-1:0] node6505;
	wire [16-1:0] node6507;
	wire [16-1:0] node6511;
	wire [16-1:0] node6513;
	wire [16-1:0] node6516;
	wire [16-1:0] node6517;
	wire [16-1:0] node6518;
	wire [16-1:0] node6519;
	wire [16-1:0] node6521;
	wire [16-1:0] node6525;
	wire [16-1:0] node6526;
	wire [16-1:0] node6528;
	wire [16-1:0] node6531;
	wire [16-1:0] node6532;
	wire [16-1:0] node6533;
	wire [16-1:0] node6536;
	wire [16-1:0] node6538;
	wire [16-1:0] node6541;
	wire [16-1:0] node6543;
	wire [16-1:0] node6546;
	wire [16-1:0] node6547;
	wire [16-1:0] node6549;
	wire [16-1:0] node6552;
	wire [16-1:0] node6553;
	wire [16-1:0] node6556;
	wire [16-1:0] node6557;
	wire [16-1:0] node6559;
	wire [16-1:0] node6563;
	wire [16-1:0] node6564;
	wire [16-1:0] node6565;
	wire [16-1:0] node6566;
	wire [16-1:0] node6568;
	wire [16-1:0] node6571;
	wire [16-1:0] node6572;
	wire [16-1:0] node6575;
	wire [16-1:0] node6577;
	wire [16-1:0] node6580;
	wire [16-1:0] node6581;
	wire [16-1:0] node6582;
	wire [16-1:0] node6585;
	wire [16-1:0] node6587;
	wire [16-1:0] node6590;
	wire [16-1:0] node6591;
	wire [16-1:0] node6594;
	wire [16-1:0] node6595;
	wire [16-1:0] node6597;
	wire [16-1:0] node6601;
	wire [16-1:0] node6602;
	wire [16-1:0] node6603;
	wire [16-1:0] node6604;
	wire [16-1:0] node6608;
	wire [16-1:0] node6609;
	wire [16-1:0] node6612;
	wire [16-1:0] node6614;
	wire [16-1:0] node6615;
	wire [16-1:0] node6619;
	wire [16-1:0] node6620;
	wire [16-1:0] node6622;
	wire [16-1:0] node6623;
	wire [16-1:0] node6625;
	wire [16-1:0] node6629;
	wire [16-1:0] node6630;
	wire [16-1:0] node6631;
	wire [16-1:0] node6632;
	wire [16-1:0] node6636;
	wire [16-1:0] node6639;
	wire [16-1:0] node6640;
	wire [16-1:0] node6644;
	wire [16-1:0] node6645;
	wire [16-1:0] node6646;
	wire [16-1:0] node6647;
	wire [16-1:0] node6648;
	wire [16-1:0] node6649;
	wire [16-1:0] node6650;
	wire [16-1:0] node6652;
	wire [16-1:0] node6654;
	wire [16-1:0] node6657;
	wire [16-1:0] node6658;
	wire [16-1:0] node6660;
	wire [16-1:0] node6663;
	wire [16-1:0] node6666;
	wire [16-1:0] node6667;
	wire [16-1:0] node6668;
	wire [16-1:0] node6669;
	wire [16-1:0] node6670;
	wire [16-1:0] node6674;
	wire [16-1:0] node6677;
	wire [16-1:0] node6678;
	wire [16-1:0] node6679;
	wire [16-1:0] node6681;
	wire [16-1:0] node6686;
	wire [16-1:0] node6687;
	wire [16-1:0] node6689;
	wire [16-1:0] node6692;
	wire [16-1:0] node6693;
	wire [16-1:0] node6697;
	wire [16-1:0] node6698;
	wire [16-1:0] node6699;
	wire [16-1:0] node6700;
	wire [16-1:0] node6701;
	wire [16-1:0] node6703;
	wire [16-1:0] node6707;
	wire [16-1:0] node6708;
	wire [16-1:0] node6712;
	wire [16-1:0] node6713;
	wire [16-1:0] node6717;
	wire [16-1:0] node6718;
	wire [16-1:0] node6719;
	wire [16-1:0] node6721;
	wire [16-1:0] node6722;
	wire [16-1:0] node6724;
	wire [16-1:0] node6728;
	wire [16-1:0] node6731;
	wire [16-1:0] node6732;
	wire [16-1:0] node6735;
	wire [16-1:0] node6736;
	wire [16-1:0] node6739;
	wire [16-1:0] node6742;
	wire [16-1:0] node6743;
	wire [16-1:0] node6744;
	wire [16-1:0] node6745;
	wire [16-1:0] node6746;
	wire [16-1:0] node6747;
	wire [16-1:0] node6750;
	wire [16-1:0] node6753;
	wire [16-1:0] node6754;
	wire [16-1:0] node6758;
	wire [16-1:0] node6760;
	wire [16-1:0] node6762;
	wire [16-1:0] node6763;
	wire [16-1:0] node6767;
	wire [16-1:0] node6768;
	wire [16-1:0] node6769;
	wire [16-1:0] node6771;
	wire [16-1:0] node6775;
	wire [16-1:0] node6776;
	wire [16-1:0] node6777;
	wire [16-1:0] node6781;
	wire [16-1:0] node6783;
	wire [16-1:0] node6785;
	wire [16-1:0] node6788;
	wire [16-1:0] node6789;
	wire [16-1:0] node6790;
	wire [16-1:0] node6791;
	wire [16-1:0] node6793;
	wire [16-1:0] node6794;
	wire [16-1:0] node6799;
	wire [16-1:0] node6800;
	wire [16-1:0] node6803;
	wire [16-1:0] node6806;
	wire [16-1:0] node6807;
	wire [16-1:0] node6810;
	wire [16-1:0] node6812;
	wire [16-1:0] node6814;
	wire [16-1:0] node6815;
	wire [16-1:0] node6819;
	wire [16-1:0] node6820;
	wire [16-1:0] node6821;
	wire [16-1:0] node6822;
	wire [16-1:0] node6823;
	wire [16-1:0] node6824;
	wire [16-1:0] node6826;
	wire [16-1:0] node6830;
	wire [16-1:0] node6831;
	wire [16-1:0] node6832;
	wire [16-1:0] node6835;
	wire [16-1:0] node6839;
	wire [16-1:0] node6840;
	wire [16-1:0] node6843;
	wire [16-1:0] node6844;
	wire [16-1:0] node6845;
	wire [16-1:0] node6847;
	wire [16-1:0] node6850;
	wire [16-1:0] node6852;
	wire [16-1:0] node6855;
	wire [16-1:0] node6856;
	wire [16-1:0] node6860;
	wire [16-1:0] node6861;
	wire [16-1:0] node6862;
	wire [16-1:0] node6863;
	wire [16-1:0] node6866;
	wire [16-1:0] node6868;
	wire [16-1:0] node6871;
	wire [16-1:0] node6873;
	wire [16-1:0] node6874;
	wire [16-1:0] node6878;
	wire [16-1:0] node6879;
	wire [16-1:0] node6880;
	wire [16-1:0] node6882;
	wire [16-1:0] node6885;
	wire [16-1:0] node6886;
	wire [16-1:0] node6890;
	wire [16-1:0] node6891;
	wire [16-1:0] node6894;
	wire [16-1:0] node6897;
	wire [16-1:0] node6898;
	wire [16-1:0] node6899;
	wire [16-1:0] node6900;
	wire [16-1:0] node6901;
	wire [16-1:0] node6903;
	wire [16-1:0] node6907;
	wire [16-1:0] node6910;
	wire [16-1:0] node6911;
	wire [16-1:0] node6912;
	wire [16-1:0] node6913;
	wire [16-1:0] node6917;
	wire [16-1:0] node6918;
	wire [16-1:0] node6919;
	wire [16-1:0] node6923;
	wire [16-1:0] node6924;
	wire [16-1:0] node6928;
	wire [16-1:0] node6929;
	wire [16-1:0] node6931;
	wire [16-1:0] node6932;
	wire [16-1:0] node6937;
	wire [16-1:0] node6938;
	wire [16-1:0] node6939;
	wire [16-1:0] node6941;
	wire [16-1:0] node6942;
	wire [16-1:0] node6946;
	wire [16-1:0] node6947;
	wire [16-1:0] node6950;
	wire [16-1:0] node6951;
	wire [16-1:0] node6953;
	wire [16-1:0] node6957;
	wire [16-1:0] node6958;
	wire [16-1:0] node6959;
	wire [16-1:0] node6960;
	wire [16-1:0] node6962;
	wire [16-1:0] node6966;
	wire [16-1:0] node6967;
	wire [16-1:0] node6970;
	wire [16-1:0] node6973;
	wire [16-1:0] node6975;
	wire [16-1:0] node6977;
	wire [16-1:0] node6978;
	wire [16-1:0] node6981;
	wire [16-1:0] node6984;
	wire [16-1:0] node6985;
	wire [16-1:0] node6986;
	wire [16-1:0] node6987;
	wire [16-1:0] node6988;
	wire [16-1:0] node6989;
	wire [16-1:0] node6990;
	wire [16-1:0] node6993;
	wire [16-1:0] node6995;
	wire [16-1:0] node6998;
	wire [16-1:0] node6999;
	wire [16-1:0] node7000;
	wire [16-1:0] node7002;
	wire [16-1:0] node7006;
	wire [16-1:0] node7009;
	wire [16-1:0] node7010;
	wire [16-1:0] node7011;
	wire [16-1:0] node7013;
	wire [16-1:0] node7014;
	wire [16-1:0] node7018;
	wire [16-1:0] node7021;
	wire [16-1:0] node7023;
	wire [16-1:0] node7026;
	wire [16-1:0] node7027;
	wire [16-1:0] node7028;
	wire [16-1:0] node7029;
	wire [16-1:0] node7030;
	wire [16-1:0] node7034;
	wire [16-1:0] node7037;
	wire [16-1:0] node7038;
	wire [16-1:0] node7039;
	wire [16-1:0] node7043;
	wire [16-1:0] node7045;
	wire [16-1:0] node7048;
	wire [16-1:0] node7049;
	wire [16-1:0] node7050;
	wire [16-1:0] node7052;
	wire [16-1:0] node7055;
	wire [16-1:0] node7056;
	wire [16-1:0] node7059;
	wire [16-1:0] node7060;
	wire [16-1:0] node7061;
	wire [16-1:0] node7066;
	wire [16-1:0] node7067;
	wire [16-1:0] node7068;
	wire [16-1:0] node7072;
	wire [16-1:0] node7075;
	wire [16-1:0] node7076;
	wire [16-1:0] node7077;
	wire [16-1:0] node7078;
	wire [16-1:0] node7079;
	wire [16-1:0] node7082;
	wire [16-1:0] node7085;
	wire [16-1:0] node7087;
	wire [16-1:0] node7090;
	wire [16-1:0] node7091;
	wire [16-1:0] node7092;
	wire [16-1:0] node7093;
	wire [16-1:0] node7095;
	wire [16-1:0] node7099;
	wire [16-1:0] node7101;
	wire [16-1:0] node7102;
	wire [16-1:0] node7106;
	wire [16-1:0] node7107;
	wire [16-1:0] node7110;
	wire [16-1:0] node7113;
	wire [16-1:0] node7114;
	wire [16-1:0] node7115;
	wire [16-1:0] node7116;
	wire [16-1:0] node7118;
	wire [16-1:0] node7120;
	wire [16-1:0] node7123;
	wire [16-1:0] node7126;
	wire [16-1:0] node7127;
	wire [16-1:0] node7131;
	wire [16-1:0] node7132;
	wire [16-1:0] node7133;
	wire [16-1:0] node7134;
	wire [16-1:0] node7138;
	wire [16-1:0] node7140;
	wire [16-1:0] node7141;
	wire [16-1:0] node7145;
	wire [16-1:0] node7146;
	wire [16-1:0] node7147;
	wire [16-1:0] node7149;
	wire [16-1:0] node7153;
	wire [16-1:0] node7156;
	wire [16-1:0] node7157;
	wire [16-1:0] node7158;
	wire [16-1:0] node7159;
	wire [16-1:0] node7160;
	wire [16-1:0] node7161;
	wire [16-1:0] node7162;
	wire [16-1:0] node7166;
	wire [16-1:0] node7167;
	wire [16-1:0] node7169;
	wire [16-1:0] node7172;
	wire [16-1:0] node7175;
	wire [16-1:0] node7176;
	wire [16-1:0] node7179;
	wire [16-1:0] node7181;
	wire [16-1:0] node7182;
	wire [16-1:0] node7183;
	wire [16-1:0] node7188;
	wire [16-1:0] node7189;
	wire [16-1:0] node7190;
	wire [16-1:0] node7193;
	wire [16-1:0] node7194;
	wire [16-1:0] node7195;
	wire [16-1:0] node7199;
	wire [16-1:0] node7200;
	wire [16-1:0] node7204;
	wire [16-1:0] node7205;
	wire [16-1:0] node7208;
	wire [16-1:0] node7211;
	wire [16-1:0] node7212;
	wire [16-1:0] node7213;
	wire [16-1:0] node7216;
	wire [16-1:0] node7217;
	wire [16-1:0] node7218;
	wire [16-1:0] node7220;
	wire [16-1:0] node7224;
	wire [16-1:0] node7226;
	wire [16-1:0] node7229;
	wire [16-1:0] node7230;
	wire [16-1:0] node7231;
	wire [16-1:0] node7232;
	wire [16-1:0] node7236;
	wire [16-1:0] node7239;
	wire [16-1:0] node7240;
	wire [16-1:0] node7241;
	wire [16-1:0] node7245;
	wire [16-1:0] node7246;
	wire [16-1:0] node7249;
	wire [16-1:0] node7251;
	wire [16-1:0] node7252;
	wire [16-1:0] node7256;
	wire [16-1:0] node7257;
	wire [16-1:0] node7258;
	wire [16-1:0] node7259;
	wire [16-1:0] node7261;
	wire [16-1:0] node7264;
	wire [16-1:0] node7265;
	wire [16-1:0] node7266;
	wire [16-1:0] node7270;
	wire [16-1:0] node7273;
	wire [16-1:0] node7274;
	wire [16-1:0] node7275;
	wire [16-1:0] node7279;
	wire [16-1:0] node7280;
	wire [16-1:0] node7282;
	wire [16-1:0] node7286;
	wire [16-1:0] node7287;
	wire [16-1:0] node7288;
	wire [16-1:0] node7289;
	wire [16-1:0] node7290;
	wire [16-1:0] node7292;
	wire [16-1:0] node7297;
	wire [16-1:0] node7298;
	wire [16-1:0] node7300;
	wire [16-1:0] node7302;
	wire [16-1:0] node7304;
	wire [16-1:0] node7307;
	wire [16-1:0] node7308;
	wire [16-1:0] node7310;
	wire [16-1:0] node7313;
	wire [16-1:0] node7316;
	wire [16-1:0] node7317;
	wire [16-1:0] node7318;
	wire [16-1:0] node7319;
	wire [16-1:0] node7322;
	wire [16-1:0] node7325;
	wire [16-1:0] node7327;
	wire [16-1:0] node7330;
	wire [16-1:0] node7331;
	wire [16-1:0] node7332;
	wire [16-1:0] node7335;
	wire [16-1:0] node7338;
	wire [16-1:0] node7340;
	wire [16-1:0] node7343;
	wire [16-1:0] node7344;
	wire [16-1:0] node7345;
	wire [16-1:0] node7346;
	wire [16-1:0] node7347;
	wire [16-1:0] node7348;
	wire [16-1:0] node7349;
	wire [16-1:0] node7350;
	wire [16-1:0] node7351;
	wire [16-1:0] node7352;
	wire [16-1:0] node7356;
	wire [16-1:0] node7358;
	wire [16-1:0] node7360;
	wire [16-1:0] node7363;
	wire [16-1:0] node7364;
	wire [16-1:0] node7365;
	wire [16-1:0] node7369;
	wire [16-1:0] node7372;
	wire [16-1:0] node7373;
	wire [16-1:0] node7374;
	wire [16-1:0] node7376;
	wire [16-1:0] node7379;
	wire [16-1:0] node7382;
	wire [16-1:0] node7383;
	wire [16-1:0] node7385;
	wire [16-1:0] node7389;
	wire [16-1:0] node7390;
	wire [16-1:0] node7391;
	wire [16-1:0] node7392;
	wire [16-1:0] node7393;
	wire [16-1:0] node7396;
	wire [16-1:0] node7397;
	wire [16-1:0] node7401;
	wire [16-1:0] node7404;
	wire [16-1:0] node7405;
	wire [16-1:0] node7407;
	wire [16-1:0] node7408;
	wire [16-1:0] node7410;
	wire [16-1:0] node7414;
	wire [16-1:0] node7417;
	wire [16-1:0] node7418;
	wire [16-1:0] node7420;
	wire [16-1:0] node7422;
	wire [16-1:0] node7425;
	wire [16-1:0] node7427;
	wire [16-1:0] node7430;
	wire [16-1:0] node7431;
	wire [16-1:0] node7432;
	wire [16-1:0] node7433;
	wire [16-1:0] node7434;
	wire [16-1:0] node7436;
	wire [16-1:0] node7439;
	wire [16-1:0] node7440;
	wire [16-1:0] node7443;
	wire [16-1:0] node7446;
	wire [16-1:0] node7447;
	wire [16-1:0] node7448;
	wire [16-1:0] node7450;
	wire [16-1:0] node7454;
	wire [16-1:0] node7455;
	wire [16-1:0] node7459;
	wire [16-1:0] node7460;
	wire [16-1:0] node7461;
	wire [16-1:0] node7465;
	wire [16-1:0] node7466;
	wire [16-1:0] node7468;
	wire [16-1:0] node7469;
	wire [16-1:0] node7474;
	wire [16-1:0] node7475;
	wire [16-1:0] node7476;
	wire [16-1:0] node7478;
	wire [16-1:0] node7481;
	wire [16-1:0] node7482;
	wire [16-1:0] node7486;
	wire [16-1:0] node7487;
	wire [16-1:0] node7488;
	wire [16-1:0] node7492;
	wire [16-1:0] node7493;
	wire [16-1:0] node7495;
	wire [16-1:0] node7498;
	wire [16-1:0] node7499;
	wire [16-1:0] node7503;
	wire [16-1:0] node7504;
	wire [16-1:0] node7505;
	wire [16-1:0] node7506;
	wire [16-1:0] node7507;
	wire [16-1:0] node7509;
	wire [16-1:0] node7512;
	wire [16-1:0] node7513;
	wire [16-1:0] node7515;
	wire [16-1:0] node7518;
	wire [16-1:0] node7519;
	wire [16-1:0] node7520;
	wire [16-1:0] node7525;
	wire [16-1:0] node7526;
	wire [16-1:0] node7528;
	wire [16-1:0] node7529;
	wire [16-1:0] node7533;
	wire [16-1:0] node7534;
	wire [16-1:0] node7537;
	wire [16-1:0] node7538;
	wire [16-1:0] node7540;
	wire [16-1:0] node7544;
	wire [16-1:0] node7545;
	wire [16-1:0] node7546;
	wire [16-1:0] node7547;
	wire [16-1:0] node7548;
	wire [16-1:0] node7553;
	wire [16-1:0] node7554;
	wire [16-1:0] node7556;
	wire [16-1:0] node7559;
	wire [16-1:0] node7560;
	wire [16-1:0] node7564;
	wire [16-1:0] node7565;
	wire [16-1:0] node7566;
	wire [16-1:0] node7567;
	wire [16-1:0] node7569;
	wire [16-1:0] node7570;
	wire [16-1:0] node7575;
	wire [16-1:0] node7576;
	wire [16-1:0] node7580;
	wire [16-1:0] node7582;
	wire [16-1:0] node7583;
	wire [16-1:0] node7585;
	wire [16-1:0] node7589;
	wire [16-1:0] node7590;
	wire [16-1:0] node7591;
	wire [16-1:0] node7592;
	wire [16-1:0] node7593;
	wire [16-1:0] node7596;
	wire [16-1:0] node7598;
	wire [16-1:0] node7601;
	wire [16-1:0] node7603;
	wire [16-1:0] node7604;
	wire [16-1:0] node7608;
	wire [16-1:0] node7609;
	wire [16-1:0] node7610;
	wire [16-1:0] node7612;
	wire [16-1:0] node7615;
	wire [16-1:0] node7616;
	wire [16-1:0] node7620;
	wire [16-1:0] node7621;
	wire [16-1:0] node7624;
	wire [16-1:0] node7626;
	wire [16-1:0] node7629;
	wire [16-1:0] node7630;
	wire [16-1:0] node7631;
	wire [16-1:0] node7632;
	wire [16-1:0] node7633;
	wire [16-1:0] node7634;
	wire [16-1:0] node7638;
	wire [16-1:0] node7641;
	wire [16-1:0] node7644;
	wire [16-1:0] node7645;
	wire [16-1:0] node7649;
	wire [16-1:0] node7650;
	wire [16-1:0] node7652;
	wire [16-1:0] node7655;
	wire [16-1:0] node7656;
	wire [16-1:0] node7658;
	wire [16-1:0] node7662;
	wire [16-1:0] node7663;
	wire [16-1:0] node7664;
	wire [16-1:0] node7665;
	wire [16-1:0] node7666;
	wire [16-1:0] node7667;
	wire [16-1:0] node7668;
	wire [16-1:0] node7670;
	wire [16-1:0] node7671;
	wire [16-1:0] node7673;
	wire [16-1:0] node7677;
	wire [16-1:0] node7678;
	wire [16-1:0] node7680;
	wire [16-1:0] node7684;
	wire [16-1:0] node7685;
	wire [16-1:0] node7689;
	wire [16-1:0] node7691;
	wire [16-1:0] node7694;
	wire [16-1:0] node7695;
	wire [16-1:0] node7696;
	wire [16-1:0] node7697;
	wire [16-1:0] node7701;
	wire [16-1:0] node7702;
	wire [16-1:0] node7705;
	wire [16-1:0] node7708;
	wire [16-1:0] node7709;
	wire [16-1:0] node7710;
	wire [16-1:0] node7711;
	wire [16-1:0] node7712;
	wire [16-1:0] node7715;
	wire [16-1:0] node7719;
	wire [16-1:0] node7722;
	wire [16-1:0] node7723;
	wire [16-1:0] node7725;
	wire [16-1:0] node7728;
	wire [16-1:0] node7730;
	wire [16-1:0] node7733;
	wire [16-1:0] node7734;
	wire [16-1:0] node7735;
	wire [16-1:0] node7736;
	wire [16-1:0] node7737;
	wire [16-1:0] node7739;
	wire [16-1:0] node7742;
	wire [16-1:0] node7743;
	wire [16-1:0] node7747;
	wire [16-1:0] node7750;
	wire [16-1:0] node7751;
	wire [16-1:0] node7754;
	wire [16-1:0] node7755;
	wire [16-1:0] node7757;
	wire [16-1:0] node7758;
	wire [16-1:0] node7763;
	wire [16-1:0] node7764;
	wire [16-1:0] node7765;
	wire [16-1:0] node7767;
	wire [16-1:0] node7768;
	wire [16-1:0] node7772;
	wire [16-1:0] node7774;
	wire [16-1:0] node7777;
	wire [16-1:0] node7778;
	wire [16-1:0] node7780;
	wire [16-1:0] node7783;
	wire [16-1:0] node7784;
	wire [16-1:0] node7786;
	wire [16-1:0] node7789;
	wire [16-1:0] node7792;
	wire [16-1:0] node7793;
	wire [16-1:0] node7794;
	wire [16-1:0] node7795;
	wire [16-1:0] node7796;
	wire [16-1:0] node7797;
	wire [16-1:0] node7800;
	wire [16-1:0] node7802;
	wire [16-1:0] node7806;
	wire [16-1:0] node7807;
	wire [16-1:0] node7809;
	wire [16-1:0] node7810;
	wire [16-1:0] node7814;
	wire [16-1:0] node7815;
	wire [16-1:0] node7816;
	wire [16-1:0] node7819;
	wire [16-1:0] node7820;
	wire [16-1:0] node7825;
	wire [16-1:0] node7826;
	wire [16-1:0] node7827;
	wire [16-1:0] node7828;
	wire [16-1:0] node7831;
	wire [16-1:0] node7834;
	wire [16-1:0] node7835;
	wire [16-1:0] node7836;
	wire [16-1:0] node7837;
	wire [16-1:0] node7842;
	wire [16-1:0] node7843;
	wire [16-1:0] node7844;
	wire [16-1:0] node7849;
	wire [16-1:0] node7850;
	wire [16-1:0] node7851;
	wire [16-1:0] node7853;
	wire [16-1:0] node7855;
	wire [16-1:0] node7859;
	wire [16-1:0] node7860;
	wire [16-1:0] node7863;
	wire [16-1:0] node7866;
	wire [16-1:0] node7867;
	wire [16-1:0] node7868;
	wire [16-1:0] node7869;
	wire [16-1:0] node7870;
	wire [16-1:0] node7871;
	wire [16-1:0] node7875;
	wire [16-1:0] node7876;
	wire [16-1:0] node7879;
	wire [16-1:0] node7883;
	wire [16-1:0] node7884;
	wire [16-1:0] node7885;
	wire [16-1:0] node7887;
	wire [16-1:0] node7890;
	wire [16-1:0] node7891;
	wire [16-1:0] node7892;
	wire [16-1:0] node7897;
	wire [16-1:0] node7899;
	wire [16-1:0] node7901;
	wire [16-1:0] node7903;
	wire [16-1:0] node7906;
	wire [16-1:0] node7907;
	wire [16-1:0] node7908;
	wire [16-1:0] node7909;
	wire [16-1:0] node7911;
	wire [16-1:0] node7914;
	wire [16-1:0] node7917;
	wire [16-1:0] node7918;
	wire [16-1:0] node7921;
	wire [16-1:0] node7923;
	wire [16-1:0] node7926;
	wire [16-1:0] node7927;
	wire [16-1:0] node7929;
	wire [16-1:0] node7930;
	wire [16-1:0] node7932;
	wire [16-1:0] node7936;
	wire [16-1:0] node7937;
	wire [16-1:0] node7940;
	wire [16-1:0] node7941;
	wire [16-1:0] node7942;
	wire [16-1:0] node7947;
	wire [16-1:0] node7948;
	wire [16-1:0] node7949;
	wire [16-1:0] node7950;
	wire [16-1:0] node7951;
	wire [16-1:0] node7952;
	wire [16-1:0] node7953;
	wire [16-1:0] node7954;
	wire [16-1:0] node7955;
	wire [16-1:0] node7956;
	wire [16-1:0] node7959;
	wire [16-1:0] node7960;
	wire [16-1:0] node7964;
	wire [16-1:0] node7967;
	wire [16-1:0] node7969;
	wire [16-1:0] node7970;
	wire [16-1:0] node7974;
	wire [16-1:0] node7977;
	wire [16-1:0] node7978;
	wire [16-1:0] node7979;
	wire [16-1:0] node7980;
	wire [16-1:0] node7984;
	wire [16-1:0] node7987;
	wire [16-1:0] node7988;
	wire [16-1:0] node7989;
	wire [16-1:0] node7992;
	wire [16-1:0] node7995;
	wire [16-1:0] node7996;
	wire [16-1:0] node7997;
	wire [16-1:0] node8002;
	wire [16-1:0] node8003;
	wire [16-1:0] node8004;
	wire [16-1:0] node8005;
	wire [16-1:0] node8006;
	wire [16-1:0] node8011;
	wire [16-1:0] node8012;
	wire [16-1:0] node8014;
	wire [16-1:0] node8017;
	wire [16-1:0] node8019;
	wire [16-1:0] node8020;
	wire [16-1:0] node8024;
	wire [16-1:0] node8025;
	wire [16-1:0] node8027;
	wire [16-1:0] node8030;
	wire [16-1:0] node8032;
	wire [16-1:0] node8035;
	wire [16-1:0] node8036;
	wire [16-1:0] node8037;
	wire [16-1:0] node8038;
	wire [16-1:0] node8039;
	wire [16-1:0] node8040;
	wire [16-1:0] node8045;
	wire [16-1:0] node8046;
	wire [16-1:0] node8049;
	wire [16-1:0] node8052;
	wire [16-1:0] node8053;
	wire [16-1:0] node8054;
	wire [16-1:0] node8055;
	wire [16-1:0] node8057;
	wire [16-1:0] node8059;
	wire [16-1:0] node8063;
	wire [16-1:0] node8065;
	wire [16-1:0] node8068;
	wire [16-1:0] node8070;
	wire [16-1:0] node8073;
	wire [16-1:0] node8074;
	wire [16-1:0] node8075;
	wire [16-1:0] node8076;
	wire [16-1:0] node8077;
	wire [16-1:0] node8078;
	wire [16-1:0] node8081;
	wire [16-1:0] node8085;
	wire [16-1:0] node8086;
	wire [16-1:0] node8090;
	wire [16-1:0] node8091;
	wire [16-1:0] node8092;
	wire [16-1:0] node8094;
	wire [16-1:0] node8098;
	wire [16-1:0] node8099;
	wire [16-1:0] node8101;
	wire [16-1:0] node8104;
	wire [16-1:0] node8106;
	wire [16-1:0] node8109;
	wire [16-1:0] node8110;
	wire [16-1:0] node8111;
	wire [16-1:0] node8114;
	wire [16-1:0] node8117;
	wire [16-1:0] node8118;
	wire [16-1:0] node8121;
	wire [16-1:0] node8123;
	wire [16-1:0] node8124;
	wire [16-1:0] node8128;
	wire [16-1:0] node8129;
	wire [16-1:0] node8130;
	wire [16-1:0] node8131;
	wire [16-1:0] node8132;
	wire [16-1:0] node8133;
	wire [16-1:0] node8136;
	wire [16-1:0] node8139;
	wire [16-1:0] node8141;
	wire [16-1:0] node8144;
	wire [16-1:0] node8145;
	wire [16-1:0] node8146;
	wire [16-1:0] node8149;
	wire [16-1:0] node8151;
	wire [16-1:0] node8154;
	wire [16-1:0] node8155;
	wire [16-1:0] node8158;
	wire [16-1:0] node8161;
	wire [16-1:0] node8162;
	wire [16-1:0] node8163;
	wire [16-1:0] node8164;
	wire [16-1:0] node8165;
	wire [16-1:0] node8166;
	wire [16-1:0] node8171;
	wire [16-1:0] node8172;
	wire [16-1:0] node8175;
	wire [16-1:0] node8176;
	wire [16-1:0] node8179;
	wire [16-1:0] node8182;
	wire [16-1:0] node8183;
	wire [16-1:0] node8185;
	wire [16-1:0] node8189;
	wire [16-1:0] node8190;
	wire [16-1:0] node8191;
	wire [16-1:0] node8194;
	wire [16-1:0] node8195;
	wire [16-1:0] node8197;
	wire [16-1:0] node8200;
	wire [16-1:0] node8201;
	wire [16-1:0] node8205;
	wire [16-1:0] node8207;
	wire [16-1:0] node8210;
	wire [16-1:0] node8211;
	wire [16-1:0] node8212;
	wire [16-1:0] node8213;
	wire [16-1:0] node8214;
	wire [16-1:0] node8217;
	wire [16-1:0] node8220;
	wire [16-1:0] node8221;
	wire [16-1:0] node8222;
	wire [16-1:0] node8224;
	wire [16-1:0] node8228;
	wire [16-1:0] node8231;
	wire [16-1:0] node8232;
	wire [16-1:0] node8233;
	wire [16-1:0] node8235;
	wire [16-1:0] node8237;
	wire [16-1:0] node8241;
	wire [16-1:0] node8243;
	wire [16-1:0] node8245;
	wire [16-1:0] node8246;
	wire [16-1:0] node8248;
	wire [16-1:0] node8252;
	wire [16-1:0] node8253;
	wire [16-1:0] node8255;
	wire [16-1:0] node8256;
	wire [16-1:0] node8259;
	wire [16-1:0] node8262;
	wire [16-1:0] node8263;
	wire [16-1:0] node8265;
	wire [16-1:0] node8266;
	wire [16-1:0] node8268;
	wire [16-1:0] node8271;
	wire [16-1:0] node8274;
	wire [16-1:0] node8275;
	wire [16-1:0] node8278;
	wire [16-1:0] node8279;
	wire [16-1:0] node8283;
	wire [16-1:0] node8284;
	wire [16-1:0] node8285;
	wire [16-1:0] node8286;
	wire [16-1:0] node8287;
	wire [16-1:0] node8288;
	wire [16-1:0] node8289;
	wire [16-1:0] node8292;
	wire [16-1:0] node8294;
	wire [16-1:0] node8297;
	wire [16-1:0] node8299;
	wire [16-1:0] node8302;
	wire [16-1:0] node8303;
	wire [16-1:0] node8304;
	wire [16-1:0] node8307;
	wire [16-1:0] node8308;
	wire [16-1:0] node8310;
	wire [16-1:0] node8314;
	wire [16-1:0] node8315;
	wire [16-1:0] node8316;
	wire [16-1:0] node8318;
	wire [16-1:0] node8322;
	wire [16-1:0] node8325;
	wire [16-1:0] node8326;
	wire [16-1:0] node8327;
	wire [16-1:0] node8331;
	wire [16-1:0] node8332;
	wire [16-1:0] node8334;
	wire [16-1:0] node8336;
	wire [16-1:0] node8339;
	wire [16-1:0] node8341;
	wire [16-1:0] node8342;
	wire [16-1:0] node8345;
	wire [16-1:0] node8348;
	wire [16-1:0] node8349;
	wire [16-1:0] node8350;
	wire [16-1:0] node8351;
	wire [16-1:0] node8352;
	wire [16-1:0] node8355;
	wire [16-1:0] node8357;
	wire [16-1:0] node8360;
	wire [16-1:0] node8361;
	wire [16-1:0] node8364;
	wire [16-1:0] node8366;
	wire [16-1:0] node8369;
	wire [16-1:0] node8370;
	wire [16-1:0] node8371;
	wire [16-1:0] node8372;
	wire [16-1:0] node8373;
	wire [16-1:0] node8378;
	wire [16-1:0] node8379;
	wire [16-1:0] node8381;
	wire [16-1:0] node8385;
	wire [16-1:0] node8386;
	wire [16-1:0] node8387;
	wire [16-1:0] node8389;
	wire [16-1:0] node8393;
	wire [16-1:0] node8396;
	wire [16-1:0] node8397;
	wire [16-1:0] node8398;
	wire [16-1:0] node8400;
	wire [16-1:0] node8401;
	wire [16-1:0] node8405;
	wire [16-1:0] node8406;
	wire [16-1:0] node8409;
	wire [16-1:0] node8411;
	wire [16-1:0] node8414;
	wire [16-1:0] node8415;
	wire [16-1:0] node8416;
	wire [16-1:0] node8418;
	wire [16-1:0] node8421;
	wire [16-1:0] node8424;
	wire [16-1:0] node8425;
	wire [16-1:0] node8426;
	wire [16-1:0] node8427;
	wire [16-1:0] node8431;
	wire [16-1:0] node8435;
	wire [16-1:0] node8436;
	wire [16-1:0] node8437;
	wire [16-1:0] node8438;
	wire [16-1:0] node8439;
	wire [16-1:0] node8440;
	wire [16-1:0] node8441;
	wire [16-1:0] node8445;
	wire [16-1:0] node8449;
	wire [16-1:0] node8450;
	wire [16-1:0] node8451;
	wire [16-1:0] node8452;
	wire [16-1:0] node8455;
	wire [16-1:0] node8459;
	wire [16-1:0] node8460;
	wire [16-1:0] node8462;
	wire [16-1:0] node8465;
	wire [16-1:0] node8468;
	wire [16-1:0] node8469;
	wire [16-1:0] node8470;
	wire [16-1:0] node8471;
	wire [16-1:0] node8472;
	wire [16-1:0] node8474;
	wire [16-1:0] node8477;
	wire [16-1:0] node8478;
	wire [16-1:0] node8482;
	wire [16-1:0] node8483;
	wire [16-1:0] node8487;
	wire [16-1:0] node8489;
	wire [16-1:0] node8490;
	wire [16-1:0] node8494;
	wire [16-1:0] node8495;
	wire [16-1:0] node8496;
	wire [16-1:0] node8499;
	wire [16-1:0] node8500;
	wire [16-1:0] node8502;
	wire [16-1:0] node8506;
	wire [16-1:0] node8507;
	wire [16-1:0] node8508;
	wire [16-1:0] node8512;
	wire [16-1:0] node8513;
	wire [16-1:0] node8517;
	wire [16-1:0] node8518;
	wire [16-1:0] node8519;
	wire [16-1:0] node8520;
	wire [16-1:0] node8521;
	wire [16-1:0] node8522;
	wire [16-1:0] node8523;
	wire [16-1:0] node8528;
	wire [16-1:0] node8531;
	wire [16-1:0] node8534;
	wire [16-1:0] node8535;
	wire [16-1:0] node8536;
	wire [16-1:0] node8537;
	wire [16-1:0] node8539;
	wire [16-1:0] node8543;
	wire [16-1:0] node8545;
	wire [16-1:0] node8547;
	wire [16-1:0] node8550;
	wire [16-1:0] node8551;
	wire [16-1:0] node8554;
	wire [16-1:0] node8555;
	wire [16-1:0] node8559;
	wire [16-1:0] node8560;
	wire [16-1:0] node8561;
	wire [16-1:0] node8562;
	wire [16-1:0] node8563;
	wire [16-1:0] node8565;
	wire [16-1:0] node8568;
	wire [16-1:0] node8569;
	wire [16-1:0] node8572;
	wire [16-1:0] node8575;
	wire [16-1:0] node8578;
	wire [16-1:0] node8580;
	wire [16-1:0] node8581;
	wire [16-1:0] node8582;
	wire [16-1:0] node8584;
	wire [16-1:0] node8589;
	wire [16-1:0] node8590;
	wire [16-1:0] node8591;
	wire [16-1:0] node8592;
	wire [16-1:0] node8597;
	wire [16-1:0] node8599;
	wire [16-1:0] node8600;
	wire [16-1:0] node8601;
	wire [16-1:0] node8604;
	wire [16-1:0] node8606;
	wire [16-1:0] node8609;
	wire [16-1:0] node8611;
	wire [16-1:0] node8614;
	wire [16-1:0] node8615;
	wire [16-1:0] node8616;
	wire [16-1:0] node8617;
	wire [16-1:0] node8618;
	wire [16-1:0] node8619;
	wire [16-1:0] node8620;
	wire [16-1:0] node8621;
	wire [16-1:0] node8622;
	wire [16-1:0] node8623;
	wire [16-1:0] node8625;
	wire [16-1:0] node8626;
	wire [16-1:0] node8630;
	wire [16-1:0] node8633;
	wire [16-1:0] node8634;
	wire [16-1:0] node8635;
	wire [16-1:0] node8638;
	wire [16-1:0] node8639;
	wire [16-1:0] node8643;
	wire [16-1:0] node8646;
	wire [16-1:0] node8647;
	wire [16-1:0] node8648;
	wire [16-1:0] node8649;
	wire [16-1:0] node8650;
	wire [16-1:0] node8655;
	wire [16-1:0] node8658;
	wire [16-1:0] node8659;
	wire [16-1:0] node8660;
	wire [16-1:0] node8664;
	wire [16-1:0] node8665;
	wire [16-1:0] node8669;
	wire [16-1:0] node8670;
	wire [16-1:0] node8671;
	wire [16-1:0] node8673;
	wire [16-1:0] node8674;
	wire [16-1:0] node8678;
	wire [16-1:0] node8679;
	wire [16-1:0] node8680;
	wire [16-1:0] node8683;
	wire [16-1:0] node8686;
	wire [16-1:0] node8687;
	wire [16-1:0] node8691;
	wire [16-1:0] node8692;
	wire [16-1:0] node8693;
	wire [16-1:0] node8696;
	wire [16-1:0] node8697;
	wire [16-1:0] node8701;
	wire [16-1:0] node8702;
	wire [16-1:0] node8705;
	wire [16-1:0] node8708;
	wire [16-1:0] node8709;
	wire [16-1:0] node8710;
	wire [16-1:0] node8711;
	wire [16-1:0] node8712;
	wire [16-1:0] node8714;
	wire [16-1:0] node8718;
	wire [16-1:0] node8719;
	wire [16-1:0] node8721;
	wire [16-1:0] node8722;
	wire [16-1:0] node8724;
	wire [16-1:0] node8728;
	wire [16-1:0] node8729;
	wire [16-1:0] node8730;
	wire [16-1:0] node8733;
	wire [16-1:0] node8737;
	wire [16-1:0] node8738;
	wire [16-1:0] node8740;
	wire [16-1:0] node8743;
	wire [16-1:0] node8744;
	wire [16-1:0] node8747;
	wire [16-1:0] node8750;
	wire [16-1:0] node8751;
	wire [16-1:0] node8752;
	wire [16-1:0] node8753;
	wire [16-1:0] node8754;
	wire [16-1:0] node8757;
	wire [16-1:0] node8758;
	wire [16-1:0] node8762;
	wire [16-1:0] node8763;
	wire [16-1:0] node8765;
	wire [16-1:0] node8769;
	wire [16-1:0] node8770;
	wire [16-1:0] node8773;
	wire [16-1:0] node8775;
	wire [16-1:0] node8778;
	wire [16-1:0] node8779;
	wire [16-1:0] node8780;
	wire [16-1:0] node8782;
	wire [16-1:0] node8783;
	wire [16-1:0] node8787;
	wire [16-1:0] node8788;
	wire [16-1:0] node8791;
	wire [16-1:0] node8793;
	wire [16-1:0] node8796;
	wire [16-1:0] node8797;
	wire [16-1:0] node8800;
	wire [16-1:0] node8802;
	wire [16-1:0] node8804;
	wire [16-1:0] node8807;
	wire [16-1:0] node8808;
	wire [16-1:0] node8809;
	wire [16-1:0] node8810;
	wire [16-1:0] node8811;
	wire [16-1:0] node8812;
	wire [16-1:0] node8815;
	wire [16-1:0] node8816;
	wire [16-1:0] node8817;
	wire [16-1:0] node8822;
	wire [16-1:0] node8823;
	wire [16-1:0] node8824;
	wire [16-1:0] node8827;
	wire [16-1:0] node8830;
	wire [16-1:0] node8832;
	wire [16-1:0] node8835;
	wire [16-1:0] node8836;
	wire [16-1:0] node8837;
	wire [16-1:0] node8838;
	wire [16-1:0] node8842;
	wire [16-1:0] node8845;
	wire [16-1:0] node8847;
	wire [16-1:0] node8850;
	wire [16-1:0] node8851;
	wire [16-1:0] node8852;
	wire [16-1:0] node8853;
	wire [16-1:0] node8855;
	wire [16-1:0] node8858;
	wire [16-1:0] node8860;
	wire [16-1:0] node8862;
	wire [16-1:0] node8865;
	wire [16-1:0] node8866;
	wire [16-1:0] node8869;
	wire [16-1:0] node8870;
	wire [16-1:0] node8874;
	wire [16-1:0] node8875;
	wire [16-1:0] node8876;
	wire [16-1:0] node8879;
	wire [16-1:0] node8880;
	wire [16-1:0] node8881;
	wire [16-1:0] node8886;
	wire [16-1:0] node8887;
	wire [16-1:0] node8888;
	wire [16-1:0] node8892;
	wire [16-1:0] node8894;
	wire [16-1:0] node8897;
	wire [16-1:0] node8898;
	wire [16-1:0] node8899;
	wire [16-1:0] node8900;
	wire [16-1:0] node8901;
	wire [16-1:0] node8903;
	wire [16-1:0] node8905;
	wire [16-1:0] node8908;
	wire [16-1:0] node8911;
	wire [16-1:0] node8912;
	wire [16-1:0] node8914;
	wire [16-1:0] node8917;
	wire [16-1:0] node8920;
	wire [16-1:0] node8921;
	wire [16-1:0] node8922;
	wire [16-1:0] node8924;
	wire [16-1:0] node8926;
	wire [16-1:0] node8929;
	wire [16-1:0] node8932;
	wire [16-1:0] node8934;
	wire [16-1:0] node8936;
	wire [16-1:0] node8939;
	wire [16-1:0] node8940;
	wire [16-1:0] node8941;
	wire [16-1:0] node8942;
	wire [16-1:0] node8945;
	wire [16-1:0] node8946;
	wire [16-1:0] node8947;
	wire [16-1:0] node8952;
	wire [16-1:0] node8953;
	wire [16-1:0] node8955;
	wire [16-1:0] node8957;
	wire [16-1:0] node8960;
	wire [16-1:0] node8963;
	wire [16-1:0] node8964;
	wire [16-1:0] node8965;
	wire [16-1:0] node8966;
	wire [16-1:0] node8969;
	wire [16-1:0] node8971;
	wire [16-1:0] node8975;
	wire [16-1:0] node8976;
	wire [16-1:0] node8977;
	wire [16-1:0] node8978;
	wire [16-1:0] node8981;
	wire [16-1:0] node8985;
	wire [16-1:0] node8987;
	wire [16-1:0] node8990;
	wire [16-1:0] node8991;
	wire [16-1:0] node8992;
	wire [16-1:0] node8993;
	wire [16-1:0] node8994;
	wire [16-1:0] node8995;
	wire [16-1:0] node8996;
	wire [16-1:0] node8998;
	wire [16-1:0] node8999;
	wire [16-1:0] node9000;
	wire [16-1:0] node9005;
	wire [16-1:0] node9007;
	wire [16-1:0] node9010;
	wire [16-1:0] node9011;
	wire [16-1:0] node9012;
	wire [16-1:0] node9015;
	wire [16-1:0] node9018;
	wire [16-1:0] node9019;
	wire [16-1:0] node9023;
	wire [16-1:0] node9024;
	wire [16-1:0] node9025;
	wire [16-1:0] node9027;
	wire [16-1:0] node9030;
	wire [16-1:0] node9033;
	wire [16-1:0] node9034;
	wire [16-1:0] node9037;
	wire [16-1:0] node9039;
	wire [16-1:0] node9042;
	wire [16-1:0] node9043;
	wire [16-1:0] node9044;
	wire [16-1:0] node9045;
	wire [16-1:0] node9047;
	wire [16-1:0] node9050;
	wire [16-1:0] node9052;
	wire [16-1:0] node9055;
	wire [16-1:0] node9057;
	wire [16-1:0] node9060;
	wire [16-1:0] node9061;
	wire [16-1:0] node9062;
	wire [16-1:0] node9065;
	wire [16-1:0] node9067;
	wire [16-1:0] node9070;
	wire [16-1:0] node9071;
	wire [16-1:0] node9073;
	wire [16-1:0] node9074;
	wire [16-1:0] node9078;
	wire [16-1:0] node9081;
	wire [16-1:0] node9082;
	wire [16-1:0] node9083;
	wire [16-1:0] node9084;
	wire [16-1:0] node9085;
	wire [16-1:0] node9086;
	wire [16-1:0] node9091;
	wire [16-1:0] node9092;
	wire [16-1:0] node9094;
	wire [16-1:0] node9097;
	wire [16-1:0] node9098;
	wire [16-1:0] node9102;
	wire [16-1:0] node9103;
	wire [16-1:0] node9104;
	wire [16-1:0] node9108;
	wire [16-1:0] node9109;
	wire [16-1:0] node9111;
	wire [16-1:0] node9112;
	wire [16-1:0] node9117;
	wire [16-1:0] node9118;
	wire [16-1:0] node9119;
	wire [16-1:0] node9120;
	wire [16-1:0] node9121;
	wire [16-1:0] node9124;
	wire [16-1:0] node9126;
	wire [16-1:0] node9130;
	wire [16-1:0] node9132;
	wire [16-1:0] node9135;
	wire [16-1:0] node9136;
	wire [16-1:0] node9138;
	wire [16-1:0] node9139;
	wire [16-1:0] node9143;
	wire [16-1:0] node9146;
	wire [16-1:0] node9147;
	wire [16-1:0] node9148;
	wire [16-1:0] node9149;
	wire [16-1:0] node9150;
	wire [16-1:0] node9151;
	wire [16-1:0] node9153;
	wire [16-1:0] node9154;
	wire [16-1:0] node9156;
	wire [16-1:0] node9160;
	wire [16-1:0] node9163;
	wire [16-1:0] node9164;
	wire [16-1:0] node9165;
	wire [16-1:0] node9166;
	wire [16-1:0] node9171;
	wire [16-1:0] node9172;
	wire [16-1:0] node9174;
	wire [16-1:0] node9177;
	wire [16-1:0] node9178;
	wire [16-1:0] node9179;
	wire [16-1:0] node9183;
	wire [16-1:0] node9186;
	wire [16-1:0] node9187;
	wire [16-1:0] node9188;
	wire [16-1:0] node9189;
	wire [16-1:0] node9192;
	wire [16-1:0] node9194;
	wire [16-1:0] node9197;
	wire [16-1:0] node9199;
	wire [16-1:0] node9202;
	wire [16-1:0] node9203;
	wire [16-1:0] node9205;
	wire [16-1:0] node9208;
	wire [16-1:0] node9211;
	wire [16-1:0] node9212;
	wire [16-1:0] node9214;
	wire [16-1:0] node9215;
	wire [16-1:0] node9217;
	wire [16-1:0] node9218;
	wire [16-1:0] node9223;
	wire [16-1:0] node9224;
	wire [16-1:0] node9225;
	wire [16-1:0] node9226;
	wire [16-1:0] node9228;
	wire [16-1:0] node9233;
	wire [16-1:0] node9234;
	wire [16-1:0] node9235;
	wire [16-1:0] node9236;
	wire [16-1:0] node9240;
	wire [16-1:0] node9242;
	wire [16-1:0] node9245;
	wire [16-1:0] node9247;
	wire [16-1:0] node9250;
	wire [16-1:0] node9251;
	wire [16-1:0] node9252;
	wire [16-1:0] node9253;
	wire [16-1:0] node9254;
	wire [16-1:0] node9255;
	wire [16-1:0] node9260;
	wire [16-1:0] node9261;
	wire [16-1:0] node9262;
	wire [16-1:0] node9265;
	wire [16-1:0] node9266;
	wire [16-1:0] node9268;
	wire [16-1:0] node9272;
	wire [16-1:0] node9274;
	wire [16-1:0] node9277;
	wire [16-1:0] node9278;
	wire [16-1:0] node9279;
	wire [16-1:0] node9280;
	wire [16-1:0] node9282;
	wire [16-1:0] node9283;
	wire [16-1:0] node9288;
	wire [16-1:0] node9291;
	wire [16-1:0] node9292;
	wire [16-1:0] node9295;
	wire [16-1:0] node9297;
	wire [16-1:0] node9299;
	wire [16-1:0] node9302;
	wire [16-1:0] node9303;
	wire [16-1:0] node9304;
	wire [16-1:0] node9306;
	wire [16-1:0] node9307;
	wire [16-1:0] node9311;
	wire [16-1:0] node9312;
	wire [16-1:0] node9315;
	wire [16-1:0] node9317;
	wire [16-1:0] node9320;
	wire [16-1:0] node9321;
	wire [16-1:0] node9322;
	wire [16-1:0] node9324;
	wire [16-1:0] node9327;
	wire [16-1:0] node9328;
	wire [16-1:0] node9330;
	wire [16-1:0] node9331;
	wire [16-1:0] node9336;
	wire [16-1:0] node9338;
	wire [16-1:0] node9340;
	wire [16-1:0] node9341;
	wire [16-1:0] node9345;
	wire [16-1:0] node9346;
	wire [16-1:0] node9347;
	wire [16-1:0] node9348;
	wire [16-1:0] node9349;
	wire [16-1:0] node9350;
	wire [16-1:0] node9351;
	wire [16-1:0] node9352;
	wire [16-1:0] node9354;
	wire [16-1:0] node9357;
	wire [16-1:0] node9358;
	wire [16-1:0] node9360;
	wire [16-1:0] node9364;
	wire [16-1:0] node9367;
	wire [16-1:0] node9369;
	wire [16-1:0] node9370;
	wire [16-1:0] node9371;
	wire [16-1:0] node9374;
	wire [16-1:0] node9376;
	wire [16-1:0] node9379;
	wire [16-1:0] node9382;
	wire [16-1:0] node9383;
	wire [16-1:0] node9384;
	wire [16-1:0] node9385;
	wire [16-1:0] node9386;
	wire [16-1:0] node9389;
	wire [16-1:0] node9390;
	wire [16-1:0] node9394;
	wire [16-1:0] node9397;
	wire [16-1:0] node9398;
	wire [16-1:0] node9400;
	wire [16-1:0] node9403;
	wire [16-1:0] node9406;
	wire [16-1:0] node9407;
	wire [16-1:0] node9408;
	wire [16-1:0] node9411;
	wire [16-1:0] node9413;
	wire [16-1:0] node9416;
	wire [16-1:0] node9417;
	wire [16-1:0] node9419;
	wire [16-1:0] node9422;
	wire [16-1:0] node9425;
	wire [16-1:0] node9426;
	wire [16-1:0] node9427;
	wire [16-1:0] node9428;
	wire [16-1:0] node9429;
	wire [16-1:0] node9430;
	wire [16-1:0] node9433;
	wire [16-1:0] node9436;
	wire [16-1:0] node9437;
	wire [16-1:0] node9441;
	wire [16-1:0] node9443;
	wire [16-1:0] node9444;
	wire [16-1:0] node9448;
	wire [16-1:0] node9449;
	wire [16-1:0] node9450;
	wire [16-1:0] node9451;
	wire [16-1:0] node9455;
	wire [16-1:0] node9458;
	wire [16-1:0] node9459;
	wire [16-1:0] node9460;
	wire [16-1:0] node9462;
	wire [16-1:0] node9466;
	wire [16-1:0] node9468;
	wire [16-1:0] node9471;
	wire [16-1:0] node9472;
	wire [16-1:0] node9473;
	wire [16-1:0] node9474;
	wire [16-1:0] node9477;
	wire [16-1:0] node9479;
	wire [16-1:0] node9480;
	wire [16-1:0] node9484;
	wire [16-1:0] node9485;
	wire [16-1:0] node9488;
	wire [16-1:0] node9491;
	wire [16-1:0] node9492;
	wire [16-1:0] node9494;
	wire [16-1:0] node9497;
	wire [16-1:0] node9498;
	wire [16-1:0] node9502;
	wire [16-1:0] node9503;
	wire [16-1:0] node9504;
	wire [16-1:0] node9505;
	wire [16-1:0] node9506;
	wire [16-1:0] node9508;
	wire [16-1:0] node9510;
	wire [16-1:0] node9511;
	wire [16-1:0] node9515;
	wire [16-1:0] node9516;
	wire [16-1:0] node9517;
	wire [16-1:0] node9519;
	wire [16-1:0] node9524;
	wire [16-1:0] node9525;
	wire [16-1:0] node9526;
	wire [16-1:0] node9527;
	wire [16-1:0] node9529;
	wire [16-1:0] node9532;
	wire [16-1:0] node9533;
	wire [16-1:0] node9537;
	wire [16-1:0] node9539;
	wire [16-1:0] node9542;
	wire [16-1:0] node9543;
	wire [16-1:0] node9546;
	wire [16-1:0] node9549;
	wire [16-1:0] node9550;
	wire [16-1:0] node9551;
	wire [16-1:0] node9552;
	wire [16-1:0] node9553;
	wire [16-1:0] node9556;
	wire [16-1:0] node9559;
	wire [16-1:0] node9561;
	wire [16-1:0] node9564;
	wire [16-1:0] node9565;
	wire [16-1:0] node9566;
	wire [16-1:0] node9570;
	wire [16-1:0] node9572;
	wire [16-1:0] node9574;
	wire [16-1:0] node9577;
	wire [16-1:0] node9578;
	wire [16-1:0] node9579;
	wire [16-1:0] node9582;
	wire [16-1:0] node9585;
	wire [16-1:0] node9586;
	wire [16-1:0] node9587;
	wire [16-1:0] node9590;
	wire [16-1:0] node9592;
	wire [16-1:0] node9595;
	wire [16-1:0] node9597;
	wire [16-1:0] node9600;
	wire [16-1:0] node9601;
	wire [16-1:0] node9602;
	wire [16-1:0] node9603;
	wire [16-1:0] node9604;
	wire [16-1:0] node9605;
	wire [16-1:0] node9607;
	wire [16-1:0] node9612;
	wire [16-1:0] node9613;
	wire [16-1:0] node9614;
	wire [16-1:0] node9618;
	wire [16-1:0] node9620;
	wire [16-1:0] node9621;
	wire [16-1:0] node9622;
	wire [16-1:0] node9627;
	wire [16-1:0] node9628;
	wire [16-1:0] node9629;
	wire [16-1:0] node9630;
	wire [16-1:0] node9634;
	wire [16-1:0] node9635;
	wire [16-1:0] node9639;
	wire [16-1:0] node9640;
	wire [16-1:0] node9643;
	wire [16-1:0] node9644;
	wire [16-1:0] node9648;
	wire [16-1:0] node9649;
	wire [16-1:0] node9650;
	wire [16-1:0] node9652;
	wire [16-1:0] node9654;
	wire [16-1:0] node9656;
	wire [16-1:0] node9659;
	wire [16-1:0] node9660;
	wire [16-1:0] node9661;
	wire [16-1:0] node9665;
	wire [16-1:0] node9668;
	wire [16-1:0] node9669;
	wire [16-1:0] node9670;
	wire [16-1:0] node9674;
	wire [16-1:0] node9676;
	wire [16-1:0] node9679;
	wire [16-1:0] node9680;
	wire [16-1:0] node9681;
	wire [16-1:0] node9682;
	wire [16-1:0] node9683;
	wire [16-1:0] node9684;
	wire [16-1:0] node9685;
	wire [16-1:0] node9686;
	wire [16-1:0] node9691;
	wire [16-1:0] node9692;
	wire [16-1:0] node9695;
	wire [16-1:0] node9698;
	wire [16-1:0] node9699;
	wire [16-1:0] node9700;
	wire [16-1:0] node9701;
	wire [16-1:0] node9704;
	wire [16-1:0] node9707;
	wire [16-1:0] node9708;
	wire [16-1:0] node9712;
	wire [16-1:0] node9713;
	wire [16-1:0] node9715;
	wire [16-1:0] node9718;
	wire [16-1:0] node9719;
	wire [16-1:0] node9721;
	wire [16-1:0] node9724;
	wire [16-1:0] node9727;
	wire [16-1:0] node9728;
	wire [16-1:0] node9729;
	wire [16-1:0] node9730;
	wire [16-1:0] node9731;
	wire [16-1:0] node9735;
	wire [16-1:0] node9738;
	wire [16-1:0] node9739;
	wire [16-1:0] node9741;
	wire [16-1:0] node9744;
	wire [16-1:0] node9745;
	wire [16-1:0] node9746;
	wire [16-1:0] node9747;
	wire [16-1:0] node9753;
	wire [16-1:0] node9754;
	wire [16-1:0] node9755;
	wire [16-1:0] node9757;
	wire [16-1:0] node9760;
	wire [16-1:0] node9761;
	wire [16-1:0] node9765;
	wire [16-1:0] node9766;
	wire [16-1:0] node9769;
	wire [16-1:0] node9770;
	wire [16-1:0] node9774;
	wire [16-1:0] node9775;
	wire [16-1:0] node9776;
	wire [16-1:0] node9777;
	wire [16-1:0] node9778;
	wire [16-1:0] node9779;
	wire [16-1:0] node9782;
	wire [16-1:0] node9786;
	wire [16-1:0] node9787;
	wire [16-1:0] node9790;
	wire [16-1:0] node9792;
	wire [16-1:0] node9793;
	wire [16-1:0] node9797;
	wire [16-1:0] node9798;
	wire [16-1:0] node9799;
	wire [16-1:0] node9801;
	wire [16-1:0] node9802;
	wire [16-1:0] node9806;
	wire [16-1:0] node9809;
	wire [16-1:0] node9810;
	wire [16-1:0] node9811;
	wire [16-1:0] node9815;
	wire [16-1:0] node9817;
	wire [16-1:0] node9820;
	wire [16-1:0] node9821;
	wire [16-1:0] node9822;
	wire [16-1:0] node9823;
	wire [16-1:0] node9827;
	wire [16-1:0] node9828;
	wire [16-1:0] node9830;
	wire [16-1:0] node9833;
	wire [16-1:0] node9835;
	wire [16-1:0] node9838;
	wire [16-1:0] node9839;
	wire [16-1:0] node9841;
	wire [16-1:0] node9842;
	wire [16-1:0] node9843;
	wire [16-1:0] node9846;
	wire [16-1:0] node9849;
	wire [16-1:0] node9852;
	wire [16-1:0] node9853;
	wire [16-1:0] node9854;
	wire [16-1:0] node9858;
	wire [16-1:0] node9860;
	wire [16-1:0] node9862;
	wire [16-1:0] node9864;
	wire [16-1:0] node9867;
	wire [16-1:0] node9868;
	wire [16-1:0] node9869;
	wire [16-1:0] node9870;
	wire [16-1:0] node9871;
	wire [16-1:0] node9872;
	wire [16-1:0] node9875;
	wire [16-1:0] node9878;
	wire [16-1:0] node9880;
	wire [16-1:0] node9883;
	wire [16-1:0] node9884;
	wire [16-1:0] node9885;
	wire [16-1:0] node9886;
	wire [16-1:0] node9891;
	wire [16-1:0] node9892;
	wire [16-1:0] node9894;
	wire [16-1:0] node9897;
	wire [16-1:0] node9900;
	wire [16-1:0] node9901;
	wire [16-1:0] node9902;
	wire [16-1:0] node9903;
	wire [16-1:0] node9906;
	wire [16-1:0] node9908;
	wire [16-1:0] node9909;
	wire [16-1:0] node9913;
	wire [16-1:0] node9914;
	wire [16-1:0] node9915;
	wire [16-1:0] node9918;
	wire [16-1:0] node9920;
	wire [16-1:0] node9924;
	wire [16-1:0] node9925;
	wire [16-1:0] node9927;
	wire [16-1:0] node9930;
	wire [16-1:0] node9931;
	wire [16-1:0] node9934;
	wire [16-1:0] node9937;
	wire [16-1:0] node9938;
	wire [16-1:0] node9939;
	wire [16-1:0] node9940;
	wire [16-1:0] node9942;
	wire [16-1:0] node9945;
	wire [16-1:0] node9946;
	wire [16-1:0] node9947;
	wire [16-1:0] node9950;
	wire [16-1:0] node9953;
	wire [16-1:0] node9954;
	wire [16-1:0] node9955;
	wire [16-1:0] node9959;
	wire [16-1:0] node9961;
	wire [16-1:0] node9964;
	wire [16-1:0] node9965;
	wire [16-1:0] node9966;
	wire [16-1:0] node9969;
	wire [16-1:0] node9970;
	wire [16-1:0] node9971;
	wire [16-1:0] node9975;
	wire [16-1:0] node9977;
	wire [16-1:0] node9980;
	wire [16-1:0] node9981;
	wire [16-1:0] node9982;
	wire [16-1:0] node9986;
	wire [16-1:0] node9987;
	wire [16-1:0] node9990;
	wire [16-1:0] node9993;
	wire [16-1:0] node9994;
	wire [16-1:0] node9995;
	wire [16-1:0] node9996;
	wire [16-1:0] node10000;
	wire [16-1:0] node10001;
	wire [16-1:0] node10002;
	wire [16-1:0] node10004;
	wire [16-1:0] node10008;
	wire [16-1:0] node10009;
	wire [16-1:0] node10013;
	wire [16-1:0] node10014;
	wire [16-1:0] node10015;
	wire [16-1:0] node10017;
	wire [16-1:0] node10021;
	wire [16-1:0] node10022;
	wire [16-1:0] node10023;
	wire [16-1:0] node10026;
	wire [16-1:0] node10028;
	wire [16-1:0] node10031;
	wire [16-1:0] node10032;
	wire [16-1:0] node10035;
	wire [16-1:0] node10037;
	wire [16-1:0] node10040;
	wire [16-1:0] node10041;
	wire [16-1:0] node10042;
	wire [16-1:0] node10043;
	wire [16-1:0] node10044;
	wire [16-1:0] node10045;
	wire [16-1:0] node10046;
	wire [16-1:0] node10047;
	wire [16-1:0] node10048;
	wire [16-1:0] node10051;
	wire [16-1:0] node10054;
	wire [16-1:0] node10056;
	wire [16-1:0] node10059;
	wire [16-1:0] node10060;
	wire [16-1:0] node10061;
	wire [16-1:0] node10064;
	wire [16-1:0] node10067;
	wire [16-1:0] node10070;
	wire [16-1:0] node10071;
	wire [16-1:0] node10072;
	wire [16-1:0] node10073;
	wire [16-1:0] node10074;
	wire [16-1:0] node10078;
	wire [16-1:0] node10079;
	wire [16-1:0] node10082;
	wire [16-1:0] node10084;
	wire [16-1:0] node10087;
	wire [16-1:0] node10088;
	wire [16-1:0] node10089;
	wire [16-1:0] node10093;
	wire [16-1:0] node10094;
	wire [16-1:0] node10095;
	wire [16-1:0] node10098;
	wire [16-1:0] node10102;
	wire [16-1:0] node10103;
	wire [16-1:0] node10106;
	wire [16-1:0] node10107;
	wire [16-1:0] node10108;
	wire [16-1:0] node10112;
	wire [16-1:0] node10115;
	wire [16-1:0] node10116;
	wire [16-1:0] node10117;
	wire [16-1:0] node10118;
	wire [16-1:0] node10119;
	wire [16-1:0] node10120;
	wire [16-1:0] node10123;
	wire [16-1:0] node10124;
	wire [16-1:0] node10127;
	wire [16-1:0] node10131;
	wire [16-1:0] node10132;
	wire [16-1:0] node10133;
	wire [16-1:0] node10138;
	wire [16-1:0] node10139;
	wire [16-1:0] node10140;
	wire [16-1:0] node10143;
	wire [16-1:0] node10145;
	wire [16-1:0] node10148;
	wire [16-1:0] node10149;
	wire [16-1:0] node10150;
	wire [16-1:0] node10153;
	wire [16-1:0] node10155;
	wire [16-1:0] node10158;
	wire [16-1:0] node10159;
	wire [16-1:0] node10161;
	wire [16-1:0] node10165;
	wire [16-1:0] node10166;
	wire [16-1:0] node10167;
	wire [16-1:0] node10168;
	wire [16-1:0] node10172;
	wire [16-1:0] node10174;
	wire [16-1:0] node10177;
	wire [16-1:0] node10178;
	wire [16-1:0] node10180;
	wire [16-1:0] node10182;
	wire [16-1:0] node10185;
	wire [16-1:0] node10186;
	wire [16-1:0] node10187;
	wire [16-1:0] node10190;
	wire [16-1:0] node10192;
	wire [16-1:0] node10195;
	wire [16-1:0] node10197;
	wire [16-1:0] node10200;
	wire [16-1:0] node10201;
	wire [16-1:0] node10202;
	wire [16-1:0] node10203;
	wire [16-1:0] node10204;
	wire [16-1:0] node10207;
	wire [16-1:0] node10209;
	wire [16-1:0] node10212;
	wire [16-1:0] node10213;
	wire [16-1:0] node10214;
	wire [16-1:0] node10215;
	wire [16-1:0] node10219;
	wire [16-1:0] node10222;
	wire [16-1:0] node10224;
	wire [16-1:0] node10225;
	wire [16-1:0] node10229;
	wire [16-1:0] node10230;
	wire [16-1:0] node10231;
	wire [16-1:0] node10232;
	wire [16-1:0] node10233;
	wire [16-1:0] node10238;
	wire [16-1:0] node10239;
	wire [16-1:0] node10241;
	wire [16-1:0] node10244;
	wire [16-1:0] node10247;
	wire [16-1:0] node10248;
	wire [16-1:0] node10249;
	wire [16-1:0] node10250;
	wire [16-1:0] node10251;
	wire [16-1:0] node10254;
	wire [16-1:0] node10258;
	wire [16-1:0] node10259;
	wire [16-1:0] node10262;
	wire [16-1:0] node10265;
	wire [16-1:0] node10266;
	wire [16-1:0] node10268;
	wire [16-1:0] node10271;
	wire [16-1:0] node10272;
	wire [16-1:0] node10273;
	wire [16-1:0] node10278;
	wire [16-1:0] node10279;
	wire [16-1:0] node10280;
	wire [16-1:0] node10281;
	wire [16-1:0] node10282;
	wire [16-1:0] node10283;
	wire [16-1:0] node10284;
	wire [16-1:0] node10290;
	wire [16-1:0] node10291;
	wire [16-1:0] node10292;
	wire [16-1:0] node10295;
	wire [16-1:0] node10298;
	wire [16-1:0] node10299;
	wire [16-1:0] node10300;
	wire [16-1:0] node10305;
	wire [16-1:0] node10306;
	wire [16-1:0] node10307;
	wire [16-1:0] node10311;
	wire [16-1:0] node10313;
	wire [16-1:0] node10314;
	wire [16-1:0] node10318;
	wire [16-1:0] node10319;
	wire [16-1:0] node10320;
	wire [16-1:0] node10321;
	wire [16-1:0] node10324;
	wire [16-1:0] node10327;
	wire [16-1:0] node10328;
	wire [16-1:0] node10329;
	wire [16-1:0] node10333;
	wire [16-1:0] node10335;
	wire [16-1:0] node10338;
	wire [16-1:0] node10339;
	wire [16-1:0] node10341;
	wire [16-1:0] node10342;
	wire [16-1:0] node10346;
	wire [16-1:0] node10347;
	wire [16-1:0] node10350;
	wire [16-1:0] node10353;
	wire [16-1:0] node10354;
	wire [16-1:0] node10355;
	wire [16-1:0] node10356;
	wire [16-1:0] node10357;
	wire [16-1:0] node10358;
	wire [16-1:0] node10359;
	wire [16-1:0] node10360;
	wire [16-1:0] node10361;
	wire [16-1:0] node10363;
	wire [16-1:0] node10368;
	wire [16-1:0] node10370;
	wire [16-1:0] node10373;
	wire [16-1:0] node10374;
	wire [16-1:0] node10377;
	wire [16-1:0] node10380;
	wire [16-1:0] node10381;
	wire [16-1:0] node10383;
	wire [16-1:0] node10386;
	wire [16-1:0] node10387;
	wire [16-1:0] node10388;
	wire [16-1:0] node10390;
	wire [16-1:0] node10394;
	wire [16-1:0] node10397;
	wire [16-1:0] node10398;
	wire [16-1:0] node10399;
	wire [16-1:0] node10400;
	wire [16-1:0] node10403;
	wire [16-1:0] node10404;
	wire [16-1:0] node10405;
	wire [16-1:0] node10408;
	wire [16-1:0] node10412;
	wire [16-1:0] node10413;
	wire [16-1:0] node10415;
	wire [16-1:0] node10417;
	wire [16-1:0] node10419;
	wire [16-1:0] node10422;
	wire [16-1:0] node10423;
	wire [16-1:0] node10424;
	wire [16-1:0] node10429;
	wire [16-1:0] node10430;
	wire [16-1:0] node10432;
	wire [16-1:0] node10434;
	wire [16-1:0] node10435;
	wire [16-1:0] node10439;
	wire [16-1:0] node10440;
	wire [16-1:0] node10441;
	wire [16-1:0] node10444;
	wire [16-1:0] node10447;
	wire [16-1:0] node10450;
	wire [16-1:0] node10451;
	wire [16-1:0] node10452;
	wire [16-1:0] node10453;
	wire [16-1:0] node10454;
	wire [16-1:0] node10456;
	wire [16-1:0] node10459;
	wire [16-1:0] node10461;
	wire [16-1:0] node10462;
	wire [16-1:0] node10463;
	wire [16-1:0] node10468;
	wire [16-1:0] node10469;
	wire [16-1:0] node10471;
	wire [16-1:0] node10474;
	wire [16-1:0] node10476;
	wire [16-1:0] node10479;
	wire [16-1:0] node10480;
	wire [16-1:0] node10482;
	wire [16-1:0] node10484;
	wire [16-1:0] node10485;
	wire [16-1:0] node10487;
	wire [16-1:0] node10491;
	wire [16-1:0] node10492;
	wire [16-1:0] node10496;
	wire [16-1:0] node10497;
	wire [16-1:0] node10498;
	wire [16-1:0] node10499;
	wire [16-1:0] node10502;
	wire [16-1:0] node10505;
	wire [16-1:0] node10506;
	wire [16-1:0] node10507;
	wire [16-1:0] node10510;
	wire [16-1:0] node10514;
	wire [16-1:0] node10515;
	wire [16-1:0] node10516;
	wire [16-1:0] node10517;
	wire [16-1:0] node10520;
	wire [16-1:0] node10522;
	wire [16-1:0] node10525;
	wire [16-1:0] node10526;
	wire [16-1:0] node10529;
	wire [16-1:0] node10532;
	wire [16-1:0] node10534;
	wire [16-1:0] node10535;
	wire [16-1:0] node10538;
	wire [16-1:0] node10541;
	wire [16-1:0] node10542;
	wire [16-1:0] node10543;
	wire [16-1:0] node10544;
	wire [16-1:0] node10545;
	wire [16-1:0] node10546;
	wire [16-1:0] node10550;
	wire [16-1:0] node10552;
	wire [16-1:0] node10554;
	wire [16-1:0] node10556;
	wire [16-1:0] node10559;
	wire [16-1:0] node10560;
	wire [16-1:0] node10561;
	wire [16-1:0] node10565;
	wire [16-1:0] node10567;
	wire [16-1:0] node10569;
	wire [16-1:0] node10572;
	wire [16-1:0] node10573;
	wire [16-1:0] node10574;
	wire [16-1:0] node10575;
	wire [16-1:0] node10576;
	wire [16-1:0] node10580;
	wire [16-1:0] node10581;
	wire [16-1:0] node10583;
	wire [16-1:0] node10587;
	wire [16-1:0] node10588;
	wire [16-1:0] node10591;
	wire [16-1:0] node10592;
	wire [16-1:0] node10593;
	wire [16-1:0] node10596;
	wire [16-1:0] node10600;
	wire [16-1:0] node10601;
	wire [16-1:0] node10603;
	wire [16-1:0] node10606;
	wire [16-1:0] node10607;
	wire [16-1:0] node10610;
	wire [16-1:0] node10613;
	wire [16-1:0] node10614;
	wire [16-1:0] node10615;
	wire [16-1:0] node10616;
	wire [16-1:0] node10617;
	wire [16-1:0] node10618;
	wire [16-1:0] node10619;
	wire [16-1:0] node10625;
	wire [16-1:0] node10626;
	wire [16-1:0] node10629;
	wire [16-1:0] node10630;
	wire [16-1:0] node10631;
	wire [16-1:0] node10632;
	wire [16-1:0] node10636;
	wire [16-1:0] node10637;
	wire [16-1:0] node10642;
	wire [16-1:0] node10643;
	wire [16-1:0] node10644;
	wire [16-1:0] node10646;
	wire [16-1:0] node10649;
	wire [16-1:0] node10650;
	wire [16-1:0] node10654;
	wire [16-1:0] node10655;
	wire [16-1:0] node10658;
	wire [16-1:0] node10659;
	wire [16-1:0] node10661;
	wire [16-1:0] node10665;
	wire [16-1:0] node10666;
	wire [16-1:0] node10667;
	wire [16-1:0] node10668;
	wire [16-1:0] node10669;
	wire [16-1:0] node10671;
	wire [16-1:0] node10675;
	wire [16-1:0] node10677;
	wire [16-1:0] node10680;
	wire [16-1:0] node10681;
	wire [16-1:0] node10682;
	wire [16-1:0] node10683;
	wire [16-1:0] node10688;
	wire [16-1:0] node10690;
	wire [16-1:0] node10691;
	wire [16-1:0] node10695;
	wire [16-1:0] node10696;
	wire [16-1:0] node10697;
	wire [16-1:0] node10698;
	wire [16-1:0] node10701;
	wire [16-1:0] node10704;
	wire [16-1:0] node10705;
	wire [16-1:0] node10708;
	wire [16-1:0] node10710;
	wire [16-1:0] node10713;
	wire [16-1:0] node10714;
	wire [16-1:0] node10717;
	wire [16-1:0] node10720;
	wire [16-1:0] node10721;
	wire [16-1:0] node10722;
	wire [16-1:0] node10723;
	wire [16-1:0] node10724;
	wire [16-1:0] node10725;
	wire [16-1:0] node10726;
	wire [16-1:0] node10728;
	wire [16-1:0] node10729;
	wire [16-1:0] node10731;
	wire [16-1:0] node10735;
	wire [16-1:0] node10736;
	wire [16-1:0] node10737;
	wire [16-1:0] node10741;
	wire [16-1:0] node10743;
	wire [16-1:0] node10744;
	wire [16-1:0] node10748;
	wire [16-1:0] node10749;
	wire [16-1:0] node10750;
	wire [16-1:0] node10751;
	wire [16-1:0] node10755;
	wire [16-1:0] node10756;
	wire [16-1:0] node10758;
	wire [16-1:0] node10760;
	wire [16-1:0] node10764;
	wire [16-1:0] node10765;
	wire [16-1:0] node10768;
	wire [16-1:0] node10771;
	wire [16-1:0] node10772;
	wire [16-1:0] node10773;
	wire [16-1:0] node10774;
	wire [16-1:0] node10776;
	wire [16-1:0] node10779;
	wire [16-1:0] node10780;
	wire [16-1:0] node10781;
	wire [16-1:0] node10784;
	wire [16-1:0] node10788;
	wire [16-1:0] node10789;
	wire [16-1:0] node10790;
	wire [16-1:0] node10791;
	wire [16-1:0] node10795;
	wire [16-1:0] node10797;
	wire [16-1:0] node10800;
	wire [16-1:0] node10803;
	wire [16-1:0] node10805;
	wire [16-1:0] node10807;
	wire [16-1:0] node10808;
	wire [16-1:0] node10810;
	wire [16-1:0] node10814;
	wire [16-1:0] node10815;
	wire [16-1:0] node10816;
	wire [16-1:0] node10817;
	wire [16-1:0] node10818;
	wire [16-1:0] node10821;
	wire [16-1:0] node10823;
	wire [16-1:0] node10826;
	wire [16-1:0] node10827;
	wire [16-1:0] node10830;
	wire [16-1:0] node10833;
	wire [16-1:0] node10834;
	wire [16-1:0] node10835;
	wire [16-1:0] node10838;
	wire [16-1:0] node10841;
	wire [16-1:0] node10842;
	wire [16-1:0] node10845;
	wire [16-1:0] node10846;
	wire [16-1:0] node10850;
	wire [16-1:0] node10851;
	wire [16-1:0] node10852;
	wire [16-1:0] node10853;
	wire [16-1:0] node10854;
	wire [16-1:0] node10856;
	wire [16-1:0] node10860;
	wire [16-1:0] node10862;
	wire [16-1:0] node10865;
	wire [16-1:0] node10866;
	wire [16-1:0] node10867;
	wire [16-1:0] node10871;
	wire [16-1:0] node10872;
	wire [16-1:0] node10875;
	wire [16-1:0] node10877;
	wire [16-1:0] node10878;
	wire [16-1:0] node10882;
	wire [16-1:0] node10883;
	wire [16-1:0] node10885;
	wire [16-1:0] node10886;
	wire [16-1:0] node10887;
	wire [16-1:0] node10890;
	wire [16-1:0] node10893;
	wire [16-1:0] node10896;
	wire [16-1:0] node10897;
	wire [16-1:0] node10900;
	wire [16-1:0] node10902;
	wire [16-1:0] node10905;
	wire [16-1:0] node10906;
	wire [16-1:0] node10907;
	wire [16-1:0] node10908;
	wire [16-1:0] node10910;
	wire [16-1:0] node10911;
	wire [16-1:0] node10912;
	wire [16-1:0] node10915;
	wire [16-1:0] node10916;
	wire [16-1:0] node10920;
	wire [16-1:0] node10921;
	wire [16-1:0] node10924;
	wire [16-1:0] node10926;
	wire [16-1:0] node10929;
	wire [16-1:0] node10930;
	wire [16-1:0] node10931;
	wire [16-1:0] node10933;
	wire [16-1:0] node10935;
	wire [16-1:0] node10939;
	wire [16-1:0] node10941;
	wire [16-1:0] node10944;
	wire [16-1:0] node10945;
	wire [16-1:0] node10946;
	wire [16-1:0] node10947;
	wire [16-1:0] node10948;
	wire [16-1:0] node10952;
	wire [16-1:0] node10953;
	wire [16-1:0] node10954;
	wire [16-1:0] node10959;
	wire [16-1:0] node10960;
	wire [16-1:0] node10962;
	wire [16-1:0] node10963;
	wire [16-1:0] node10967;
	wire [16-1:0] node10970;
	wire [16-1:0] node10971;
	wire [16-1:0] node10972;
	wire [16-1:0] node10973;
	wire [16-1:0] node10974;
	wire [16-1:0] node10977;
	wire [16-1:0] node10981;
	wire [16-1:0] node10982;
	wire [16-1:0] node10984;
	wire [16-1:0] node10988;
	wire [16-1:0] node10989;
	wire [16-1:0] node10991;
	wire [16-1:0] node10992;
	wire [16-1:0] node10997;
	wire [16-1:0] node10998;
	wire [16-1:0] node10999;
	wire [16-1:0] node11000;
	wire [16-1:0] node11001;
	wire [16-1:0] node11004;
	wire [16-1:0] node11007;
	wire [16-1:0] node11009;
	wire [16-1:0] node11011;
	wire [16-1:0] node11014;
	wire [16-1:0] node11015;
	wire [16-1:0] node11016;
	wire [16-1:0] node11018;
	wire [16-1:0] node11019;
	wire [16-1:0] node11023;
	wire [16-1:0] node11024;
	wire [16-1:0] node11025;
	wire [16-1:0] node11028;
	wire [16-1:0] node11031;
	wire [16-1:0] node11034;
	wire [16-1:0] node11035;
	wire [16-1:0] node11036;
	wire [16-1:0] node11037;
	wire [16-1:0] node11041;
	wire [16-1:0] node11044;
	wire [16-1:0] node11046;
	wire [16-1:0] node11049;
	wire [16-1:0] node11050;
	wire [16-1:0] node11051;
	wire [16-1:0] node11052;
	wire [16-1:0] node11055;
	wire [16-1:0] node11058;
	wire [16-1:0] node11059;
	wire [16-1:0] node11060;
	wire [16-1:0] node11064;
	wire [16-1:0] node11067;
	wire [16-1:0] node11068;
	wire [16-1:0] node11069;
	wire [16-1:0] node11073;
	wire [16-1:0] node11074;
	wire [16-1:0] node11077;
	wire [16-1:0] node11079;
	wire [16-1:0] node11082;
	wire [16-1:0] node11083;
	wire [16-1:0] node11084;
	wire [16-1:0] node11085;
	wire [16-1:0] node11086;
	wire [16-1:0] node11087;
	wire [16-1:0] node11088;
	wire [16-1:0] node11091;
	wire [16-1:0] node11092;
	wire [16-1:0] node11094;
	wire [16-1:0] node11098;
	wire [16-1:0] node11101;
	wire [16-1:0] node11102;
	wire [16-1:0] node11104;
	wire [16-1:0] node11107;
	wire [16-1:0] node11108;
	wire [16-1:0] node11110;
	wire [16-1:0] node11113;
	wire [16-1:0] node11114;
	wire [16-1:0] node11116;
	wire [16-1:0] node11119;
	wire [16-1:0] node11120;
	wire [16-1:0] node11124;
	wire [16-1:0] node11125;
	wire [16-1:0] node11126;
	wire [16-1:0] node11127;
	wire [16-1:0] node11128;
	wire [16-1:0] node11129;
	wire [16-1:0] node11133;
	wire [16-1:0] node11134;
	wire [16-1:0] node11138;
	wire [16-1:0] node11139;
	wire [16-1:0] node11141;
	wire [16-1:0] node11145;
	wire [16-1:0] node11146;
	wire [16-1:0] node11147;
	wire [16-1:0] node11148;
	wire [16-1:0] node11152;
	wire [16-1:0] node11153;
	wire [16-1:0] node11157;
	wire [16-1:0] node11160;
	wire [16-1:0] node11161;
	wire [16-1:0] node11162;
	wire [16-1:0] node11163;
	wire [16-1:0] node11167;
	wire [16-1:0] node11170;
	wire [16-1:0] node11171;
	wire [16-1:0] node11173;
	wire [16-1:0] node11176;
	wire [16-1:0] node11178;
	wire [16-1:0] node11181;
	wire [16-1:0] node11182;
	wire [16-1:0] node11183;
	wire [16-1:0] node11184;
	wire [16-1:0] node11185;
	wire [16-1:0] node11188;
	wire [16-1:0] node11191;
	wire [16-1:0] node11192;
	wire [16-1:0] node11194;
	wire [16-1:0] node11198;
	wire [16-1:0] node11199;
	wire [16-1:0] node11200;
	wire [16-1:0] node11202;
	wire [16-1:0] node11203;
	wire [16-1:0] node11207;
	wire [16-1:0] node11210;
	wire [16-1:0] node11211;
	wire [16-1:0] node11214;
	wire [16-1:0] node11215;
	wire [16-1:0] node11217;
	wire [16-1:0] node11219;
	wire [16-1:0] node11223;
	wire [16-1:0] node11224;
	wire [16-1:0] node11225;
	wire [16-1:0] node11227;
	wire [16-1:0] node11230;
	wire [16-1:0] node11231;
	wire [16-1:0] node11233;
	wire [16-1:0] node11236;
	wire [16-1:0] node11238;
	wire [16-1:0] node11239;
	wire [16-1:0] node11243;
	wire [16-1:0] node11244;
	wire [16-1:0] node11246;
	wire [16-1:0] node11247;
	wire [16-1:0] node11251;
	wire [16-1:0] node11252;
	wire [16-1:0] node11254;
	wire [16-1:0] node11255;
	wire [16-1:0] node11256;
	wire [16-1:0] node11261;
	wire [16-1:0] node11263;
	wire [16-1:0] node11266;
	wire [16-1:0] node11267;
	wire [16-1:0] node11268;
	wire [16-1:0] node11269;
	wire [16-1:0] node11270;
	wire [16-1:0] node11271;
	wire [16-1:0] node11273;
	wire [16-1:0] node11276;
	wire [16-1:0] node11277;
	wire [16-1:0] node11278;
	wire [16-1:0] node11283;
	wire [16-1:0] node11284;
	wire [16-1:0] node11287;
	wire [16-1:0] node11288;
	wire [16-1:0] node11290;
	wire [16-1:0] node11294;
	wire [16-1:0] node11295;
	wire [16-1:0] node11296;
	wire [16-1:0] node11297;
	wire [16-1:0] node11302;
	wire [16-1:0] node11303;
	wire [16-1:0] node11304;
	wire [16-1:0] node11309;
	wire [16-1:0] node11310;
	wire [16-1:0] node11311;
	wire [16-1:0] node11312;
	wire [16-1:0] node11314;
	wire [16-1:0] node11317;
	wire [16-1:0] node11318;
	wire [16-1:0] node11319;
	wire [16-1:0] node11324;
	wire [16-1:0] node11325;
	wire [16-1:0] node11326;
	wire [16-1:0] node11328;
	wire [16-1:0] node11333;
	wire [16-1:0] node11334;
	wire [16-1:0] node11335;
	wire [16-1:0] node11337;
	wire [16-1:0] node11340;
	wire [16-1:0] node11341;
	wire [16-1:0] node11343;
	wire [16-1:0] node11344;
	wire [16-1:0] node11348;
	wire [16-1:0] node11351;
	wire [16-1:0] node11352;
	wire [16-1:0] node11355;
	wire [16-1:0] node11357;
	wire [16-1:0] node11360;
	wire [16-1:0] node11361;
	wire [16-1:0] node11362;
	wire [16-1:0] node11363;
	wire [16-1:0] node11365;
	wire [16-1:0] node11366;
	wire [16-1:0] node11370;
	wire [16-1:0] node11371;
	wire [16-1:0] node11373;
	wire [16-1:0] node11376;
	wire [16-1:0] node11378;
	wire [16-1:0] node11379;
	wire [16-1:0] node11383;
	wire [16-1:0] node11384;
	wire [16-1:0] node11385;
	wire [16-1:0] node11387;
	wire [16-1:0] node11390;
	wire [16-1:0] node11391;
	wire [16-1:0] node11392;
	wire [16-1:0] node11395;
	wire [16-1:0] node11399;
	wire [16-1:0] node11400;
	wire [16-1:0] node11401;
	wire [16-1:0] node11405;
	wire [16-1:0] node11406;
	wire [16-1:0] node11408;
	wire [16-1:0] node11411;
	wire [16-1:0] node11414;
	wire [16-1:0] node11415;
	wire [16-1:0] node11416;
	wire [16-1:0] node11417;
	wire [16-1:0] node11418;
	wire [16-1:0] node11421;
	wire [16-1:0] node11422;
	wire [16-1:0] node11425;
	wire [16-1:0] node11428;
	wire [16-1:0] node11430;
	wire [16-1:0] node11431;
	wire [16-1:0] node11435;
	wire [16-1:0] node11436;
	wire [16-1:0] node11437;
	wire [16-1:0] node11438;
	wire [16-1:0] node11441;
	wire [16-1:0] node11444;
	wire [16-1:0] node11447;
	wire [16-1:0] node11450;
	wire [16-1:0] node11451;
	wire [16-1:0] node11452;
	wire [16-1:0] node11454;
	wire [16-1:0] node11457;
	wire [16-1:0] node11458;
	wire [16-1:0] node11462;
	wire [16-1:0] node11463;
	wire [16-1:0] node11464;
	wire [16-1:0] node11466;
	wire [16-1:0] node11470;
	wire [16-1:0] node11471;
	wire [16-1:0] node11474;
	wire [16-1:0] node11475;

	assign outp = (inp[6]) ? node5960 : node1;
		assign node1 = (inp[12]) ? node2989 : node2;
			assign node2 = (inp[0]) ? node1482 : node3;
				assign node3 = (inp[3]) ? node705 : node4;
					assign node4 = (inp[7]) ? node348 : node5;
						assign node5 = (inp[5]) ? node189 : node6;
							assign node6 = (inp[13]) ? node98 : node7;
								assign node7 = (inp[14]) ? node49 : node8;
									assign node8 = (inp[8]) ? node30 : node9;
										assign node9 = (inp[11]) ? node21 : node10;
											assign node10 = (inp[9]) ? node12 : 16'b0011111111111111;
												assign node12 = (inp[1]) ? 16'b0000111111111111 : node13;
													assign node13 = (inp[2]) ? 16'b0001111111111111 : node14;
														assign node14 = (inp[10]) ? node16 : 16'b0111111111111111;
															assign node16 = (inp[4]) ? 16'b0001111111111111 : 16'b0011111111111111;
											assign node21 = (inp[15]) ? node23 : 16'b0001111111111111;
												assign node23 = (inp[1]) ? 16'b0000011111111111 : node24;
													assign node24 = (inp[2]) ? 16'b0000111111111111 : node25;
														assign node25 = (inp[9]) ? 16'b0000111111111111 : 16'b0001111111111111;
										assign node30 = (inp[10]) ? node44 : node31;
											assign node31 = (inp[15]) ? node37 : node32;
												assign node32 = (inp[4]) ? 16'b0000111111111111 : node33;
													assign node33 = (inp[11]) ? 16'b0001111111111111 : 16'b0011111111111111;
												assign node37 = (inp[11]) ? node39 : 16'b0000011111111111;
													assign node39 = (inp[9]) ? node41 : 16'b0000111111111111;
														assign node41 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node44 = (inp[11]) ? node46 : 16'b0000111111111111;
												assign node46 = (inp[1]) ? 16'b0000001111111111 : 16'b0000000111111111;
									assign node49 = (inp[1]) ? node83 : node50;
										assign node50 = (inp[4]) ? node70 : node51;
											assign node51 = (inp[15]) ? node59 : node52;
												assign node52 = (inp[8]) ? 16'b0000111111111111 : node53;
													assign node53 = (inp[2]) ? 16'b0001111111111111 : node54;
														assign node54 = (inp[9]) ? 16'b0001111111111111 : 16'b0011111111111111;
												assign node59 = (inp[9]) ? node65 : node60;
													assign node60 = (inp[10]) ? 16'b0000111111111111 : node61;
														assign node61 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node65 = (inp[2]) ? 16'b0000011111111111 : node66;
														assign node66 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node70 = (inp[9]) ? node78 : node71;
												assign node71 = (inp[10]) ? 16'b0000011111111111 : node72;
													assign node72 = (inp[8]) ? node74 : 16'b0000111111111111;
														assign node74 = (inp[2]) ? 16'b0000111111111111 : 16'b0000011111111111;
												assign node78 = (inp[2]) ? 16'b0000011111111111 : node79;
													assign node79 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node83 = (inp[10]) ? node93 : node84;
											assign node84 = (inp[2]) ? 16'b0000011111111111 : node85;
												assign node85 = (inp[8]) ? node87 : 16'b0000111111111111;
													assign node87 = (inp[11]) ? 16'b0000011111111111 : node88;
														assign node88 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node93 = (inp[2]) ? node95 : 16'b0000001111111111;
												assign node95 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
								assign node98 = (inp[15]) ? node148 : node99;
									assign node99 = (inp[8]) ? node119 : node100;
										assign node100 = (inp[4]) ? node110 : node101;
											assign node101 = (inp[2]) ? 16'b0000111111111111 : node102;
												assign node102 = (inp[1]) ? node104 : 16'b0001111111111111;
													assign node104 = (inp[10]) ? 16'b0000111111111111 : node105;
														assign node105 = (inp[14]) ? 16'b0000111111111111 : 16'b0011111111111111;
											assign node110 = (inp[1]) ? node114 : node111;
												assign node111 = (inp[2]) ? 16'b0000011111111111 : 16'b0001111111111111;
												assign node114 = (inp[11]) ? node116 : 16'b0000011111111111;
													assign node116 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node119 = (inp[2]) ? node133 : node120;
											assign node120 = (inp[9]) ? node124 : node121;
												assign node121 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node124 = (inp[11]) ? node128 : node125;
													assign node125 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node128 = (inp[4]) ? 16'b0000001111111111 : node129;
														assign node129 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node133 = (inp[11]) ? node139 : node134;
												assign node134 = (inp[14]) ? 16'b0000001111111111 : node135;
													assign node135 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node139 = (inp[4]) ? node145 : node140;
													assign node140 = (inp[1]) ? 16'b0000001111111111 : node141;
														assign node141 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node145 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node148 = (inp[11]) ? node168 : node149;
										assign node149 = (inp[4]) ? node159 : node150;
											assign node150 = (inp[14]) ? node154 : node151;
												assign node151 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node154 = (inp[1]) ? node156 : 16'b0000011111111111;
													assign node156 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node159 = (inp[1]) ? node163 : node160;
												assign node160 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node163 = (inp[2]) ? node165 : 16'b0000001111111111;
													assign node165 = (inp[9]) ? 16'b0000001111111111 : 16'b0000000011111111;
										assign node168 = (inp[9]) ? node180 : node169;
											assign node169 = (inp[14]) ? node175 : node170;
												assign node170 = (inp[4]) ? 16'b0000001111111111 : node171;
													assign node171 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node175 = (inp[8]) ? 16'b0000001111111111 : node176;
													assign node176 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node180 = (inp[1]) ? node186 : node181;
												assign node181 = (inp[2]) ? 16'b0000000111111111 : node182;
													assign node182 = (inp[8]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node186 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node189 = (inp[13]) ? node265 : node190;
								assign node190 = (inp[14]) ? node230 : node191;
									assign node191 = (inp[2]) ? node209 : node192;
										assign node192 = (inp[11]) ? node198 : node193;
											assign node193 = (inp[1]) ? node195 : 16'b0001111111111111;
												assign node195 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node198 = (inp[4]) ? node206 : node199;
												assign node199 = (inp[9]) ? node201 : 16'b0000111111111111;
													assign node201 = (inp[1]) ? 16'b0000011111111111 : node202;
														assign node202 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node206 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node209 = (inp[10]) ? node221 : node210;
											assign node210 = (inp[4]) ? node214 : node211;
												assign node211 = (inp[1]) ? 16'b0000111111111111 : 16'b0000011111111111;
												assign node214 = (inp[15]) ? 16'b0000001111111111 : node215;
													assign node215 = (inp[9]) ? node217 : 16'b0000011111111111;
														assign node217 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node221 = (inp[11]) ? node227 : node222;
												assign node222 = (inp[4]) ? node224 : 16'b0000001111111111;
													assign node224 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node227 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node230 = (inp[15]) ? node250 : node231;
										assign node231 = (inp[4]) ? node241 : node232;
											assign node232 = (inp[11]) ? 16'b0000001111111111 : node233;
												assign node233 = (inp[10]) ? node235 : 16'b0000111111111111;
													assign node235 = (inp[9]) ? node237 : 16'b0000011111111111;
														assign node237 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node241 = (inp[1]) ? node247 : node242;
												assign node242 = (inp[11]) ? node244 : 16'b0000001111111111;
													assign node244 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node247 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node250 = (inp[10]) ? node258 : node251;
											assign node251 = (inp[9]) ? node255 : node252;
												assign node252 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node255 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node258 = (inp[4]) ? node262 : node259;
												assign node259 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node262 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node265 = (inp[9]) ? node309 : node266;
									assign node266 = (inp[4]) ? node286 : node267;
										assign node267 = (inp[11]) ? node273 : node268;
											assign node268 = (inp[15]) ? 16'b0000011111111111 : node269;
												assign node269 = (inp[1]) ? 16'b0001111111111111 : 16'b0000111111111111;
											assign node273 = (inp[10]) ? node281 : node274;
												assign node274 = (inp[14]) ? 16'b0000001111111111 : node275;
													assign node275 = (inp[2]) ? 16'b0000001111111111 : node276;
														assign node276 = (inp[15]) ? 16'b0000111111111111 : 16'b0000011111111111;
												assign node281 = (inp[1]) ? node283 : 16'b0000001111111111;
													assign node283 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node286 = (inp[2]) ? node300 : node287;
											assign node287 = (inp[15]) ? node295 : node288;
												assign node288 = (inp[8]) ? 16'b0000000111111111 : node289;
													assign node289 = (inp[14]) ? 16'b0000011111111111 : node290;
														assign node290 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node295 = (inp[1]) ? node297 : 16'b0000001111111111;
													assign node297 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node300 = (inp[11]) ? node306 : node301;
												assign node301 = (inp[15]) ? node303 : 16'b0000001111111111;
													assign node303 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node306 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
									assign node309 = (inp[10]) ? node329 : node310;
										assign node310 = (inp[2]) ? node318 : node311;
											assign node311 = (inp[8]) ? node315 : node312;
												assign node312 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node315 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node318 = (inp[1]) ? node326 : node319;
												assign node319 = (inp[11]) ? node321 : 16'b0000001111111111;
													assign node321 = (inp[14]) ? node323 : 16'b0000000111111111;
														assign node323 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node326 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node329 = (inp[4]) ? node339 : node330;
											assign node330 = (inp[11]) ? node332 : 16'b0000000111111111;
												assign node332 = (inp[2]) ? node334 : 16'b0000000001111111;
													assign node334 = (inp[15]) ? 16'b0000000011111111 : node335;
														assign node335 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node339 = (inp[11]) ? 16'b0000000000111111 : node340;
												assign node340 = (inp[8]) ? node342 : 16'b0000000011111111;
													assign node342 = (inp[14]) ? 16'b0000000001111111 : node343;
														assign node343 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
						assign node348 = (inp[14]) ? node534 : node349;
							assign node349 = (inp[5]) ? node439 : node350;
								assign node350 = (inp[8]) ? node390 : node351;
									assign node351 = (inp[4]) ? node363 : node352;
										assign node352 = (inp[15]) ? node358 : node353;
											assign node353 = (inp[11]) ? 16'b0000111111111111 : node354;
												assign node354 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
											assign node358 = (inp[9]) ? 16'b0000001111111111 : node359;
												assign node359 = (inp[10]) ? 16'b0000011111111111 : 16'b0001111111111111;
										assign node363 = (inp[13]) ? node373 : node364;
											assign node364 = (inp[15]) ? node368 : node365;
												assign node365 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node368 = (inp[9]) ? 16'b0000011111111111 : node369;
													assign node369 = (inp[1]) ? 16'b0000011111111111 : 16'b0001111111111111;
											assign node373 = (inp[9]) ? node385 : node374;
												assign node374 = (inp[1]) ? node378 : node375;
													assign node375 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node378 = (inp[2]) ? 16'b0000001111111111 : node379;
														assign node379 = (inp[10]) ? node381 : 16'b0000011111111111;
															assign node381 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node385 = (inp[10]) ? node387 : 16'b0000001111111111;
													assign node387 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node390 = (inp[1]) ? node416 : node391;
										assign node391 = (inp[15]) ? node405 : node392;
											assign node392 = (inp[4]) ? node396 : node393;
												assign node393 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node396 = (inp[11]) ? node398 : 16'b0000011111111111;
													assign node398 = (inp[2]) ? node400 : 16'b0000011111111111;
														assign node400 = (inp[9]) ? 16'b0000001111111111 : node401;
															assign node401 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node405 = (inp[4]) ? node413 : node406;
												assign node406 = (inp[9]) ? 16'b0000001111111111 : node407;
													assign node407 = (inp[13]) ? node409 : 16'b0000011111111111;
														assign node409 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node413 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node416 = (inp[2]) ? node430 : node417;
											assign node417 = (inp[10]) ? node423 : node418;
												assign node418 = (inp[13]) ? node420 : 16'b0000011111111111;
													assign node420 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node423 = (inp[13]) ? 16'b0000000011111111 : node424;
													assign node424 = (inp[15]) ? node426 : 16'b0000001111111111;
														assign node426 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node430 = (inp[11]) ? node432 : 16'b0000000111111111;
												assign node432 = (inp[15]) ? node434 : 16'b0000000111111111;
													assign node434 = (inp[9]) ? 16'b0000000011111111 : node435;
														assign node435 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node439 = (inp[13]) ? node481 : node440;
									assign node440 = (inp[15]) ? node464 : node441;
										assign node441 = (inp[10]) ? node451 : node442;
											assign node442 = (inp[2]) ? node446 : node443;
												assign node443 = (inp[1]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node446 = (inp[9]) ? 16'b0000000011111111 : node447;
													assign node447 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node451 = (inp[4]) ? 16'b0000001111111111 : node452;
												assign node452 = (inp[11]) ? node458 : node453;
													assign node453 = (inp[2]) ? node455 : 16'b0000011111111111;
														assign node455 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node458 = (inp[2]) ? 16'b0000001111111111 : node459;
														assign node459 = (inp[8]) ? 16'b0000001111111111 : 16'b0000111111111111;
										assign node464 = (inp[10]) ? node470 : node465;
											assign node465 = (inp[9]) ? 16'b0000000111111111 : node466;
												assign node466 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node470 = (inp[11]) ? node474 : node471;
												assign node471 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node474 = (inp[1]) ? 16'b0000000011111111 : node475;
													assign node475 = (inp[9]) ? node477 : 16'b0000000111111111;
														assign node477 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node481 = (inp[2]) ? node513 : node482;
										assign node482 = (inp[1]) ? node500 : node483;
											assign node483 = (inp[4]) ? node487 : node484;
												assign node484 = (inp[11]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node487 = (inp[11]) ? node495 : node488;
													assign node488 = (inp[9]) ? node492 : node489;
														assign node489 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node492 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node495 = (inp[15]) ? 16'b0000000111111111 : node496;
														assign node496 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node500 = (inp[8]) ? node508 : node501;
												assign node501 = (inp[10]) ? node505 : node502;
													assign node502 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node505 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node508 = (inp[10]) ? 16'b0000000000111111 : node509;
													assign node509 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node513 = (inp[11]) ? node525 : node514;
											assign node514 = (inp[8]) ? node518 : node515;
												assign node515 = (inp[15]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node518 = (inp[4]) ? node520 : 16'b0000000011111111;
													assign node520 = (inp[9]) ? 16'b0000000011111111 : node521;
														assign node521 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node525 = (inp[1]) ? node527 : 16'b0000000111111111;
												assign node527 = (inp[8]) ? node529 : 16'b0000000000111111;
													assign node529 = (inp[15]) ? node531 : 16'b0000000001111111;
														assign node531 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node534 = (inp[10]) ? node626 : node535;
								assign node535 = (inp[8]) ? node573 : node536;
									assign node536 = (inp[13]) ? node556 : node537;
										assign node537 = (inp[15]) ? node549 : node538;
											assign node538 = (inp[4]) ? node544 : node539;
												assign node539 = (inp[9]) ? 16'b0000011111111111 : node540;
													assign node540 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node544 = (inp[5]) ? node546 : 16'b0000011111111111;
													assign node546 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node549 = (inp[2]) ? 16'b0000000111111111 : node550;
												assign node550 = (inp[4]) ? node552 : 16'b0000011111111111;
													assign node552 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node556 = (inp[15]) ? node566 : node557;
											assign node557 = (inp[5]) ? node559 : 16'b0000111111111111;
												assign node559 = (inp[1]) ? 16'b0000000111111111 : node560;
													assign node560 = (inp[4]) ? 16'b0000001111111111 : node561;
														assign node561 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node566 = (inp[1]) ? 16'b0000000011111111 : node567;
												assign node567 = (inp[9]) ? 16'b0000000111111111 : node568;
													assign node568 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node573 = (inp[9]) ? node599 : node574;
										assign node574 = (inp[4]) ? node588 : node575;
											assign node575 = (inp[15]) ? node583 : node576;
												assign node576 = (inp[1]) ? node578 : 16'b0000011111111111;
													assign node578 = (inp[13]) ? 16'b0000001111111111 : node579;
														assign node579 = (inp[11]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node583 = (inp[13]) ? node585 : 16'b0000001111111111;
													assign node585 = (inp[2]) ? 16'b0000000111111111 : 16'b0000011111111111;
											assign node588 = (inp[2]) ? node594 : node589;
												assign node589 = (inp[15]) ? 16'b0000000111111111 : node590;
													assign node590 = (inp[13]) ? 16'b0000011111111111 : 16'b0000001111111111;
												assign node594 = (inp[5]) ? node596 : 16'b0000000111111111;
													assign node596 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node599 = (inp[13]) ? node615 : node600;
											assign node600 = (inp[2]) ? node610 : node601;
												assign node601 = (inp[15]) ? node605 : node602;
													assign node602 = (inp[1]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node605 = (inp[1]) ? 16'b0000000111111111 : node606;
														assign node606 = (inp[11]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node610 = (inp[11]) ? node612 : 16'b0000000111111111;
													assign node612 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node615 = (inp[15]) ? node621 : node616;
												assign node616 = (inp[1]) ? 16'b0000000011111111 : node617;
													assign node617 = (inp[4]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node621 = (inp[5]) ? node623 : 16'b0000000011111111;
													assign node623 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000001111111;
								assign node626 = (inp[11]) ? node668 : node627;
									assign node627 = (inp[8]) ? node647 : node628;
										assign node628 = (inp[4]) ? node636 : node629;
											assign node629 = (inp[1]) ? 16'b0000001111111111 : node630;
												assign node630 = (inp[13]) ? node632 : 16'b0001111111111111;
													assign node632 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node636 = (inp[15]) ? node644 : node637;
												assign node637 = (inp[2]) ? 16'b0000000111111111 : node638;
													assign node638 = (inp[13]) ? 16'b0000001111111111 : node639;
														assign node639 = (inp[1]) ? 16'b0000011111111111 : 16'b0000001111111111;
												assign node644 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node647 = (inp[1]) ? node655 : node648;
											assign node648 = (inp[4]) ? node650 : 16'b0000001111111111;
												assign node650 = (inp[15]) ? node652 : 16'b0000000111111111;
													assign node652 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node655 = (inp[5]) ? node661 : node656;
												assign node656 = (inp[4]) ? 16'b0000000001111111 : node657;
													assign node657 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node661 = (inp[15]) ? node663 : 16'b0000000011111111;
													assign node663 = (inp[9]) ? 16'b0000000001111111 : node664;
														assign node664 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node668 = (inp[2]) ? node686 : node669;
										assign node669 = (inp[4]) ? node675 : node670;
											assign node670 = (inp[8]) ? node672 : 16'b0000000111111111;
												assign node672 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node675 = (inp[5]) ? 16'b0000000001111111 : node676;
												assign node676 = (inp[9]) ? node678 : 16'b0000000111111111;
													assign node678 = (inp[1]) ? node682 : node679;
														assign node679 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node682 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node686 = (inp[9]) ? node692 : node687;
											assign node687 = (inp[15]) ? 16'b0000000011111111 : node688;
												assign node688 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node692 = (inp[5]) ? node696 : node693;
												assign node693 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node696 = (inp[1]) ? node702 : node697;
													assign node697 = (inp[8]) ? node699 : 16'b0000000111111111;
														assign node699 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node702 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
					assign node705 = (inp[8]) ? node1075 : node706;
						assign node706 = (inp[2]) ? node886 : node707;
							assign node707 = (inp[13]) ? node799 : node708;
								assign node708 = (inp[14]) ? node756 : node709;
									assign node709 = (inp[7]) ? node729 : node710;
										assign node710 = (inp[1]) ? node724 : node711;
											assign node711 = (inp[10]) ? node717 : node712;
												assign node712 = (inp[15]) ? node714 : 16'b0001111111111111;
													assign node714 = (inp[11]) ? 16'b0000011111111111 : 16'b0001111111111111;
												assign node717 = (inp[5]) ? 16'b0000011111111111 : node718;
													assign node718 = (inp[9]) ? node720 : 16'b0000111111111111;
														assign node720 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
											assign node724 = (inp[5]) ? 16'b0000000111111111 : node725;
												assign node725 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node729 = (inp[10]) ? node739 : node730;
											assign node730 = (inp[15]) ? node734 : node731;
												assign node731 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node734 = (inp[4]) ? node736 : 16'b0000111111111111;
													assign node736 = (inp[1]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node739 = (inp[11]) ? node751 : node740;
												assign node740 = (inp[1]) ? node746 : node741;
													assign node741 = (inp[9]) ? node743 : 16'b0000111111111111;
														assign node743 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node746 = (inp[9]) ? node748 : 16'b0000011111111111;
														assign node748 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node751 = (inp[4]) ? node753 : 16'b0000011111111111;
													assign node753 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node756 = (inp[9]) ? node778 : node757;
										assign node757 = (inp[1]) ? node765 : node758;
											assign node758 = (inp[11]) ? 16'b0000011111111111 : node759;
												assign node759 = (inp[15]) ? node761 : 16'b0000011111111111;
													assign node761 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node765 = (inp[11]) ? node771 : node766;
												assign node766 = (inp[7]) ? node768 : 16'b0000111111111111;
													assign node768 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node771 = (inp[4]) ? node773 : 16'b0000001111111111;
													assign node773 = (inp[15]) ? 16'b0000000011111111 : node774;
														assign node774 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node778 = (inp[10]) ? node788 : node779;
											assign node779 = (inp[7]) ? node785 : node780;
												assign node780 = (inp[11]) ? node782 : 16'b0000011111111111;
													assign node782 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node785 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node788 = (inp[15]) ? node792 : node789;
												assign node789 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node792 = (inp[1]) ? node794 : 16'b0000000001111111;
													assign node794 = (inp[4]) ? 16'b0000000011111111 : node795;
														assign node795 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node799 = (inp[10]) ? node849 : node800;
									assign node800 = (inp[4]) ? node826 : node801;
										assign node801 = (inp[15]) ? node815 : node802;
											assign node802 = (inp[1]) ? node812 : node803;
												assign node803 = (inp[5]) ? node809 : node804;
													assign node804 = (inp[14]) ? node806 : 16'b0000111111111111;
														assign node806 = (inp[9]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node809 = (inp[14]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node812 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node815 = (inp[14]) ? node823 : node816;
												assign node816 = (inp[5]) ? node818 : 16'b0000011111111111;
													assign node818 = (inp[7]) ? node820 : 16'b0000001111111111;
														assign node820 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node823 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node826 = (inp[5]) ? node834 : node827;
											assign node827 = (inp[14]) ? 16'b0000000111111111 : node828;
												assign node828 = (inp[7]) ? node830 : 16'b0000011111111111;
													assign node830 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node834 = (inp[15]) ? node840 : node835;
												assign node835 = (inp[9]) ? node837 : 16'b0000001111111111;
													assign node837 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node840 = (inp[7]) ? node846 : node841;
													assign node841 = (inp[11]) ? 16'b0000000111111111 : node842;
														assign node842 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node846 = (inp[9]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node849 = (inp[15]) ? node877 : node850;
										assign node850 = (inp[11]) ? node870 : node851;
											assign node851 = (inp[5]) ? node859 : node852;
												assign node852 = (inp[1]) ? 16'b0000001111111111 : node853;
													assign node853 = (inp[9]) ? node855 : 16'b0000011111111111;
														assign node855 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node859 = (inp[14]) ? node865 : node860;
													assign node860 = (inp[9]) ? 16'b0000011111111111 : node861;
														assign node861 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node865 = (inp[9]) ? 16'b0000000111111111 : node866;
														assign node866 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node870 = (inp[4]) ? node874 : node871;
												assign node871 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node874 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node877 = (inp[5]) ? node879 : 16'b0000000111111111;
											assign node879 = (inp[7]) ? 16'b0000000011111111 : node880;
												assign node880 = (inp[14]) ? node882 : 16'b0000000111111111;
													assign node882 = (inp[9]) ? 16'b0000000111111111 : 16'b0000000011111111;
							assign node886 = (inp[1]) ? node978 : node887;
								assign node887 = (inp[11]) ? node927 : node888;
									assign node888 = (inp[15]) ? node908 : node889;
										assign node889 = (inp[13]) ? node903 : node890;
											assign node890 = (inp[5]) ? node900 : node891;
												assign node891 = (inp[7]) ? node893 : 16'b0000111111111111;
													assign node893 = (inp[14]) ? 16'b0000001111111111 : node894;
														assign node894 = (inp[10]) ? node896 : 16'b0000111111111111;
															assign node896 = (inp[9]) ? 16'b0000011111111111 : 16'b0000011111111111;
												assign node900 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node903 = (inp[4]) ? 16'b0000001111111111 : node904;
												assign node904 = (inp[9]) ? 16'b0000011111111111 : 16'b0000001111111111;
										assign node908 = (inp[10]) ? node920 : node909;
											assign node909 = (inp[7]) ? node915 : node910;
												assign node910 = (inp[9]) ? 16'b0000011111111111 : node911;
													assign node911 = (inp[13]) ? 16'b0000011111111111 : 16'b0001111111111111;
												assign node915 = (inp[14]) ? 16'b0000000111111111 : node916;
													assign node916 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node920 = (inp[13]) ? node922 : 16'b0000000111111111;
												assign node922 = (inp[7]) ? 16'b0000000111111111 : node923;
													assign node923 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node927 = (inp[9]) ? node951 : node928;
										assign node928 = (inp[10]) ? node938 : node929;
											assign node929 = (inp[13]) ? node931 : 16'b0000001111111111;
												assign node931 = (inp[5]) ? node933 : 16'b0000001111111111;
													assign node933 = (inp[4]) ? 16'b0000000111111111 : node934;
														assign node934 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node938 = (inp[15]) ? node946 : node939;
												assign node939 = (inp[5]) ? 16'b0000000111111111 : node940;
													assign node940 = (inp[14]) ? 16'b0000001111111111 : node941;
														assign node941 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node946 = (inp[14]) ? node948 : 16'b0000000111111111;
													assign node948 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node951 = (inp[14]) ? node967 : node952;
											assign node952 = (inp[7]) ? node960 : node953;
												assign node953 = (inp[5]) ? node955 : 16'b0000011111111111;
													assign node955 = (inp[4]) ? 16'b0000001111111111 : node956;
														assign node956 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node960 = (inp[15]) ? node964 : node961;
													assign node961 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node964 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node967 = (inp[4]) ? node971 : node968;
												assign node968 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node971 = (inp[7]) ? node975 : node972;
													assign node972 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node975 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
								assign node978 = (inp[11]) ? node1016 : node979;
									assign node979 = (inp[7]) ? node997 : node980;
										assign node980 = (inp[9]) ? node990 : node981;
											assign node981 = (inp[13]) ? node985 : node982;
												assign node982 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node985 = (inp[10]) ? node987 : 16'b0000001111111111;
													assign node987 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node990 = (inp[5]) ? node994 : node991;
												assign node991 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node994 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node997 = (inp[5]) ? node1003 : node998;
											assign node998 = (inp[9]) ? 16'b0000000011111111 : node999;
												assign node999 = (inp[13]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node1003 = (inp[4]) ? node1009 : node1004;
												assign node1004 = (inp[13]) ? node1006 : 16'b0000000111111111;
													assign node1006 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1009 = (inp[13]) ? node1013 : node1010;
													assign node1010 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node1013 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000000111111;
									assign node1016 = (inp[15]) ? node1042 : node1017;
										assign node1017 = (inp[9]) ? node1025 : node1018;
											assign node1018 = (inp[4]) ? 16'b0000000111111111 : node1019;
												assign node1019 = (inp[14]) ? 16'b0000000111111111 : node1020;
													assign node1020 = (inp[7]) ? 16'b0000000111111111 : 16'b0000011111111111;
											assign node1025 = (inp[4]) ? node1033 : node1026;
												assign node1026 = (inp[14]) ? 16'b0000000011111111 : node1027;
													assign node1027 = (inp[5]) ? node1029 : 16'b0000000111111111;
														assign node1029 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1033 = (inp[5]) ? 16'b0000000000111111 : node1034;
													assign node1034 = (inp[13]) ? 16'b0000000001111111 : node1035;
														assign node1035 = (inp[7]) ? node1037 : 16'b0000000011111111;
															assign node1037 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1042 = (inp[10]) ? node1052 : node1043;
											assign node1043 = (inp[7]) ? node1047 : node1044;
												assign node1044 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1047 = (inp[5]) ? 16'b0000000000111111 : node1048;
													assign node1048 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1052 = (inp[13]) ? node1060 : node1053;
												assign node1053 = (inp[7]) ? 16'b0000000001111111 : node1054;
													assign node1054 = (inp[4]) ? node1056 : 16'b0000000011111111;
														assign node1056 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1060 = (inp[14]) ? node1068 : node1061;
													assign node1061 = (inp[4]) ? node1065 : node1062;
														assign node1062 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node1065 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node1068 = (inp[9]) ? node1072 : node1069;
														assign node1069 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node1072 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node1075 = (inp[9]) ? node1289 : node1076;
							assign node1076 = (inp[1]) ? node1162 : node1077;
								assign node1077 = (inp[15]) ? node1127 : node1078;
									assign node1078 = (inp[11]) ? node1106 : node1079;
										assign node1079 = (inp[14]) ? node1097 : node1080;
											assign node1080 = (inp[13]) ? node1088 : node1081;
												assign node1081 = (inp[2]) ? node1085 : node1082;
													assign node1082 = (inp[5]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node1085 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1088 = (inp[10]) ? node1094 : node1089;
													assign node1089 = (inp[2]) ? 16'b0000011111111111 : node1090;
														assign node1090 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1094 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1097 = (inp[5]) ? node1101 : node1098;
												assign node1098 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1101 = (inp[4]) ? node1103 : 16'b0000001111111111;
													assign node1103 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1106 = (inp[7]) ? node1120 : node1107;
											assign node1107 = (inp[13]) ? node1115 : node1108;
												assign node1108 = (inp[14]) ? 16'b0000001111111111 : node1109;
													assign node1109 = (inp[10]) ? 16'b0000001111111111 : node1110;
														assign node1110 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1115 = (inp[5]) ? node1117 : 16'b0000001111111111;
													assign node1117 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1120 = (inp[2]) ? node1124 : node1121;
												assign node1121 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1124 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1127 = (inp[7]) ? node1149 : node1128;
										assign node1128 = (inp[11]) ? node1144 : node1129;
											assign node1129 = (inp[4]) ? node1139 : node1130;
												assign node1130 = (inp[10]) ? node1132 : 16'b0000011111111111;
													assign node1132 = (inp[5]) ? node1136 : node1133;
														assign node1133 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1136 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1139 = (inp[10]) ? 16'b0000000111111111 : node1140;
													assign node1140 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1144 = (inp[10]) ? node1146 : 16'b0000000111111111;
												assign node1146 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node1149 = (inp[13]) ? node1155 : node1150;
											assign node1150 = (inp[10]) ? node1152 : 16'b0000000011111111;
												assign node1152 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1155 = (inp[14]) ? node1157 : 16'b0000000111111111;
												assign node1157 = (inp[11]) ? 16'b0000000001111111 : node1158;
													assign node1158 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1162 = (inp[14]) ? node1230 : node1163;
									assign node1163 = (inp[10]) ? node1195 : node1164;
										assign node1164 = (inp[4]) ? node1180 : node1165;
											assign node1165 = (inp[15]) ? node1173 : node1166;
												assign node1166 = (inp[7]) ? 16'b0000011111111111 : node1167;
													assign node1167 = (inp[2]) ? 16'b0000011111111111 : node1168;
														assign node1168 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1173 = (inp[13]) ? node1177 : node1174;
													assign node1174 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1177 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1180 = (inp[5]) ? node1192 : node1181;
												assign node1181 = (inp[11]) ? node1185 : node1182;
													assign node1182 = (inp[15]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node1185 = (inp[13]) ? 16'b0000000111111111 : node1186;
														assign node1186 = (inp[7]) ? 16'b0000000111111111 : node1187;
															assign node1187 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1192 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1195 = (inp[13]) ? node1207 : node1196;
											assign node1196 = (inp[5]) ? node1204 : node1197;
												assign node1197 = (inp[2]) ? 16'b0000000111111111 : node1198;
													assign node1198 = (inp[7]) ? node1200 : 16'b0000001111111111;
														assign node1200 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1204 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1207 = (inp[11]) ? node1217 : node1208;
												assign node1208 = (inp[2]) ? node1210 : 16'b0000000111111111;
													assign node1210 = (inp[15]) ? node1212 : 16'b0000000111111111;
														assign node1212 = (inp[4]) ? 16'b0000000011111111 : node1213;
															assign node1213 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1217 = (inp[5]) ? node1223 : node1218;
													assign node1218 = (inp[2]) ? 16'b0000000011111111 : node1219;
														assign node1219 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node1223 = (inp[2]) ? node1225 : 16'b0000000001111111;
														assign node1225 = (inp[7]) ? node1227 : 16'b0000000000111111;
															assign node1227 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node1230 = (inp[7]) ? node1262 : node1231;
										assign node1231 = (inp[10]) ? node1247 : node1232;
											assign node1232 = (inp[4]) ? node1240 : node1233;
												assign node1233 = (inp[5]) ? 16'b0000000111111111 : node1234;
													assign node1234 = (inp[15]) ? 16'b0000001111111111 : node1235;
														assign node1235 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1240 = (inp[13]) ? node1244 : node1241;
													assign node1241 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1244 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1247 = (inp[11]) ? node1255 : node1248;
												assign node1248 = (inp[13]) ? node1250 : 16'b0000000111111111;
													assign node1250 = (inp[5]) ? node1252 : 16'b0000000011111111;
														assign node1252 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1255 = (inp[5]) ? 16'b0000000000111111 : node1256;
													assign node1256 = (inp[2]) ? 16'b0000000001111111 : node1257;
														assign node1257 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1262 = (inp[15]) ? node1274 : node1263;
											assign node1263 = (inp[5]) ? node1271 : node1264;
												assign node1264 = (inp[13]) ? node1266 : 16'b0000000011111111;
													assign node1266 = (inp[4]) ? node1268 : 16'b0000000011111111;
														assign node1268 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1271 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1274 = (inp[5]) ? node1280 : node1275;
												assign node1275 = (inp[11]) ? 16'b0000000001111111 : node1276;
													assign node1276 = (inp[10]) ? 16'b0000000001111111 : 16'b0000001111111111;
												assign node1280 = (inp[2]) ? node1286 : node1281;
													assign node1281 = (inp[13]) ? node1283 : 16'b0000000001111111;
														assign node1283 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node1286 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node1289 = (inp[7]) ? node1395 : node1290;
								assign node1290 = (inp[10]) ? node1334 : node1291;
									assign node1291 = (inp[5]) ? node1317 : node1292;
										assign node1292 = (inp[13]) ? node1306 : node1293;
											assign node1293 = (inp[14]) ? node1301 : node1294;
												assign node1294 = (inp[2]) ? node1296 : 16'b0000011111111111;
													assign node1296 = (inp[4]) ? 16'b0000001111111111 : node1297;
														assign node1297 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1301 = (inp[11]) ? node1303 : 16'b0000001111111111;
													assign node1303 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1306 = (inp[4]) ? node1310 : node1307;
												assign node1307 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1310 = (inp[2]) ? node1312 : 16'b0000000111111111;
													assign node1312 = (inp[15]) ? 16'b0000000011111111 : node1313;
														assign node1313 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1317 = (inp[2]) ? node1327 : node1318;
											assign node1318 = (inp[11]) ? node1322 : node1319;
												assign node1319 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1322 = (inp[13]) ? node1324 : 16'b0000000111111111;
													assign node1324 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1327 = (inp[1]) ? node1331 : node1328;
												assign node1328 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1331 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1334 = (inp[4]) ? node1350 : node1335;
										assign node1335 = (inp[11]) ? node1347 : node1336;
											assign node1336 = (inp[13]) ? node1342 : node1337;
												assign node1337 = (inp[2]) ? node1339 : 16'b0000011111111111;
													assign node1339 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1342 = (inp[2]) ? 16'b0000000111111111 : node1343;
													assign node1343 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1347 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node1350 = (inp[13]) ? node1368 : node1351;
											assign node1351 = (inp[1]) ? node1361 : node1352;
												assign node1352 = (inp[5]) ? node1356 : node1353;
													assign node1353 = (inp[14]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node1356 = (inp[2]) ? 16'b0000000011111111 : node1357;
														assign node1357 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1361 = (inp[5]) ? node1363 : 16'b0000000011111111;
													assign node1363 = (inp[2]) ? node1365 : 16'b0000000001111111;
														assign node1365 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node1368 = (inp[2]) ? node1382 : node1369;
												assign node1369 = (inp[5]) ? node1377 : node1370;
													assign node1370 = (inp[15]) ? 16'b0000000001111111 : node1371;
														assign node1371 = (inp[1]) ? 16'b0000000011111111 : node1372;
															assign node1372 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node1377 = (inp[1]) ? 16'b0000000000111111 : node1378;
														assign node1378 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1382 = (inp[5]) ? node1390 : node1383;
													assign node1383 = (inp[15]) ? node1385 : 16'b0000000001111111;
														assign node1385 = (inp[1]) ? 16'b0000000000111111 : node1386;
															assign node1386 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node1390 = (inp[11]) ? 16'b0000000000011111 : node1391;
														assign node1391 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000001111111;
								assign node1395 = (inp[14]) ? node1451 : node1396;
									assign node1396 = (inp[1]) ? node1428 : node1397;
										assign node1397 = (inp[5]) ? node1417 : node1398;
											assign node1398 = (inp[13]) ? node1406 : node1399;
												assign node1399 = (inp[15]) ? node1401 : 16'b0000011111111111;
													assign node1401 = (inp[2]) ? 16'b0000000111111111 : node1402;
														assign node1402 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1406 = (inp[11]) ? node1410 : node1407;
													assign node1407 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1410 = (inp[2]) ? node1412 : 16'b0000000011111111;
														assign node1412 = (inp[15]) ? 16'b0000000001111111 : node1413;
															assign node1413 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1417 = (inp[11]) ? node1419 : 16'b0000000011111111;
												assign node1419 = (inp[2]) ? 16'b0000000001111111 : node1420;
													assign node1420 = (inp[10]) ? node1422 : 16'b0000000111111111;
														assign node1422 = (inp[13]) ? node1424 : 16'b0000000011111111;
															assign node1424 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1428 = (inp[2]) ? node1438 : node1429;
											assign node1429 = (inp[15]) ? node1431 : 16'b0000000011111111;
												assign node1431 = (inp[4]) ? 16'b0000000000111111 : node1432;
													assign node1432 = (inp[10]) ? node1434 : 16'b0000000011111111;
														assign node1434 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1438 = (inp[11]) ? node1444 : node1439;
												assign node1439 = (inp[15]) ? node1441 : 16'b0000000001111111;
													assign node1441 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node1444 = (inp[13]) ? 16'b0000000000001111 : node1445;
													assign node1445 = (inp[15]) ? node1447 : 16'b0000000000111111;
														assign node1447 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node1451 = (inp[15]) ? node1465 : node1452;
										assign node1452 = (inp[11]) ? node1456 : node1453;
											assign node1453 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node1456 = (inp[2]) ? node1458 : 16'b0000000001111111;
												assign node1458 = (inp[10]) ? 16'b0000000000111111 : node1459;
													assign node1459 = (inp[1]) ? node1461 : 16'b0000000001111111;
														assign node1461 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1465 = (inp[4]) ? node1467 : 16'b0000000001111111;
											assign node1467 = (inp[11]) ? node1475 : node1468;
												assign node1468 = (inp[1]) ? node1472 : node1469;
													assign node1469 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1472 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node1475 = (inp[2]) ? 16'b0000000000011111 : node1476;
													assign node1476 = (inp[13]) ? node1478 : 16'b0000000000111111;
														assign node1478 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
				assign node1482 = (inp[7]) ? node2256 : node1483;
					assign node1483 = (inp[9]) ? node1843 : node1484;
						assign node1484 = (inp[13]) ? node1672 : node1485;
							assign node1485 = (inp[14]) ? node1565 : node1486;
								assign node1486 = (inp[10]) ? node1522 : node1487;
									assign node1487 = (inp[8]) ? node1505 : node1488;
										assign node1488 = (inp[4]) ? node1498 : node1489;
											assign node1489 = (inp[15]) ? node1495 : node1490;
												assign node1490 = (inp[5]) ? node1492 : 16'b0001111111111111;
													assign node1492 = (inp[3]) ? 16'b0001111111111111 : 16'b0000111111111111;
												assign node1495 = (inp[5]) ? 16'b0000111111111111 : 16'b0000011111111111;
											assign node1498 = (inp[15]) ? node1500 : 16'b0000011111111111;
												assign node1500 = (inp[2]) ? 16'b0000000111111111 : node1501;
													assign node1501 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node1505 = (inp[4]) ? node1511 : node1506;
											assign node1506 = (inp[3]) ? node1508 : 16'b0000011111111111;
												assign node1508 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1511 = (inp[15]) ? node1515 : node1512;
												assign node1512 = (inp[2]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node1515 = (inp[5]) ? node1519 : node1516;
													assign node1516 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1519 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node1522 = (inp[15]) ? node1542 : node1523;
										assign node1523 = (inp[5]) ? node1533 : node1524;
											assign node1524 = (inp[11]) ? node1530 : node1525;
												assign node1525 = (inp[3]) ? 16'b0000011111111111 : node1526;
													assign node1526 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1530 = (inp[4]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node1533 = (inp[4]) ? node1539 : node1534;
												assign node1534 = (inp[3]) ? 16'b0000001111111111 : node1535;
													assign node1535 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1539 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1542 = (inp[2]) ? node1554 : node1543;
											assign node1543 = (inp[3]) ? node1547 : node1544;
												assign node1544 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1547 = (inp[8]) ? node1549 : 16'b0000011111111111;
													assign node1549 = (inp[1]) ? node1551 : 16'b0000000111111111;
														assign node1551 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1554 = (inp[11]) ? node1556 : 16'b0000000111111111;
												assign node1556 = (inp[8]) ? node1558 : 16'b0000001111111111;
													assign node1558 = (inp[5]) ? 16'b0000000011111111 : node1559;
														assign node1559 = (inp[3]) ? node1561 : 16'b0000001111111111;
															assign node1561 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node1565 = (inp[8]) ? node1615 : node1566;
									assign node1566 = (inp[2]) ? node1594 : node1567;
										assign node1567 = (inp[1]) ? node1581 : node1568;
											assign node1568 = (inp[11]) ? node1574 : node1569;
												assign node1569 = (inp[5]) ? 16'b0000011111111111 : node1570;
													assign node1570 = (inp[15]) ? 16'b0000011111111111 : 16'b0001111111111111;
												assign node1574 = (inp[5]) ? 16'b0000001111111111 : node1575;
													assign node1575 = (inp[4]) ? node1577 : 16'b0000011111111111;
														assign node1577 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1581 = (inp[15]) ? node1587 : node1582;
												assign node1582 = (inp[5]) ? 16'b0000001111111111 : node1583;
													assign node1583 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1587 = (inp[11]) ? 16'b0000000111111111 : node1588;
													assign node1588 = (inp[5]) ? node1590 : 16'b0000001111111111;
														assign node1590 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1594 = (inp[4]) ? node1604 : node1595;
											assign node1595 = (inp[1]) ? node1601 : node1596;
												assign node1596 = (inp[15]) ? node1598 : 16'b0000111111111111;
													assign node1598 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1601 = (inp[11]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node1604 = (inp[10]) ? node1612 : node1605;
												assign node1605 = (inp[1]) ? 16'b0000000111111111 : node1606;
													assign node1606 = (inp[5]) ? node1608 : 16'b0000000111111111;
														assign node1608 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1612 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1615 = (inp[4]) ? node1649 : node1616;
										assign node1616 = (inp[1]) ? node1634 : node1617;
											assign node1617 = (inp[5]) ? 16'b0000000011111111 : node1618;
												assign node1618 = (inp[3]) ? node1624 : node1619;
													assign node1619 = (inp[15]) ? node1621 : 16'b0000011111111111;
														assign node1621 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1624 = (inp[2]) ? node1628 : node1625;
														assign node1625 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1628 = (inp[10]) ? node1630 : 16'b0000001111111111;
															assign node1630 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1634 = (inp[11]) ? node1644 : node1635;
												assign node1635 = (inp[5]) ? node1637 : 16'b0000001111111111;
													assign node1637 = (inp[10]) ? 16'b0000000111111111 : node1638;
														assign node1638 = (inp[2]) ? 16'b0000000111111111 : node1639;
															assign node1639 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1644 = (inp[3]) ? node1646 : 16'b0000000111111111;
													assign node1646 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1649 = (inp[15]) ? node1665 : node1650;
											assign node1650 = (inp[11]) ? node1654 : node1651;
												assign node1651 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1654 = (inp[1]) ? node1658 : node1655;
													assign node1655 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1658 = (inp[2]) ? 16'b0000000011111111 : node1659;
														assign node1659 = (inp[10]) ? node1661 : 16'b0000000111111111;
															assign node1661 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1665 = (inp[2]) ? 16'b0000000001111111 : node1666;
												assign node1666 = (inp[10]) ? node1668 : 16'b0000000111111111;
													assign node1668 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node1672 = (inp[3]) ? node1754 : node1673;
								assign node1673 = (inp[1]) ? node1719 : node1674;
									assign node1674 = (inp[4]) ? node1690 : node1675;
										assign node1675 = (inp[15]) ? node1681 : node1676;
											assign node1676 = (inp[2]) ? node1678 : 16'b0000011111111111;
												assign node1678 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node1681 = (inp[11]) ? node1687 : node1682;
												assign node1682 = (inp[14]) ? 16'b0000001111111111 : node1683;
													assign node1683 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1687 = (inp[2]) ? 16'b0000001111111111 : 16'b0000000111111111;
										assign node1690 = (inp[11]) ? node1704 : node1691;
											assign node1691 = (inp[8]) ? node1695 : node1692;
												assign node1692 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node1695 = (inp[14]) ? node1699 : node1696;
													assign node1696 = (inp[5]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node1699 = (inp[10]) ? 16'b0000000011111111 : node1700;
														assign node1700 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1704 = (inp[8]) ? node1712 : node1705;
												assign node1705 = (inp[15]) ? node1707 : 16'b0000000111111111;
													assign node1707 = (inp[2]) ? node1709 : 16'b0000001111111111;
														assign node1709 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1712 = (inp[14]) ? node1714 : 16'b0000000111111111;
													assign node1714 = (inp[15]) ? node1716 : 16'b0000001111111111;
														assign node1716 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1719 = (inp[15]) ? node1733 : node1720;
										assign node1720 = (inp[14]) ? node1728 : node1721;
											assign node1721 = (inp[4]) ? node1723 : 16'b0000001111111111;
												assign node1723 = (inp[10]) ? node1725 : 16'b0000001111111111;
													assign node1725 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1728 = (inp[5]) ? 16'b0000000111111111 : node1729;
												assign node1729 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1733 = (inp[5]) ? node1745 : node1734;
											assign node1734 = (inp[8]) ? node1738 : node1735;
												assign node1735 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1738 = (inp[10]) ? node1740 : 16'b0000000111111111;
													assign node1740 = (inp[11]) ? 16'b0000000011111111 : node1741;
														assign node1741 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1745 = (inp[11]) ? node1751 : node1746;
												assign node1746 = (inp[4]) ? 16'b0000000001111111 : node1747;
													assign node1747 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1751 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
								assign node1754 = (inp[8]) ? node1802 : node1755;
									assign node1755 = (inp[4]) ? node1787 : node1756;
										assign node1756 = (inp[10]) ? node1766 : node1757;
											assign node1757 = (inp[11]) ? 16'b0000001111111111 : node1758;
												assign node1758 = (inp[2]) ? 16'b0000001111111111 : node1759;
													assign node1759 = (inp[5]) ? node1761 : 16'b0000011111111111;
														assign node1761 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node1766 = (inp[14]) ? node1778 : node1767;
												assign node1767 = (inp[5]) ? node1773 : node1768;
													assign node1768 = (inp[2]) ? 16'b0000001111111111 : node1769;
														assign node1769 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1773 = (inp[11]) ? node1775 : 16'b0000001111111111;
														assign node1775 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1778 = (inp[5]) ? node1782 : node1779;
													assign node1779 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1782 = (inp[2]) ? 16'b0000000011111111 : node1783;
														assign node1783 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1787 = (inp[15]) ? node1795 : node1788;
											assign node1788 = (inp[2]) ? node1792 : node1789;
												assign node1789 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1792 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node1795 = (inp[2]) ? node1797 : 16'b0000000011111111;
												assign node1797 = (inp[5]) ? node1799 : 16'b0000000111111111;
													assign node1799 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node1802 = (inp[14]) ? node1826 : node1803;
										assign node1803 = (inp[2]) ? node1819 : node1804;
											assign node1804 = (inp[1]) ? node1814 : node1805;
												assign node1805 = (inp[15]) ? node1807 : 16'b0000011111111111;
													assign node1807 = (inp[5]) ? 16'b0000000111111111 : node1808;
														assign node1808 = (inp[11]) ? node1810 : 16'b0000001111111111;
															assign node1810 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1814 = (inp[11]) ? node1816 : 16'b0000000111111111;
													assign node1816 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node1819 = (inp[11]) ? node1821 : 16'b0000000011111111;
												assign node1821 = (inp[15]) ? 16'b0000000001111111 : node1822;
													assign node1822 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000001111111;
										assign node1826 = (inp[4]) ? node1836 : node1827;
											assign node1827 = (inp[10]) ? node1829 : 16'b0000000011111111;
												assign node1829 = (inp[11]) ? 16'b0000000001111111 : node1830;
													assign node1830 = (inp[1]) ? 16'b0000000001111111 : node1831;
														assign node1831 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1836 = (inp[10]) ? node1840 : node1837;
												assign node1837 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node1840 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node1843 = (inp[3]) ? node2063 : node1844;
							assign node1844 = (inp[2]) ? node1954 : node1845;
								assign node1845 = (inp[14]) ? node1903 : node1846;
									assign node1846 = (inp[8]) ? node1870 : node1847;
										assign node1847 = (inp[15]) ? node1857 : node1848;
											assign node1848 = (inp[11]) ? node1854 : node1849;
												assign node1849 = (inp[5]) ? 16'b0000111111111111 : node1850;
													assign node1850 = (inp[1]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node1854 = (inp[5]) ? 16'b0000001111111111 : 16'b0000111111111111;
											assign node1857 = (inp[5]) ? node1865 : node1858;
												assign node1858 = (inp[13]) ? node1862 : node1859;
													assign node1859 = (inp[4]) ? 16'b0000111111111111 : 16'b0000011111111111;
													assign node1862 = (inp[1]) ? 16'b0000011111111111 : 16'b0000001111111111;
												assign node1865 = (inp[13]) ? 16'b0000000111111111 : node1866;
													assign node1866 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node1870 = (inp[1]) ? node1882 : node1871;
											assign node1871 = (inp[10]) ? node1879 : node1872;
												assign node1872 = (inp[13]) ? node1874 : 16'b0000111111111111;
													assign node1874 = (inp[5]) ? node1876 : 16'b0000011111111111;
														assign node1876 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1879 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1882 = (inp[15]) ? node1894 : node1883;
												assign node1883 = (inp[11]) ? node1889 : node1884;
													assign node1884 = (inp[4]) ? 16'b0000001111111111 : node1885;
														assign node1885 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1889 = (inp[5]) ? 16'b0000000011111111 : node1890;
														assign node1890 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1894 = (inp[4]) ? node1898 : node1895;
													assign node1895 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1898 = (inp[10]) ? node1900 : 16'b0000000111111111;
														assign node1900 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node1903 = (inp[15]) ? node1933 : node1904;
										assign node1904 = (inp[4]) ? node1918 : node1905;
											assign node1905 = (inp[10]) ? node1915 : node1906;
												assign node1906 = (inp[13]) ? node1910 : node1907;
													assign node1907 = (inp[11]) ? 16'b0000011111111111 : 16'b0001111111111111;
													assign node1910 = (inp[8]) ? node1912 : 16'b0000001111111111;
														assign node1912 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1915 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node1918 = (inp[10]) ? node1928 : node1919;
												assign node1919 = (inp[8]) ? node1925 : node1920;
													assign node1920 = (inp[5]) ? node1922 : 16'b0000001111111111;
														assign node1922 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1925 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1928 = (inp[13]) ? node1930 : 16'b0000000111111111;
													assign node1930 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1933 = (inp[5]) ? node1947 : node1934;
											assign node1934 = (inp[8]) ? node1942 : node1935;
												assign node1935 = (inp[4]) ? node1937 : 16'b0000001111111111;
													assign node1937 = (inp[13]) ? node1939 : 16'b0000000111111111;
														assign node1939 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1942 = (inp[1]) ? 16'b0000000011111111 : node1943;
													assign node1943 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1947 = (inp[11]) ? node1951 : node1948;
												assign node1948 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node1951 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1954 = (inp[11]) ? node2008 : node1955;
									assign node1955 = (inp[4]) ? node1973 : node1956;
										assign node1956 = (inp[1]) ? node1968 : node1957;
											assign node1957 = (inp[5]) ? node1963 : node1958;
												assign node1958 = (inp[13]) ? node1960 : 16'b0000011111111111;
													assign node1960 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1963 = (inp[14]) ? 16'b0000000111111111 : node1964;
													assign node1964 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1968 = (inp[8]) ? 16'b0000000000111111 : node1969;
												assign node1969 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1973 = (inp[14]) ? node1989 : node1974;
											assign node1974 = (inp[5]) ? node1982 : node1975;
												assign node1975 = (inp[13]) ? node1979 : node1976;
													assign node1976 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1979 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1982 = (inp[8]) ? node1984 : 16'b0000000111111111;
													assign node1984 = (inp[1]) ? node1986 : 16'b0000000011111111;
														assign node1986 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1989 = (inp[13]) ? node1999 : node1990;
												assign node1990 = (inp[15]) ? node1992 : 16'b0000000111111111;
													assign node1992 = (inp[8]) ? node1996 : node1993;
														assign node1993 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1996 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node1999 = (inp[5]) ? 16'b0000000000111111 : node2000;
													assign node2000 = (inp[1]) ? node2004 : node2001;
														assign node2001 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2004 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2008 = (inp[10]) ? node2036 : node2009;
										assign node2009 = (inp[14]) ? node2021 : node2010;
											assign node2010 = (inp[8]) ? node2016 : node2011;
												assign node2011 = (inp[4]) ? node2013 : 16'b0000001111111111;
													assign node2013 = (inp[1]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node2016 = (inp[4]) ? node2018 : 16'b0000000111111111;
													assign node2018 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node2021 = (inp[5]) ? node2031 : node2022;
												assign node2022 = (inp[1]) ? node2028 : node2023;
													assign node2023 = (inp[4]) ? node2025 : 16'b0000000111111111;
														assign node2025 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2028 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node2031 = (inp[13]) ? node2033 : 16'b0000000011111111;
													assign node2033 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2036 = (inp[8]) ? node2044 : node2037;
											assign node2037 = (inp[15]) ? node2039 : 16'b0000000011111111;
												assign node2039 = (inp[5]) ? 16'b0000000001111111 : node2040;
													assign node2040 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2044 = (inp[13]) ? node2052 : node2045;
												assign node2045 = (inp[1]) ? node2047 : 16'b0000000011111111;
													assign node2047 = (inp[15]) ? 16'b0000000001111111 : node2048;
														assign node2048 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2052 = (inp[5]) ? node2056 : node2053;
													assign node2053 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node2056 = (inp[14]) ? node2058 : 16'b0000000000111111;
														assign node2058 = (inp[15]) ? 16'b0000000000011111 : node2059;
															assign node2059 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node2063 = (inp[15]) ? node2157 : node2064;
								assign node2064 = (inp[8]) ? node2106 : node2065;
									assign node2065 = (inp[11]) ? node2089 : node2066;
										assign node2066 = (inp[4]) ? node2076 : node2067;
											assign node2067 = (inp[2]) ? node2071 : node2068;
												assign node2068 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2071 = (inp[5]) ? 16'b0000001111111111 : node2072;
													assign node2072 = (inp[10]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node2076 = (inp[1]) ? node2078 : 16'b0000001111111111;
												assign node2078 = (inp[13]) ? node2082 : node2079;
													assign node2079 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2082 = (inp[14]) ? node2084 : 16'b0000000011111111;
														assign node2084 = (inp[10]) ? node2086 : 16'b0000000011111111;
															assign node2086 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2089 = (inp[2]) ? node2095 : node2090;
											assign node2090 = (inp[5]) ? 16'b0000000111111111 : node2091;
												assign node2091 = (inp[1]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node2095 = (inp[4]) ? node2103 : node2096;
												assign node2096 = (inp[1]) ? node2098 : 16'b0000000111111111;
													assign node2098 = (inp[5]) ? 16'b0000000011111111 : node2099;
														assign node2099 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2103 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2106 = (inp[10]) ? node2136 : node2107;
										assign node2107 = (inp[5]) ? node2121 : node2108;
											assign node2108 = (inp[1]) ? node2114 : node2109;
												assign node2109 = (inp[2]) ? 16'b0000000111111111 : node2110;
													assign node2110 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2114 = (inp[13]) ? 16'b0000000011111111 : node2115;
													assign node2115 = (inp[2]) ? 16'b0000000111111111 : node2116;
														assign node2116 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2121 = (inp[4]) ? node2133 : node2122;
												assign node2122 = (inp[13]) ? node2124 : 16'b0000000111111111;
													assign node2124 = (inp[1]) ? node2130 : node2125;
														assign node2125 = (inp[14]) ? node2127 : 16'b0000000111111111;
															assign node2127 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2130 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2133 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2136 = (inp[2]) ? node2148 : node2137;
											assign node2137 = (inp[4]) ? node2143 : node2138;
												assign node2138 = (inp[11]) ? node2140 : 16'b0000011111111111;
													assign node2140 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2143 = (inp[13]) ? node2145 : 16'b0000000011111111;
													assign node2145 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2148 = (inp[11]) ? node2154 : node2149;
												assign node2149 = (inp[13]) ? 16'b0000000001111111 : node2150;
													assign node2150 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2154 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000111111;
								assign node2157 = (inp[11]) ? node2199 : node2158;
									assign node2158 = (inp[5]) ? node2178 : node2159;
										assign node2159 = (inp[10]) ? node2169 : node2160;
											assign node2160 = (inp[4]) ? 16'b0000000111111111 : node2161;
												assign node2161 = (inp[1]) ? node2165 : node2162;
													assign node2162 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2165 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2169 = (inp[4]) ? node2175 : node2170;
												assign node2170 = (inp[13]) ? 16'b0000000011111111 : node2171;
													assign node2171 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2175 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2178 = (inp[8]) ? node2190 : node2179;
											assign node2179 = (inp[2]) ? node2183 : node2180;
												assign node2180 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2183 = (inp[13]) ? node2185 : 16'b0000000011111111;
													assign node2185 = (inp[10]) ? 16'b0000000001111111 : node2186;
														assign node2186 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2190 = (inp[13]) ? node2192 : 16'b0000000011111111;
												assign node2192 = (inp[14]) ? node2194 : 16'b0000000001111111;
													assign node2194 = (inp[2]) ? 16'b0000000000111111 : node2195;
														assign node2195 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node2199 = (inp[5]) ? node2231 : node2200;
										assign node2200 = (inp[10]) ? node2214 : node2201;
											assign node2201 = (inp[2]) ? 16'b0000000011111111 : node2202;
												assign node2202 = (inp[1]) ? node2210 : node2203;
													assign node2203 = (inp[8]) ? 16'b0000000011111111 : node2204;
														assign node2204 = (inp[13]) ? node2206 : 16'b0000000111111111;
															assign node2206 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2210 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2214 = (inp[14]) ? node2224 : node2215;
												assign node2215 = (inp[2]) ? node2219 : node2216;
													assign node2216 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node2219 = (inp[8]) ? node2221 : 16'b0000000001111111;
														assign node2221 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node2224 = (inp[4]) ? 16'b0000000000111111 : node2225;
													assign node2225 = (inp[13]) ? node2227 : 16'b0000000001111111;
														assign node2227 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2231 = (inp[1]) ? node2243 : node2232;
											assign node2232 = (inp[8]) ? node2240 : node2233;
												assign node2233 = (inp[2]) ? node2235 : 16'b0000000011111111;
													assign node2235 = (inp[14]) ? 16'b0000000000111111 : node2236;
														assign node2236 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2240 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2243 = (inp[8]) ? node2249 : node2244;
												assign node2244 = (inp[2]) ? node2246 : 16'b0000000000111111;
													assign node2246 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node2249 = (inp[2]) ? node2251 : 16'b0000000000011111;
													assign node2251 = (inp[4]) ? node2253 : 16'b0000000000011111;
														assign node2253 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node2256 = (inp[1]) ? node2636 : node2257;
						assign node2257 = (inp[2]) ? node2459 : node2258;
							assign node2258 = (inp[15]) ? node2354 : node2259;
								assign node2259 = (inp[14]) ? node2307 : node2260;
									assign node2260 = (inp[3]) ? node2286 : node2261;
										assign node2261 = (inp[8]) ? node2273 : node2262;
											assign node2262 = (inp[9]) ? node2270 : node2263;
												assign node2263 = (inp[11]) ? node2265 : 16'b0000111111111111;
													assign node2265 = (inp[5]) ? 16'b0000011111111111 : node2266;
														assign node2266 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2270 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2273 = (inp[10]) ? 16'b0000000111111111 : node2274;
												assign node2274 = (inp[4]) ? node2282 : node2275;
													assign node2275 = (inp[9]) ? node2277 : 16'b0000011111111111;
														assign node2277 = (inp[5]) ? 16'b0000001111111111 : node2278;
															assign node2278 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2282 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2286 = (inp[8]) ? node2298 : node2287;
											assign node2287 = (inp[10]) ? node2293 : node2288;
												assign node2288 = (inp[4]) ? 16'b0000001111111111 : node2289;
													assign node2289 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2293 = (inp[5]) ? node2295 : 16'b0000001111111111;
													assign node2295 = (inp[9]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node2298 = (inp[13]) ? node2304 : node2299;
												assign node2299 = (inp[5]) ? 16'b0000000111111111 : node2300;
													assign node2300 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2304 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node2307 = (inp[4]) ? node2335 : node2308;
										assign node2308 = (inp[9]) ? node2322 : node2309;
											assign node2309 = (inp[5]) ? node2319 : node2310;
												assign node2310 = (inp[13]) ? 16'b0000001111111111 : node2311;
													assign node2311 = (inp[10]) ? node2313 : 16'b0000111111111111;
														assign node2313 = (inp[11]) ? 16'b0000011111111111 : node2314;
															assign node2314 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2319 = (inp[8]) ? 16'b0000000111111111 : 16'b0000011111111111;
											assign node2322 = (inp[8]) ? node2330 : node2323;
												assign node2323 = (inp[13]) ? node2327 : node2324;
													assign node2324 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2327 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node2330 = (inp[5]) ? 16'b0000000011111111 : node2331;
													assign node2331 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2335 = (inp[11]) ? node2347 : node2336;
											assign node2336 = (inp[8]) ? node2344 : node2337;
												assign node2337 = (inp[9]) ? node2341 : node2338;
													assign node2338 = (inp[5]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node2341 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2344 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2347 = (inp[9]) ? node2349 : 16'b0000000011111111;
												assign node2349 = (inp[5]) ? node2351 : 16'b0000000001111111;
													assign node2351 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node2354 = (inp[11]) ? node2404 : node2355;
									assign node2355 = (inp[10]) ? node2379 : node2356;
										assign node2356 = (inp[5]) ? node2368 : node2357;
											assign node2357 = (inp[9]) ? node2365 : node2358;
												assign node2358 = (inp[8]) ? 16'b0000001111111111 : node2359;
													assign node2359 = (inp[14]) ? 16'b0000011111111111 : node2360;
														assign node2360 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2365 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2368 = (inp[4]) ? 16'b0000000011111111 : node2369;
												assign node2369 = (inp[8]) ? node2371 : 16'b0000001111111111;
													assign node2371 = (inp[14]) ? 16'b0000000001111111 : node2372;
														assign node2372 = (inp[3]) ? node2374 : 16'b0000001111111111;
															assign node2374 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2379 = (inp[4]) ? node2385 : node2380;
											assign node2380 = (inp[14]) ? node2382 : 16'b0000000111111111;
												assign node2382 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2385 = (inp[5]) ? node2395 : node2386;
												assign node2386 = (inp[8]) ? node2388 : 16'b0000001111111111;
													assign node2388 = (inp[9]) ? 16'b0000000011111111 : node2389;
														assign node2389 = (inp[3]) ? node2391 : 16'b0000000111111111;
															assign node2391 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node2395 = (inp[8]) ? node2399 : node2396;
													assign node2396 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2399 = (inp[3]) ? node2401 : 16'b0000000001111111;
														assign node2401 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node2404 = (inp[8]) ? node2434 : node2405;
										assign node2405 = (inp[13]) ? node2421 : node2406;
											assign node2406 = (inp[10]) ? node2412 : node2407;
												assign node2407 = (inp[3]) ? node2409 : 16'b0000001111111111;
													assign node2409 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2412 = (inp[5]) ? node2418 : node2413;
													assign node2413 = (inp[3]) ? 16'b0000000111111111 : node2414;
														assign node2414 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2418 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000111111111;
											assign node2421 = (inp[14]) ? node2425 : node2422;
												assign node2422 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2425 = (inp[10]) ? node2429 : node2426;
													assign node2426 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node2429 = (inp[9]) ? node2431 : 16'b0000000001111111;
														assign node2431 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2434 = (inp[3]) ? node2450 : node2435;
											assign node2435 = (inp[5]) ? node2441 : node2436;
												assign node2436 = (inp[4]) ? node2438 : 16'b0000000111111111;
													assign node2438 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2441 = (inp[10]) ? node2447 : node2442;
													assign node2442 = (inp[4]) ? node2444 : 16'b0000000011111111;
														assign node2444 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2447 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2450 = (inp[10]) ? node2454 : node2451;
												assign node2451 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2454 = (inp[14]) ? node2456 : 16'b0000000000111111;
													assign node2456 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node2459 = (inp[11]) ? node2551 : node2460;
								assign node2460 = (inp[9]) ? node2502 : node2461;
									assign node2461 = (inp[15]) ? node2483 : node2462;
										assign node2462 = (inp[14]) ? node2470 : node2463;
											assign node2463 = (inp[3]) ? node2467 : node2464;
												assign node2464 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2467 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2470 = (inp[4]) ? node2476 : node2471;
												assign node2471 = (inp[5]) ? 16'b0000000111111111 : node2472;
													assign node2472 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2476 = (inp[5]) ? 16'b0000000011111111 : node2477;
													assign node2477 = (inp[10]) ? node2479 : 16'b0000000111111111;
														assign node2479 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2483 = (inp[3]) ? node2489 : node2484;
											assign node2484 = (inp[10]) ? 16'b0000000011111111 : node2485;
												assign node2485 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2489 = (inp[13]) ? node2491 : 16'b0000001111111111;
												assign node2491 = (inp[4]) ? node2497 : node2492;
													assign node2492 = (inp[5]) ? 16'b0000000011111111 : node2493;
														assign node2493 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2497 = (inp[5]) ? 16'b0000000001111111 : node2498;
														assign node2498 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2502 = (inp[3]) ? node2526 : node2503;
										assign node2503 = (inp[5]) ? node2515 : node2504;
											assign node2504 = (inp[15]) ? node2512 : node2505;
												assign node2505 = (inp[10]) ? node2507 : 16'b0000011111111111;
													assign node2507 = (inp[14]) ? 16'b0000000111111111 : node2508;
														assign node2508 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2512 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2515 = (inp[13]) ? node2519 : node2516;
												assign node2516 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2519 = (inp[4]) ? node2521 : 16'b0000000011111111;
													assign node2521 = (inp[10]) ? 16'b0000000000111111 : node2522;
														assign node2522 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2526 = (inp[10]) ? node2538 : node2527;
											assign node2527 = (inp[8]) ? node2531 : node2528;
												assign node2528 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2531 = (inp[5]) ? 16'b0000000001111111 : node2532;
													assign node2532 = (inp[4]) ? node2534 : 16'b0000000011111111;
														assign node2534 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2538 = (inp[4]) ? node2546 : node2539;
												assign node2539 = (inp[14]) ? node2541 : 16'b0000000011111111;
													assign node2541 = (inp[8]) ? 16'b0000000001111111 : node2542;
														assign node2542 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2546 = (inp[13]) ? node2548 : 16'b0000000001111111;
													assign node2548 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node2551 = (inp[8]) ? node2593 : node2552;
									assign node2552 = (inp[3]) ? node2574 : node2553;
										assign node2553 = (inp[4]) ? node2567 : node2554;
											assign node2554 = (inp[13]) ? node2558 : node2555;
												assign node2555 = (inp[9]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node2558 = (inp[15]) ? node2562 : node2559;
													assign node2559 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2562 = (inp[5]) ? node2564 : 16'b0000000111111111;
														assign node2564 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2567 = (inp[13]) ? node2569 : 16'b0000000111111111;
												assign node2569 = (inp[14]) ? node2571 : 16'b0000000011111111;
													assign node2571 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2574 = (inp[5]) ? node2582 : node2575;
											assign node2575 = (inp[15]) ? node2579 : node2576;
												assign node2576 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2579 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2582 = (inp[10]) ? node2588 : node2583;
												assign node2583 = (inp[15]) ? node2585 : 16'b0000000011111111;
													assign node2585 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2588 = (inp[9]) ? node2590 : 16'b0000000001111111;
													assign node2590 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node2593 = (inp[15]) ? node2621 : node2594;
										assign node2594 = (inp[13]) ? node2610 : node2595;
											assign node2595 = (inp[3]) ? node2601 : node2596;
												assign node2596 = (inp[10]) ? node2598 : 16'b0000000111111111;
													assign node2598 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node2601 = (inp[14]) ? node2603 : 16'b0000000011111111;
													assign node2603 = (inp[5]) ? node2607 : node2604;
														assign node2604 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node2607 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node2610 = (inp[4]) ? node2614 : node2611;
												assign node2611 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2614 = (inp[3]) ? 16'b0000000000111111 : node2615;
													assign node2615 = (inp[5]) ? 16'b0000000000111111 : node2616;
														assign node2616 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2621 = (inp[14]) ? node2631 : node2622;
											assign node2622 = (inp[5]) ? node2626 : node2623;
												assign node2623 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2626 = (inp[4]) ? node2628 : 16'b0000000000011111;
													assign node2628 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2631 = (inp[3]) ? 16'b0000000000011111 : node2632;
												assign node2632 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node2636 = (inp[10]) ? node2810 : node2637;
							assign node2637 = (inp[14]) ? node2719 : node2638;
								assign node2638 = (inp[15]) ? node2688 : node2639;
									assign node2639 = (inp[11]) ? node2661 : node2640;
										assign node2640 = (inp[2]) ? node2654 : node2641;
											assign node2641 = (inp[8]) ? node2651 : node2642;
												assign node2642 = (inp[13]) ? 16'b0000001111111111 : node2643;
													assign node2643 = (inp[9]) ? 16'b0000011111111111 : node2644;
														assign node2644 = (inp[4]) ? node2646 : 16'b0001111111111111;
															assign node2646 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2651 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2654 = (inp[3]) ? node2658 : node2655;
												assign node2655 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2658 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node2661 = (inp[5]) ? node2673 : node2662;
											assign node2662 = (inp[9]) ? node2670 : node2663;
												assign node2663 = (inp[13]) ? 16'b0000000111111111 : node2664;
													assign node2664 = (inp[2]) ? node2666 : 16'b0000011111111111;
														assign node2666 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2670 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node2673 = (inp[4]) ? node2681 : node2674;
												assign node2674 = (inp[9]) ? 16'b0000000011111111 : node2675;
													assign node2675 = (inp[13]) ? node2677 : 16'b0000000111111111;
														assign node2677 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2681 = (inp[3]) ? 16'b0000000001111111 : node2682;
													assign node2682 = (inp[13]) ? node2684 : 16'b0000000011111111;
														assign node2684 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2688 = (inp[9]) ? node2708 : node2689;
										assign node2689 = (inp[2]) ? node2699 : node2690;
											assign node2690 = (inp[4]) ? node2694 : node2691;
												assign node2691 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node2694 = (inp[11]) ? node2696 : 16'b0000000111111111;
													assign node2696 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2699 = (inp[4]) ? node2705 : node2700;
												assign node2700 = (inp[3]) ? 16'b0000000011111111 : node2701;
													assign node2701 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2705 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2708 = (inp[3]) ? node2710 : 16'b0000000011111111;
											assign node2710 = (inp[13]) ? node2714 : node2711;
												assign node2711 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node2714 = (inp[5]) ? node2716 : 16'b0000000000111111;
													assign node2716 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node2719 = (inp[8]) ? node2759 : node2720;
									assign node2720 = (inp[5]) ? node2740 : node2721;
										assign node2721 = (inp[2]) ? node2729 : node2722;
											assign node2722 = (inp[11]) ? 16'b0000000011111111 : node2723;
												assign node2723 = (inp[15]) ? 16'b0000000111111111 : node2724;
													assign node2724 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2729 = (inp[9]) ? node2733 : node2730;
												assign node2730 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2733 = (inp[15]) ? node2735 : 16'b0000000011111111;
													assign node2735 = (inp[3]) ? 16'b0000000001111111 : node2736;
														assign node2736 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2740 = (inp[13]) ? node2752 : node2741;
											assign node2741 = (inp[11]) ? node2747 : node2742;
												assign node2742 = (inp[4]) ? 16'b0000000011111111 : node2743;
													assign node2743 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2747 = (inp[2]) ? 16'b0000000001111111 : node2748;
													assign node2748 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node2752 = (inp[3]) ? node2756 : node2753;
												assign node2753 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2756 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000000011111;
									assign node2759 = (inp[4]) ? node2781 : node2760;
										assign node2760 = (inp[5]) ? node2774 : node2761;
											assign node2761 = (inp[2]) ? node2769 : node2762;
												assign node2762 = (inp[11]) ? 16'b0000000011111111 : node2763;
													assign node2763 = (inp[15]) ? 16'b0000000111111111 : node2764;
														assign node2764 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2769 = (inp[15]) ? node2771 : 16'b0000000011111111;
													assign node2771 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2774 = (inp[2]) ? node2778 : node2775;
												assign node2775 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2778 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000011111;
										assign node2781 = (inp[5]) ? node2791 : node2782;
											assign node2782 = (inp[15]) ? node2784 : 16'b0000000001111111;
												assign node2784 = (inp[11]) ? node2788 : node2785;
													assign node2785 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node2788 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2791 = (inp[9]) ? node2801 : node2792;
												assign node2792 = (inp[11]) ? 16'b0000000000111111 : node2793;
													assign node2793 = (inp[2]) ? node2795 : 16'b0000000001111111;
														assign node2795 = (inp[15]) ? 16'b0000000000011111 : node2796;
															assign node2796 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2801 = (inp[11]) ? node2803 : 16'b0000000000111111;
													assign node2803 = (inp[3]) ? 16'b0000000000001111 : node2804;
														assign node2804 = (inp[15]) ? node2806 : 16'b0000000000011111;
															assign node2806 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node2810 = (inp[15]) ? node2904 : node2811;
								assign node2811 = (inp[2]) ? node2853 : node2812;
									assign node2812 = (inp[9]) ? node2830 : node2813;
										assign node2813 = (inp[11]) ? node2821 : node2814;
											assign node2814 = (inp[5]) ? 16'b0000000111111111 : node2815;
												assign node2815 = (inp[14]) ? node2817 : 16'b0000011111111111;
													assign node2817 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2821 = (inp[14]) ? node2827 : node2822;
												assign node2822 = (inp[8]) ? node2824 : 16'b0000000111111111;
													assign node2824 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2827 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2830 = (inp[8]) ? node2842 : node2831;
											assign node2831 = (inp[3]) ? node2837 : node2832;
												assign node2832 = (inp[11]) ? 16'b0000000011111111 : node2833;
													assign node2833 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2837 = (inp[11]) ? 16'b0000000011111111 : node2838;
													assign node2838 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2842 = (inp[3]) ? node2846 : node2843;
												assign node2843 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2846 = (inp[13]) ? node2848 : 16'b0000000111111111;
													assign node2848 = (inp[5]) ? node2850 : 16'b0000000000111111;
														assign node2850 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node2853 = (inp[13]) ? node2879 : node2854;
										assign node2854 = (inp[11]) ? node2872 : node2855;
											assign node2855 = (inp[8]) ? node2867 : node2856;
												assign node2856 = (inp[5]) ? node2860 : node2857;
													assign node2857 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2860 = (inp[3]) ? node2862 : 16'b0000000011111111;
														assign node2862 = (inp[9]) ? node2864 : 16'b0000000011111111;
															assign node2864 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2867 = (inp[14]) ? 16'b0000000001111111 : node2868;
													assign node2868 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node2872 = (inp[9]) ? node2874 : 16'b0000000001111111;
												assign node2874 = (inp[14]) ? 16'b0000000000111111 : node2875;
													assign node2875 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2879 = (inp[9]) ? node2889 : node2880;
											assign node2880 = (inp[4]) ? node2886 : node2881;
												assign node2881 = (inp[3]) ? 16'b0000000001111111 : node2882;
													assign node2882 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2886 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node2889 = (inp[5]) ? node2897 : node2890;
												assign node2890 = (inp[3]) ? 16'b0000000001111111 : node2891;
													assign node2891 = (inp[4]) ? node2893 : 16'b0000000000111111;
														assign node2893 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node2897 = (inp[8]) ? node2899 : 16'b0000000000111111;
													assign node2899 = (inp[11]) ? node2901 : 16'b0000000000011111;
														assign node2901 = (inp[3]) ? 16'b0000000000000111 : 16'b0000000000011111;
								assign node2904 = (inp[9]) ? node2942 : node2905;
									assign node2905 = (inp[2]) ? node2927 : node2906;
										assign node2906 = (inp[8]) ? node2916 : node2907;
											assign node2907 = (inp[3]) ? node2909 : 16'b0000000011111111;
												assign node2909 = (inp[14]) ? 16'b0000000001111111 : node2910;
													assign node2910 = (inp[4]) ? 16'b0000000001111111 : node2911;
														assign node2911 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node2916 = (inp[13]) ? 16'b0000000000111111 : node2917;
												assign node2917 = (inp[4]) ? node2921 : node2918;
													assign node2918 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2921 = (inp[3]) ? node2923 : 16'b0000000001111111;
														assign node2923 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000000111111;
										assign node2927 = (inp[3]) ? node2931 : node2928;
											assign node2928 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2931 = (inp[11]) ? node2937 : node2932;
												assign node2932 = (inp[5]) ? node2934 : 16'b0000000000111111;
													assign node2934 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2937 = (inp[14]) ? 16'b0000000000001111 : node2938;
													assign node2938 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node2942 = (inp[3]) ? node2964 : node2943;
										assign node2943 = (inp[11]) ? node2953 : node2944;
											assign node2944 = (inp[8]) ? node2950 : node2945;
												assign node2945 = (inp[5]) ? 16'b0000000001111111 : node2946;
													assign node2946 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2950 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node2953 = (inp[8]) ? node2959 : node2954;
												assign node2954 = (inp[14]) ? 16'b0000000000011111 : node2955;
													assign node2955 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2959 = (inp[13]) ? 16'b0000000000001111 : node2960;
													assign node2960 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node2964 = (inp[4]) ? node2976 : node2965;
											assign node2965 = (inp[13]) ? node2971 : node2966;
												assign node2966 = (inp[14]) ? 16'b0000000000111111 : node2967;
													assign node2967 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node2971 = (inp[5]) ? node2973 : 16'b0000000000111111;
													assign node2973 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node2976 = (inp[13]) ? node2984 : node2977;
												assign node2977 = (inp[14]) ? node2979 : 16'b0000000000011111;
													assign node2979 = (inp[5]) ? node2981 : 16'b0000000000111111;
														assign node2981 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node2984 = (inp[8]) ? node2986 : 16'b0000000000011111;
													assign node2986 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
			assign node2989 = (inp[10]) ? node4451 : node2990;
				assign node2990 = (inp[13]) ? node3708 : node2991;
					assign node2991 = (inp[11]) ? node3349 : node2992;
						assign node2992 = (inp[14]) ? node3190 : node2993;
							assign node2993 = (inp[4]) ? node3095 : node2994;
								assign node2994 = (inp[0]) ? node3040 : node2995;
									assign node2995 = (inp[8]) ? node3019 : node2996;
										assign node2996 = (inp[7]) ? node3010 : node2997;
											assign node2997 = (inp[5]) ? 16'b0000111111111111 : node2998;
												assign node2998 = (inp[9]) ? node3006 : node2999;
													assign node2999 = (inp[15]) ? 16'b0001111111111111 : node3000;
														assign node3000 = (inp[3]) ? node3002 : 16'b0011111111111111;
															assign node3002 = (inp[2]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node3006 = (inp[15]) ? 16'b0000111111111111 : 16'b0001111111111111;
											assign node3010 = (inp[3]) ? 16'b0000001111111111 : node3011;
												assign node3011 = (inp[5]) ? node3013 : 16'b0000111111111111;
													assign node3013 = (inp[1]) ? 16'b0000011111111111 : node3014;
														assign node3014 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node3019 = (inp[9]) ? node3037 : node3020;
											assign node3020 = (inp[15]) ? node3030 : node3021;
												assign node3021 = (inp[7]) ? node3027 : node3022;
													assign node3022 = (inp[3]) ? 16'b0000111111111111 : node3023;
														assign node3023 = (inp[2]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node3027 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node3030 = (inp[1]) ? node3032 : 16'b0000011111111111;
													assign node3032 = (inp[3]) ? 16'b0000001111111111 : node3033;
														assign node3033 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3037 = (inp[5]) ? 16'b0000000111111111 : 16'b0000011111111111;
									assign node3040 = (inp[1]) ? node3066 : node3041;
										assign node3041 = (inp[15]) ? node3053 : node3042;
											assign node3042 = (inp[7]) ? node3046 : node3043;
												assign node3043 = (inp[5]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node3046 = (inp[3]) ? 16'b0000001111111111 : node3047;
													assign node3047 = (inp[9]) ? 16'b0000011111111111 : node3048;
														assign node3048 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node3053 = (inp[8]) ? node3061 : node3054;
												assign node3054 = (inp[2]) ? node3058 : node3055;
													assign node3055 = (inp[7]) ? 16'b0000111111111111 : 16'b0000011111111111;
													assign node3058 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3061 = (inp[2]) ? node3063 : 16'b0000001111111111;
													assign node3063 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node3066 = (inp[3]) ? node3082 : node3067;
											assign node3067 = (inp[2]) ? node3079 : node3068;
												assign node3068 = (inp[15]) ? node3074 : node3069;
													assign node3069 = (inp[9]) ? node3071 : 16'b0000011111111111;
														assign node3071 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3074 = (inp[7]) ? node3076 : 16'b0000001111111111;
														assign node3076 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3079 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3082 = (inp[15]) ? node3092 : node3083;
												assign node3083 = (inp[8]) ? node3087 : node3084;
													assign node3084 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3087 = (inp[7]) ? 16'b0000000111111111 : node3088;
														assign node3088 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3092 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node3095 = (inp[7]) ? node3137 : node3096;
									assign node3096 = (inp[1]) ? node3116 : node3097;
										assign node3097 = (inp[0]) ? node3107 : node3098;
											assign node3098 = (inp[9]) ? node3102 : node3099;
												assign node3099 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node3102 = (inp[15]) ? 16'b0000011111111111 : node3103;
													assign node3103 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node3107 = (inp[2]) ? node3113 : node3108;
												assign node3108 = (inp[9]) ? node3110 : 16'b0000011111111111;
													assign node3110 = (inp[5]) ? 16'b0000011111111111 : 16'b0000001111111111;
												assign node3113 = (inp[9]) ? 16'b0000001111111111 : 16'b0000000111111111;
										assign node3116 = (inp[15]) ? node3130 : node3117;
											assign node3117 = (inp[0]) ? node3127 : node3118;
												assign node3118 = (inp[3]) ? node3122 : node3119;
													assign node3119 = (inp[8]) ? 16'b0000111111111111 : 16'b0000011111111111;
													assign node3122 = (inp[9]) ? 16'b0000001111111111 : node3123;
														assign node3123 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3127 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3130 = (inp[5]) ? node3134 : node3131;
												assign node3131 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3134 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
									assign node3137 = (inp[5]) ? node3163 : node3138;
										assign node3138 = (inp[9]) ? node3150 : node3139;
											assign node3139 = (inp[0]) ? node3147 : node3140;
												assign node3140 = (inp[3]) ? node3142 : 16'b0000111111111111;
													assign node3142 = (inp[2]) ? 16'b0000001111111111 : node3143;
														assign node3143 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3147 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3150 = (inp[15]) ? node3158 : node3151;
												assign node3151 = (inp[2]) ? 16'b0000000111111111 : node3152;
													assign node3152 = (inp[3]) ? node3154 : 16'b0000001111111111;
														assign node3154 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3158 = (inp[3]) ? node3160 : 16'b0000001111111111;
													assign node3160 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3163 = (inp[9]) ? node3179 : node3164;
											assign node3164 = (inp[3]) ? node3170 : node3165;
												assign node3165 = (inp[8]) ? node3167 : 16'b0000001111111111;
													assign node3167 = (inp[1]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node3170 = (inp[1]) ? node3174 : node3171;
													assign node3171 = (inp[2]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node3174 = (inp[15]) ? 16'b0000000011111111 : node3175;
														assign node3175 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node3179 = (inp[2]) ? node3185 : node3180;
												assign node3180 = (inp[0]) ? 16'b0000000011111111 : node3181;
													assign node3181 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3185 = (inp[0]) ? node3187 : 16'b0000000011111111;
													assign node3187 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node3190 = (inp[7]) ? node3274 : node3191;
								assign node3191 = (inp[8]) ? node3241 : node3192;
									assign node3192 = (inp[1]) ? node3214 : node3193;
										assign node3193 = (inp[2]) ? node3201 : node3194;
											assign node3194 = (inp[4]) ? 16'b0000011111111111 : node3195;
												assign node3195 = (inp[0]) ? node3197 : 16'b0000111111111111;
													assign node3197 = (inp[9]) ? 16'b0000111111111111 : 16'b0000011111111111;
											assign node3201 = (inp[5]) ? node3203 : 16'b0000011111111111;
												assign node3203 = (inp[9]) ? node3211 : node3204;
													assign node3204 = (inp[0]) ? 16'b0000000111111111 : node3205;
														assign node3205 = (inp[3]) ? 16'b0000011111111111 : node3206;
															assign node3206 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3211 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node3214 = (inp[9]) ? node3232 : node3215;
											assign node3215 = (inp[15]) ? node3225 : node3216;
												assign node3216 = (inp[5]) ? node3220 : node3217;
													assign node3217 = (inp[4]) ? 16'b0000111111111111 : 16'b0000011111111111;
													assign node3220 = (inp[3]) ? 16'b0000001111111111 : node3221;
														assign node3221 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3225 = (inp[5]) ? node3227 : 16'b0000001111111111;
													assign node3227 = (inp[2]) ? 16'b0000000111111111 : node3228;
														assign node3228 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3232 = (inp[4]) ? node3236 : node3233;
												assign node3233 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3236 = (inp[2]) ? 16'b0000000000111111 : node3237;
													assign node3237 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node3241 = (inp[0]) ? node3259 : node3242;
										assign node3242 = (inp[3]) ? node3246 : node3243;
											assign node3243 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3246 = (inp[5]) ? node3254 : node3247;
												assign node3247 = (inp[2]) ? 16'b0000000111111111 : node3248;
													assign node3248 = (inp[1]) ? node3250 : 16'b0000011111111111;
														assign node3250 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3254 = (inp[4]) ? 16'b0000000011111111 : node3255;
													assign node3255 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3259 = (inp[15]) ? node3267 : node3260;
											assign node3260 = (inp[2]) ? node3264 : node3261;
												assign node3261 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3264 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3267 = (inp[4]) ? 16'b0000000011111111 : node3268;
												assign node3268 = (inp[5]) ? 16'b0000000001111111 : node3269;
													assign node3269 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node3274 = (inp[4]) ? node3316 : node3275;
									assign node3275 = (inp[2]) ? node3297 : node3276;
										assign node3276 = (inp[1]) ? node3284 : node3277;
											assign node3277 = (inp[15]) ? node3279 : 16'b0000011111111111;
												assign node3279 = (inp[3]) ? 16'b0000001111111111 : node3280;
													assign node3280 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3284 = (inp[8]) ? node3294 : node3285;
												assign node3285 = (inp[15]) ? node3291 : node3286;
													assign node3286 = (inp[0]) ? 16'b0000001111111111 : node3287;
														assign node3287 = (inp[9]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node3291 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3294 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3297 = (inp[3]) ? node3307 : node3298;
											assign node3298 = (inp[9]) ? node3302 : node3299;
												assign node3299 = (inp[8]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node3302 = (inp[0]) ? node3304 : 16'b0000000111111111;
													assign node3304 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3307 = (inp[9]) ? node3311 : node3308;
												assign node3308 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3311 = (inp[5]) ? 16'b0000000001111111 : node3312;
													assign node3312 = (inp[8]) ? 16'b0000000001111111 : 16'b0000001111111111;
									assign node3316 = (inp[3]) ? node3328 : node3317;
										assign node3317 = (inp[0]) ? node3325 : node3318;
											assign node3318 = (inp[15]) ? node3320 : 16'b0000000111111111;
												assign node3320 = (inp[5]) ? node3322 : 16'b0000001111111111;
													assign node3322 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3325 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3328 = (inp[5]) ? node3338 : node3329;
											assign node3329 = (inp[0]) ? node3333 : node3330;
												assign node3330 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3333 = (inp[9]) ? node3335 : 16'b0000000011111111;
													assign node3335 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3338 = (inp[1]) ? 16'b0000000001111111 : node3339;
												assign node3339 = (inp[15]) ? node3343 : node3340;
													assign node3340 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node3343 = (inp[9]) ? 16'b0000000001111111 : node3344;
														assign node3344 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
						assign node3349 = (inp[8]) ? node3541 : node3350;
							assign node3350 = (inp[3]) ? node3430 : node3351;
								assign node3351 = (inp[7]) ? node3379 : node3352;
									assign node3352 = (inp[0]) ? node3366 : node3353;
										assign node3353 = (inp[1]) ? node3361 : node3354;
											assign node3354 = (inp[4]) ? node3358 : node3355;
												assign node3355 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node3358 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node3361 = (inp[14]) ? node3363 : 16'b0000011111111111;
												assign node3363 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node3366 = (inp[14]) ? node3374 : node3367;
											assign node3367 = (inp[5]) ? node3371 : node3368;
												assign node3368 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3371 = (inp[15]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node3374 = (inp[1]) ? 16'b0000000111111111 : node3375;
												assign node3375 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node3379 = (inp[9]) ? node3407 : node3380;
										assign node3380 = (inp[2]) ? node3396 : node3381;
											assign node3381 = (inp[4]) ? node3387 : node3382;
												assign node3382 = (inp[0]) ? node3384 : 16'b0000011111111111;
													assign node3384 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3387 = (inp[15]) ? node3391 : node3388;
													assign node3388 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3391 = (inp[0]) ? 16'b0000000111111111 : node3392;
														assign node3392 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3396 = (inp[4]) ? node3400 : node3397;
												assign node3397 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3400 = (inp[5]) ? 16'b0000000011111111 : node3401;
													assign node3401 = (inp[15]) ? 16'b0000001111111111 : node3402;
														assign node3402 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3407 = (inp[5]) ? node3411 : node3408;
											assign node3408 = (inp[0]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node3411 = (inp[14]) ? 16'b0000000011111111 : node3412;
												assign node3412 = (inp[1]) ? node3420 : node3413;
													assign node3413 = (inp[0]) ? node3415 : 16'b0000000111111111;
														assign node3415 = (inp[4]) ? node3417 : 16'b0000000111111111;
															assign node3417 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3420 = (inp[0]) ? 16'b0000000011111111 : node3421;
														assign node3421 = (inp[15]) ? node3425 : node3422;
															assign node3422 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
															assign node3425 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000011111111;
								assign node3430 = (inp[15]) ? node3486 : node3431;
									assign node3431 = (inp[0]) ? node3459 : node3432;
										assign node3432 = (inp[9]) ? node3450 : node3433;
											assign node3433 = (inp[1]) ? node3447 : node3434;
												assign node3434 = (inp[7]) ? node3440 : node3435;
													assign node3435 = (inp[2]) ? node3437 : 16'b0000011111111111;
														assign node3437 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3440 = (inp[5]) ? node3442 : 16'b0000011111111111;
														assign node3442 = (inp[14]) ? node3444 : 16'b0000001111111111;
															assign node3444 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3447 = (inp[14]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node3450 = (inp[4]) ? 16'b0000000111111111 : node3451;
												assign node3451 = (inp[2]) ? node3453 : 16'b0000001111111111;
													assign node3453 = (inp[14]) ? 16'b0000000011111111 : node3454;
														assign node3454 = (inp[1]) ? 16'b0000001111111111 : 16'b0000000111111111;
										assign node3459 = (inp[5]) ? node3471 : node3460;
											assign node3460 = (inp[2]) ? node3464 : node3461;
												assign node3461 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3464 = (inp[1]) ? 16'b0000000011111111 : node3465;
													assign node3465 = (inp[7]) ? node3467 : 16'b0000000111111111;
														assign node3467 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3471 = (inp[14]) ? node3479 : node3472;
												assign node3472 = (inp[2]) ? 16'b0000000011111111 : node3473;
													assign node3473 = (inp[1]) ? 16'b0000000111111111 : node3474;
														assign node3474 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3479 = (inp[1]) ? node3481 : 16'b0000000011111111;
													assign node3481 = (inp[7]) ? node3483 : 16'b0000000000111111;
														assign node3483 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node3486 = (inp[1]) ? node3518 : node3487;
										assign node3487 = (inp[14]) ? node3501 : node3488;
											assign node3488 = (inp[2]) ? node3492 : node3489;
												assign node3489 = (inp[5]) ? 16'b0000000011111111 : 16'b0000011111111111;
												assign node3492 = (inp[0]) ? node3498 : node3493;
													assign node3493 = (inp[7]) ? 16'b0000000111111111 : node3494;
														assign node3494 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3498 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3501 = (inp[0]) ? node3511 : node3502;
												assign node3502 = (inp[9]) ? 16'b0000000011111111 : node3503;
													assign node3503 = (inp[7]) ? node3505 : 16'b0000000111111111;
														assign node3505 = (inp[2]) ? 16'b0000000011111111 : node3506;
															assign node3506 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3511 = (inp[2]) ? node3513 : 16'b0000000011111111;
													assign node3513 = (inp[7]) ? 16'b0000000001111111 : node3514;
														assign node3514 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node3518 = (inp[14]) ? node3534 : node3519;
											assign node3519 = (inp[2]) ? node3531 : node3520;
												assign node3520 = (inp[0]) ? node3526 : node3521;
													assign node3521 = (inp[4]) ? 16'b0000000111111111 : node3522;
														assign node3522 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3526 = (inp[9]) ? node3528 : 16'b0000000011111111;
														assign node3528 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node3531 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3534 = (inp[7]) ? node3536 : 16'b0000000011111111;
												assign node3536 = (inp[0]) ? node3538 : 16'b0000000000011111;
													assign node3538 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node3541 = (inp[0]) ? node3623 : node3542;
								assign node3542 = (inp[1]) ? node3580 : node3543;
									assign node3543 = (inp[7]) ? node3557 : node3544;
										assign node3544 = (inp[9]) ? node3548 : node3545;
											assign node3545 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node3548 = (inp[5]) ? node3552 : node3549;
												assign node3549 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3552 = (inp[2]) ? node3554 : 16'b0000000111111111;
													assign node3554 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node3557 = (inp[5]) ? node3571 : node3558;
											assign node3558 = (inp[3]) ? node3566 : node3559;
												assign node3559 = (inp[15]) ? 16'b0000000111111111 : node3560;
													assign node3560 = (inp[4]) ? 16'b0000001111111111 : node3561;
														assign node3561 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3566 = (inp[4]) ? node3568 : 16'b0000000111111111;
													assign node3568 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3571 = (inp[2]) ? 16'b0000000001111111 : node3572;
												assign node3572 = (inp[9]) ? node3576 : node3573;
													assign node3573 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3576 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node3580 = (inp[3]) ? node3594 : node3581;
										assign node3581 = (inp[4]) ? node3589 : node3582;
											assign node3582 = (inp[15]) ? node3586 : node3583;
												assign node3583 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3586 = (inp[2]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node3589 = (inp[2]) ? 16'b0000000111111111 : node3590;
												assign node3590 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3594 = (inp[5]) ? node3604 : node3595;
											assign node3595 = (inp[14]) ? node3597 : 16'b0000000111111111;
												assign node3597 = (inp[7]) ? node3601 : node3598;
													assign node3598 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3601 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node3604 = (inp[9]) ? node3616 : node3605;
												assign node3605 = (inp[2]) ? node3613 : node3606;
													assign node3606 = (inp[7]) ? node3608 : 16'b0000000011111111;
														assign node3608 = (inp[15]) ? node3610 : 16'b0000000011111111;
															assign node3610 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3613 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3616 = (inp[4]) ? node3620 : node3617;
													assign node3617 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3620 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node3623 = (inp[14]) ? node3661 : node3624;
									assign node3624 = (inp[4]) ? node3642 : node3625;
										assign node3625 = (inp[2]) ? node3631 : node3626;
											assign node3626 = (inp[7]) ? 16'b0000000111111111 : node3627;
												assign node3627 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3631 = (inp[5]) ? node3637 : node3632;
												assign node3632 = (inp[1]) ? 16'b0000000011111111 : node3633;
													assign node3633 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3637 = (inp[15]) ? node3639 : 16'b0000000011111111;
													assign node3639 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3642 = (inp[2]) ? node3654 : node3643;
											assign node3643 = (inp[9]) ? node3647 : node3644;
												assign node3644 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3647 = (inp[7]) ? node3651 : node3648;
													assign node3648 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3651 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3654 = (inp[15]) ? 16'b0000000001111111 : node3655;
												assign node3655 = (inp[7]) ? node3657 : 16'b0000000001111111;
													assign node3657 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3661 = (inp[2]) ? node3689 : node3662;
										assign node3662 = (inp[7]) ? node3674 : node3663;
											assign node3663 = (inp[9]) ? node3669 : node3664;
												assign node3664 = (inp[5]) ? 16'b0000000011111111 : node3665;
													assign node3665 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node3669 = (inp[1]) ? 16'b0000000001111111 : node3670;
													assign node3670 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3674 = (inp[1]) ? node3684 : node3675;
												assign node3675 = (inp[15]) ? node3677 : 16'b0000000011111111;
													assign node3677 = (inp[5]) ? 16'b0000000000011111 : node3678;
														assign node3678 = (inp[4]) ? node3680 : 16'b0000000011111111;
															assign node3680 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3684 = (inp[9]) ? 16'b0000000000111111 : node3685;
													assign node3685 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3689 = (inp[9]) ? node3695 : node3690;
											assign node3690 = (inp[7]) ? node3692 : 16'b0000000001111111;
												assign node3692 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node3695 = (inp[4]) ? node3705 : node3696;
												assign node3696 = (inp[5]) ? 16'b0000000000111111 : node3697;
													assign node3697 = (inp[1]) ? node3699 : 16'b0000000000111111;
														assign node3699 = (inp[7]) ? node3701 : 16'b0000000000111111;
															assign node3701 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node3705 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000001111111;
					assign node3708 = (inp[2]) ? node4090 : node3709;
						assign node3709 = (inp[3]) ? node3893 : node3710;
							assign node3710 = (inp[5]) ? node3808 : node3711;
								assign node3711 = (inp[15]) ? node3743 : node3712;
									assign node3712 = (inp[8]) ? node3730 : node3713;
										assign node3713 = (inp[0]) ? node3721 : node3714;
											assign node3714 = (inp[7]) ? 16'b0000001111111111 : node3715;
												assign node3715 = (inp[4]) ? 16'b0000011111111111 : node3716;
													assign node3716 = (inp[1]) ? 16'b0000111111111111 : 16'b0001111111111111;
											assign node3721 = (inp[1]) ? node3727 : node3722;
												assign node3722 = (inp[14]) ? 16'b0000001111111111 : node3723;
													assign node3723 = (inp[9]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node3727 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node3730 = (inp[1]) ? node3732 : 16'b0000001111111111;
											assign node3732 = (inp[11]) ? node3740 : node3733;
												assign node3733 = (inp[7]) ? 16'b0000000111111111 : node3734;
													assign node3734 = (inp[9]) ? node3736 : 16'b0000001111111111;
														assign node3736 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3740 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node3743 = (inp[0]) ? node3777 : node3744;
										assign node3744 = (inp[8]) ? node3754 : node3745;
											assign node3745 = (inp[4]) ? node3751 : node3746;
												assign node3746 = (inp[1]) ? 16'b0000001111111111 : node3747;
													assign node3747 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node3751 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3754 = (inp[7]) ? node3762 : node3755;
												assign node3755 = (inp[11]) ? 16'b0000000111111111 : node3756;
													assign node3756 = (inp[14]) ? 16'b0000000111111111 : node3757;
														assign node3757 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3762 = (inp[1]) ? node3770 : node3763;
													assign node3763 = (inp[4]) ? 16'b0000000111111111 : node3764;
														assign node3764 = (inp[11]) ? 16'b0000000111111111 : node3765;
															assign node3765 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3770 = (inp[9]) ? 16'b0000000011111111 : node3771;
														assign node3771 = (inp[4]) ? node3773 : 16'b0000000111111111;
															assign node3773 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node3777 = (inp[11]) ? node3791 : node3778;
											assign node3778 = (inp[8]) ? node3788 : node3779;
												assign node3779 = (inp[1]) ? node3781 : 16'b0000000111111111;
													assign node3781 = (inp[14]) ? 16'b0000000011111111 : node3782;
														assign node3782 = (inp[7]) ? node3784 : 16'b0000000111111111;
															assign node3784 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3788 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3791 = (inp[1]) ? node3799 : node3792;
												assign node3792 = (inp[7]) ? node3794 : 16'b0000000111111111;
													assign node3794 = (inp[8]) ? 16'b0000000001111111 : node3795;
														assign node3795 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3799 = (inp[4]) ? node3801 : 16'b0000000011111111;
													assign node3801 = (inp[9]) ? node3803 : 16'b0000000011111111;
														assign node3803 = (inp[14]) ? 16'b0000000001111111 : node3804;
															assign node3804 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node3808 = (inp[8]) ? node3858 : node3809;
									assign node3809 = (inp[9]) ? node3833 : node3810;
										assign node3810 = (inp[11]) ? node3826 : node3811;
											assign node3811 = (inp[14]) ? node3821 : node3812;
												assign node3812 = (inp[0]) ? node3814 : 16'b0000011111111111;
													assign node3814 = (inp[1]) ? 16'b0000000111111111 : node3815;
														assign node3815 = (inp[4]) ? node3817 : 16'b0000011111111111;
															assign node3817 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3821 = (inp[15]) ? node3823 : 16'b0000001111111111;
													assign node3823 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3826 = (inp[7]) ? 16'b0000000011111111 : node3827;
												assign node3827 = (inp[1]) ? 16'b0000000111111111 : node3828;
													assign node3828 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node3833 = (inp[11]) ? node3849 : node3834;
											assign node3834 = (inp[0]) ? node3844 : node3835;
												assign node3835 = (inp[14]) ? node3839 : node3836;
													assign node3836 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3839 = (inp[4]) ? 16'b0000000111111111 : node3840;
														assign node3840 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3844 = (inp[15]) ? 16'b0000000001111111 : node3845;
													assign node3845 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3849 = (inp[7]) ? node3851 : 16'b0000000011111111;
												assign node3851 = (inp[14]) ? node3855 : node3852;
													assign node3852 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3855 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3858 = (inp[9]) ? node3880 : node3859;
										assign node3859 = (inp[4]) ? node3875 : node3860;
											assign node3860 = (inp[11]) ? node3866 : node3861;
												assign node3861 = (inp[15]) ? 16'b0000000011111111 : node3862;
													assign node3862 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3866 = (inp[1]) ? 16'b0000000011111111 : node3867;
													assign node3867 = (inp[7]) ? node3869 : 16'b0000000111111111;
														assign node3869 = (inp[15]) ? 16'b0000000001111111 : node3870;
															assign node3870 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3875 = (inp[11]) ? node3877 : 16'b0000000011111111;
												assign node3877 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3880 = (inp[15]) ? node3882 : 16'b0000000011111111;
											assign node3882 = (inp[0]) ? node3886 : node3883;
												assign node3883 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node3886 = (inp[7]) ? 16'b0000000000111111 : node3887;
													assign node3887 = (inp[14]) ? node3889 : 16'b0000000001111111;
														assign node3889 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node3893 = (inp[0]) ? node3983 : node3894;
								assign node3894 = (inp[7]) ? node3944 : node3895;
									assign node3895 = (inp[1]) ? node3917 : node3896;
										assign node3896 = (inp[4]) ? node3908 : node3897;
											assign node3897 = (inp[5]) ? 16'b0000011111111111 : node3898;
												assign node3898 = (inp[15]) ? node3904 : node3899;
													assign node3899 = (inp[9]) ? node3901 : 16'b0000111111111111;
														assign node3901 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3904 = (inp[14]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node3908 = (inp[8]) ? node3914 : node3909;
												assign node3909 = (inp[11]) ? node3911 : 16'b0000001111111111;
													assign node3911 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3914 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000001111111;
										assign node3917 = (inp[8]) ? node3927 : node3918;
											assign node3918 = (inp[15]) ? node3922 : node3919;
												assign node3919 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node3922 = (inp[9]) ? node3924 : 16'b0000000111111111;
													assign node3924 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3927 = (inp[11]) ? node3937 : node3928;
												assign node3928 = (inp[9]) ? node3930 : 16'b0000001111111111;
													assign node3930 = (inp[14]) ? 16'b0000000011111111 : node3931;
														assign node3931 = (inp[4]) ? node3933 : 16'b0000000111111111;
															assign node3933 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3937 = (inp[9]) ? node3939 : 16'b0000000011111111;
													assign node3939 = (inp[15]) ? 16'b0000000000111111 : node3940;
														assign node3940 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000001111111;
									assign node3944 = (inp[14]) ? node3966 : node3945;
										assign node3945 = (inp[15]) ? node3955 : node3946;
											assign node3946 = (inp[1]) ? node3948 : 16'b0000001111111111;
												assign node3948 = (inp[4]) ? node3950 : 16'b0000001111111111;
													assign node3950 = (inp[11]) ? 16'b0000000011111111 : node3951;
														assign node3951 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3955 = (inp[4]) ? node3963 : node3956;
												assign node3956 = (inp[11]) ? 16'b0000000111111111 : node3957;
													assign node3957 = (inp[8]) ? 16'b0000000011111111 : node3958;
														assign node3958 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3963 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3966 = (inp[5]) ? node3974 : node3967;
											assign node3967 = (inp[8]) ? node3971 : node3968;
												assign node3968 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3971 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node3974 = (inp[9]) ? node3980 : node3975;
												assign node3975 = (inp[11]) ? 16'b0000000001111111 : node3976;
													assign node3976 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3980 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
								assign node3983 = (inp[9]) ? node4033 : node3984;
									assign node3984 = (inp[8]) ? node4014 : node3985;
										assign node3985 = (inp[5]) ? node4005 : node3986;
											assign node3986 = (inp[7]) ? node3996 : node3987;
												assign node3987 = (inp[1]) ? node3991 : node3988;
													assign node3988 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3991 = (inp[15]) ? node3993 : 16'b0000001111111111;
														assign node3993 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3996 = (inp[15]) ? node3998 : 16'b0000000111111111;
													assign node3998 = (inp[1]) ? 16'b0000000011111111 : node3999;
														assign node3999 = (inp[14]) ? node4001 : 16'b0000000111111111;
															assign node4001 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4005 = (inp[7]) ? 16'b0000000001111111 : node4006;
												assign node4006 = (inp[1]) ? node4008 : 16'b0000000111111111;
													assign node4008 = (inp[15]) ? 16'b0000000011111111 : node4009;
														assign node4009 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4014 = (inp[11]) ? node4018 : node4015;
											assign node4015 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4018 = (inp[1]) ? node4024 : node4019;
												assign node4019 = (inp[5]) ? node4021 : 16'b0000000011111111;
													assign node4021 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4024 = (inp[7]) ? node4028 : node4025;
													assign node4025 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node4028 = (inp[15]) ? 16'b0000000000111111 : node4029;
														assign node4029 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node4033 = (inp[1]) ? node4059 : node4034;
										assign node4034 = (inp[4]) ? node4046 : node4035;
											assign node4035 = (inp[15]) ? node4043 : node4036;
												assign node4036 = (inp[7]) ? 16'b0000000011111111 : node4037;
													assign node4037 = (inp[11]) ? node4039 : 16'b0000000111111111;
														assign node4039 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4043 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node4046 = (inp[14]) ? node4050 : node4047;
												assign node4047 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4050 = (inp[5]) ? node4054 : node4051;
													assign node4051 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node4054 = (inp[8]) ? 16'b0000000000111111 : node4055;
														assign node4055 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node4059 = (inp[5]) ? node4071 : node4060;
											assign node4060 = (inp[11]) ? node4064 : node4061;
												assign node4061 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4064 = (inp[15]) ? node4066 : 16'b0000000001111111;
													assign node4066 = (inp[8]) ? 16'b0000000000111111 : node4067;
														assign node4067 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node4071 = (inp[14]) ? node4081 : node4072;
												assign node4072 = (inp[4]) ? node4074 : 16'b0000000001111111;
													assign node4074 = (inp[7]) ? 16'b0000000000111111 : node4075;
														assign node4075 = (inp[8]) ? 16'b0000000000111111 : node4076;
															assign node4076 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4081 = (inp[11]) ? node4083 : 16'b0000000000111111;
													assign node4083 = (inp[8]) ? 16'b0000000000011111 : node4084;
														assign node4084 = (inp[4]) ? 16'b0000000000011111 : node4085;
															assign node4085 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node4090 = (inp[7]) ? node4262 : node4091;
							assign node4091 = (inp[8]) ? node4193 : node4092;
								assign node4092 = (inp[4]) ? node4154 : node4093;
									assign node4093 = (inp[5]) ? node4129 : node4094;
										assign node4094 = (inp[9]) ? node4112 : node4095;
											assign node4095 = (inp[14]) ? node4105 : node4096;
												assign node4096 = (inp[15]) ? node4098 : 16'b0000011111111111;
													assign node4098 = (inp[11]) ? 16'b0000001111111111 : node4099;
														assign node4099 = (inp[1]) ? node4101 : 16'b0000011111111111;
															assign node4101 = (inp[0]) ? 16'b0000001111111111 : 16'b0000001111111111;
												assign node4105 = (inp[0]) ? 16'b0000000111111111 : node4106;
													assign node4106 = (inp[11]) ? node4108 : 16'b0000001111111111;
														assign node4108 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4112 = (inp[11]) ? node4120 : node4113;
												assign node4113 = (inp[15]) ? 16'b0000000111111111 : node4114;
													assign node4114 = (inp[14]) ? node4116 : 16'b0000011111111111;
														assign node4116 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4120 = (inp[3]) ? node4126 : node4121;
													assign node4121 = (inp[15]) ? node4123 : 16'b0000000111111111;
														assign node4123 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4126 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4129 = (inp[3]) ? node4145 : node4130;
											assign node4130 = (inp[14]) ? node4134 : node4131;
												assign node4131 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4134 = (inp[1]) ? node4140 : node4135;
													assign node4135 = (inp[0]) ? 16'b0000000011111111 : node4136;
														assign node4136 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4140 = (inp[0]) ? node4142 : 16'b0000000011111111;
														assign node4142 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4145 = (inp[14]) ? node4151 : node4146;
												assign node4146 = (inp[0]) ? 16'b0000000011111111 : node4147;
													assign node4147 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4151 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000001111111;
									assign node4154 = (inp[11]) ? node4174 : node4155;
										assign node4155 = (inp[0]) ? node4161 : node4156;
											assign node4156 = (inp[1]) ? node4158 : 16'b0000011111111111;
												assign node4158 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4161 = (inp[9]) ? node4167 : node4162;
												assign node4162 = (inp[15]) ? node4164 : 16'b0000000111111111;
													assign node4164 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4167 = (inp[5]) ? node4169 : 16'b0000000011111111;
													assign node4169 = (inp[3]) ? 16'b0000000001111111 : node4170;
														assign node4170 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4174 = (inp[9]) ? node4182 : node4175;
											assign node4175 = (inp[14]) ? node4177 : 16'b0000000011111111;
												assign node4177 = (inp[3]) ? 16'b0000000000111111 : node4178;
													assign node4178 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4182 = (inp[3]) ? node4186 : node4183;
												assign node4183 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4186 = (inp[14]) ? node4188 : 16'b0000000001111111;
													assign node4188 = (inp[5]) ? 16'b0000000000111111 : node4189;
														assign node4189 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node4193 = (inp[5]) ? node4229 : node4194;
									assign node4194 = (inp[0]) ? node4208 : node4195;
										assign node4195 = (inp[14]) ? node4203 : node4196;
											assign node4196 = (inp[9]) ? node4198 : 16'b0000000011111111;
												assign node4198 = (inp[15]) ? 16'b0000000111111111 : node4199;
													assign node4199 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4203 = (inp[3]) ? 16'b0000000001111111 : node4204;
												assign node4204 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node4208 = (inp[15]) ? node4220 : node4209;
											assign node4209 = (inp[3]) ? node4211 : 16'b0000000011111111;
												assign node4211 = (inp[11]) ? node4215 : node4212;
													assign node4212 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4215 = (inp[4]) ? 16'b0000000001111111 : node4216;
														assign node4216 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4220 = (inp[14]) ? node4226 : node4221;
												assign node4221 = (inp[4]) ? 16'b0000000001111111 : node4222;
													assign node4222 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4226 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node4229 = (inp[1]) ? node4241 : node4230;
										assign node4230 = (inp[4]) ? node4236 : node4231;
											assign node4231 = (inp[9]) ? node4233 : 16'b0000000011111111;
												assign node4233 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4236 = (inp[0]) ? 16'b0000000000111111 : node4237;
												assign node4237 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4241 = (inp[3]) ? node4249 : node4242;
											assign node4242 = (inp[15]) ? 16'b0000000000111111 : node4243;
												assign node4243 = (inp[4]) ? 16'b0000000011111111 : node4244;
													assign node4244 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4249 = (inp[11]) ? node4255 : node4250;
												assign node4250 = (inp[9]) ? 16'b0000000000111111 : node4251;
													assign node4251 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4255 = (inp[15]) ? 16'b0000000000011111 : node4256;
													assign node4256 = (inp[14]) ? 16'b0000000000111111 : node4257;
														assign node4257 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node4262 = (inp[1]) ? node4354 : node4263;
								assign node4263 = (inp[15]) ? node4317 : node4264;
									assign node4264 = (inp[4]) ? node4294 : node4265;
										assign node4265 = (inp[8]) ? node4279 : node4266;
											assign node4266 = (inp[9]) ? node4270 : node4267;
												assign node4267 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4270 = (inp[0]) ? node4276 : node4271;
													assign node4271 = (inp[5]) ? node4273 : 16'b0000000111111111;
														assign node4273 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4276 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4279 = (inp[11]) ? node4287 : node4280;
												assign node4280 = (inp[5]) ? node4282 : 16'b0000000111111111;
													assign node4282 = (inp[9]) ? 16'b0000000011111111 : node4283;
														assign node4283 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4287 = (inp[9]) ? node4291 : node4288;
													assign node4288 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4291 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000001111111;
										assign node4294 = (inp[5]) ? node4306 : node4295;
											assign node4295 = (inp[14]) ? node4301 : node4296;
												assign node4296 = (inp[8]) ? node4298 : 16'b0000000111111111;
													assign node4298 = (inp[9]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node4301 = (inp[8]) ? node4303 : 16'b0000000011111111;
													assign node4303 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000111111111;
											assign node4306 = (inp[11]) ? node4312 : node4307;
												assign node4307 = (inp[3]) ? node4309 : 16'b0000000011111111;
													assign node4309 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4312 = (inp[14]) ? node4314 : 16'b0000000000111111;
													assign node4314 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node4317 = (inp[5]) ? node4333 : node4318;
										assign node4318 = (inp[3]) ? node4328 : node4319;
											assign node4319 = (inp[14]) ? node4325 : node4320;
												assign node4320 = (inp[11]) ? 16'b0000000111111111 : node4321;
													assign node4321 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4325 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node4328 = (inp[0]) ? 16'b0000000001111111 : node4329;
												assign node4329 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000000111111;
										assign node4333 = (inp[8]) ? node4343 : node4334;
											assign node4334 = (inp[14]) ? node4338 : node4335;
												assign node4335 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4338 = (inp[3]) ? node4340 : 16'b0000000001111111;
													assign node4340 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node4343 = (inp[9]) ? node4347 : node4344;
												assign node4344 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4347 = (inp[11]) ? 16'b0000000000011111 : node4348;
													assign node4348 = (inp[0]) ? node4350 : 16'b0000000000111111;
														assign node4350 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node4354 = (inp[0]) ? node4398 : node4355;
									assign node4355 = (inp[4]) ? node4375 : node4356;
										assign node4356 = (inp[5]) ? node4366 : node4357;
											assign node4357 = (inp[11]) ? node4363 : node4358;
												assign node4358 = (inp[3]) ? node4360 : 16'b0000000111111111;
													assign node4360 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4363 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node4366 = (inp[9]) ? node4370 : node4367;
												assign node4367 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4370 = (inp[15]) ? node4372 : 16'b0000000001111111;
													assign node4372 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node4375 = (inp[11]) ? node4385 : node4376;
											assign node4376 = (inp[15]) ? 16'b0000000001111111 : node4377;
												assign node4377 = (inp[5]) ? 16'b0000000000011111 : node4378;
													assign node4378 = (inp[3]) ? node4380 : 16'b0000000011111111;
														assign node4380 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4385 = (inp[14]) ? node4393 : node4386;
												assign node4386 = (inp[3]) ? 16'b0000000000111111 : node4387;
													assign node4387 = (inp[9]) ? node4389 : 16'b0000000011111111;
														assign node4389 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4393 = (inp[3]) ? 16'b0000000000001111 : node4394;
													assign node4394 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node4398 = (inp[3]) ? node4418 : node4399;
										assign node4399 = (inp[15]) ? node4405 : node4400;
											assign node4400 = (inp[5]) ? 16'b0000000000111111 : node4401;
												assign node4401 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4405 = (inp[11]) ? node4407 : 16'b0000000000111111;
												assign node4407 = (inp[9]) ? 16'b0000000000011111 : node4408;
													assign node4408 = (inp[5]) ? node4414 : node4409;
														assign node4409 = (inp[8]) ? 16'b0000000000111111 : node4410;
															assign node4410 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node4414 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node4418 = (inp[9]) ? node4432 : node4419;
											assign node4419 = (inp[5]) ? node4423 : node4420;
												assign node4420 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4423 = (inp[8]) ? node4429 : node4424;
													assign node4424 = (inp[11]) ? node4426 : 16'b0000000000111111;
														assign node4426 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node4429 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node4432 = (inp[14]) ? node4442 : node4433;
												assign node4433 = (inp[11]) ? node4437 : node4434;
													assign node4434 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node4437 = (inp[15]) ? node4439 : 16'b0000000000011111;
														assign node4439 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node4442 = (inp[4]) ? node4446 : node4443;
													assign node4443 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node4446 = (inp[11]) ? node4448 : 16'b0000000000001111;
														assign node4448 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
				assign node4451 = (inp[1]) ? node5171 : node4452;
					assign node4452 = (inp[5]) ? node4830 : node4453;
						assign node4453 = (inp[4]) ? node4649 : node4454;
							assign node4454 = (inp[7]) ? node4554 : node4455;
								assign node4455 = (inp[13]) ? node4509 : node4456;
									assign node4456 = (inp[8]) ? node4482 : node4457;
										assign node4457 = (inp[3]) ? node4467 : node4458;
											assign node4458 = (inp[11]) ? 16'b0000011111111111 : node4459;
												assign node4459 = (inp[9]) ? 16'b0000011111111111 : node4460;
													assign node4460 = (inp[14]) ? node4462 : 16'b0001111111111111;
														assign node4462 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node4467 = (inp[15]) ? node4477 : node4468;
												assign node4468 = (inp[0]) ? node4474 : node4469;
													assign node4469 = (inp[11]) ? 16'b0000011111111111 : node4470;
														assign node4470 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4474 = (inp[2]) ? 16'b0000011111111111 : 16'b0000001111111111;
												assign node4477 = (inp[9]) ? 16'b0000000111111111 : node4478;
													assign node4478 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node4482 = (inp[0]) ? node4496 : node4483;
											assign node4483 = (inp[11]) ? node4493 : node4484;
												assign node4484 = (inp[2]) ? node4486 : 16'b0000111111111111;
													assign node4486 = (inp[3]) ? 16'b0000001111111111 : node4487;
														assign node4487 = (inp[14]) ? node4489 : 16'b0000111111111111;
															assign node4489 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4493 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4496 = (inp[14]) ? 16'b0000000011111111 : node4497;
												assign node4497 = (inp[9]) ? node4503 : node4498;
													assign node4498 = (inp[15]) ? 16'b0000001111111111 : node4499;
														assign node4499 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4503 = (inp[2]) ? node4505 : 16'b0000000111111111;
														assign node4505 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node4509 = (inp[14]) ? node4529 : node4510;
										assign node4510 = (inp[9]) ? node4518 : node4511;
											assign node4511 = (inp[0]) ? node4515 : node4512;
												assign node4512 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node4515 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4518 = (inp[11]) ? node4524 : node4519;
												assign node4519 = (inp[2]) ? 16'b0000000111111111 : node4520;
													assign node4520 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4524 = (inp[15]) ? 16'b0000000011111111 : node4525;
													assign node4525 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4529 = (inp[11]) ? node4543 : node4530;
											assign node4530 = (inp[9]) ? node4538 : node4531;
												assign node4531 = (inp[8]) ? node4533 : 16'b0000001111111111;
													assign node4533 = (inp[3]) ? node4535 : 16'b0000000111111111;
														assign node4535 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node4538 = (inp[2]) ? 16'b0000000011111111 : node4539;
													assign node4539 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node4543 = (inp[9]) ? 16'b0000000111111111 : node4544;
												assign node4544 = (inp[15]) ? node4546 : 16'b0000000011111111;
													assign node4546 = (inp[2]) ? node4548 : 16'b0000000011111111;
														assign node4548 = (inp[3]) ? 16'b0000000001111111 : node4549;
															assign node4549 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node4554 = (inp[8]) ? node4606 : node4555;
									assign node4555 = (inp[9]) ? node4581 : node4556;
										assign node4556 = (inp[0]) ? node4568 : node4557;
											assign node4557 = (inp[2]) ? node4565 : node4558;
												assign node4558 = (inp[14]) ? node4560 : 16'b0000111111111111;
													assign node4560 = (inp[15]) ? node4562 : 16'b0000001111111111;
														assign node4562 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4565 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4568 = (inp[14]) ? node4572 : node4569;
												assign node4569 = (inp[15]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node4572 = (inp[3]) ? node4576 : node4573;
													assign node4573 = (inp[11]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node4576 = (inp[15]) ? node4578 : 16'b0000000111111111;
														assign node4578 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4581 = (inp[15]) ? node4593 : node4582;
											assign node4582 = (inp[13]) ? node4588 : node4583;
												assign node4583 = (inp[0]) ? 16'b0000000111111111 : node4584;
													assign node4584 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4588 = (inp[11]) ? node4590 : 16'b0000000111111111;
													assign node4590 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4593 = (inp[11]) ? node4601 : node4594;
												assign node4594 = (inp[3]) ? node4596 : 16'b0000000111111111;
													assign node4596 = (inp[0]) ? 16'b0000000011111111 : node4597;
														assign node4597 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4601 = (inp[2]) ? node4603 : 16'b0000000011111111;
													assign node4603 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node4606 = (inp[2]) ? node4628 : node4607;
										assign node4607 = (inp[9]) ? node4619 : node4608;
											assign node4608 = (inp[0]) ? node4614 : node4609;
												assign node4609 = (inp[11]) ? node4611 : 16'b0000011111111111;
													assign node4611 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4614 = (inp[13]) ? node4616 : 16'b0000000111111111;
													assign node4616 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node4619 = (inp[15]) ? node4621 : 16'b0000000111111111;
												assign node4621 = (inp[3]) ? 16'b0000000001111111 : node4622;
													assign node4622 = (inp[14]) ? 16'b0000000011111111 : node4623;
														assign node4623 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4628 = (inp[0]) ? node4640 : node4629;
											assign node4629 = (inp[13]) ? node4635 : node4630;
												assign node4630 = (inp[15]) ? 16'b0000000011111111 : node4631;
													assign node4631 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4635 = (inp[9]) ? 16'b0000000000111111 : node4636;
													assign node4636 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4640 = (inp[14]) ? node4644 : node4641;
												assign node4641 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node4644 = (inp[9]) ? 16'b0000000000011111 : node4645;
													assign node4645 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node4649 = (inp[2]) ? node4731 : node4650;
								assign node4650 = (inp[11]) ? node4682 : node4651;
									assign node4651 = (inp[3]) ? node4671 : node4652;
										assign node4652 = (inp[0]) ? node4660 : node4653;
											assign node4653 = (inp[14]) ? node4657 : node4654;
												assign node4654 = (inp[13]) ? 16'b0000011111111111 : 16'b0000001111111111;
												assign node4657 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4660 = (inp[15]) ? node4664 : node4661;
												assign node4661 = (inp[8]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node4664 = (inp[9]) ? 16'b0000000011111111 : node4665;
													assign node4665 = (inp[8]) ? node4667 : 16'b0000000111111111;
														assign node4667 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4671 = (inp[15]) ? node4677 : node4672;
											assign node4672 = (inp[7]) ? 16'b0000000111111111 : node4673;
												assign node4673 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4677 = (inp[7]) ? 16'b0000000001111111 : node4678;
												assign node4678 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node4682 = (inp[9]) ? node4700 : node4683;
										assign node4683 = (inp[7]) ? node4693 : node4684;
											assign node4684 = (inp[15]) ? 16'b0000000011111111 : node4685;
												assign node4685 = (inp[3]) ? node4687 : 16'b0000001111111111;
													assign node4687 = (inp[14]) ? 16'b0000000111111111 : node4688;
														assign node4688 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4693 = (inp[13]) ? node4697 : node4694;
												assign node4694 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4697 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4700 = (inp[8]) ? node4716 : node4701;
											assign node4701 = (inp[14]) ? node4709 : node4702;
												assign node4702 = (inp[13]) ? node4704 : 16'b0000000111111111;
													assign node4704 = (inp[3]) ? 16'b0000000011111111 : node4705;
														assign node4705 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4709 = (inp[15]) ? 16'b0000000011111111 : node4710;
													assign node4710 = (inp[3]) ? node4712 : 16'b0000000011111111;
														assign node4712 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4716 = (inp[13]) ? node4722 : node4717;
												assign node4717 = (inp[0]) ? node4719 : 16'b0000000111111111;
													assign node4719 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4722 = (inp[0]) ? node4728 : node4723;
													assign node4723 = (inp[15]) ? 16'b0000000001111111 : node4724;
														assign node4724 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4728 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000011111;
								assign node4731 = (inp[13]) ? node4771 : node4732;
									assign node4732 = (inp[0]) ? node4748 : node4733;
										assign node4733 = (inp[3]) ? node4743 : node4734;
											assign node4734 = (inp[9]) ? node4738 : node4735;
												assign node4735 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4738 = (inp[8]) ? 16'b0000000011111111 : node4739;
													assign node4739 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4743 = (inp[9]) ? 16'b0000000011111111 : node4744;
												assign node4744 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4748 = (inp[11]) ? node4766 : node4749;
											assign node4749 = (inp[14]) ? node4759 : node4750;
												assign node4750 = (inp[3]) ? node4756 : node4751;
													assign node4751 = (inp[9]) ? 16'b0000000011111111 : node4752;
														assign node4752 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4756 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4759 = (inp[15]) ? node4763 : node4760;
													assign node4760 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4763 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node4766 = (inp[7]) ? node4768 : 16'b0000000001111111;
												assign node4768 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node4771 = (inp[15]) ? node4799 : node4772;
										assign node4772 = (inp[11]) ? node4782 : node4773;
											assign node4773 = (inp[9]) ? node4779 : node4774;
												assign node4774 = (inp[0]) ? node4776 : 16'b0000011111111111;
													assign node4776 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4779 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4782 = (inp[9]) ? node4794 : node4783;
												assign node4783 = (inp[8]) ? node4789 : node4784;
													assign node4784 = (inp[7]) ? node4786 : 16'b0000001111111111;
														assign node4786 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4789 = (inp[7]) ? node4791 : 16'b0000000001111111;
														assign node4791 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node4794 = (inp[8]) ? 16'b0000000000111111 : node4795;
													assign node4795 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node4799 = (inp[7]) ? node4815 : node4800;
											assign node4800 = (inp[9]) ? node4804 : node4801;
												assign node4801 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node4804 = (inp[3]) ? node4812 : node4805;
													assign node4805 = (inp[11]) ? node4807 : 16'b0000000001111111;
														assign node4807 = (inp[8]) ? 16'b0000000000111111 : node4808;
															assign node4808 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node4812 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node4815 = (inp[8]) ? node4819 : node4816;
												assign node4816 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4819 = (inp[9]) ? node4825 : node4820;
													assign node4820 = (inp[0]) ? 16'b0000000000011111 : node4821;
														assign node4821 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node4825 = (inp[3]) ? node4827 : 16'b0000000000011111;
														assign node4827 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000011111;
						assign node4830 = (inp[3]) ? node5008 : node4831;
							assign node4831 = (inp[2]) ? node4921 : node4832;
								assign node4832 = (inp[15]) ? node4868 : node4833;
									assign node4833 = (inp[4]) ? node4851 : node4834;
										assign node4834 = (inp[14]) ? node4842 : node4835;
											assign node4835 = (inp[9]) ? node4837 : 16'b0000011111111111;
												assign node4837 = (inp[8]) ? node4839 : 16'b0000001111111111;
													assign node4839 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4842 = (inp[7]) ? node4848 : node4843;
												assign node4843 = (inp[9]) ? 16'b0000000111111111 : node4844;
													assign node4844 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4848 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node4851 = (inp[14]) ? node4863 : node4852;
											assign node4852 = (inp[9]) ? node4858 : node4853;
												assign node4853 = (inp[8]) ? 16'b0000000111111111 : node4854;
													assign node4854 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4858 = (inp[7]) ? 16'b0000000001111111 : node4859;
													assign node4859 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node4863 = (inp[13]) ? 16'b0000000001111111 : node4864;
												assign node4864 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node4868 = (inp[8]) ? node4886 : node4869;
										assign node4869 = (inp[0]) ? node4875 : node4870;
											assign node4870 = (inp[14]) ? 16'b0000000111111111 : node4871;
												assign node4871 = (inp[7]) ? 16'b0000000111111111 : 16'b0000011111111111;
											assign node4875 = (inp[11]) ? node4883 : node4876;
												assign node4876 = (inp[9]) ? node4878 : 16'b0000000111111111;
													assign node4878 = (inp[14]) ? 16'b0000000011111111 : node4879;
														assign node4879 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4883 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4886 = (inp[4]) ? node4902 : node4887;
											assign node4887 = (inp[14]) ? node4895 : node4888;
												assign node4888 = (inp[7]) ? 16'b0000000011111111 : node4889;
													assign node4889 = (inp[0]) ? node4891 : 16'b0000000111111111;
														assign node4891 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4895 = (inp[13]) ? node4897 : 16'b0000000011111111;
													assign node4897 = (inp[7]) ? 16'b0000000001111111 : node4898;
														assign node4898 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4902 = (inp[14]) ? node4916 : node4903;
												assign node4903 = (inp[11]) ? node4909 : node4904;
													assign node4904 = (inp[13]) ? node4906 : 16'b0000000011111111;
														assign node4906 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4909 = (inp[9]) ? node4913 : node4910;
														assign node4910 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node4913 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4916 = (inp[11]) ? 16'b0000000000111111 : node4917;
													assign node4917 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000000111111;
								assign node4921 = (inp[13]) ? node4959 : node4922;
									assign node4922 = (inp[11]) ? node4946 : node4923;
										assign node4923 = (inp[14]) ? node4933 : node4924;
											assign node4924 = (inp[15]) ? node4930 : node4925;
												assign node4925 = (inp[9]) ? 16'b0000000111111111 : node4926;
													assign node4926 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4930 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4933 = (inp[9]) ? node4939 : node4934;
												assign node4934 = (inp[15]) ? 16'b0000000011111111 : node4935;
													assign node4935 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4939 = (inp[4]) ? node4943 : node4940;
													assign node4940 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node4943 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node4946 = (inp[8]) ? node4954 : node4947;
											assign node4947 = (inp[4]) ? node4951 : node4948;
												assign node4948 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4951 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4954 = (inp[15]) ? 16'b0000000001111111 : node4955;
												assign node4955 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000001111111;
									assign node4959 = (inp[15]) ? node4985 : node4960;
										assign node4960 = (inp[7]) ? node4968 : node4961;
											assign node4961 = (inp[9]) ? 16'b0000000011111111 : node4962;
												assign node4962 = (inp[11]) ? node4964 : 16'b0000000111111111;
													assign node4964 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4968 = (inp[0]) ? node4976 : node4969;
												assign node4969 = (inp[9]) ? 16'b0000000001111111 : node4970;
													assign node4970 = (inp[4]) ? 16'b0000000001111111 : node4971;
														assign node4971 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4976 = (inp[8]) ? node4980 : node4977;
													assign node4977 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4980 = (inp[9]) ? node4982 : 16'b0000000000111111;
														assign node4982 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node4985 = (inp[4]) ? node4999 : node4986;
											assign node4986 = (inp[11]) ? node4992 : node4987;
												assign node4987 = (inp[8]) ? node4989 : 16'b0000000011111111;
													assign node4989 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4992 = (inp[8]) ? 16'b0000000000011111 : node4993;
													assign node4993 = (inp[7]) ? node4995 : 16'b0000000001111111;
														assign node4995 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node4999 = (inp[11]) ? node5001 : 16'b0000000000111111;
												assign node5001 = (inp[14]) ? node5003 : 16'b0000000000111111;
													assign node5003 = (inp[9]) ? 16'b0000000000011111 : node5004;
														assign node5004 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node5008 = (inp[8]) ? node5086 : node5009;
								assign node5009 = (inp[15]) ? node5041 : node5010;
									assign node5010 = (inp[13]) ? node5022 : node5011;
										assign node5011 = (inp[4]) ? node5017 : node5012;
											assign node5012 = (inp[2]) ? 16'b0000000111111111 : node5013;
												assign node5013 = (inp[11]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node5017 = (inp[7]) ? 16'b0000000011111111 : node5018;
												assign node5018 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node5022 = (inp[0]) ? node5030 : node5023;
											assign node5023 = (inp[7]) ? 16'b0000000011111111 : node5024;
												assign node5024 = (inp[2]) ? node5026 : 16'b0000000111111111;
													assign node5026 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node5030 = (inp[7]) ? node5034 : node5031;
												assign node5031 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5034 = (inp[2]) ? node5036 : 16'b0000000000111111;
													assign node5036 = (inp[9]) ? node5038 : 16'b0000000001111111;
														assign node5038 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node5041 = (inp[4]) ? node5065 : node5042;
										assign node5042 = (inp[14]) ? node5056 : node5043;
											assign node5043 = (inp[7]) ? node5051 : node5044;
												assign node5044 = (inp[9]) ? node5046 : 16'b0000001111111111;
													assign node5046 = (inp[11]) ? 16'b0000000011111111 : node5047;
														assign node5047 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node5051 = (inp[9]) ? node5053 : 16'b0000000011111111;
													assign node5053 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5056 = (inp[0]) ? node5062 : node5057;
												assign node5057 = (inp[11]) ? 16'b0000000001111111 : node5058;
													assign node5058 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5062 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5065 = (inp[11]) ? node5075 : node5066;
											assign node5066 = (inp[13]) ? node5068 : 16'b0000000001111111;
												assign node5068 = (inp[9]) ? 16'b0000000000111111 : node5069;
													assign node5069 = (inp[7]) ? node5071 : 16'b0000000111111111;
														assign node5071 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node5075 = (inp[7]) ? node5077 : 16'b0000000001111111;
												assign node5077 = (inp[13]) ? node5083 : node5078;
													assign node5078 = (inp[2]) ? node5080 : 16'b0000000001111111;
														assign node5080 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node5083 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node5086 = (inp[13]) ? node5130 : node5087;
									assign node5087 = (inp[11]) ? node5107 : node5088;
										assign node5088 = (inp[0]) ? node5094 : node5089;
											assign node5089 = (inp[2]) ? node5091 : 16'b0000000111111111;
												assign node5091 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5094 = (inp[7]) ? node5102 : node5095;
												assign node5095 = (inp[4]) ? node5099 : node5096;
													assign node5096 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node5099 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node5102 = (inp[9]) ? 16'b0000000000001111 : node5103;
													assign node5103 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5107 = (inp[14]) ? node5121 : node5108;
											assign node5108 = (inp[0]) ? node5112 : node5109;
												assign node5109 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5112 = (inp[7]) ? node5114 : 16'b0000000011111111;
													assign node5114 = (inp[9]) ? node5118 : node5115;
														assign node5115 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5118 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node5121 = (inp[2]) ? node5125 : node5122;
												assign node5122 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5125 = (inp[4]) ? 16'b0000000000011111 : node5126;
													assign node5126 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node5130 = (inp[9]) ? node5150 : node5131;
										assign node5131 = (inp[15]) ? node5137 : node5132;
											assign node5132 = (inp[14]) ? 16'b0000000000011111 : node5133;
												assign node5133 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5137 = (inp[4]) ? node5145 : node5138;
												assign node5138 = (inp[7]) ? 16'b0000000000011111 : node5139;
													assign node5139 = (inp[11]) ? node5141 : 16'b0000000001111111;
														assign node5141 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5145 = (inp[0]) ? node5147 : 16'b0000000000011111;
													assign node5147 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node5150 = (inp[2]) ? node5160 : node5151;
											assign node5151 = (inp[15]) ? node5153 : 16'b0000000000111111;
												assign node5153 = (inp[7]) ? 16'b0000000000001111 : node5154;
													assign node5154 = (inp[11]) ? 16'b0000000000011111 : node5155;
														assign node5155 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node5160 = (inp[14]) ? node5168 : node5161;
												assign node5161 = (inp[15]) ? node5163 : 16'b0000000000011111;
													assign node5163 = (inp[0]) ? node5165 : 16'b0000000000011111;
														assign node5165 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node5168 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000011111;
					assign node5171 = (inp[11]) ? node5535 : node5172;
						assign node5172 = (inp[15]) ? node5346 : node5173;
							assign node5173 = (inp[14]) ? node5259 : node5174;
								assign node5174 = (inp[7]) ? node5216 : node5175;
									assign node5175 = (inp[4]) ? node5195 : node5176;
										assign node5176 = (inp[8]) ? node5186 : node5177;
											assign node5177 = (inp[13]) ? node5181 : node5178;
												assign node5178 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5181 = (inp[2]) ? node5183 : 16'b0000001111111111;
													assign node5183 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node5186 = (inp[2]) ? node5190 : node5187;
												assign node5187 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5190 = (inp[9]) ? node5192 : 16'b0000000111111111;
													assign node5192 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node5195 = (inp[2]) ? node5209 : node5196;
											assign node5196 = (inp[13]) ? node5204 : node5197;
												assign node5197 = (inp[3]) ? 16'b0000000011111111 : node5198;
													assign node5198 = (inp[8]) ? 16'b0000001111111111 : node5199;
														assign node5199 = (inp[0]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node5204 = (inp[8]) ? node5206 : 16'b0000000111111111;
													assign node5206 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node5209 = (inp[0]) ? node5213 : node5210;
												assign node5210 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5213 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node5216 = (inp[5]) ? node5232 : node5217;
										assign node5217 = (inp[8]) ? node5223 : node5218;
											assign node5218 = (inp[9]) ? node5220 : 16'b0000001111111111;
												assign node5220 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5223 = (inp[0]) ? node5225 : 16'b0000000011111111;
												assign node5225 = (inp[2]) ? 16'b0000000001111111 : node5226;
													assign node5226 = (inp[3]) ? node5228 : 16'b0000000111111111;
														assign node5228 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5232 = (inp[13]) ? node5244 : node5233;
											assign node5233 = (inp[9]) ? node5237 : node5234;
												assign node5234 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5237 = (inp[0]) ? node5239 : 16'b0000000011111111;
													assign node5239 = (inp[2]) ? 16'b0000000000111111 : node5240;
														assign node5240 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5244 = (inp[0]) ? node5256 : node5245;
												assign node5245 = (inp[3]) ? node5251 : node5246;
													assign node5246 = (inp[4]) ? node5248 : 16'b0000000001111111;
														assign node5248 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5251 = (inp[4]) ? node5253 : 16'b0000000001111111;
														assign node5253 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5256 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000011111;
								assign node5259 = (inp[5]) ? node5283 : node5260;
									assign node5260 = (inp[4]) ? node5276 : node5261;
										assign node5261 = (inp[8]) ? node5269 : node5262;
											assign node5262 = (inp[13]) ? node5264 : 16'b0000000111111111;
												assign node5264 = (inp[9]) ? 16'b0000000011111111 : node5265;
													assign node5265 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5269 = (inp[0]) ? node5273 : node5270;
												assign node5270 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5273 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000000111111;
										assign node5276 = (inp[2]) ? 16'b0000000001111111 : node5277;
											assign node5277 = (inp[3]) ? 16'b0000000011111111 : node5278;
												assign node5278 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node5283 = (inp[13]) ? node5313 : node5284;
										assign node5284 = (inp[2]) ? node5296 : node5285;
											assign node5285 = (inp[9]) ? node5287 : 16'b0000000111111111;
												assign node5287 = (inp[7]) ? node5293 : node5288;
													assign node5288 = (inp[8]) ? node5290 : 16'b0000000011111111;
														assign node5290 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5293 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5296 = (inp[3]) ? node5304 : node5297;
												assign node5297 = (inp[4]) ? 16'b0000000001111111 : node5298;
													assign node5298 = (inp[9]) ? node5300 : 16'b0000000111111111;
														assign node5300 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5304 = (inp[9]) ? node5306 : 16'b0000000011111111;
													assign node5306 = (inp[4]) ? node5310 : node5307;
														assign node5307 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5310 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node5313 = (inp[7]) ? node5327 : node5314;
											assign node5314 = (inp[3]) ? node5324 : node5315;
												assign node5315 = (inp[8]) ? 16'b0000000001111111 : node5316;
													assign node5316 = (inp[2]) ? node5318 : 16'b0000000011111111;
														assign node5318 = (inp[0]) ? 16'b0000000001111111 : node5319;
															assign node5319 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5324 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5327 = (inp[0]) ? node5335 : node5328;
												assign node5328 = (inp[4]) ? node5332 : node5329;
													assign node5329 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5332 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5335 = (inp[3]) ? node5343 : node5336;
													assign node5336 = (inp[9]) ? node5340 : node5337;
														assign node5337 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5340 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node5343 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node5346 = (inp[2]) ? node5438 : node5347;
								assign node5347 = (inp[9]) ? node5395 : node5348;
									assign node5348 = (inp[3]) ? node5366 : node5349;
										assign node5349 = (inp[0]) ? node5363 : node5350;
											assign node5350 = (inp[13]) ? node5358 : node5351;
												assign node5351 = (inp[7]) ? 16'b0000000111111111 : node5352;
													assign node5352 = (inp[5]) ? 16'b0000001111111111 : node5353;
														assign node5353 = (inp[8]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node5358 = (inp[7]) ? 16'b0000000111111111 : node5359;
													assign node5359 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5363 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5366 = (inp[7]) ? node5386 : node5367;
											assign node5367 = (inp[4]) ? node5381 : node5368;
												assign node5368 = (inp[14]) ? node5372 : node5369;
													assign node5369 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5372 = (inp[13]) ? node5378 : node5373;
														assign node5373 = (inp[0]) ? node5375 : 16'b0000000111111111;
															assign node5375 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5378 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5381 = (inp[13]) ? 16'b0000000001111111 : node5382;
													assign node5382 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5386 = (inp[5]) ? node5390 : node5387;
												assign node5387 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5390 = (inp[4]) ? node5392 : 16'b0000000000111111;
													assign node5392 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node5395 = (inp[7]) ? node5419 : node5396;
										assign node5396 = (inp[4]) ? node5402 : node5397;
											assign node5397 = (inp[8]) ? 16'b0000000011111111 : node5398;
												assign node5398 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5402 = (inp[14]) ? node5410 : node5403;
												assign node5403 = (inp[0]) ? 16'b0000000001111111 : node5404;
													assign node5404 = (inp[8]) ? node5406 : 16'b0000000011111111;
														assign node5406 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5410 = (inp[13]) ? node5416 : node5411;
													assign node5411 = (inp[3]) ? node5413 : 16'b0000000001111111;
														assign node5413 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5416 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node5419 = (inp[5]) ? node5433 : node5420;
											assign node5420 = (inp[4]) ? node5424 : node5421;
												assign node5421 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5424 = (inp[0]) ? 16'b0000000000111111 : node5425;
													assign node5425 = (inp[8]) ? node5427 : 16'b0000000001111111;
														assign node5427 = (inp[3]) ? node5429 : 16'b0000000001111111;
															assign node5429 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5433 = (inp[3]) ? 16'b0000000000111111 : node5434;
												assign node5434 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node5438 = (inp[4]) ? node5496 : node5439;
									assign node5439 = (inp[13]) ? node5459 : node5440;
										assign node5440 = (inp[7]) ? node5452 : node5441;
											assign node5441 = (inp[14]) ? node5449 : node5442;
												assign node5442 = (inp[8]) ? 16'b0000000011111111 : node5443;
													assign node5443 = (inp[3]) ? 16'b0000000111111111 : node5444;
														assign node5444 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node5449 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node5452 = (inp[9]) ? node5456 : node5453;
												assign node5453 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node5456 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5459 = (inp[3]) ? node5471 : node5460;
											assign node5460 = (inp[7]) ? node5464 : node5461;
												assign node5461 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5464 = (inp[8]) ? node5466 : 16'b0000000001111111;
													assign node5466 = (inp[5]) ? 16'b0000000000111111 : node5467;
														assign node5467 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5471 = (inp[14]) ? node5483 : node5472;
												assign node5472 = (inp[7]) ? 16'b0000000000111111 : node5473;
													assign node5473 = (inp[0]) ? node5479 : node5474;
														assign node5474 = (inp[9]) ? node5476 : 16'b0000000001111111;
															assign node5476 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5479 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5483 = (inp[8]) ? node5487 : node5484;
													assign node5484 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5487 = (inp[0]) ? node5493 : node5488;
														assign node5488 = (inp[5]) ? node5490 : 16'b0000000000111111;
															assign node5490 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node5493 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node5496 = (inp[14]) ? node5518 : node5497;
										assign node5497 = (inp[5]) ? node5509 : node5498;
											assign node5498 = (inp[9]) ? node5504 : node5499;
												assign node5499 = (inp[13]) ? 16'b0000000001111111 : node5500;
													assign node5500 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5504 = (inp[7]) ? 16'b0000000000001111 : node5505;
													assign node5505 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5509 = (inp[13]) ? node5515 : node5510;
												assign node5510 = (inp[7]) ? 16'b0000000000111111 : node5511;
													assign node5511 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5515 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node5518 = (inp[7]) ? node5530 : node5519;
											assign node5519 = (inp[5]) ? node5527 : node5520;
												assign node5520 = (inp[0]) ? node5522 : 16'b0000000001111111;
													assign node5522 = (inp[9]) ? node5524 : 16'b0000000000111111;
														assign node5524 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node5527 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node5530 = (inp[8]) ? node5532 : 16'b0000000000011111;
												assign node5532 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node5535 = (inp[8]) ? node5723 : node5536;
							assign node5536 = (inp[5]) ? node5634 : node5537;
								assign node5537 = (inp[4]) ? node5581 : node5538;
									assign node5538 = (inp[2]) ? node5568 : node5539;
										assign node5539 = (inp[0]) ? node5559 : node5540;
											assign node5540 = (inp[14]) ? node5552 : node5541;
												assign node5541 = (inp[7]) ? node5549 : node5542;
													assign node5542 = (inp[3]) ? 16'b0000001111111111 : node5543;
														assign node5543 = (inp[9]) ? 16'b0000001111111111 : node5544;
															assign node5544 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node5549 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5552 = (inp[3]) ? node5556 : node5553;
													assign node5553 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5556 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5559 = (inp[15]) ? node5565 : node5560;
												assign node5560 = (inp[14]) ? node5562 : 16'b0000000111111111;
													assign node5562 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5565 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node5568 = (inp[14]) ? node5574 : node5569;
											assign node5569 = (inp[7]) ? node5571 : 16'b0000000111111111;
												assign node5571 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5574 = (inp[13]) ? node5578 : node5575;
												assign node5575 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5578 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node5581 = (inp[15]) ? node5613 : node5582;
										assign node5582 = (inp[14]) ? node5596 : node5583;
											assign node5583 = (inp[13]) ? node5591 : node5584;
												assign node5584 = (inp[0]) ? node5586 : 16'b0000000111111111;
													assign node5586 = (inp[9]) ? 16'b0000000011111111 : node5587;
														assign node5587 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5591 = (inp[7]) ? node5593 : 16'b0000000011111111;
													assign node5593 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5596 = (inp[9]) ? node5608 : node5597;
												assign node5597 = (inp[7]) ? 16'b0000000001111111 : node5598;
													assign node5598 = (inp[0]) ? node5604 : node5599;
														assign node5599 = (inp[13]) ? 16'b0000000011111111 : node5600;
															assign node5600 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5604 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5608 = (inp[2]) ? node5610 : 16'b0000000001111111;
													assign node5610 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000000011111;
										assign node5613 = (inp[7]) ? node5621 : node5614;
											assign node5614 = (inp[13]) ? node5616 : 16'b0000000001111111;
												assign node5616 = (inp[2]) ? node5618 : 16'b0000000001111111;
													assign node5618 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5621 = (inp[9]) ? node5625 : node5622;
												assign node5622 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5625 = (inp[0]) ? node5629 : node5626;
													assign node5626 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000000011111;
													assign node5629 = (inp[3]) ? node5631 : 16'b0000000000011111;
														assign node5631 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node5634 = (inp[7]) ? node5676 : node5635;
									assign node5635 = (inp[15]) ? node5657 : node5636;
										assign node5636 = (inp[3]) ? node5644 : node5637;
											assign node5637 = (inp[4]) ? node5641 : node5638;
												assign node5638 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5641 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5644 = (inp[14]) ? node5652 : node5645;
												assign node5645 = (inp[9]) ? 16'b0000000001111111 : node5646;
													assign node5646 = (inp[0]) ? 16'b0000000001111111 : node5647;
														assign node5647 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5652 = (inp[4]) ? 16'b0000000000011111 : node5653;
													assign node5653 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5657 = (inp[4]) ? node5673 : node5658;
											assign node5658 = (inp[14]) ? node5662 : node5659;
												assign node5659 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5662 = (inp[13]) ? node5664 : 16'b0000000001111111;
													assign node5664 = (inp[3]) ? node5668 : node5665;
														assign node5665 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5668 = (inp[2]) ? node5670 : 16'b0000000000111111;
															assign node5670 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node5673 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node5676 = (inp[4]) ? node5696 : node5677;
										assign node5677 = (inp[14]) ? node5685 : node5678;
											assign node5678 = (inp[13]) ? node5680 : 16'b0000000011111111;
												assign node5680 = (inp[3]) ? node5682 : 16'b0000000001111111;
													assign node5682 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5685 = (inp[13]) ? 16'b0000000000111111 : node5686;
												assign node5686 = (inp[3]) ? node5688 : 16'b0000000001111111;
													assign node5688 = (inp[15]) ? node5692 : node5689;
														assign node5689 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5692 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node5696 = (inp[13]) ? node5708 : node5697;
											assign node5697 = (inp[3]) ? node5703 : node5698;
												assign node5698 = (inp[15]) ? 16'b0000000000111111 : node5699;
													assign node5699 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5703 = (inp[9]) ? node5705 : 16'b0000000000111111;
													assign node5705 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node5708 = (inp[14]) ? node5716 : node5709;
												assign node5709 = (inp[0]) ? 16'b0000000000011111 : node5710;
													assign node5710 = (inp[3]) ? node5712 : 16'b0000000001111111;
														assign node5712 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5716 = (inp[15]) ? 16'b0000000000001111 : node5717;
													assign node5717 = (inp[3]) ? node5719 : 16'b0000000000111111;
														assign node5719 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node5723 = (inp[0]) ? node5845 : node5724;
								assign node5724 = (inp[4]) ? node5786 : node5725;
									assign node5725 = (inp[7]) ? node5757 : node5726;
										assign node5726 = (inp[15]) ? node5736 : node5727;
											assign node5727 = (inp[9]) ? node5733 : node5728;
												assign node5728 = (inp[5]) ? 16'b0000000000111111 : node5729;
													assign node5729 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5733 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5736 = (inp[3]) ? node5744 : node5737;
												assign node5737 = (inp[5]) ? node5741 : node5738;
													assign node5738 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5741 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node5744 = (inp[2]) ? node5750 : node5745;
													assign node5745 = (inp[13]) ? 16'b0000000001111111 : node5746;
														assign node5746 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5750 = (inp[9]) ? node5754 : node5751;
														assign node5751 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5754 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node5757 = (inp[14]) ? node5777 : node5758;
											assign node5758 = (inp[3]) ? node5772 : node5759;
												assign node5759 = (inp[2]) ? node5767 : node5760;
													assign node5760 = (inp[15]) ? node5762 : 16'b0000000001111111;
														assign node5762 = (inp[9]) ? node5764 : 16'b0000000011111111;
															assign node5764 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5767 = (inp[15]) ? node5769 : 16'b0000000001111111;
														assign node5769 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5772 = (inp[2]) ? node5774 : 16'b0000000000111111;
													assign node5774 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5777 = (inp[3]) ? node5783 : node5778;
												assign node5778 = (inp[15]) ? 16'b0000000000111111 : node5779;
													assign node5779 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node5783 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node5786 = (inp[13]) ? node5820 : node5787;
										assign node5787 = (inp[7]) ? node5807 : node5788;
											assign node5788 = (inp[2]) ? node5798 : node5789;
												assign node5789 = (inp[9]) ? node5793 : node5790;
													assign node5790 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5793 = (inp[3]) ? node5795 : 16'b0000000001111111;
														assign node5795 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5798 = (inp[9]) ? 16'b0000000000111111 : node5799;
													assign node5799 = (inp[3]) ? node5801 : 16'b0000000001111111;
														assign node5801 = (inp[5]) ? 16'b0000000000111111 : node5802;
															assign node5802 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5807 = (inp[5]) ? node5813 : node5808;
												assign node5808 = (inp[15]) ? node5810 : 16'b0000000001111111;
													assign node5810 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5813 = (inp[2]) ? node5815 : 16'b0000000000111111;
													assign node5815 = (inp[9]) ? node5817 : 16'b0000000000011111;
														assign node5817 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node5820 = (inp[9]) ? node5834 : node5821;
											assign node5821 = (inp[15]) ? node5829 : node5822;
												assign node5822 = (inp[7]) ? node5824 : 16'b0000000011111111;
													assign node5824 = (inp[3]) ? node5826 : 16'b0000000000111111;
														assign node5826 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node5829 = (inp[2]) ? 16'b0000000000011111 : node5830;
													assign node5830 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node5834 = (inp[7]) ? node5842 : node5835;
												assign node5835 = (inp[14]) ? node5837 : 16'b0000000000111111;
													assign node5837 = (inp[5]) ? node5839 : 16'b0000000000011111;
														assign node5839 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000011111;
												assign node5842 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node5845 = (inp[3]) ? node5897 : node5846;
									assign node5846 = (inp[13]) ? node5872 : node5847;
										assign node5847 = (inp[4]) ? node5861 : node5848;
											assign node5848 = (inp[2]) ? node5856 : node5849;
												assign node5849 = (inp[9]) ? 16'b0000000001111111 : node5850;
													assign node5850 = (inp[14]) ? 16'b0000000011111111 : node5851;
														assign node5851 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5856 = (inp[15]) ? 16'b0000000000111111 : node5857;
													assign node5857 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5861 = (inp[5]) ? node5865 : node5862;
												assign node5862 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5865 = (inp[7]) ? node5867 : 16'b0000000011111111;
													assign node5867 = (inp[2]) ? node5869 : 16'b0000000000011111;
														assign node5869 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000011111;
										assign node5872 = (inp[5]) ? node5882 : node5873;
											assign node5873 = (inp[4]) ? node5879 : node5874;
												assign node5874 = (inp[14]) ? 16'b0000000000111111 : node5875;
													assign node5875 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5879 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node5882 = (inp[2]) ? node5890 : node5883;
												assign node5883 = (inp[9]) ? node5887 : node5884;
													assign node5884 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5887 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000000011111;
												assign node5890 = (inp[9]) ? node5894 : node5891;
													assign node5891 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node5894 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node5897 = (inp[7]) ? node5925 : node5898;
										assign node5898 = (inp[15]) ? node5912 : node5899;
											assign node5899 = (inp[14]) ? node5905 : node5900;
												assign node5900 = (inp[4]) ? 16'b0000000000111111 : node5901;
													assign node5901 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5905 = (inp[2]) ? node5907 : 16'b0000000000111111;
													assign node5907 = (inp[13]) ? 16'b0000000000011111 : node5908;
														assign node5908 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node5912 = (inp[5]) ? 16'b0000000000011111 : node5913;
												assign node5913 = (inp[9]) ? node5919 : node5914;
													assign node5914 = (inp[2]) ? node5916 : 16'b0000000000111111;
														assign node5916 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node5919 = (inp[13]) ? node5921 : 16'b0000000000011111;
														assign node5921 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node5925 = (inp[2]) ? node5941 : node5926;
											assign node5926 = (inp[5]) ? node5930 : node5927;
												assign node5927 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node5930 = (inp[14]) ? node5938 : node5931;
													assign node5931 = (inp[15]) ? node5935 : node5932;
														assign node5932 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node5935 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node5938 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node5941 = (inp[4]) ? node5951 : node5942;
												assign node5942 = (inp[13]) ? 16'b0000000000001111 : node5943;
													assign node5943 = (inp[14]) ? 16'b0000000000111111 : node5944;
														assign node5944 = (inp[5]) ? node5946 : 16'b0000000000011111;
															assign node5946 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node5951 = (inp[9]) ? node5957 : node5952;
													assign node5952 = (inp[14]) ? node5954 : 16'b0000000000001111;
														assign node5954 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node5957 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000000011;
		assign node5960 = (inp[2]) ? node8614 : node5961;
			assign node5961 = (inp[11]) ? node7343 : node5962;
				assign node5962 = (inp[4]) ? node6644 : node5963;
					assign node5963 = (inp[12]) ? node6317 : node5964;
						assign node5964 = (inp[1]) ? node6118 : node5965;
							assign node5965 = (inp[0]) ? node6037 : node5966;
								assign node5966 = (inp[9]) ? node6002 : node5967;
									assign node5967 = (inp[5]) ? node5987 : node5968;
										assign node5968 = (inp[13]) ? node5972 : node5969;
											assign node5969 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
											assign node5972 = (inp[8]) ? node5982 : node5973;
												assign node5973 = (inp[7]) ? node5975 : 16'b0000111111111111;
													assign node5975 = (inp[3]) ? node5979 : node5976;
														assign node5976 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node5979 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5982 = (inp[14]) ? node5984 : 16'b0000011111111111;
													assign node5984 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node5987 = (inp[10]) ? node5997 : node5988;
											assign node5988 = (inp[3]) ? node5992 : node5989;
												assign node5989 = (inp[15]) ? 16'b0000111111111111 : 16'b0000011111111111;
												assign node5992 = (inp[8]) ? node5994 : 16'b0000011111111111;
													assign node5994 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node5997 = (inp[7]) ? 16'b0000001111111111 : node5998;
												assign node5998 = (inp[13]) ? 16'b0000000111111111 : 16'b0000011111111111;
									assign node6002 = (inp[14]) ? node6018 : node6003;
										assign node6003 = (inp[13]) ? node6013 : node6004;
											assign node6004 = (inp[7]) ? 16'b0000011111111111 : node6005;
												assign node6005 = (inp[10]) ? node6007 : 16'b0000111111111111;
													assign node6007 = (inp[3]) ? 16'b0000011111111111 : node6008;
														assign node6008 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node6013 = (inp[7]) ? 16'b0000000111111111 : node6014;
												assign node6014 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
										assign node6018 = (inp[8]) ? node6024 : node6019;
											assign node6019 = (inp[15]) ? 16'b0000001111111111 : node6020;
												assign node6020 = (inp[10]) ? 16'b0000001111111111 : 16'b0000111111111111;
											assign node6024 = (inp[15]) ? node6030 : node6025;
												assign node6025 = (inp[13]) ? 16'b0000000111111111 : node6026;
													assign node6026 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6030 = (inp[10]) ? node6032 : 16'b0000000111111111;
													assign node6032 = (inp[7]) ? 16'b0000000011111111 : node6033;
														assign node6033 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node6037 = (inp[7]) ? node6077 : node6038;
									assign node6038 = (inp[14]) ? node6056 : node6039;
										assign node6039 = (inp[10]) ? 16'b0000001111111111 : node6040;
											assign node6040 = (inp[15]) ? node6048 : node6041;
												assign node6041 = (inp[3]) ? node6043 : 16'b0000111111111111;
													assign node6043 = (inp[8]) ? node6045 : 16'b0000111111111111;
														assign node6045 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6048 = (inp[5]) ? node6050 : 16'b0000011111111111;
													assign node6050 = (inp[9]) ? 16'b0000000011111111 : node6051;
														assign node6051 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node6056 = (inp[8]) ? node6068 : node6057;
											assign node6057 = (inp[10]) ? node6061 : node6058;
												assign node6058 = (inp[9]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node6061 = (inp[3]) ? node6063 : 16'b0000001111111111;
													assign node6063 = (inp[5]) ? 16'b0000000111111111 : node6064;
														assign node6064 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6068 = (inp[5]) ? node6072 : node6069;
												assign node6069 = (inp[3]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node6072 = (inp[9]) ? node6074 : 16'b0000000111111111;
													assign node6074 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node6077 = (inp[8]) ? node6097 : node6078;
										assign node6078 = (inp[13]) ? node6084 : node6079;
											assign node6079 = (inp[14]) ? node6081 : 16'b0000011111111111;
												assign node6081 = (inp[15]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node6084 = (inp[3]) ? node6094 : node6085;
												assign node6085 = (inp[15]) ? node6087 : 16'b0000011111111111;
													assign node6087 = (inp[10]) ? 16'b0000000111111111 : node6088;
														assign node6088 = (inp[9]) ? node6090 : 16'b0000001111111111;
															assign node6090 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6094 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node6097 = (inp[14]) ? node6111 : node6098;
											assign node6098 = (inp[5]) ? node6104 : node6099;
												assign node6099 = (inp[13]) ? node6101 : 16'b0000001111111111;
													assign node6101 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6104 = (inp[15]) ? node6106 : 16'b0000000111111111;
													assign node6106 = (inp[3]) ? 16'b0000000011111111 : node6107;
														assign node6107 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6111 = (inp[3]) ? node6115 : node6112;
												assign node6112 = (inp[9]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node6115 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node6118 = (inp[0]) ? node6224 : node6119;
								assign node6119 = (inp[15]) ? node6179 : node6120;
									assign node6120 = (inp[3]) ? node6144 : node6121;
										assign node6121 = (inp[10]) ? node6133 : node6122;
											assign node6122 = (inp[14]) ? node6128 : node6123;
												assign node6123 = (inp[13]) ? node6125 : 16'b0000111111111111;
													assign node6125 = (inp[7]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node6128 = (inp[5]) ? 16'b0000001111111111 : node6129;
													assign node6129 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node6133 = (inp[5]) ? node6141 : node6134;
												assign node6134 = (inp[7]) ? 16'b0000001111111111 : node6135;
													assign node6135 = (inp[8]) ? node6137 : 16'b0000011111111111;
														assign node6137 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6141 = (inp[14]) ? 16'b0000001111111111 : 16'b0000000111111111;
										assign node6144 = (inp[13]) ? node6160 : node6145;
											assign node6145 = (inp[14]) ? node6155 : node6146;
												assign node6146 = (inp[5]) ? node6148 : 16'b0000011111111111;
													assign node6148 = (inp[9]) ? 16'b0000001111111111 : node6149;
														assign node6149 = (inp[10]) ? 16'b0000001111111111 : node6150;
															assign node6150 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6155 = (inp[8]) ? node6157 : 16'b0000001111111111;
													assign node6157 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6160 = (inp[9]) ? node6174 : node6161;
												assign node6161 = (inp[14]) ? node6167 : node6162;
													assign node6162 = (inp[5]) ? node6164 : 16'b0000001111111111;
														assign node6164 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6167 = (inp[10]) ? node6171 : node6168;
														assign node6168 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6171 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node6174 = (inp[8]) ? node6176 : 16'b0000000111111111;
													assign node6176 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node6179 = (inp[10]) ? node6205 : node6180;
										assign node6180 = (inp[13]) ? node6188 : node6181;
											assign node6181 = (inp[7]) ? 16'b0000001111111111 : node6182;
												assign node6182 = (inp[5]) ? node6184 : 16'b0000011111111111;
													assign node6184 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node6188 = (inp[14]) ? node6196 : node6189;
												assign node6189 = (inp[5]) ? 16'b0000000111111111 : node6190;
													assign node6190 = (inp[8]) ? 16'b0000000111111111 : node6191;
														assign node6191 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6196 = (inp[8]) ? node6202 : node6197;
													assign node6197 = (inp[9]) ? node6199 : 16'b0000001111111111;
														assign node6199 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6202 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6205 = (inp[9]) ? node6217 : node6206;
											assign node6206 = (inp[5]) ? node6212 : node6207;
												assign node6207 = (inp[8]) ? 16'b0000000111111111 : node6208;
													assign node6208 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6212 = (inp[13]) ? node6214 : 16'b0000000111111111;
													assign node6214 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node6217 = (inp[8]) ? 16'b0000000001111111 : node6218;
												assign node6218 = (inp[5]) ? node6220 : 16'b0000000011111111;
													assign node6220 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node6224 = (inp[7]) ? node6270 : node6225;
									assign node6225 = (inp[5]) ? node6243 : node6226;
										assign node6226 = (inp[8]) ? 16'b0000000011111111 : node6227;
											assign node6227 = (inp[9]) ? node6233 : node6228;
												assign node6228 = (inp[13]) ? 16'b0000001111111111 : node6229;
													assign node6229 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node6233 = (inp[3]) ? node6237 : node6234;
													assign node6234 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6237 = (inp[10]) ? 16'b0000001111111111 : node6238;
														assign node6238 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node6243 = (inp[10]) ? node6261 : node6244;
											assign node6244 = (inp[13]) ? node6256 : node6245;
												assign node6245 = (inp[14]) ? node6251 : node6246;
													assign node6246 = (inp[8]) ? node6248 : 16'b0000011111111111;
														assign node6248 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6251 = (inp[3]) ? 16'b0000000111111111 : node6252;
														assign node6252 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6256 = (inp[3]) ? node6258 : 16'b0000000111111111;
													assign node6258 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6261 = (inp[9]) ? node6265 : node6262;
												assign node6262 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node6265 = (inp[3]) ? node6267 : 16'b0000000011111111;
													assign node6267 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000001111111;
									assign node6270 = (inp[9]) ? node6294 : node6271;
										assign node6271 = (inp[13]) ? node6281 : node6272;
											assign node6272 = (inp[14]) ? node6276 : node6273;
												assign node6273 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node6276 = (inp[15]) ? node6278 : 16'b0000000111111111;
													assign node6278 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6281 = (inp[15]) ? node6289 : node6282;
												assign node6282 = (inp[8]) ? 16'b0000000011111111 : node6283;
													assign node6283 = (inp[5]) ? node6285 : 16'b0000000111111111;
														assign node6285 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node6289 = (inp[3]) ? node6291 : 16'b0000000011111111;
													assign node6291 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node6294 = (inp[13]) ? node6308 : node6295;
											assign node6295 = (inp[14]) ? node6301 : node6296;
												assign node6296 = (inp[8]) ? 16'b0000000011111111 : node6297;
													assign node6297 = (inp[10]) ? 16'b0000001111111111 : 16'b0000000011111111;
												assign node6301 = (inp[8]) ? node6303 : 16'b0000000011111111;
													assign node6303 = (inp[15]) ? 16'b0000000000111111 : node6304;
														assign node6304 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6308 = (inp[5]) ? node6312 : node6309;
												assign node6309 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6312 = (inp[10]) ? node6314 : 16'b0000000001111111;
													assign node6314 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
						assign node6317 = (inp[13]) ? node6465 : node6318;
							assign node6318 = (inp[14]) ? node6384 : node6319;
								assign node6319 = (inp[9]) ? node6351 : node6320;
									assign node6320 = (inp[5]) ? node6340 : node6321;
										assign node6321 = (inp[3]) ? node6333 : node6322;
											assign node6322 = (inp[0]) ? node6328 : node6323;
												assign node6323 = (inp[15]) ? 16'b0000011111111111 : node6324;
													assign node6324 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node6328 = (inp[7]) ? 16'b0000001111111111 : node6329;
													assign node6329 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node6333 = (inp[10]) ? node6337 : node6334;
												assign node6334 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6337 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node6340 = (inp[10]) ? node6344 : node6341;
											assign node6341 = (inp[15]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node6344 = (inp[0]) ? 16'b0000000011111111 : node6345;
												assign node6345 = (inp[1]) ? node6347 : 16'b0000001111111111;
													assign node6347 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node6351 = (inp[10]) ? node6367 : node6352;
										assign node6352 = (inp[0]) ? node6362 : node6353;
											assign node6353 = (inp[5]) ? node6357 : node6354;
												assign node6354 = (inp[8]) ? 16'b0000011111111111 : 16'b0000001111111111;
												assign node6357 = (inp[1]) ? node6359 : 16'b0000001111111111;
													assign node6359 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node6362 = (inp[1]) ? 16'b0000000111111111 : node6363;
												assign node6363 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node6367 = (inp[5]) ? node6379 : node6368;
											assign node6368 = (inp[15]) ? node6374 : node6369;
												assign node6369 = (inp[7]) ? node6371 : 16'b0000011111111111;
													assign node6371 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6374 = (inp[1]) ? node6376 : 16'b0000000111111111;
													assign node6376 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6379 = (inp[0]) ? 16'b0000000001111111 : node6380;
												assign node6380 = (inp[1]) ? 16'b0000000111111111 : 16'b0000000011111111;
								assign node6384 = (inp[7]) ? node6426 : node6385;
									assign node6385 = (inp[5]) ? node6403 : node6386;
										assign node6386 = (inp[10]) ? node6392 : node6387;
											assign node6387 = (inp[9]) ? 16'b0000001111111111 : node6388;
												assign node6388 = (inp[3]) ? 16'b0000001111111111 : 16'b0000111111111111;
											assign node6392 = (inp[3]) ? node6396 : node6393;
												assign node6393 = (inp[8]) ? 16'b0000011111111111 : 16'b0000001111111111;
												assign node6396 = (inp[0]) ? node6398 : 16'b0000000111111111;
													assign node6398 = (inp[9]) ? node6400 : 16'b0000000111111111;
														assign node6400 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6403 = (inp[10]) ? node6419 : node6404;
											assign node6404 = (inp[15]) ? node6412 : node6405;
												assign node6405 = (inp[3]) ? node6407 : 16'b0000001111111111;
													assign node6407 = (inp[9]) ? 16'b0000000111111111 : node6408;
														assign node6408 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6412 = (inp[1]) ? node6414 : 16'b0000000111111111;
													assign node6414 = (inp[0]) ? 16'b0000000011111111 : node6415;
														assign node6415 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6419 = (inp[1]) ? node6423 : node6420;
												assign node6420 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6423 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node6426 = (inp[9]) ? node6440 : node6427;
										assign node6427 = (inp[5]) ? node6437 : node6428;
											assign node6428 = (inp[8]) ? node6434 : node6429;
												assign node6429 = (inp[1]) ? 16'b0000000111111111 : node6430;
													assign node6430 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6434 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6437 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node6440 = (inp[1]) ? node6458 : node6441;
											assign node6441 = (inp[0]) ? node6453 : node6442;
												assign node6442 = (inp[8]) ? node6450 : node6443;
													assign node6443 = (inp[15]) ? 16'b0000000011111111 : node6444;
														assign node6444 = (inp[5]) ? node6446 : 16'b0000000111111111;
															assign node6446 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6450 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6453 = (inp[15]) ? node6455 : 16'b0000000011111111;
													assign node6455 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6458 = (inp[10]) ? node6462 : node6459;
												assign node6459 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6462 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node6465 = (inp[0]) ? node6563 : node6466;
								assign node6466 = (inp[10]) ? node6516 : node6467;
									assign node6467 = (inp[5]) ? node6495 : node6468;
										assign node6468 = (inp[14]) ? node6490 : node6469;
											assign node6469 = (inp[8]) ? node6479 : node6470;
												assign node6470 = (inp[15]) ? node6474 : node6471;
													assign node6471 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node6474 = (inp[3]) ? node6476 : 16'b0000001111111111;
														assign node6476 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6479 = (inp[3]) ? node6485 : node6480;
													assign node6480 = (inp[1]) ? 16'b0000001111111111 : node6481;
														assign node6481 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6485 = (inp[15]) ? 16'b0000000011111111 : node6486;
														assign node6486 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6490 = (inp[9]) ? node6492 : 16'b0000001111111111;
												assign node6492 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6495 = (inp[7]) ? node6511 : node6496;
											assign node6496 = (inp[3]) ? node6502 : node6497;
												assign node6497 = (inp[9]) ? 16'b0000000111111111 : node6498;
													assign node6498 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6502 = (inp[15]) ? 16'b0000000011111111 : node6503;
													assign node6503 = (inp[8]) ? node6505 : 16'b0000001111111111;
														assign node6505 = (inp[9]) ? node6507 : 16'b0000000111111111;
															assign node6507 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000011111111;
											assign node6511 = (inp[1]) ? node6513 : 16'b0000000001111111;
												assign node6513 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node6516 = (inp[7]) ? node6546 : node6517;
										assign node6517 = (inp[9]) ? node6525 : node6518;
											assign node6518 = (inp[15]) ? 16'b0000000111111111 : node6519;
												assign node6519 = (inp[14]) ? node6521 : 16'b0000001111111111;
													assign node6521 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6525 = (inp[8]) ? node6531 : node6526;
												assign node6526 = (inp[1]) ? node6528 : 16'b0000000111111111;
													assign node6528 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6531 = (inp[14]) ? node6541 : node6532;
													assign node6532 = (inp[5]) ? node6536 : node6533;
														assign node6533 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6536 = (inp[1]) ? node6538 : 16'b0000000011111111;
															assign node6538 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6541 = (inp[1]) ? node6543 : 16'b0000000001111111;
														assign node6543 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6546 = (inp[1]) ? node6552 : node6547;
											assign node6547 = (inp[3]) ? node6549 : 16'b0000000111111111;
												assign node6549 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node6552 = (inp[5]) ? node6556 : node6553;
												assign node6553 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6556 = (inp[8]) ? 16'b0000000000011111 : node6557;
													assign node6557 = (inp[15]) ? node6559 : 16'b0000000001111111;
														assign node6559 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node6563 = (inp[8]) ? node6601 : node6564;
									assign node6564 = (inp[14]) ? node6580 : node6565;
										assign node6565 = (inp[15]) ? node6571 : node6566;
											assign node6566 = (inp[3]) ? node6568 : 16'b0000001111111111;
												assign node6568 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6571 = (inp[5]) ? node6575 : node6572;
												assign node6572 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6575 = (inp[7]) ? node6577 : 16'b0000000011111111;
													assign node6577 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6580 = (inp[10]) ? node6590 : node6581;
											assign node6581 = (inp[3]) ? node6585 : node6582;
												assign node6582 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6585 = (inp[7]) ? node6587 : 16'b0000000011111111;
													assign node6587 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6590 = (inp[7]) ? node6594 : node6591;
												assign node6591 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6594 = (inp[3]) ? 16'b0000000000111111 : node6595;
													assign node6595 = (inp[5]) ? node6597 : 16'b0000000001111111;
														assign node6597 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node6601 = (inp[7]) ? node6619 : node6602;
										assign node6602 = (inp[10]) ? node6608 : node6603;
											assign node6603 = (inp[5]) ? 16'b0000000001111111 : node6604;
												assign node6604 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6608 = (inp[9]) ? node6612 : node6609;
												assign node6609 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6612 = (inp[3]) ? node6614 : 16'b0000000001111111;
													assign node6614 = (inp[15]) ? 16'b0000000000111111 : node6615;
														assign node6615 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node6619 = (inp[9]) ? node6629 : node6620;
											assign node6620 = (inp[1]) ? node6622 : 16'b0000000001111111;
												assign node6622 = (inp[3]) ? 16'b0000000000111111 : node6623;
													assign node6623 = (inp[15]) ? node6625 : 16'b0000000011111111;
														assign node6625 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6629 = (inp[5]) ? node6639 : node6630;
												assign node6630 = (inp[10]) ? node6636 : node6631;
													assign node6631 = (inp[1]) ? 16'b0000000001111111 : node6632;
														assign node6632 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node6636 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000011111;
												assign node6639 = (inp[1]) ? 16'b0000000000001111 : node6640;
													assign node6640 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000000011111;
					assign node6644 = (inp[1]) ? node6984 : node6645;
						assign node6645 = (inp[8]) ? node6819 : node6646;
							assign node6646 = (inp[0]) ? node6742 : node6647;
								assign node6647 = (inp[13]) ? node6697 : node6648;
									assign node6648 = (inp[14]) ? node6666 : node6649;
										assign node6649 = (inp[15]) ? node6657 : node6650;
											assign node6650 = (inp[12]) ? node6652 : 16'b0000111111111111;
												assign node6652 = (inp[3]) ? node6654 : 16'b0000111111111111;
													assign node6654 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node6657 = (inp[3]) ? node6663 : node6658;
												assign node6658 = (inp[9]) ? node6660 : 16'b0001111111111111;
													assign node6660 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6663 = (inp[9]) ? 16'b0000001111111111 : 16'b0000000111111111;
										assign node6666 = (inp[7]) ? node6686 : node6667;
											assign node6667 = (inp[9]) ? node6677 : node6668;
												assign node6668 = (inp[3]) ? node6674 : node6669;
													assign node6669 = (inp[10]) ? 16'b0000011111111111 : node6670;
														assign node6670 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node6674 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6677 = (inp[10]) ? 16'b0000000111111111 : node6678;
													assign node6678 = (inp[5]) ? 16'b0000001111111111 : node6679;
														assign node6679 = (inp[15]) ? node6681 : 16'b0000011111111111;
															assign node6681 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node6686 = (inp[9]) ? node6692 : node6687;
												assign node6687 = (inp[12]) ? node6689 : 16'b0000001111111111;
													assign node6689 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node6692 = (inp[3]) ? 16'b0000000000111111 : node6693;
													assign node6693 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node6697 = (inp[12]) ? node6717 : node6698;
										assign node6698 = (inp[9]) ? node6712 : node6699;
											assign node6699 = (inp[10]) ? node6707 : node6700;
												assign node6700 = (inp[14]) ? 16'b0000111111111111 : node6701;
													assign node6701 = (inp[5]) ? node6703 : 16'b0000011111111111;
														assign node6703 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6707 = (inp[14]) ? 16'b0000001111111111 : node6708;
													assign node6708 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node6712 = (inp[5]) ? 16'b0000001111111111 : node6713;
												assign node6713 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6717 = (inp[3]) ? node6731 : node6718;
											assign node6718 = (inp[5]) ? node6728 : node6719;
												assign node6719 = (inp[10]) ? node6721 : 16'b0000001111111111;
													assign node6721 = (inp[7]) ? 16'b0000000111111111 : node6722;
														assign node6722 = (inp[9]) ? node6724 : 16'b0000001111111111;
															assign node6724 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6728 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6731 = (inp[10]) ? node6735 : node6732;
												assign node6732 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6735 = (inp[9]) ? node6739 : node6736;
													assign node6736 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6739 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node6742 = (inp[7]) ? node6788 : node6743;
									assign node6743 = (inp[13]) ? node6767 : node6744;
										assign node6744 = (inp[5]) ? node6758 : node6745;
											assign node6745 = (inp[9]) ? node6753 : node6746;
												assign node6746 = (inp[15]) ? node6750 : node6747;
													assign node6747 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node6750 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6753 = (inp[10]) ? 16'b0000000011111111 : node6754;
													assign node6754 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6758 = (inp[15]) ? node6760 : 16'b0000001111111111;
												assign node6760 = (inp[10]) ? node6762 : 16'b0000000111111111;
													assign node6762 = (inp[3]) ? 16'b0000000111111111 : node6763;
														assign node6763 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node6767 = (inp[10]) ? node6775 : node6768;
											assign node6768 = (inp[9]) ? 16'b0000000111111111 : node6769;
												assign node6769 = (inp[3]) ? node6771 : 16'b0000001111111111;
													assign node6771 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node6775 = (inp[15]) ? node6781 : node6776;
												assign node6776 = (inp[12]) ? 16'b0000000011111111 : node6777;
													assign node6777 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6781 = (inp[5]) ? node6783 : 16'b0000000011111111;
													assign node6783 = (inp[9]) ? node6785 : 16'b0000000001111111;
														assign node6785 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000001111111;
									assign node6788 = (inp[14]) ? node6806 : node6789;
										assign node6789 = (inp[10]) ? node6799 : node6790;
											assign node6790 = (inp[5]) ? 16'b0000000111111111 : node6791;
												assign node6791 = (inp[9]) ? node6793 : 16'b0000001111111111;
													assign node6793 = (inp[12]) ? 16'b0000000111111111 : node6794;
														assign node6794 = (inp[3]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node6799 = (inp[13]) ? node6803 : node6800;
												assign node6800 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6803 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6806 = (inp[9]) ? node6810 : node6807;
											assign node6807 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6810 = (inp[12]) ? node6812 : 16'b0000000001111111;
												assign node6812 = (inp[5]) ? node6814 : 16'b0000000001111111;
													assign node6814 = (inp[13]) ? 16'b0000000000011111 : node6815;
														assign node6815 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node6819 = (inp[0]) ? node6897 : node6820;
								assign node6820 = (inp[12]) ? node6860 : node6821;
									assign node6821 = (inp[13]) ? node6839 : node6822;
										assign node6822 = (inp[9]) ? node6830 : node6823;
											assign node6823 = (inp[14]) ? 16'b0000001111111111 : node6824;
												assign node6824 = (inp[3]) ? node6826 : 16'b0000001111111111;
													assign node6826 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6830 = (inp[7]) ? 16'b0000000011111111 : node6831;
												assign node6831 = (inp[3]) ? node6835 : node6832;
													assign node6832 = (inp[10]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node6835 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node6839 = (inp[5]) ? node6843 : node6840;
											assign node6840 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node6843 = (inp[15]) ? node6855 : node6844;
												assign node6844 = (inp[10]) ? node6850 : node6845;
													assign node6845 = (inp[14]) ? node6847 : 16'b0000000111111111;
														assign node6847 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6850 = (inp[7]) ? node6852 : 16'b0000000011111111;
														assign node6852 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6855 = (inp[9]) ? 16'b0000000001111111 : node6856;
													assign node6856 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node6860 = (inp[14]) ? node6878 : node6861;
										assign node6861 = (inp[5]) ? node6871 : node6862;
											assign node6862 = (inp[10]) ? node6866 : node6863;
												assign node6863 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6866 = (inp[9]) ? node6868 : 16'b0000000111111111;
													assign node6868 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node6871 = (inp[7]) ? node6873 : 16'b0000000001111111;
												assign node6873 = (inp[3]) ? 16'b0000000011111111 : node6874;
													assign node6874 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node6878 = (inp[15]) ? node6890 : node6879;
											assign node6879 = (inp[10]) ? node6885 : node6880;
												assign node6880 = (inp[9]) ? node6882 : 16'b0000000111111111;
													assign node6882 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node6885 = (inp[13]) ? 16'b0000000001111111 : node6886;
													assign node6886 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6890 = (inp[10]) ? node6894 : node6891;
												assign node6891 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6894 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000000111111;
								assign node6897 = (inp[14]) ? node6937 : node6898;
									assign node6898 = (inp[5]) ? node6910 : node6899;
										assign node6899 = (inp[10]) ? node6907 : node6900;
											assign node6900 = (inp[3]) ? 16'b0000000111111111 : node6901;
												assign node6901 = (inp[15]) ? node6903 : 16'b0000011111111111;
													assign node6903 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6907 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node6910 = (inp[9]) ? node6928 : node6911;
											assign node6911 = (inp[12]) ? node6917 : node6912;
												assign node6912 = (inp[13]) ? 16'b0000000011111111 : node6913;
													assign node6913 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6917 = (inp[15]) ? node6923 : node6918;
													assign node6918 = (inp[7]) ? 16'b0000000011111111 : node6919;
														assign node6919 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6923 = (inp[10]) ? 16'b0000000001111111 : node6924;
														assign node6924 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6928 = (inp[12]) ? 16'b0000000000111111 : node6929;
												assign node6929 = (inp[7]) ? node6931 : 16'b0000000011111111;
													assign node6931 = (inp[15]) ? 16'b0000000001111111 : node6932;
														assign node6932 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000001111111;
									assign node6937 = (inp[3]) ? node6957 : node6938;
										assign node6938 = (inp[7]) ? node6946 : node6939;
											assign node6939 = (inp[9]) ? node6941 : 16'b0000000111111111;
												assign node6941 = (inp[12]) ? 16'b0000000011111111 : node6942;
													assign node6942 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node6946 = (inp[9]) ? node6950 : node6947;
												assign node6947 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node6950 = (inp[5]) ? 16'b0000000000011111 : node6951;
													assign node6951 = (inp[10]) ? node6953 : 16'b0000000001111111;
														assign node6953 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6957 = (inp[7]) ? node6973 : node6958;
											assign node6958 = (inp[12]) ? node6966 : node6959;
												assign node6959 = (inp[10]) ? 16'b0000000001111111 : node6960;
													assign node6960 = (inp[15]) ? node6962 : 16'b0000000011111111;
														assign node6962 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node6966 = (inp[5]) ? node6970 : node6967;
													assign node6967 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node6970 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node6973 = (inp[12]) ? node6975 : 16'b0000000000011111;
												assign node6975 = (inp[15]) ? node6977 : 16'b0000000000011111;
													assign node6977 = (inp[5]) ? node6981 : node6978;
														assign node6978 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node6981 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
						assign node6984 = (inp[13]) ? node7156 : node6985;
							assign node6985 = (inp[3]) ? node7075 : node6986;
								assign node6986 = (inp[15]) ? node7026 : node6987;
									assign node6987 = (inp[0]) ? node7009 : node6988;
										assign node6988 = (inp[9]) ? node6998 : node6989;
											assign node6989 = (inp[5]) ? node6993 : node6990;
												assign node6990 = (inp[12]) ? 16'b0000001111111111 : 16'b0000111111111111;
												assign node6993 = (inp[14]) ? node6995 : 16'b0000001111111111;
													assign node6995 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6998 = (inp[14]) ? node7006 : node6999;
												assign node6999 = (inp[8]) ? 16'b0000000111111111 : node7000;
													assign node7000 = (inp[12]) ? node7002 : 16'b0000001111111111;
														assign node7002 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7006 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node7009 = (inp[14]) ? node7021 : node7010;
											assign node7010 = (inp[8]) ? node7018 : node7011;
												assign node7011 = (inp[5]) ? node7013 : 16'b0000011111111111;
													assign node7013 = (inp[9]) ? 16'b0000000111111111 : node7014;
														assign node7014 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7018 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7021 = (inp[10]) ? node7023 : 16'b0000000011111111;
												assign node7023 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node7026 = (inp[7]) ? node7048 : node7027;
										assign node7027 = (inp[14]) ? node7037 : node7028;
											assign node7028 = (inp[5]) ? node7034 : node7029;
												assign node7029 = (inp[12]) ? 16'b0000000111111111 : node7030;
													assign node7030 = (inp[0]) ? 16'b0000011111111111 : 16'b0000001111111111;
												assign node7034 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7037 = (inp[9]) ? node7043 : node7038;
												assign node7038 = (inp[0]) ? 16'b0000000011111111 : node7039;
													assign node7039 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7043 = (inp[12]) ? node7045 : 16'b0000000011111111;
													assign node7045 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000000111111;
										assign node7048 = (inp[12]) ? node7066 : node7049;
											assign node7049 = (inp[5]) ? node7055 : node7050;
												assign node7050 = (inp[14]) ? node7052 : 16'b0000000111111111;
													assign node7052 = (inp[9]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node7055 = (inp[8]) ? node7059 : node7056;
													assign node7056 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7059 = (inp[10]) ? 16'b0000000000111111 : node7060;
														assign node7060 = (inp[14]) ? 16'b0000000001111111 : node7061;
															assign node7061 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7066 = (inp[5]) ? node7072 : node7067;
												assign node7067 = (inp[10]) ? 16'b0000000001111111 : node7068;
													assign node7068 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7072 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node7075 = (inp[14]) ? node7113 : node7076;
									assign node7076 = (inp[10]) ? node7090 : node7077;
										assign node7077 = (inp[9]) ? node7085 : node7078;
											assign node7078 = (inp[5]) ? node7082 : node7079;
												assign node7079 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7082 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node7085 = (inp[5]) ? node7087 : 16'b0000000011111111;
												assign node7087 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node7090 = (inp[9]) ? node7106 : node7091;
											assign node7091 = (inp[0]) ? node7099 : node7092;
												assign node7092 = (inp[7]) ? 16'b0000000011111111 : node7093;
													assign node7093 = (inp[12]) ? node7095 : 16'b0000001111111111;
														assign node7095 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node7099 = (inp[12]) ? node7101 : 16'b0000000011111111;
													assign node7101 = (inp[8]) ? 16'b0000000000011111 : node7102;
														assign node7102 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7106 = (inp[7]) ? node7110 : node7107;
												assign node7107 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7110 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node7113 = (inp[8]) ? node7131 : node7114;
										assign node7114 = (inp[9]) ? node7126 : node7115;
											assign node7115 = (inp[10]) ? node7123 : node7116;
												assign node7116 = (inp[5]) ? node7118 : 16'b0000000111111111;
													assign node7118 = (inp[0]) ? node7120 : 16'b0000000011111111;
														assign node7120 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7123 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7126 = (inp[12]) ? 16'b0000000000111111 : node7127;
												assign node7127 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node7131 = (inp[5]) ? node7145 : node7132;
											assign node7132 = (inp[10]) ? node7138 : node7133;
												assign node7133 = (inp[9]) ? 16'b0000000001111111 : node7134;
													assign node7134 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7138 = (inp[0]) ? node7140 : 16'b0000000001111111;
													assign node7140 = (inp[7]) ? 16'b0000000000111111 : node7141;
														assign node7141 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7145 = (inp[0]) ? node7153 : node7146;
												assign node7146 = (inp[12]) ? 16'b0000000000111111 : node7147;
													assign node7147 = (inp[15]) ? node7149 : 16'b0000000011111111;
														assign node7149 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7153 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node7156 = (inp[10]) ? node7256 : node7157;
								assign node7157 = (inp[15]) ? node7211 : node7158;
									assign node7158 = (inp[12]) ? node7188 : node7159;
										assign node7159 = (inp[3]) ? node7175 : node7160;
											assign node7160 = (inp[8]) ? node7166 : node7161;
												assign node7161 = (inp[14]) ? 16'b0000000111111111 : node7162;
													assign node7162 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7166 = (inp[0]) ? node7172 : node7167;
													assign node7167 = (inp[7]) ? node7169 : 16'b0000000111111111;
														assign node7169 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7172 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7175 = (inp[0]) ? node7179 : node7176;
												assign node7176 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node7179 = (inp[9]) ? node7181 : 16'b0000000111111111;
													assign node7181 = (inp[5]) ? 16'b0000000001111111 : node7182;
														assign node7182 = (inp[8]) ? 16'b0000000001111111 : node7183;
															assign node7183 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node7188 = (inp[9]) ? node7204 : node7189;
											assign node7189 = (inp[0]) ? node7193 : node7190;
												assign node7190 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7193 = (inp[8]) ? node7199 : node7194;
													assign node7194 = (inp[7]) ? 16'b0000000011111111 : node7195;
														assign node7195 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7199 = (inp[3]) ? 16'b0000000001111111 : node7200;
														assign node7200 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7204 = (inp[8]) ? node7208 : node7205;
												assign node7205 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7208 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000000011111;
									assign node7211 = (inp[14]) ? node7229 : node7212;
										assign node7212 = (inp[8]) ? node7216 : node7213;
											assign node7213 = (inp[9]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node7216 = (inp[9]) ? node7224 : node7217;
												assign node7217 = (inp[5]) ? 16'b0000000001111111 : node7218;
													assign node7218 = (inp[12]) ? node7220 : 16'b0000000011111111;
														assign node7220 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7224 = (inp[5]) ? node7226 : 16'b0000000000111111;
													assign node7226 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7229 = (inp[3]) ? node7239 : node7230;
											assign node7230 = (inp[0]) ? node7236 : node7231;
												assign node7231 = (inp[12]) ? 16'b0000000001111111 : node7232;
													assign node7232 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7236 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7239 = (inp[5]) ? node7245 : node7240;
												assign node7240 = (inp[7]) ? 16'b0000000000111111 : node7241;
													assign node7241 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7245 = (inp[12]) ? node7249 : node7246;
													assign node7246 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node7249 = (inp[9]) ? node7251 : 16'b0000000000011111;
														assign node7251 = (inp[7]) ? 16'b0000000000001111 : node7252;
															assign node7252 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node7256 = (inp[7]) ? node7286 : node7257;
									assign node7257 = (inp[0]) ? node7273 : node7258;
										assign node7258 = (inp[9]) ? node7264 : node7259;
											assign node7259 = (inp[12]) ? node7261 : 16'b0000000011111111;
												assign node7261 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7264 = (inp[8]) ? node7270 : node7265;
												assign node7265 = (inp[14]) ? 16'b0000000011111111 : node7266;
													assign node7266 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7270 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7273 = (inp[5]) ? node7279 : node7274;
											assign node7274 = (inp[15]) ? 16'b0000000000111111 : node7275;
												assign node7275 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node7279 = (inp[14]) ? 16'b0000000000011111 : node7280;
												assign node7280 = (inp[12]) ? node7282 : 16'b0000000011111111;
													assign node7282 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node7286 = (inp[5]) ? node7316 : node7287;
										assign node7287 = (inp[0]) ? node7297 : node7288;
											assign node7288 = (inp[15]) ? 16'b0000000000111111 : node7289;
												assign node7289 = (inp[8]) ? 16'b0000000001111111 : node7290;
													assign node7290 = (inp[12]) ? node7292 : 16'b0000000011111111;
														assign node7292 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7297 = (inp[12]) ? node7307 : node7298;
												assign node7298 = (inp[8]) ? node7300 : 16'b0000000001111111;
													assign node7300 = (inp[14]) ? node7302 : 16'b0000000000111111;
														assign node7302 = (inp[15]) ? node7304 : 16'b0000000000111111;
															assign node7304 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7307 = (inp[14]) ? node7313 : node7308;
													assign node7308 = (inp[8]) ? node7310 : 16'b0000000000111111;
														assign node7310 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node7313 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node7316 = (inp[15]) ? node7330 : node7317;
											assign node7317 = (inp[14]) ? node7325 : node7318;
												assign node7318 = (inp[8]) ? node7322 : node7319;
													assign node7319 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7322 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7325 = (inp[3]) ? node7327 : 16'b0000000000111111;
													assign node7327 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node7330 = (inp[12]) ? node7338 : node7331;
												assign node7331 = (inp[0]) ? node7335 : node7332;
													assign node7332 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node7335 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7338 = (inp[14]) ? node7340 : 16'b0000000000001111;
													assign node7340 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
				assign node7343 = (inp[9]) ? node7947 : node7344;
					assign node7344 = (inp[3]) ? node7662 : node7345;
						assign node7345 = (inp[0]) ? node7503 : node7346;
							assign node7346 = (inp[15]) ? node7430 : node7347;
								assign node7347 = (inp[7]) ? node7389 : node7348;
									assign node7348 = (inp[14]) ? node7372 : node7349;
										assign node7349 = (inp[4]) ? node7363 : node7350;
											assign node7350 = (inp[8]) ? node7356 : node7351;
												assign node7351 = (inp[12]) ? 16'b0000011111111111 : node7352;
													assign node7352 = (inp[5]) ? 16'b0001111111111111 : 16'b0000111111111111;
												assign node7356 = (inp[5]) ? node7358 : 16'b0000011111111111;
													assign node7358 = (inp[1]) ? node7360 : 16'b0000011111111111;
														assign node7360 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node7363 = (inp[10]) ? node7369 : node7364;
												assign node7364 = (inp[8]) ? 16'b0000001111111111 : node7365;
													assign node7365 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node7369 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node7372 = (inp[5]) ? node7382 : node7373;
											assign node7373 = (inp[13]) ? node7379 : node7374;
												assign node7374 = (inp[10]) ? node7376 : 16'b0000011111111111;
													assign node7376 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node7379 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node7382 = (inp[12]) ? 16'b0000000111111111 : node7383;
												assign node7383 = (inp[10]) ? node7385 : 16'b0000111111111111;
													assign node7385 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
									assign node7389 = (inp[13]) ? node7417 : node7390;
										assign node7390 = (inp[10]) ? node7404 : node7391;
											assign node7391 = (inp[8]) ? node7401 : node7392;
												assign node7392 = (inp[5]) ? node7396 : node7393;
													assign node7393 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node7396 = (inp[14]) ? 16'b0000001111111111 : node7397;
														assign node7397 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node7401 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
											assign node7404 = (inp[1]) ? node7414 : node7405;
												assign node7405 = (inp[12]) ? node7407 : 16'b0000001111111111;
													assign node7407 = (inp[4]) ? 16'b0000000111111111 : node7408;
														assign node7408 = (inp[8]) ? node7410 : 16'b0000001111111111;
															assign node7410 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7414 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node7417 = (inp[4]) ? node7425 : node7418;
											assign node7418 = (inp[1]) ? node7420 : 16'b0000000111111111;
												assign node7420 = (inp[12]) ? node7422 : 16'b0000000011111111;
													assign node7422 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7425 = (inp[1]) ? node7427 : 16'b0000000011111111;
												assign node7427 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node7430 = (inp[1]) ? node7474 : node7431;
									assign node7431 = (inp[4]) ? node7459 : node7432;
										assign node7432 = (inp[8]) ? node7446 : node7433;
											assign node7433 = (inp[13]) ? node7439 : node7434;
												assign node7434 = (inp[5]) ? node7436 : 16'b0000111111111111;
													assign node7436 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node7439 = (inp[10]) ? node7443 : node7440;
													assign node7440 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7443 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7446 = (inp[10]) ? node7454 : node7447;
												assign node7447 = (inp[5]) ? 16'b0000000111111111 : node7448;
													assign node7448 = (inp[14]) ? node7450 : 16'b0000001111111111;
														assign node7450 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7454 = (inp[14]) ? 16'b0000000011111111 : node7455;
													assign node7455 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node7459 = (inp[7]) ? node7465 : node7460;
											assign node7460 = (inp[13]) ? 16'b0000000111111111 : node7461;
												assign node7461 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node7465 = (inp[14]) ? 16'b0000000001111111 : node7466;
												assign node7466 = (inp[13]) ? node7468 : 16'b0000001111111111;
													assign node7468 = (inp[10]) ? 16'b0000000011111111 : node7469;
														assign node7469 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node7474 = (inp[13]) ? node7486 : node7475;
										assign node7475 = (inp[4]) ? node7481 : node7476;
											assign node7476 = (inp[7]) ? node7478 : 16'b0000001111111111;
												assign node7478 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node7481 = (inp[12]) ? 16'b0000000011111111 : node7482;
												assign node7482 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node7486 = (inp[5]) ? node7492 : node7487;
											assign node7487 = (inp[10]) ? 16'b0000000011111111 : node7488;
												assign node7488 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7492 = (inp[10]) ? node7498 : node7493;
												assign node7493 = (inp[14]) ? node7495 : 16'b0000000011111111;
													assign node7495 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7498 = (inp[14]) ? 16'b0000000000011111 : node7499;
													assign node7499 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node7503 = (inp[7]) ? node7589 : node7504;
								assign node7504 = (inp[10]) ? node7544 : node7505;
									assign node7505 = (inp[5]) ? node7525 : node7506;
										assign node7506 = (inp[14]) ? node7512 : node7507;
											assign node7507 = (inp[1]) ? node7509 : 16'b0000011111111111;
												assign node7509 = (inp[8]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node7512 = (inp[15]) ? node7518 : node7513;
												assign node7513 = (inp[4]) ? node7515 : 16'b0000001111111111;
													assign node7515 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7518 = (inp[1]) ? 16'b0000000011111111 : node7519;
													assign node7519 = (inp[12]) ? 16'b0000000111111111 : node7520;
														assign node7520 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node7525 = (inp[12]) ? node7533 : node7526;
											assign node7526 = (inp[4]) ? node7528 : 16'b0000001111111111;
												assign node7528 = (inp[13]) ? 16'b0000000111111111 : node7529;
													assign node7529 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7533 = (inp[14]) ? node7537 : node7534;
												assign node7534 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7537 = (inp[15]) ? 16'b0000000001111111 : node7538;
													assign node7538 = (inp[13]) ? node7540 : 16'b0000000011111111;
														assign node7540 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node7544 = (inp[4]) ? node7564 : node7545;
										assign node7545 = (inp[14]) ? node7553 : node7546;
											assign node7546 = (inp[13]) ? 16'b0000000111111111 : node7547;
												assign node7547 = (inp[5]) ? 16'b0000001111111111 : node7548;
													assign node7548 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node7553 = (inp[8]) ? node7559 : node7554;
												assign node7554 = (inp[13]) ? node7556 : 16'b0000000111111111;
													assign node7556 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7559 = (inp[5]) ? 16'b0000000001111111 : node7560;
													assign node7560 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node7564 = (inp[13]) ? node7580 : node7565;
											assign node7565 = (inp[5]) ? node7575 : node7566;
												assign node7566 = (inp[8]) ? 16'b0000000011111111 : node7567;
													assign node7567 = (inp[15]) ? node7569 : 16'b0000001111111111;
														assign node7569 = (inp[1]) ? 16'b0000000011111111 : node7570;
															assign node7570 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7575 = (inp[15]) ? 16'b0000000000011111 : node7576;
													assign node7576 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7580 = (inp[8]) ? node7582 : 16'b0000000001111111;
												assign node7582 = (inp[15]) ? 16'b0000000000111111 : node7583;
													assign node7583 = (inp[12]) ? node7585 : 16'b0000000001111111;
														assign node7585 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node7589 = (inp[8]) ? node7629 : node7590;
									assign node7590 = (inp[15]) ? node7608 : node7591;
										assign node7591 = (inp[5]) ? node7601 : node7592;
											assign node7592 = (inp[13]) ? node7596 : node7593;
												assign node7593 = (inp[10]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node7596 = (inp[10]) ? node7598 : 16'b0000000111111111;
													assign node7598 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7601 = (inp[1]) ? node7603 : 16'b0000000011111111;
												assign node7603 = (inp[10]) ? 16'b0000000011111111 : node7604;
													assign node7604 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000011111111;
										assign node7608 = (inp[1]) ? node7620 : node7609;
											assign node7609 = (inp[13]) ? node7615 : node7610;
												assign node7610 = (inp[4]) ? node7612 : 16'b0000000111111111;
													assign node7612 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7615 = (inp[12]) ? 16'b0000000001111111 : node7616;
													assign node7616 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node7620 = (inp[13]) ? node7624 : node7621;
												assign node7621 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7624 = (inp[14]) ? node7626 : 16'b0000000001111111;
													assign node7626 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node7629 = (inp[14]) ? node7649 : node7630;
										assign node7630 = (inp[12]) ? node7644 : node7631;
											assign node7631 = (inp[5]) ? node7641 : node7632;
												assign node7632 = (inp[4]) ? node7638 : node7633;
													assign node7633 = (inp[15]) ? 16'b0000000111111111 : node7634;
														assign node7634 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7638 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7641 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7644 = (inp[13]) ? 16'b0000000000111111 : node7645;
												assign node7645 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node7649 = (inp[10]) ? node7655 : node7650;
											assign node7650 = (inp[1]) ? node7652 : 16'b0000000001111111;
												assign node7652 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7655 = (inp[12]) ? 16'b0000000000111111 : node7656;
												assign node7656 = (inp[1]) ? node7658 : 16'b0000000001111111;
													assign node7658 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node7662 = (inp[1]) ? node7792 : node7663;
							assign node7663 = (inp[4]) ? node7733 : node7664;
								assign node7664 = (inp[14]) ? node7694 : node7665;
									assign node7665 = (inp[8]) ? node7689 : node7666;
										assign node7666 = (inp[15]) ? node7684 : node7667;
											assign node7667 = (inp[13]) ? node7677 : node7668;
												assign node7668 = (inp[10]) ? node7670 : 16'b0001111111111111;
													assign node7670 = (inp[0]) ? 16'b0000001111111111 : node7671;
														assign node7671 = (inp[12]) ? node7673 : 16'b0000011111111111;
															assign node7673 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node7677 = (inp[10]) ? 16'b0000000111111111 : node7678;
													assign node7678 = (inp[0]) ? node7680 : 16'b0000001111111111;
														assign node7680 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node7684 = (inp[5]) ? 16'b0000000011111111 : node7685;
												assign node7685 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
										assign node7689 = (inp[10]) ? node7691 : 16'b0000000111111111;
											assign node7691 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000001111111;
									assign node7694 = (inp[0]) ? node7708 : node7695;
										assign node7695 = (inp[7]) ? node7701 : node7696;
											assign node7696 = (inp[15]) ? 16'b0000000111111111 : node7697;
												assign node7697 = (inp[8]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node7701 = (inp[10]) ? node7705 : node7702;
												assign node7702 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node7705 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node7708 = (inp[12]) ? node7722 : node7709;
											assign node7709 = (inp[10]) ? node7719 : node7710;
												assign node7710 = (inp[7]) ? 16'b0000000011111111 : node7711;
													assign node7711 = (inp[15]) ? node7715 : node7712;
														assign node7712 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7715 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7719 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7722 = (inp[5]) ? node7728 : node7723;
												assign node7723 = (inp[15]) ? node7725 : 16'b0000000011111111;
													assign node7725 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7728 = (inp[15]) ? node7730 : 16'b0000000001111111;
													assign node7730 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node7733 = (inp[5]) ? node7763 : node7734;
									assign node7734 = (inp[15]) ? node7750 : node7735;
										assign node7735 = (inp[10]) ? node7747 : node7736;
											assign node7736 = (inp[8]) ? node7742 : node7737;
												assign node7737 = (inp[14]) ? node7739 : 16'b0000001111111111;
													assign node7739 = (inp[12]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node7742 = (inp[7]) ? 16'b0000000011111111 : node7743;
													assign node7743 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node7747 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000001111111;
										assign node7750 = (inp[13]) ? node7754 : node7751;
											assign node7751 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node7754 = (inp[0]) ? 16'b0000000001111111 : node7755;
												assign node7755 = (inp[14]) ? node7757 : 16'b0000000011111111;
													assign node7757 = (inp[12]) ? 16'b0000000001111111 : node7758;
														assign node7758 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node7763 = (inp[8]) ? node7777 : node7764;
										assign node7764 = (inp[15]) ? node7772 : node7765;
											assign node7765 = (inp[14]) ? node7767 : 16'b0000000111111111;
												assign node7767 = (inp[12]) ? 16'b0000000001111111 : node7768;
													assign node7768 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7772 = (inp[0]) ? node7774 : 16'b0000000011111111;
												assign node7774 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7777 = (inp[0]) ? node7783 : node7778;
											assign node7778 = (inp[15]) ? node7780 : 16'b0000000001111111;
												assign node7780 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7783 = (inp[15]) ? node7789 : node7784;
												assign node7784 = (inp[14]) ? node7786 : 16'b0000000001111111;
													assign node7786 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7789 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node7792 = (inp[0]) ? node7866 : node7793;
								assign node7793 = (inp[4]) ? node7825 : node7794;
									assign node7794 = (inp[13]) ? node7806 : node7795;
										assign node7795 = (inp[8]) ? 16'b0000000001111111 : node7796;
											assign node7796 = (inp[12]) ? node7800 : node7797;
												assign node7797 = (inp[5]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node7800 = (inp[5]) ? node7802 : 16'b0000000111111111;
													assign node7802 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node7806 = (inp[10]) ? node7814 : node7807;
											assign node7807 = (inp[15]) ? node7809 : 16'b0000000011111111;
												assign node7809 = (inp[8]) ? 16'b0000000000111111 : node7810;
													assign node7810 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7814 = (inp[7]) ? 16'b0000000001111111 : node7815;
												assign node7815 = (inp[5]) ? node7819 : node7816;
													assign node7816 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7819 = (inp[14]) ? 16'b0000000000111111 : node7820;
														assign node7820 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node7825 = (inp[10]) ? node7849 : node7826;
										assign node7826 = (inp[13]) ? node7834 : node7827;
											assign node7827 = (inp[8]) ? node7831 : node7828;
												assign node7828 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7831 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node7834 = (inp[5]) ? node7842 : node7835;
												assign node7835 = (inp[14]) ? 16'b0000000001111111 : node7836;
													assign node7836 = (inp[7]) ? 16'b0000000001111111 : node7837;
														assign node7837 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7842 = (inp[12]) ? 16'b0000000000111111 : node7843;
													assign node7843 = (inp[14]) ? 16'b0000000000111111 : node7844;
														assign node7844 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node7849 = (inp[15]) ? node7859 : node7850;
											assign node7850 = (inp[5]) ? 16'b0000000000111111 : node7851;
												assign node7851 = (inp[8]) ? node7853 : 16'b0000000011111111;
													assign node7853 = (inp[13]) ? node7855 : 16'b0000000001111111;
														assign node7855 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7859 = (inp[13]) ? node7863 : node7860;
												assign node7860 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7863 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node7866 = (inp[10]) ? node7906 : node7867;
									assign node7867 = (inp[8]) ? node7883 : node7868;
										assign node7868 = (inp[15]) ? 16'b0000000001111111 : node7869;
											assign node7869 = (inp[13]) ? node7875 : node7870;
												assign node7870 = (inp[4]) ? 16'b0000000111111111 : node7871;
													assign node7871 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7875 = (inp[14]) ? node7879 : node7876;
													assign node7876 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7879 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node7883 = (inp[5]) ? node7897 : node7884;
											assign node7884 = (inp[12]) ? node7890 : node7885;
												assign node7885 = (inp[7]) ? node7887 : 16'b0000000111111111;
													assign node7887 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7890 = (inp[7]) ? 16'b0000000000111111 : node7891;
													assign node7891 = (inp[13]) ? 16'b0000000001111111 : node7892;
														assign node7892 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7897 = (inp[13]) ? node7899 : 16'b0000000000111111;
												assign node7899 = (inp[14]) ? node7901 : 16'b0000000000111111;
													assign node7901 = (inp[4]) ? node7903 : 16'b0000000000011111;
														assign node7903 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node7906 = (inp[13]) ? node7926 : node7907;
										assign node7907 = (inp[14]) ? node7917 : node7908;
											assign node7908 = (inp[7]) ? node7914 : node7909;
												assign node7909 = (inp[8]) ? node7911 : 16'b0000000011111111;
													assign node7911 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7914 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node7917 = (inp[4]) ? node7921 : node7918;
												assign node7918 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7921 = (inp[15]) ? node7923 : 16'b0000000000011111;
													assign node7923 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node7926 = (inp[4]) ? node7936 : node7927;
											assign node7927 = (inp[14]) ? node7929 : 16'b0000000000111111;
												assign node7929 = (inp[7]) ? 16'b0000000000001111 : node7930;
													assign node7930 = (inp[12]) ? node7932 : 16'b0000000000111111;
														assign node7932 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node7936 = (inp[14]) ? node7940 : node7937;
												assign node7937 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node7940 = (inp[8]) ? 16'b0000000000000111 : node7941;
													assign node7941 = (inp[12]) ? 16'b0000000000000111 : node7942;
														assign node7942 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node7947 = (inp[14]) ? node8283 : node7948;
						assign node7948 = (inp[15]) ? node8128 : node7949;
							assign node7949 = (inp[5]) ? node8035 : node7950;
								assign node7950 = (inp[7]) ? node8002 : node7951;
									assign node7951 = (inp[13]) ? node7977 : node7952;
										assign node7952 = (inp[8]) ? node7974 : node7953;
											assign node7953 = (inp[4]) ? node7967 : node7954;
												assign node7954 = (inp[1]) ? node7964 : node7955;
													assign node7955 = (inp[0]) ? node7959 : node7956;
														assign node7956 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node7959 = (inp[10]) ? 16'b0000001111111111 : node7960;
															assign node7960 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node7964 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7967 = (inp[10]) ? node7969 : 16'b0000001111111111;
													assign node7969 = (inp[12]) ? 16'b0000000011111111 : node7970;
														assign node7970 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node7974 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node7977 = (inp[10]) ? node7987 : node7978;
											assign node7978 = (inp[12]) ? node7984 : node7979;
												assign node7979 = (inp[3]) ? 16'b0000000111111111 : node7980;
													assign node7980 = (inp[4]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node7984 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7987 = (inp[4]) ? node7995 : node7988;
												assign node7988 = (inp[8]) ? node7992 : node7989;
													assign node7989 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7992 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node7995 = (inp[3]) ? 16'b0000000001111111 : node7996;
													assign node7996 = (inp[0]) ? 16'b0000000011111111 : node7997;
														assign node7997 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node8002 = (inp[13]) ? node8024 : node8003;
										assign node8003 = (inp[1]) ? node8011 : node8004;
											assign node8004 = (inp[8]) ? 16'b0000000111111111 : node8005;
												assign node8005 = (inp[10]) ? 16'b0000000111111111 : node8006;
													assign node8006 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node8011 = (inp[0]) ? node8017 : node8012;
												assign node8012 = (inp[12]) ? node8014 : 16'b0000000111111111;
													assign node8014 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8017 = (inp[12]) ? node8019 : 16'b0000000011111111;
													assign node8019 = (inp[3]) ? 16'b0000000000111111 : node8020;
														assign node8020 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node8024 = (inp[3]) ? node8030 : node8025;
											assign node8025 = (inp[10]) ? node8027 : 16'b0000000111111111;
												assign node8027 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8030 = (inp[8]) ? node8032 : 16'b0000000001111111;
												assign node8032 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node8035 = (inp[12]) ? node8073 : node8036;
									assign node8036 = (inp[13]) ? node8052 : node8037;
										assign node8037 = (inp[3]) ? node8045 : node8038;
											assign node8038 = (inp[8]) ? 16'b0000000111111111 : node8039;
												assign node8039 = (inp[1]) ? 16'b0000001111111111 : node8040;
													assign node8040 = (inp[7]) ? 16'b0000001111111111 : 16'b0000111111111111;
											assign node8045 = (inp[0]) ? node8049 : node8046;
												assign node8046 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node8049 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node8052 = (inp[4]) ? node8068 : node8053;
											assign node8053 = (inp[7]) ? node8063 : node8054;
												assign node8054 = (inp[1]) ? 16'b0000000001111111 : node8055;
													assign node8055 = (inp[3]) ? node8057 : 16'b0000001111111111;
														assign node8057 = (inp[0]) ? node8059 : 16'b0000000111111111;
															assign node8059 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8063 = (inp[10]) ? node8065 : 16'b0000000011111111;
													assign node8065 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8068 = (inp[0]) ? node8070 : 16'b0000000001111111;
												assign node8070 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node8073 = (inp[0]) ? node8109 : node8074;
										assign node8074 = (inp[10]) ? node8090 : node8075;
											assign node8075 = (inp[8]) ? node8085 : node8076;
												assign node8076 = (inp[4]) ? 16'b0000000001111111 : node8077;
													assign node8077 = (inp[7]) ? node8081 : node8078;
														assign node8078 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8081 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8085 = (inp[1]) ? 16'b0000000001111111 : node8086;
													assign node8086 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8090 = (inp[1]) ? node8098 : node8091;
												assign node8091 = (inp[3]) ? 16'b0000000001111111 : node8092;
													assign node8092 = (inp[7]) ? node8094 : 16'b0000000011111111;
														assign node8094 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8098 = (inp[4]) ? node8104 : node8099;
													assign node8099 = (inp[13]) ? node8101 : 16'b0000000001111111;
														assign node8101 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node8104 = (inp[7]) ? node8106 : 16'b0000000000111111;
														assign node8106 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node8109 = (inp[3]) ? node8117 : node8110;
											assign node8110 = (inp[8]) ? node8114 : node8111;
												assign node8111 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8114 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8117 = (inp[7]) ? node8121 : node8118;
												assign node8118 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node8121 = (inp[13]) ? node8123 : 16'b0000000000001111;
													assign node8123 = (inp[10]) ? 16'b0000000000011111 : node8124;
														assign node8124 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node8128 = (inp[10]) ? node8210 : node8129;
								assign node8129 = (inp[5]) ? node8161 : node8130;
									assign node8130 = (inp[4]) ? node8144 : node8131;
										assign node8131 = (inp[3]) ? node8139 : node8132;
											assign node8132 = (inp[0]) ? node8136 : node8133;
												assign node8133 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8136 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8139 = (inp[12]) ? node8141 : 16'b0000000011111111;
												assign node8141 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node8144 = (inp[7]) ? node8154 : node8145;
											assign node8145 = (inp[0]) ? node8149 : node8146;
												assign node8146 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8149 = (inp[12]) ? node8151 : 16'b0000000011111111;
													assign node8151 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000011111111;
											assign node8154 = (inp[1]) ? node8158 : node8155;
												assign node8155 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8158 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
									assign node8161 = (inp[4]) ? node8189 : node8162;
										assign node8162 = (inp[7]) ? node8182 : node8163;
											assign node8163 = (inp[1]) ? node8171 : node8164;
												assign node8164 = (inp[8]) ? 16'b0000000011111111 : node8165;
													assign node8165 = (inp[0]) ? 16'b0000000111111111 : node8166;
														assign node8166 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8171 = (inp[13]) ? node8175 : node8172;
													assign node8172 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8175 = (inp[12]) ? node8179 : node8176;
														assign node8176 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8179 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8182 = (inp[0]) ? 16'b0000000000111111 : node8183;
												assign node8183 = (inp[8]) ? node8185 : 16'b0000000011111111;
													assign node8185 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000000111111;
										assign node8189 = (inp[1]) ? node8205 : node8190;
											assign node8190 = (inp[3]) ? node8194 : node8191;
												assign node8191 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8194 = (inp[0]) ? node8200 : node8195;
													assign node8195 = (inp[12]) ? node8197 : 16'b0000000001111111;
														assign node8197 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node8200 = (inp[13]) ? 16'b0000000000111111 : node8201;
														assign node8201 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8205 = (inp[12]) ? node8207 : 16'b0000000000111111;
												assign node8207 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node8210 = (inp[13]) ? node8252 : node8211;
									assign node8211 = (inp[1]) ? node8231 : node8212;
										assign node8212 = (inp[7]) ? node8220 : node8213;
											assign node8213 = (inp[0]) ? node8217 : node8214;
												assign node8214 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8217 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8220 = (inp[0]) ? node8228 : node8221;
												assign node8221 = (inp[4]) ? 16'b0000000001111111 : node8222;
													assign node8222 = (inp[8]) ? node8224 : 16'b0000000011111111;
														assign node8224 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8228 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node8231 = (inp[5]) ? node8241 : node8232;
											assign node8232 = (inp[4]) ? 16'b0000000000111111 : node8233;
												assign node8233 = (inp[7]) ? node8235 : 16'b0000001111111111;
													assign node8235 = (inp[3]) ? node8237 : 16'b0000000001111111;
														assign node8237 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8241 = (inp[3]) ? node8243 : 16'b0000000000111111;
												assign node8243 = (inp[12]) ? node8245 : 16'b0000000000001111;
													assign node8245 = (inp[7]) ? 16'b0000000000011111 : node8246;
														assign node8246 = (inp[4]) ? node8248 : 16'b0000000000111111;
															assign node8248 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node8252 = (inp[8]) ? node8262 : node8253;
										assign node8253 = (inp[4]) ? node8255 : 16'b0000000001111111;
											assign node8255 = (inp[3]) ? node8259 : node8256;
												assign node8256 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8259 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node8262 = (inp[7]) ? node8274 : node8263;
											assign node8263 = (inp[3]) ? node8265 : 16'b0000000001111111;
												assign node8265 = (inp[5]) ? node8271 : node8266;
													assign node8266 = (inp[1]) ? node8268 : 16'b0000000000111111;
														assign node8268 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node8271 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000001111;
											assign node8274 = (inp[0]) ? node8278 : node8275;
												assign node8275 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8278 = (inp[12]) ? 16'b0000000000001111 : node8279;
													assign node8279 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node8283 = (inp[5]) ? node8435 : node8284;
							assign node8284 = (inp[3]) ? node8348 : node8285;
								assign node8285 = (inp[0]) ? node8325 : node8286;
									assign node8286 = (inp[8]) ? node8302 : node8287;
										assign node8287 = (inp[1]) ? node8297 : node8288;
											assign node8288 = (inp[13]) ? node8292 : node8289;
												assign node8289 = (inp[12]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node8292 = (inp[15]) ? node8294 : 16'b0000000111111111;
													assign node8294 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8297 = (inp[12]) ? node8299 : 16'b0000000011111111;
												assign node8299 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node8302 = (inp[13]) ? node8314 : node8303;
											assign node8303 = (inp[12]) ? node8307 : node8304;
												assign node8304 = (inp[10]) ? 16'b0000000001111111 : 16'b0000001111111111;
												assign node8307 = (inp[1]) ? 16'b0000000001111111 : node8308;
													assign node8308 = (inp[4]) ? node8310 : 16'b0000000011111111;
														assign node8310 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8314 = (inp[7]) ? node8322 : node8315;
												assign node8315 = (inp[12]) ? 16'b0000000001111111 : node8316;
													assign node8316 = (inp[15]) ? node8318 : 16'b0000000011111111;
														assign node8318 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8322 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node8325 = (inp[7]) ? node8331 : node8326;
										assign node8326 = (inp[12]) ? 16'b0000000001111111 : node8327;
											assign node8327 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node8331 = (inp[8]) ? node8339 : node8332;
											assign node8332 = (inp[15]) ? node8334 : 16'b0000000011111111;
												assign node8334 = (inp[1]) ? node8336 : 16'b0000000001111111;
													assign node8336 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8339 = (inp[10]) ? node8341 : 16'b0000000001111111;
												assign node8341 = (inp[1]) ? node8345 : node8342;
													assign node8342 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node8345 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node8348 = (inp[8]) ? node8396 : node8349;
									assign node8349 = (inp[0]) ? node8369 : node8350;
										assign node8350 = (inp[7]) ? node8360 : node8351;
											assign node8351 = (inp[4]) ? node8355 : node8352;
												assign node8352 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8355 = (inp[13]) ? node8357 : 16'b0000000011111111;
													assign node8357 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8360 = (inp[1]) ? node8364 : node8361;
												assign node8361 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8364 = (inp[13]) ? node8366 : 16'b0000000001111111;
													assign node8366 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node8369 = (inp[10]) ? node8385 : node8370;
											assign node8370 = (inp[4]) ? node8378 : node8371;
												assign node8371 = (inp[15]) ? 16'b0000000001111111 : node8372;
													assign node8372 = (inp[1]) ? 16'b0000000011111111 : node8373;
														assign node8373 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8378 = (inp[1]) ? 16'b0000000000111111 : node8379;
													assign node8379 = (inp[13]) ? node8381 : 16'b0000000011111111;
														assign node8381 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8385 = (inp[4]) ? node8393 : node8386;
												assign node8386 = (inp[7]) ? 16'b0000000000011111 : node8387;
													assign node8387 = (inp[12]) ? node8389 : 16'b0000000001111111;
														assign node8389 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8393 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node8396 = (inp[12]) ? node8414 : node8397;
										assign node8397 = (inp[10]) ? node8405 : node8398;
											assign node8398 = (inp[7]) ? node8400 : 16'b0000000011111111;
												assign node8400 = (inp[13]) ? 16'b0000000000111111 : node8401;
													assign node8401 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8405 = (inp[13]) ? node8409 : node8406;
												assign node8406 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node8409 = (inp[7]) ? node8411 : 16'b0000000000111111;
													assign node8411 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node8414 = (inp[15]) ? node8424 : node8415;
											assign node8415 = (inp[0]) ? node8421 : node8416;
												assign node8416 = (inp[4]) ? node8418 : 16'b0000000001111111;
													assign node8418 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8421 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node8424 = (inp[0]) ? 16'b0000000000001111 : node8425;
												assign node8425 = (inp[1]) ? node8431 : node8426;
													assign node8426 = (inp[7]) ? 16'b0000000000111111 : node8427;
														assign node8427 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node8431 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000011111;
							assign node8435 = (inp[4]) ? node8517 : node8436;
								assign node8436 = (inp[7]) ? node8468 : node8437;
									assign node8437 = (inp[8]) ? node8449 : node8438;
										assign node8438 = (inp[0]) ? 16'b0000000000111111 : node8439;
											assign node8439 = (inp[15]) ? node8445 : node8440;
												assign node8440 = (inp[12]) ? 16'b0000000011111111 : node8441;
													assign node8441 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8445 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node8449 = (inp[1]) ? node8459 : node8450;
											assign node8450 = (inp[3]) ? 16'b0000000001111111 : node8451;
												assign node8451 = (inp[13]) ? node8455 : node8452;
													assign node8452 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node8455 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8459 = (inp[10]) ? node8465 : node8460;
												assign node8460 = (inp[12]) ? node8462 : 16'b0000000111111111;
													assign node8462 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8465 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node8468 = (inp[10]) ? node8494 : node8469;
										assign node8469 = (inp[12]) ? node8487 : node8470;
											assign node8470 = (inp[0]) ? node8482 : node8471;
												assign node8471 = (inp[1]) ? node8477 : node8472;
													assign node8472 = (inp[13]) ? node8474 : 16'b0000000011111111;
														assign node8474 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8477 = (inp[8]) ? 16'b0000000001111111 : node8478;
														assign node8478 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8482 = (inp[1]) ? 16'b0000000000111111 : node8483;
													assign node8483 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8487 = (inp[13]) ? node8489 : 16'b0000000000111111;
												assign node8489 = (inp[1]) ? 16'b0000000000011111 : node8490;
													assign node8490 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000011111;
										assign node8494 = (inp[8]) ? node8506 : node8495;
											assign node8495 = (inp[0]) ? node8499 : node8496;
												assign node8496 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8499 = (inp[12]) ? 16'b0000000000011111 : node8500;
													assign node8500 = (inp[3]) ? node8502 : 16'b0000000000111111;
														assign node8502 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node8506 = (inp[13]) ? node8512 : node8507;
												assign node8507 = (inp[1]) ? 16'b0000000000001111 : node8508;
													assign node8508 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8512 = (inp[12]) ? 16'b0000000000001111 : node8513;
													assign node8513 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node8517 = (inp[15]) ? node8559 : node8518;
									assign node8518 = (inp[3]) ? node8534 : node8519;
										assign node8519 = (inp[1]) ? node8531 : node8520;
											assign node8520 = (inp[7]) ? node8528 : node8521;
												assign node8521 = (inp[8]) ? 16'b0000000000111111 : node8522;
													assign node8522 = (inp[10]) ? 16'b0000000011111111 : node8523;
														assign node8523 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8528 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8531 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000000011111;
										assign node8534 = (inp[0]) ? node8550 : node8535;
											assign node8535 = (inp[7]) ? node8543 : node8536;
												assign node8536 = (inp[12]) ? 16'b0000000000111111 : node8537;
													assign node8537 = (inp[10]) ? node8539 : 16'b0000000001111111;
														assign node8539 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8543 = (inp[1]) ? node8545 : 16'b0000000001111111;
													assign node8545 = (inp[13]) ? node8547 : 16'b0000000000011111;
														assign node8547 = (inp[8]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node8550 = (inp[8]) ? node8554 : node8551;
												assign node8551 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000011111;
												assign node8554 = (inp[13]) ? 16'b0000000000001111 : node8555;
													assign node8555 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node8559 = (inp[1]) ? node8589 : node8560;
										assign node8560 = (inp[3]) ? node8578 : node8561;
											assign node8561 = (inp[13]) ? node8575 : node8562;
												assign node8562 = (inp[12]) ? node8568 : node8563;
													assign node8563 = (inp[7]) ? node8565 : 16'b0000000011111111;
														assign node8565 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node8568 = (inp[7]) ? node8572 : node8569;
														assign node8569 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node8572 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node8575 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node8578 = (inp[10]) ? node8580 : 16'b0000000000011111;
												assign node8580 = (inp[12]) ? 16'b0000000000000111 : node8581;
													assign node8581 = (inp[7]) ? 16'b0000000000001111 : node8582;
														assign node8582 = (inp[13]) ? node8584 : 16'b0000000000011111;
															assign node8584 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node8589 = (inp[12]) ? node8597 : node8590;
											assign node8590 = (inp[0]) ? 16'b0000000000001111 : node8591;
												assign node8591 = (inp[7]) ? 16'b0000000000011111 : node8592;
													assign node8592 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node8597 = (inp[13]) ? node8599 : 16'b0000000000001111;
												assign node8599 = (inp[0]) ? node8609 : node8600;
													assign node8600 = (inp[7]) ? node8604 : node8601;
														assign node8601 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node8604 = (inp[8]) ? node8606 : 16'b0000000000011111;
															assign node8606 = (inp[3]) ? 16'b0000000000000111 : 16'b0000000000000111;
													assign node8609 = (inp[10]) ? node8611 : 16'b0000000000000111;
														assign node8611 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000001111;
			assign node8614 = (inp[3]) ? node10040 : node8615;
				assign node8615 = (inp[15]) ? node9345 : node8616;
					assign node8616 = (inp[10]) ? node8990 : node8617;
						assign node8617 = (inp[12]) ? node8807 : node8618;
							assign node8618 = (inp[13]) ? node8708 : node8619;
								assign node8619 = (inp[11]) ? node8669 : node8620;
									assign node8620 = (inp[7]) ? node8646 : node8621;
										assign node8621 = (inp[5]) ? node8633 : node8622;
											assign node8622 = (inp[1]) ? node8630 : node8623;
												assign node8623 = (inp[4]) ? node8625 : 16'b0000111111111111;
													assign node8625 = (inp[14]) ? 16'b0000011111111111 : node8626;
														assign node8626 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node8630 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node8633 = (inp[8]) ? node8643 : node8634;
												assign node8634 = (inp[1]) ? node8638 : node8635;
													assign node8635 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node8638 = (inp[14]) ? 16'b0000001111111111 : node8639;
														assign node8639 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8643 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node8646 = (inp[14]) ? node8658 : node8647;
											assign node8647 = (inp[1]) ? node8655 : node8648;
												assign node8648 = (inp[8]) ? 16'b0000001111111111 : node8649;
													assign node8649 = (inp[5]) ? 16'b0000011111111111 : node8650;
														assign node8650 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node8655 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node8658 = (inp[4]) ? node8664 : node8659;
												assign node8659 = (inp[8]) ? 16'b0000000111111111 : node8660;
													assign node8660 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8664 = (inp[5]) ? 16'b0000000011111111 : node8665;
													assign node8665 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node8669 = (inp[0]) ? node8691 : node8670;
										assign node8670 = (inp[4]) ? node8678 : node8671;
											assign node8671 = (inp[1]) ? node8673 : 16'b0000011111111111;
												assign node8673 = (inp[9]) ? 16'b0000001111111111 : node8674;
													assign node8674 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node8678 = (inp[5]) ? node8686 : node8679;
												assign node8679 = (inp[8]) ? node8683 : node8680;
													assign node8680 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8683 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8686 = (inp[9]) ? 16'b0000000011111111 : node8687;
													assign node8687 = (inp[1]) ? 16'b0000000011111111 : 16'b0000001111111111;
										assign node8691 = (inp[9]) ? node8701 : node8692;
											assign node8692 = (inp[14]) ? node8696 : node8693;
												assign node8693 = (inp[1]) ? 16'b0000001111111111 : 16'b0000000111111111;
												assign node8696 = (inp[8]) ? 16'b0000000011111111 : node8697;
													assign node8697 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node8701 = (inp[14]) ? node8705 : node8702;
												assign node8702 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8705 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
								assign node8708 = (inp[1]) ? node8750 : node8709;
									assign node8709 = (inp[7]) ? node8737 : node8710;
										assign node8710 = (inp[5]) ? node8718 : node8711;
											assign node8711 = (inp[4]) ? 16'b0000001111111111 : node8712;
												assign node8712 = (inp[0]) ? node8714 : 16'b0000111111111111;
													assign node8714 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node8718 = (inp[4]) ? node8728 : node8719;
												assign node8719 = (inp[9]) ? node8721 : 16'b0000001111111111;
													assign node8721 = (inp[14]) ? 16'b0000000111111111 : node8722;
														assign node8722 = (inp[8]) ? node8724 : 16'b0000011111111111;
															assign node8724 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8728 = (inp[11]) ? 16'b0000000011111111 : node8729;
													assign node8729 = (inp[14]) ? node8733 : node8730;
														assign node8730 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8733 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node8737 = (inp[14]) ? node8743 : node8738;
											assign node8738 = (inp[11]) ? node8740 : 16'b0000001111111111;
												assign node8740 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8743 = (inp[11]) ? node8747 : node8744;
												assign node8744 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8747 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node8750 = (inp[9]) ? node8778 : node8751;
										assign node8751 = (inp[11]) ? node8769 : node8752;
											assign node8752 = (inp[14]) ? node8762 : node8753;
												assign node8753 = (inp[4]) ? node8757 : node8754;
													assign node8754 = (inp[7]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node8757 = (inp[0]) ? 16'b0000000111111111 : node8758;
														assign node8758 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8762 = (inp[5]) ? 16'b0000000001111111 : node8763;
													assign node8763 = (inp[8]) ? node8765 : 16'b0000001111111111;
														assign node8765 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8769 = (inp[8]) ? node8773 : node8770;
												assign node8770 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8773 = (inp[0]) ? node8775 : 16'b0000000011111111;
													assign node8775 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node8778 = (inp[5]) ? node8796 : node8779;
											assign node8779 = (inp[11]) ? node8787 : node8780;
												assign node8780 = (inp[7]) ? node8782 : 16'b0000000111111111;
													assign node8782 = (inp[14]) ? 16'b0000000001111111 : node8783;
														assign node8783 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8787 = (inp[7]) ? node8791 : node8788;
													assign node8788 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8791 = (inp[14]) ? node8793 : 16'b0000000001111111;
														assign node8793 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node8796 = (inp[4]) ? node8800 : node8797;
												assign node8797 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8800 = (inp[14]) ? node8802 : 16'b0000000000111111;
													assign node8802 = (inp[0]) ? node8804 : 16'b0000000000111111;
														assign node8804 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node8807 = (inp[4]) ? node8897 : node8808;
								assign node8808 = (inp[1]) ? node8850 : node8809;
									assign node8809 = (inp[14]) ? node8835 : node8810;
										assign node8810 = (inp[8]) ? node8822 : node8811;
											assign node8811 = (inp[5]) ? node8815 : node8812;
												assign node8812 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node8815 = (inp[0]) ? 16'b0000000111111111 : node8816;
													assign node8816 = (inp[11]) ? 16'b0000001111111111 : node8817;
														assign node8817 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node8822 = (inp[13]) ? node8830 : node8823;
												assign node8823 = (inp[11]) ? node8827 : node8824;
													assign node8824 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8827 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node8830 = (inp[0]) ? node8832 : 16'b0000000111111111;
													assign node8832 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node8835 = (inp[8]) ? node8845 : node8836;
											assign node8836 = (inp[11]) ? node8842 : node8837;
												assign node8837 = (inp[7]) ? 16'b0000000111111111 : node8838;
													assign node8838 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8842 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8845 = (inp[11]) ? node8847 : 16'b0000000011111111;
												assign node8847 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node8850 = (inp[7]) ? node8874 : node8851;
										assign node8851 = (inp[13]) ? node8865 : node8852;
											assign node8852 = (inp[8]) ? node8858 : node8853;
												assign node8853 = (inp[11]) ? node8855 : 16'b0000001111111111;
													assign node8855 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node8858 = (inp[9]) ? node8860 : 16'b0000000111111111;
													assign node8860 = (inp[5]) ? node8862 : 16'b0000000111111111;
														assign node8862 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8865 = (inp[11]) ? node8869 : node8866;
												assign node8866 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node8869 = (inp[5]) ? 16'b0000000011111111 : node8870;
													assign node8870 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node8874 = (inp[5]) ? node8886 : node8875;
											assign node8875 = (inp[11]) ? node8879 : node8876;
												assign node8876 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8879 = (inp[14]) ? 16'b0000000011111111 : node8880;
													assign node8880 = (inp[0]) ? 16'b0000000011111111 : node8881;
														assign node8881 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8886 = (inp[11]) ? node8892 : node8887;
												assign node8887 = (inp[0]) ? 16'b0000000001111111 : node8888;
													assign node8888 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8892 = (inp[14]) ? node8894 : 16'b0000000001111111;
													assign node8894 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node8897 = (inp[11]) ? node8939 : node8898;
									assign node8898 = (inp[5]) ? node8920 : node8899;
										assign node8899 = (inp[9]) ? node8911 : node8900;
											assign node8900 = (inp[0]) ? node8908 : node8901;
												assign node8901 = (inp[1]) ? node8903 : 16'b0000001111111111;
													assign node8903 = (inp[8]) ? node8905 : 16'b0000000111111111;
														assign node8905 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8908 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8911 = (inp[1]) ? node8917 : node8912;
												assign node8912 = (inp[7]) ? node8914 : 16'b0000000111111111;
													assign node8914 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8917 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node8920 = (inp[0]) ? node8932 : node8921;
											assign node8921 = (inp[13]) ? node8929 : node8922;
												assign node8922 = (inp[14]) ? node8924 : 16'b0000000111111111;
													assign node8924 = (inp[7]) ? node8926 : 16'b0000000111111111;
														assign node8926 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8929 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8932 = (inp[8]) ? node8934 : 16'b0000000011111111;
												assign node8934 = (inp[14]) ? node8936 : 16'b0000000001111111;
													assign node8936 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node8939 = (inp[7]) ? node8963 : node8940;
										assign node8940 = (inp[8]) ? node8952 : node8941;
											assign node8941 = (inp[9]) ? node8945 : node8942;
												assign node8942 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8945 = (inp[5]) ? 16'b0000000001111111 : node8946;
													assign node8946 = (inp[13]) ? 16'b0000000011111111 : node8947;
														assign node8947 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8952 = (inp[9]) ? node8960 : node8953;
												assign node8953 = (inp[13]) ? node8955 : 16'b0000000011111111;
													assign node8955 = (inp[1]) ? node8957 : 16'b0000000001111111;
														assign node8957 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8960 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node8963 = (inp[14]) ? node8975 : node8964;
											assign node8964 = (inp[13]) ? 16'b0000000000111111 : node8965;
												assign node8965 = (inp[0]) ? node8969 : node8966;
													assign node8966 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8969 = (inp[5]) ? node8971 : 16'b0000000001111111;
														assign node8971 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8975 = (inp[8]) ? node8985 : node8976;
												assign node8976 = (inp[5]) ? 16'b0000000000111111 : node8977;
													assign node8977 = (inp[1]) ? node8981 : node8978;
														assign node8978 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8981 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8985 = (inp[1]) ? node8987 : 16'b0000000000111111;
													assign node8987 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node8990 = (inp[5]) ? node9146 : node8991;
							assign node8991 = (inp[7]) ? node9081 : node8992;
								assign node8992 = (inp[4]) ? node9042 : node8993;
									assign node8993 = (inp[9]) ? node9023 : node8994;
										assign node8994 = (inp[0]) ? node9010 : node8995;
											assign node8995 = (inp[8]) ? node9005 : node8996;
												assign node8996 = (inp[13]) ? node8998 : 16'b0000011111111111;
													assign node8998 = (inp[11]) ? 16'b0000001111111111 : node8999;
														assign node8999 = (inp[14]) ? 16'b0000001111111111 : node9000;
															assign node9000 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node9005 = (inp[11]) ? node9007 : 16'b0000000111111111;
													assign node9007 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node9010 = (inp[12]) ? node9018 : node9011;
												assign node9011 = (inp[14]) ? node9015 : node9012;
													assign node9012 = (inp[8]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node9015 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9018 = (inp[14]) ? 16'b0000000011111111 : node9019;
													assign node9019 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node9023 = (inp[13]) ? node9033 : node9024;
											assign node9024 = (inp[14]) ? node9030 : node9025;
												assign node9025 = (inp[11]) ? node9027 : 16'b0000011111111111;
													assign node9027 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9030 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9033 = (inp[12]) ? node9037 : node9034;
												assign node9034 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9037 = (inp[14]) ? node9039 : 16'b0000000011111111;
													assign node9039 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node9042 = (inp[11]) ? node9060 : node9043;
										assign node9043 = (inp[1]) ? node9055 : node9044;
											assign node9044 = (inp[14]) ? node9050 : node9045;
												assign node9045 = (inp[9]) ? node9047 : 16'b0000001111111111;
													assign node9047 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9050 = (inp[9]) ? node9052 : 16'b0000000111111111;
													assign node9052 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node9055 = (inp[14]) ? node9057 : 16'b0000000111111111;
												assign node9057 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node9060 = (inp[0]) ? node9070 : node9061;
											assign node9061 = (inp[9]) ? node9065 : node9062;
												assign node9062 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9065 = (inp[8]) ? node9067 : 16'b0000000011111111;
													assign node9067 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9070 = (inp[9]) ? node9078 : node9071;
												assign node9071 = (inp[13]) ? node9073 : 16'b0000000011111111;
													assign node9073 = (inp[12]) ? 16'b0000000001111111 : node9074;
														assign node9074 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9078 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node9081 = (inp[13]) ? node9117 : node9082;
									assign node9082 = (inp[12]) ? node9102 : node9083;
										assign node9083 = (inp[14]) ? node9091 : node9084;
											assign node9084 = (inp[11]) ? 16'b0000000111111111 : node9085;
												assign node9085 = (inp[1]) ? 16'b0000001111111111 : node9086;
													assign node9086 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node9091 = (inp[8]) ? node9097 : node9092;
												assign node9092 = (inp[0]) ? node9094 : 16'b0000000111111111;
													assign node9094 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9097 = (inp[9]) ? 16'b0000000011111111 : node9098;
													assign node9098 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node9102 = (inp[8]) ? node9108 : node9103;
											assign node9103 = (inp[14]) ? 16'b0000000001111111 : node9104;
												assign node9104 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node9108 = (inp[9]) ? 16'b0000000000111111 : node9109;
												assign node9109 = (inp[1]) ? node9111 : 16'b0000000111111111;
													assign node9111 = (inp[0]) ? 16'b0000000001111111 : node9112;
														assign node9112 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node9117 = (inp[9]) ? node9135 : node9118;
										assign node9118 = (inp[1]) ? node9130 : node9119;
											assign node9119 = (inp[0]) ? 16'b0000000001111111 : node9120;
												assign node9120 = (inp[12]) ? node9124 : node9121;
													assign node9121 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9124 = (inp[11]) ? node9126 : 16'b0000000011111111;
														assign node9126 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9130 = (inp[12]) ? node9132 : 16'b0000000011111111;
												assign node9132 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node9135 = (inp[11]) ? node9143 : node9136;
											assign node9136 = (inp[1]) ? node9138 : 16'b0000000001111111;
												assign node9138 = (inp[14]) ? 16'b0000000000111111 : node9139;
													assign node9139 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9143 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node9146 = (inp[0]) ? node9250 : node9147;
								assign node9147 = (inp[12]) ? node9211 : node9148;
									assign node9148 = (inp[14]) ? node9186 : node9149;
										assign node9149 = (inp[4]) ? node9163 : node9150;
											assign node9150 = (inp[8]) ? node9160 : node9151;
												assign node9151 = (inp[1]) ? node9153 : 16'b0000011111111111;
													assign node9153 = (inp[7]) ? 16'b0000000111111111 : node9154;
														assign node9154 = (inp[9]) ? node9156 : 16'b0000001111111111;
															assign node9156 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9160 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9163 = (inp[11]) ? node9171 : node9164;
												assign node9164 = (inp[13]) ? 16'b0000000011111111 : node9165;
													assign node9165 = (inp[7]) ? 16'b0000000111111111 : node9166;
														assign node9166 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9171 = (inp[8]) ? node9177 : node9172;
													assign node9172 = (inp[1]) ? node9174 : 16'b0000000011111111;
														assign node9174 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9177 = (inp[13]) ? node9183 : node9178;
														assign node9178 = (inp[7]) ? 16'b0000000001111111 : node9179;
															assign node9179 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node9183 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node9186 = (inp[1]) ? node9202 : node9187;
											assign node9187 = (inp[8]) ? node9197 : node9188;
												assign node9188 = (inp[11]) ? node9192 : node9189;
													assign node9189 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9192 = (inp[9]) ? node9194 : 16'b0000000011111111;
														assign node9194 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9197 = (inp[7]) ? node9199 : 16'b0000000001111111;
													assign node9199 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9202 = (inp[9]) ? node9208 : node9203;
												assign node9203 = (inp[13]) ? node9205 : 16'b0000000011111111;
													assign node9205 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9208 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node9211 = (inp[4]) ? node9223 : node9212;
										assign node9212 = (inp[7]) ? node9214 : 16'b0000000011111111;
											assign node9214 = (inp[11]) ? 16'b0000000000111111 : node9215;
												assign node9215 = (inp[13]) ? node9217 : 16'b0000000011111111;
													assign node9217 = (inp[8]) ? 16'b0000000001111111 : node9218;
														assign node9218 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node9223 = (inp[11]) ? node9233 : node9224;
											assign node9224 = (inp[7]) ? 16'b0000000000111111 : node9225;
												assign node9225 = (inp[1]) ? 16'b0000000001111111 : node9226;
													assign node9226 = (inp[8]) ? node9228 : 16'b0000000011111111;
														assign node9228 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9233 = (inp[14]) ? node9245 : node9234;
												assign node9234 = (inp[8]) ? node9240 : node9235;
													assign node9235 = (inp[1]) ? 16'b0000000001111111 : node9236;
														assign node9236 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9240 = (inp[7]) ? node9242 : 16'b0000000001111111;
														assign node9242 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node9245 = (inp[7]) ? node9247 : 16'b0000000000111111;
													assign node9247 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000000011111;
								assign node9250 = (inp[14]) ? node9302 : node9251;
									assign node9251 = (inp[1]) ? node9277 : node9252;
										assign node9252 = (inp[8]) ? node9260 : node9253;
											assign node9253 = (inp[11]) ? 16'b0000000011111111 : node9254;
												assign node9254 = (inp[12]) ? 16'b0000000011111111 : node9255;
													assign node9255 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9260 = (inp[4]) ? node9272 : node9261;
												assign node9261 = (inp[11]) ? node9265 : node9262;
													assign node9262 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9265 = (inp[13]) ? 16'b0000000001111111 : node9266;
														assign node9266 = (inp[9]) ? node9268 : 16'b0000000111111111;
															assign node9268 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9272 = (inp[11]) ? node9274 : 16'b0000000001111111;
													assign node9274 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node9277 = (inp[8]) ? node9291 : node9278;
											assign node9278 = (inp[11]) ? node9288 : node9279;
												assign node9279 = (inp[4]) ? 16'b0000000001111111 : node9280;
													assign node9280 = (inp[12]) ? node9282 : 16'b0000000011111111;
														assign node9282 = (inp[9]) ? 16'b0000000001111111 : node9283;
															assign node9283 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9288 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000011111111;
											assign node9291 = (inp[7]) ? node9295 : node9292;
												assign node9292 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9295 = (inp[12]) ? node9297 : 16'b0000000000111111;
													assign node9297 = (inp[13]) ? node9299 : 16'b0000000000001111;
														assign node9299 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node9302 = (inp[4]) ? node9320 : node9303;
										assign node9303 = (inp[1]) ? node9311 : node9304;
											assign node9304 = (inp[9]) ? node9306 : 16'b0000000011111111;
												assign node9306 = (inp[7]) ? 16'b0000000000111111 : node9307;
													assign node9307 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9311 = (inp[11]) ? node9315 : node9312;
												assign node9312 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9315 = (inp[7]) ? node9317 : 16'b0000000000111111;
													assign node9317 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000001111;
										assign node9320 = (inp[8]) ? node9336 : node9321;
											assign node9321 = (inp[13]) ? node9327 : node9322;
												assign node9322 = (inp[11]) ? node9324 : 16'b0000000001111111;
													assign node9324 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node9327 = (inp[9]) ? 16'b0000000000011111 : node9328;
													assign node9328 = (inp[1]) ? node9330 : 16'b0000000000111111;
														assign node9330 = (inp[12]) ? 16'b0000000000011111 : node9331;
															assign node9331 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node9336 = (inp[13]) ? node9338 : 16'b0000000000011111;
												assign node9338 = (inp[7]) ? node9340 : 16'b0000000000011111;
													assign node9340 = (inp[11]) ? 16'b0000000000001111 : node9341;
														assign node9341 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node9345 = (inp[11]) ? node9679 : node9346;
						assign node9346 = (inp[8]) ? node9502 : node9347;
							assign node9347 = (inp[14]) ? node9425 : node9348;
								assign node9348 = (inp[13]) ? node9382 : node9349;
									assign node9349 = (inp[12]) ? node9367 : node9350;
										assign node9350 = (inp[0]) ? node9364 : node9351;
											assign node9351 = (inp[9]) ? node9357 : node9352;
												assign node9352 = (inp[5]) ? node9354 : 16'b0000111111111111;
													assign node9354 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node9357 = (inp[5]) ? 16'b0000000111111111 : node9358;
													assign node9358 = (inp[4]) ? node9360 : 16'b0000001111111111;
														assign node9360 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node9364 = (inp[7]) ? 16'b0000001111111111 : 16'b0000000111111111;
										assign node9367 = (inp[1]) ? node9369 : 16'b0000000111111111;
											assign node9369 = (inp[9]) ? node9379 : node9370;
												assign node9370 = (inp[5]) ? node9374 : node9371;
													assign node9371 = (inp[0]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node9374 = (inp[7]) ? node9376 : 16'b0000000011111111;
														assign node9376 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9379 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node9382 = (inp[0]) ? node9406 : node9383;
										assign node9383 = (inp[7]) ? node9397 : node9384;
											assign node9384 = (inp[4]) ? node9394 : node9385;
												assign node9385 = (inp[12]) ? node9389 : node9386;
													assign node9386 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9389 = (inp[10]) ? 16'b0000000011111111 : node9390;
														assign node9390 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9394 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9397 = (inp[4]) ? node9403 : node9398;
												assign node9398 = (inp[1]) ? node9400 : 16'b0000000011111111;
													assign node9400 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9403 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node9406 = (inp[12]) ? node9416 : node9407;
											assign node9407 = (inp[9]) ? node9411 : node9408;
												assign node9408 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node9411 = (inp[5]) ? node9413 : 16'b0000000011111111;
													assign node9413 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9416 = (inp[9]) ? node9422 : node9417;
												assign node9417 = (inp[7]) ? node9419 : 16'b0000000001111111;
													assign node9419 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node9422 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000001111111;
								assign node9425 = (inp[10]) ? node9471 : node9426;
									assign node9426 = (inp[12]) ? node9448 : node9427;
										assign node9427 = (inp[9]) ? node9441 : node9428;
											assign node9428 = (inp[7]) ? node9436 : node9429;
												assign node9429 = (inp[5]) ? node9433 : node9430;
													assign node9430 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9433 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9436 = (inp[1]) ? 16'b0000000011111111 : node9437;
													assign node9437 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node9441 = (inp[0]) ? node9443 : 16'b0000000111111111;
												assign node9443 = (inp[4]) ? 16'b0000000001111111 : node9444;
													assign node9444 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node9448 = (inp[7]) ? node9458 : node9449;
											assign node9449 = (inp[9]) ? node9455 : node9450;
												assign node9450 = (inp[13]) ? 16'b0000000011111111 : node9451;
													assign node9451 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9455 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9458 = (inp[5]) ? node9466 : node9459;
												assign node9459 = (inp[9]) ? 16'b0000000001111111 : node9460;
													assign node9460 = (inp[1]) ? node9462 : 16'b0000000011111111;
														assign node9462 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9466 = (inp[1]) ? node9468 : 16'b0000000001111111;
													assign node9468 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node9471 = (inp[5]) ? node9491 : node9472;
										assign node9472 = (inp[13]) ? node9484 : node9473;
											assign node9473 = (inp[1]) ? node9477 : node9474;
												assign node9474 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9477 = (inp[7]) ? node9479 : 16'b0000000011111111;
													assign node9479 = (inp[12]) ? 16'b0000000001111111 : node9480;
														assign node9480 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9484 = (inp[0]) ? node9488 : node9485;
												assign node9485 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9488 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node9491 = (inp[9]) ? node9497 : node9492;
											assign node9492 = (inp[0]) ? node9494 : 16'b0000000001111111;
												assign node9494 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000011111;
											assign node9497 = (inp[0]) ? 16'b0000000000011111 : node9498;
												assign node9498 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node9502 = (inp[5]) ? node9600 : node9503;
								assign node9503 = (inp[10]) ? node9549 : node9504;
									assign node9504 = (inp[9]) ? node9524 : node9505;
										assign node9505 = (inp[0]) ? node9515 : node9506;
											assign node9506 = (inp[12]) ? node9508 : 16'b0000001111111111;
												assign node9508 = (inp[4]) ? node9510 : 16'b0000001111111111;
													assign node9510 = (inp[13]) ? 16'b0000000011111111 : node9511;
														assign node9511 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9515 = (inp[1]) ? 16'b0000000001111111 : node9516;
												assign node9516 = (inp[7]) ? 16'b0000000011111111 : node9517;
													assign node9517 = (inp[14]) ? node9519 : 16'b0000000111111111;
														assign node9519 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node9524 = (inp[12]) ? node9542 : node9525;
											assign node9525 = (inp[13]) ? node9537 : node9526;
												assign node9526 = (inp[4]) ? node9532 : node9527;
													assign node9527 = (inp[1]) ? node9529 : 16'b0000000111111111;
														assign node9529 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9532 = (inp[1]) ? 16'b0000000011111111 : node9533;
														assign node9533 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9537 = (inp[4]) ? node9539 : 16'b0000000011111111;
													assign node9539 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9542 = (inp[4]) ? node9546 : node9543;
												assign node9543 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9546 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000001111111;
									assign node9549 = (inp[13]) ? node9577 : node9550;
										assign node9550 = (inp[12]) ? node9564 : node9551;
											assign node9551 = (inp[9]) ? node9559 : node9552;
												assign node9552 = (inp[7]) ? node9556 : node9553;
													assign node9553 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node9556 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node9559 = (inp[14]) ? node9561 : 16'b0000000011111111;
													assign node9561 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9564 = (inp[1]) ? node9570 : node9565;
												assign node9565 = (inp[0]) ? 16'b0000000001111111 : node9566;
													assign node9566 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9570 = (inp[4]) ? node9572 : 16'b0000000111111111;
													assign node9572 = (inp[14]) ? node9574 : 16'b0000000001111111;
														assign node9574 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node9577 = (inp[14]) ? node9585 : node9578;
											assign node9578 = (inp[9]) ? node9582 : node9579;
												assign node9579 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9582 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9585 = (inp[7]) ? node9595 : node9586;
												assign node9586 = (inp[4]) ? node9590 : node9587;
													assign node9587 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node9590 = (inp[0]) ? node9592 : 16'b0000000000111111;
														assign node9592 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node9595 = (inp[0]) ? node9597 : 16'b0000000000011111;
													assign node9597 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node9600 = (inp[12]) ? node9648 : node9601;
									assign node9601 = (inp[1]) ? node9627 : node9602;
										assign node9602 = (inp[9]) ? node9612 : node9603;
											assign node9603 = (inp[0]) ? 16'b0000000011111111 : node9604;
												assign node9604 = (inp[7]) ? 16'b0000000011111111 : node9605;
													assign node9605 = (inp[10]) ? node9607 : 16'b0000000111111111;
														assign node9607 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node9612 = (inp[4]) ? node9618 : node9613;
												assign node9613 = (inp[0]) ? 16'b0000000001111111 : node9614;
													assign node9614 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9618 = (inp[14]) ? node9620 : 16'b0000000011111111;
													assign node9620 = (inp[10]) ? 16'b0000000000011111 : node9621;
														assign node9621 = (inp[7]) ? 16'b0000000000111111 : node9622;
															assign node9622 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node9627 = (inp[0]) ? node9639 : node9628;
											assign node9628 = (inp[9]) ? node9634 : node9629;
												assign node9629 = (inp[13]) ? 16'b0000000001111111 : node9630;
													assign node9630 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node9634 = (inp[7]) ? 16'b0000000000011111 : node9635;
													assign node9635 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9639 = (inp[4]) ? node9643 : node9640;
												assign node9640 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node9643 = (inp[14]) ? 16'b0000000000001111 : node9644;
													assign node9644 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node9648 = (inp[0]) ? node9668 : node9649;
										assign node9649 = (inp[14]) ? node9659 : node9650;
											assign node9650 = (inp[10]) ? node9652 : 16'b0000000011111111;
												assign node9652 = (inp[7]) ? node9654 : 16'b0000000001111111;
													assign node9654 = (inp[13]) ? node9656 : 16'b0000000001111111;
														assign node9656 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node9659 = (inp[13]) ? node9665 : node9660;
												assign node9660 = (inp[10]) ? 16'b0000000000111111 : node9661;
													assign node9661 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9665 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node9668 = (inp[1]) ? node9674 : node9669;
											assign node9669 = (inp[14]) ? 16'b0000000000001111 : node9670;
												assign node9670 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9674 = (inp[10]) ? node9676 : 16'b0000000000111111;
												assign node9676 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node9679 = (inp[8]) ? node9867 : node9680;
							assign node9680 = (inp[7]) ? node9774 : node9681;
								assign node9681 = (inp[0]) ? node9727 : node9682;
									assign node9682 = (inp[9]) ? node9698 : node9683;
										assign node9683 = (inp[1]) ? node9691 : node9684;
											assign node9684 = (inp[12]) ? 16'b0000000111111111 : node9685;
												assign node9685 = (inp[14]) ? 16'b0000001111111111 : node9686;
													assign node9686 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node9691 = (inp[12]) ? node9695 : node9692;
												assign node9692 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9695 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node9698 = (inp[5]) ? node9712 : node9699;
											assign node9699 = (inp[4]) ? node9707 : node9700;
												assign node9700 = (inp[12]) ? node9704 : node9701;
													assign node9701 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9704 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node9707 = (inp[12]) ? 16'b0000000001111111 : node9708;
													assign node9708 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node9712 = (inp[13]) ? node9718 : node9713;
												assign node9713 = (inp[1]) ? node9715 : 16'b0000000011111111;
													assign node9715 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9718 = (inp[1]) ? node9724 : node9719;
													assign node9719 = (inp[4]) ? node9721 : 16'b0000000001111111;
														assign node9721 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9724 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000001111111;
									assign node9727 = (inp[14]) ? node9753 : node9728;
										assign node9728 = (inp[1]) ? node9738 : node9729;
											assign node9729 = (inp[13]) ? node9735 : node9730;
												assign node9730 = (inp[12]) ? 16'b0000000011111111 : node9731;
													assign node9731 = (inp[9]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node9735 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node9738 = (inp[10]) ? node9744 : node9739;
												assign node9739 = (inp[5]) ? node9741 : 16'b0000000001111111;
													assign node9741 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node9744 = (inp[9]) ? 16'b0000000001111111 : node9745;
													assign node9745 = (inp[4]) ? 16'b0000000001111111 : node9746;
														assign node9746 = (inp[13]) ? 16'b0000000001111111 : node9747;
															assign node9747 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node9753 = (inp[10]) ? node9765 : node9754;
											assign node9754 = (inp[9]) ? node9760 : node9755;
												assign node9755 = (inp[13]) ? node9757 : 16'b0000000011111111;
													assign node9757 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9760 = (inp[12]) ? 16'b0000000000111111 : node9761;
													assign node9761 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node9765 = (inp[5]) ? node9769 : node9766;
												assign node9766 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9769 = (inp[9]) ? 16'b0000000000001111 : node9770;
													assign node9770 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node9774 = (inp[0]) ? node9820 : node9775;
									assign node9775 = (inp[4]) ? node9797 : node9776;
										assign node9776 = (inp[14]) ? node9786 : node9777;
											assign node9777 = (inp[10]) ? 16'b0000000001111111 : node9778;
												assign node9778 = (inp[12]) ? node9782 : node9779;
													assign node9779 = (inp[13]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node9782 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node9786 = (inp[9]) ? node9790 : node9787;
												assign node9787 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node9790 = (inp[5]) ? node9792 : 16'b0000000001111111;
													assign node9792 = (inp[10]) ? 16'b0000000000011111 : node9793;
														assign node9793 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node9797 = (inp[13]) ? node9809 : node9798;
											assign node9798 = (inp[14]) ? node9806 : node9799;
												assign node9799 = (inp[5]) ? node9801 : 16'b0000000111111111;
													assign node9801 = (inp[12]) ? 16'b0000000001111111 : node9802;
														assign node9802 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9806 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9809 = (inp[12]) ? node9815 : node9810;
												assign node9810 = (inp[10]) ? 16'b0000000000111111 : node9811;
													assign node9811 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9815 = (inp[5]) ? node9817 : 16'b0000000000111111;
													assign node9817 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node9820 = (inp[5]) ? node9838 : node9821;
										assign node9821 = (inp[1]) ? node9827 : node9822;
											assign node9822 = (inp[9]) ? 16'b0000000001111111 : node9823;
												assign node9823 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9827 = (inp[13]) ? node9833 : node9828;
												assign node9828 = (inp[10]) ? node9830 : 16'b0000000011111111;
													assign node9830 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9833 = (inp[9]) ? node9835 : 16'b0000000000111111;
													assign node9835 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000111111;
										assign node9838 = (inp[1]) ? node9852 : node9839;
											assign node9839 = (inp[14]) ? node9841 : 16'b0000000000111111;
												assign node9841 = (inp[10]) ? node9849 : node9842;
													assign node9842 = (inp[4]) ? node9846 : node9843;
														assign node9843 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node9846 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node9849 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000001111;
											assign node9852 = (inp[13]) ? node9858 : node9853;
												assign node9853 = (inp[14]) ? 16'b0000000000000111 : node9854;
													assign node9854 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node9858 = (inp[4]) ? node9860 : 16'b0000000000001111;
													assign node9860 = (inp[10]) ? node9862 : 16'b0000000000000111;
														assign node9862 = (inp[9]) ? node9864 : 16'b0000000000001111;
															assign node9864 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node9867 = (inp[14]) ? node9937 : node9868;
								assign node9868 = (inp[10]) ? node9900 : node9869;
									assign node9869 = (inp[4]) ? node9883 : node9870;
										assign node9870 = (inp[12]) ? node9878 : node9871;
											assign node9871 = (inp[9]) ? node9875 : node9872;
												assign node9872 = (inp[0]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node9875 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node9878 = (inp[9]) ? node9880 : 16'b0000000011111111;
												assign node9880 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node9883 = (inp[1]) ? node9891 : node9884;
											assign node9884 = (inp[13]) ? 16'b0000000001111111 : node9885;
												assign node9885 = (inp[9]) ? 16'b0000000001111111 : node9886;
													assign node9886 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9891 = (inp[9]) ? node9897 : node9892;
												assign node9892 = (inp[5]) ? node9894 : 16'b0000000001111111;
													assign node9894 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node9897 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000111111;
									assign node9900 = (inp[13]) ? node9924 : node9901;
										assign node9901 = (inp[0]) ? node9913 : node9902;
											assign node9902 = (inp[12]) ? node9906 : node9903;
												assign node9903 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9906 = (inp[7]) ? node9908 : 16'b0000000001111111;
													assign node9908 = (inp[9]) ? 16'b0000000000011111 : node9909;
														assign node9909 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9913 = (inp[5]) ? 16'b0000000000011111 : node9914;
												assign node9914 = (inp[7]) ? node9918 : node9915;
													assign node9915 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9918 = (inp[1]) ? node9920 : 16'b0000000001111111;
														assign node9920 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node9924 = (inp[9]) ? node9930 : node9925;
											assign node9925 = (inp[4]) ? node9927 : 16'b0000000000111111;
												assign node9927 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node9930 = (inp[7]) ? node9934 : node9931;
												assign node9931 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node9934 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000011111;
								assign node9937 = (inp[4]) ? node9993 : node9938;
									assign node9938 = (inp[13]) ? node9964 : node9939;
										assign node9939 = (inp[1]) ? node9945 : node9940;
											assign node9940 = (inp[9]) ? node9942 : 16'b0000000001111111;
												assign node9942 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000111111111;
											assign node9945 = (inp[5]) ? node9953 : node9946;
												assign node9946 = (inp[7]) ? node9950 : node9947;
													assign node9947 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node9950 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node9953 = (inp[7]) ? node9959 : node9954;
													assign node9954 = (inp[12]) ? 16'b0000000000011111 : node9955;
														assign node9955 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node9959 = (inp[0]) ? node9961 : 16'b0000000000011111;
														assign node9961 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node9964 = (inp[12]) ? node9980 : node9965;
											assign node9965 = (inp[10]) ? node9969 : node9966;
												assign node9966 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9969 = (inp[0]) ? node9975 : node9970;
													assign node9970 = (inp[7]) ? 16'b0000000000011111 : node9971;
														assign node9971 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node9975 = (inp[7]) ? node9977 : 16'b0000000000011111;
														assign node9977 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node9980 = (inp[9]) ? node9986 : node9981;
												assign node9981 = (inp[1]) ? 16'b0000000000011111 : node9982;
													assign node9982 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node9986 = (inp[10]) ? node9990 : node9987;
													assign node9987 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node9990 = (inp[7]) ? 16'b0000000000000011 : 16'b0000000000000111;
									assign node9993 = (inp[7]) ? node10013 : node9994;
										assign node9994 = (inp[1]) ? node10000 : node9995;
											assign node9995 = (inp[9]) ? 16'b0000000000111111 : node9996;
												assign node9996 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node10000 = (inp[5]) ? node10008 : node10001;
												assign node10001 = (inp[10]) ? 16'b0000000000011111 : node10002;
													assign node10002 = (inp[0]) ? node10004 : 16'b0000000000111111;
														assign node10004 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10008 = (inp[9]) ? 16'b0000000000001111 : node10009;
													assign node10009 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000001111;
										assign node10013 = (inp[12]) ? node10021 : node10014;
											assign node10014 = (inp[5]) ? 16'b0000000000111111 : node10015;
												assign node10015 = (inp[0]) ? node10017 : 16'b0000000000011111;
													assign node10017 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node10021 = (inp[13]) ? node10031 : node10022;
												assign node10022 = (inp[1]) ? node10026 : node10023;
													assign node10023 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node10026 = (inp[9]) ? node10028 : 16'b0000000000001111;
														assign node10028 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node10031 = (inp[5]) ? node10035 : node10032;
													assign node10032 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node10035 = (inp[0]) ? node10037 : 16'b0000000000000111;
														assign node10037 = (inp[10]) ? 16'b0000000000000011 : 16'b0000000000000111;
				assign node10040 = (inp[4]) ? node10720 : node10041;
					assign node10041 = (inp[13]) ? node10353 : node10042;
						assign node10042 = (inp[10]) ? node10200 : node10043;
							assign node10043 = (inp[8]) ? node10115 : node10044;
								assign node10044 = (inp[0]) ? node10070 : node10045;
									assign node10045 = (inp[5]) ? node10059 : node10046;
										assign node10046 = (inp[1]) ? node10054 : node10047;
											assign node10047 = (inp[14]) ? node10051 : node10048;
												assign node10048 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node10051 = (inp[15]) ? 16'b0000001111111111 : 16'b0000000111111111;
											assign node10054 = (inp[15]) ? node10056 : 16'b0000001111111111;
												assign node10056 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
										assign node10059 = (inp[11]) ? node10067 : node10060;
											assign node10060 = (inp[9]) ? node10064 : node10061;
												assign node10061 = (inp[7]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node10064 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node10067 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node10070 = (inp[15]) ? node10102 : node10071;
										assign node10071 = (inp[9]) ? node10087 : node10072;
											assign node10072 = (inp[12]) ? node10078 : node10073;
												assign node10073 = (inp[11]) ? 16'b0000000111111111 : node10074;
													assign node10074 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node10078 = (inp[1]) ? node10082 : node10079;
													assign node10079 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10082 = (inp[7]) ? node10084 : 16'b0000000011111111;
														assign node10084 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node10087 = (inp[14]) ? node10093 : node10088;
												assign node10088 = (inp[5]) ? 16'b0000000011111111 : node10089;
													assign node10089 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10093 = (inp[11]) ? 16'b0000000001111111 : node10094;
													assign node10094 = (inp[7]) ? node10098 : node10095;
														assign node10095 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10098 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node10102 = (inp[7]) ? node10106 : node10103;
											assign node10103 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10106 = (inp[12]) ? node10112 : node10107;
												assign node10107 = (inp[5]) ? 16'b0000000001111111 : node10108;
													assign node10108 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10112 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node10115 = (inp[0]) ? node10165 : node10116;
									assign node10116 = (inp[14]) ? node10138 : node10117;
										assign node10117 = (inp[12]) ? node10131 : node10118;
											assign node10118 = (inp[7]) ? 16'b0000000011111111 : node10119;
												assign node10119 = (inp[1]) ? node10123 : node10120;
													assign node10120 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node10123 = (inp[9]) ? node10127 : node10124;
														assign node10124 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10127 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node10131 = (inp[1]) ? 16'b0000000001111111 : node10132;
												assign node10132 = (inp[11]) ? 16'b0000000011111111 : node10133;
													assign node10133 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node10138 = (inp[15]) ? node10148 : node10139;
											assign node10139 = (inp[7]) ? node10143 : node10140;
												assign node10140 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10143 = (inp[9]) ? node10145 : 16'b0000000011111111;
													assign node10145 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10148 = (inp[7]) ? node10158 : node10149;
												assign node10149 = (inp[12]) ? node10153 : node10150;
													assign node10150 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10153 = (inp[11]) ? node10155 : 16'b0000000001111111;
														assign node10155 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10158 = (inp[1]) ? 16'b0000000000011111 : node10159;
													assign node10159 = (inp[12]) ? node10161 : 16'b0000000000111111;
														assign node10161 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node10165 = (inp[1]) ? node10177 : node10166;
										assign node10166 = (inp[7]) ? node10172 : node10167;
											assign node10167 = (inp[9]) ? 16'b0000000011111111 : node10168;
												assign node10168 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node10172 = (inp[9]) ? node10174 : 16'b0000000001111111;
												assign node10174 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node10177 = (inp[14]) ? node10185 : node10178;
											assign node10178 = (inp[5]) ? node10180 : 16'b0000000001111111;
												assign node10180 = (inp[12]) ? node10182 : 16'b0000000001111111;
													assign node10182 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10185 = (inp[12]) ? node10195 : node10186;
												assign node10186 = (inp[5]) ? node10190 : node10187;
													assign node10187 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10190 = (inp[7]) ? node10192 : 16'b0000000000111111;
														assign node10192 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10195 = (inp[11]) ? node10197 : 16'b0000000000111111;
													assign node10197 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node10200 = (inp[12]) ? node10278 : node10201;
								assign node10201 = (inp[0]) ? node10229 : node10202;
									assign node10202 = (inp[8]) ? node10212 : node10203;
										assign node10203 = (inp[15]) ? node10207 : node10204;
											assign node10204 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node10207 = (inp[9]) ? node10209 : 16'b0000000111111111;
												assign node10209 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node10212 = (inp[1]) ? node10222 : node10213;
											assign node10213 = (inp[5]) ? node10219 : node10214;
												assign node10214 = (inp[9]) ? 16'b0000000011111111 : node10215;
													assign node10215 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10219 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node10222 = (inp[15]) ? node10224 : 16'b0000000011111111;
												assign node10224 = (inp[14]) ? 16'b0000000001111111 : node10225;
													assign node10225 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node10229 = (inp[11]) ? node10247 : node10230;
										assign node10230 = (inp[15]) ? node10238 : node10231;
											assign node10231 = (inp[14]) ? 16'b0000000001111111 : node10232;
												assign node10232 = (inp[5]) ? 16'b0000000011111111 : node10233;
													assign node10233 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node10238 = (inp[5]) ? node10244 : node10239;
												assign node10239 = (inp[1]) ? node10241 : 16'b0000000011111111;
													assign node10241 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node10244 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node10247 = (inp[8]) ? node10265 : node10248;
											assign node10248 = (inp[7]) ? node10258 : node10249;
												assign node10249 = (inp[9]) ? 16'b0000000001111111 : node10250;
													assign node10250 = (inp[5]) ? node10254 : node10251;
														assign node10251 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10254 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10258 = (inp[5]) ? node10262 : node10259;
													assign node10259 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10262 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10265 = (inp[7]) ? node10271 : node10266;
												assign node10266 = (inp[9]) ? node10268 : 16'b0000000001111111;
													assign node10268 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10271 = (inp[5]) ? 16'b0000000000111111 : node10272;
													assign node10272 = (inp[14]) ? 16'b0000000000111111 : node10273;
														assign node10273 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node10278 = (inp[9]) ? node10318 : node10279;
									assign node10279 = (inp[0]) ? node10305 : node10280;
										assign node10280 = (inp[1]) ? node10290 : node10281;
											assign node10281 = (inp[11]) ? 16'b0000000011111111 : node10282;
												assign node10282 = (inp[8]) ? 16'b0000000011111111 : node10283;
													assign node10283 = (inp[15]) ? 16'b0000000111111111 : node10284;
														assign node10284 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node10290 = (inp[8]) ? node10298 : node10291;
												assign node10291 = (inp[5]) ? node10295 : node10292;
													assign node10292 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10295 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10298 = (inp[7]) ? 16'b0000000000111111 : node10299;
													assign node10299 = (inp[5]) ? 16'b0000000000111111 : node10300;
														assign node10300 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node10305 = (inp[8]) ? node10311 : node10306;
											assign node10306 = (inp[7]) ? 16'b0000000000111111 : node10307;
												assign node10307 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10311 = (inp[7]) ? node10313 : 16'b0000000000111111;
												assign node10313 = (inp[5]) ? 16'b0000000000011111 : node10314;
													assign node10314 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node10318 = (inp[8]) ? node10338 : node10319;
										assign node10319 = (inp[11]) ? node10327 : node10320;
											assign node10320 = (inp[0]) ? node10324 : node10321;
												assign node10321 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node10324 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10327 = (inp[1]) ? node10333 : node10328;
												assign node10328 = (inp[14]) ? 16'b0000000000111111 : node10329;
													assign node10329 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node10333 = (inp[5]) ? node10335 : 16'b0000000000111111;
													assign node10335 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node10338 = (inp[15]) ? node10346 : node10339;
											assign node10339 = (inp[0]) ? node10341 : 16'b0000000000111111;
												assign node10341 = (inp[1]) ? 16'b0000000000011111 : node10342;
													assign node10342 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000011111;
											assign node10346 = (inp[14]) ? node10350 : node10347;
												assign node10347 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10350 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node10353 = (inp[14]) ? node10541 : node10354;
							assign node10354 = (inp[11]) ? node10450 : node10355;
								assign node10355 = (inp[10]) ? node10397 : node10356;
									assign node10356 = (inp[12]) ? node10380 : node10357;
										assign node10357 = (inp[1]) ? node10373 : node10358;
											assign node10358 = (inp[0]) ? node10368 : node10359;
												assign node10359 = (inp[9]) ? 16'b0000000111111111 : node10360;
													assign node10360 = (inp[7]) ? 16'b0000001111111111 : node10361;
														assign node10361 = (inp[15]) ? node10363 : 16'b0000011111111111;
															assign node10363 = (inp[5]) ? 16'b0000001111111111 : 16'b0000001111111111;
												assign node10368 = (inp[15]) ? node10370 : 16'b0000001111111111;
													assign node10370 = (inp[7]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node10373 = (inp[15]) ? node10377 : node10374;
												assign node10374 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node10377 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node10380 = (inp[5]) ? node10386 : node10381;
											assign node10381 = (inp[15]) ? node10383 : 16'b0000000111111111;
												assign node10383 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10386 = (inp[9]) ? node10394 : node10387;
												assign node10387 = (inp[0]) ? 16'b0000000001111111 : node10388;
													assign node10388 = (inp[1]) ? node10390 : 16'b0000000011111111;
														assign node10390 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10394 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node10397 = (inp[5]) ? node10429 : node10398;
										assign node10398 = (inp[0]) ? node10412 : node10399;
											assign node10399 = (inp[7]) ? node10403 : node10400;
												assign node10400 = (inp[9]) ? 16'b0000001111111111 : 16'b0000000011111111;
												assign node10403 = (inp[1]) ? 16'b0000000001111111 : node10404;
													assign node10404 = (inp[15]) ? node10408 : node10405;
														assign node10405 = (inp[9]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node10408 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10412 = (inp[15]) ? node10422 : node10413;
												assign node10413 = (inp[8]) ? node10415 : 16'b0000000011111111;
													assign node10415 = (inp[7]) ? node10417 : 16'b0000000011111111;
														assign node10417 = (inp[12]) ? node10419 : 16'b0000000001111111;
															assign node10419 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10422 = (inp[1]) ? 16'b0000000000011111 : node10423;
													assign node10423 = (inp[12]) ? 16'b0000000001111111 : node10424;
														assign node10424 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node10429 = (inp[0]) ? node10439 : node10430;
											assign node10430 = (inp[9]) ? node10432 : 16'b0000000111111111;
												assign node10432 = (inp[15]) ? node10434 : 16'b0000000001111111;
													assign node10434 = (inp[1]) ? 16'b0000000000111111 : node10435;
														assign node10435 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10439 = (inp[12]) ? node10447 : node10440;
												assign node10440 = (inp[8]) ? node10444 : node10441;
													assign node10441 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node10444 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10447 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node10450 = (inp[7]) ? node10496 : node10451;
									assign node10451 = (inp[15]) ? node10479 : node10452;
										assign node10452 = (inp[10]) ? node10468 : node10453;
											assign node10453 = (inp[8]) ? node10459 : node10454;
												assign node10454 = (inp[9]) ? node10456 : 16'b0000001111111111;
													assign node10456 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10459 = (inp[1]) ? node10461 : 16'b0000000011111111;
													assign node10461 = (inp[0]) ? 16'b0000000000111111 : node10462;
														assign node10462 = (inp[5]) ? 16'b0000000001111111 : node10463;
															assign node10463 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10468 = (inp[8]) ? node10474 : node10469;
												assign node10469 = (inp[5]) ? node10471 : 16'b0000000011111111;
													assign node10471 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10474 = (inp[1]) ? node10476 : 16'b0000000001111111;
													assign node10476 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node10479 = (inp[9]) ? node10491 : node10480;
											assign node10480 = (inp[12]) ? node10482 : 16'b0000000001111111;
												assign node10482 = (inp[8]) ? node10484 : 16'b0000000001111111;
													assign node10484 = (inp[1]) ? 16'b0000000000111111 : node10485;
														assign node10485 = (inp[0]) ? node10487 : 16'b0000000001111111;
															assign node10487 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10491 = (inp[8]) ? 16'b0000000000011111 : node10492;
												assign node10492 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node10496 = (inp[15]) ? node10514 : node10497;
										assign node10497 = (inp[5]) ? node10505 : node10498;
											assign node10498 = (inp[1]) ? node10502 : node10499;
												assign node10499 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10502 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10505 = (inp[8]) ? 16'b0000000000111111 : node10506;
												assign node10506 = (inp[9]) ? node10510 : node10507;
													assign node10507 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node10510 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node10514 = (inp[9]) ? node10532 : node10515;
											assign node10515 = (inp[10]) ? node10525 : node10516;
												assign node10516 = (inp[8]) ? node10520 : node10517;
													assign node10517 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10520 = (inp[0]) ? node10522 : 16'b0000000000111111;
														assign node10522 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10525 = (inp[5]) ? node10529 : node10526;
													assign node10526 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000000011111;
													assign node10529 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node10532 = (inp[1]) ? node10534 : 16'b0000000000011111;
												assign node10534 = (inp[5]) ? node10538 : node10535;
													assign node10535 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000001111;
													assign node10538 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node10541 = (inp[1]) ? node10613 : node10542;
								assign node10542 = (inp[12]) ? node10572 : node10543;
									assign node10543 = (inp[5]) ? node10559 : node10544;
										assign node10544 = (inp[11]) ? node10550 : node10545;
											assign node10545 = (inp[10]) ? 16'b0000000011111111 : node10546;
												assign node10546 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node10550 = (inp[7]) ? node10552 : 16'b0000000011111111;
												assign node10552 = (inp[8]) ? node10554 : 16'b0000000001111111;
													assign node10554 = (inp[0]) ? node10556 : 16'b0000000000111111;
														assign node10556 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node10559 = (inp[0]) ? node10565 : node10560;
											assign node10560 = (inp[7]) ? 16'b0000000001111111 : node10561;
												assign node10561 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node10565 = (inp[11]) ? node10567 : 16'b0000000000111111;
												assign node10567 = (inp[7]) ? node10569 : 16'b0000000001111111;
													assign node10569 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node10572 = (inp[0]) ? node10600 : node10573;
										assign node10573 = (inp[9]) ? node10587 : node10574;
											assign node10574 = (inp[7]) ? node10580 : node10575;
												assign node10575 = (inp[8]) ? 16'b0000000001111111 : node10576;
													assign node10576 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node10580 = (inp[5]) ? 16'b0000000000111111 : node10581;
													assign node10581 = (inp[15]) ? node10583 : 16'b0000000001111111;
														assign node10583 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10587 = (inp[15]) ? node10591 : node10588;
												assign node10588 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node10591 = (inp[11]) ? 16'b0000000000011111 : node10592;
													assign node10592 = (inp[10]) ? node10596 : node10593;
														assign node10593 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10596 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000111111;
										assign node10600 = (inp[11]) ? node10606 : node10601;
											assign node10601 = (inp[7]) ? node10603 : 16'b0000000000111111;
												assign node10603 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node10606 = (inp[7]) ? node10610 : node10607;
												assign node10607 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10610 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node10613 = (inp[12]) ? node10665 : node10614;
									assign node10614 = (inp[8]) ? node10642 : node10615;
										assign node10615 = (inp[11]) ? node10625 : node10616;
											assign node10616 = (inp[7]) ? 16'b0000000001111111 : node10617;
												assign node10617 = (inp[5]) ? 16'b0000000001111111 : node10618;
													assign node10618 = (inp[9]) ? 16'b0000000011111111 : node10619;
														assign node10619 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10625 = (inp[9]) ? node10629 : node10626;
												assign node10626 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10629 = (inp[5]) ? 16'b0000000000001111 : node10630;
													assign node10630 = (inp[0]) ? node10636 : node10631;
														assign node10631 = (inp[15]) ? 16'b0000000000111111 : node10632;
															assign node10632 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10636 = (inp[10]) ? 16'b0000000000011111 : node10637;
															assign node10637 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node10642 = (inp[10]) ? node10654 : node10643;
											assign node10643 = (inp[15]) ? node10649 : node10644;
												assign node10644 = (inp[11]) ? node10646 : 16'b0000000001111111;
													assign node10646 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node10649 = (inp[5]) ? 16'b0000000000011111 : node10650;
													assign node10650 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000011111;
											assign node10654 = (inp[0]) ? node10658 : node10655;
												assign node10655 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10658 = (inp[9]) ? 16'b0000000000001111 : node10659;
													assign node10659 = (inp[7]) ? node10661 : 16'b0000000000011111;
														assign node10661 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node10665 = (inp[9]) ? node10695 : node10666;
										assign node10666 = (inp[15]) ? node10680 : node10667;
											assign node10667 = (inp[0]) ? node10675 : node10668;
												assign node10668 = (inp[10]) ? 16'b0000000000111111 : node10669;
													assign node10669 = (inp[7]) ? node10671 : 16'b0000000001111111;
														assign node10671 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10675 = (inp[8]) ? node10677 : 16'b0000000000111111;
													assign node10677 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node10680 = (inp[7]) ? node10688 : node10681;
												assign node10681 = (inp[5]) ? 16'b0000000000011111 : node10682;
													assign node10682 = (inp[8]) ? 16'b0000000000011111 : node10683;
														assign node10683 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node10688 = (inp[10]) ? node10690 : 16'b0000000000011111;
													assign node10690 = (inp[11]) ? 16'b0000000000000111 : node10691;
														assign node10691 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node10695 = (inp[7]) ? node10713 : node10696;
											assign node10696 = (inp[10]) ? node10704 : node10697;
												assign node10697 = (inp[8]) ? node10701 : node10698;
													assign node10698 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10701 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node10704 = (inp[8]) ? node10708 : node10705;
													assign node10705 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node10708 = (inp[5]) ? node10710 : 16'b0000000000001111;
														assign node10710 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node10713 = (inp[10]) ? node10717 : node10714;
												assign node10714 = (inp[8]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node10717 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000001111;
					assign node10720 = (inp[9]) ? node11082 : node10721;
						assign node10721 = (inp[10]) ? node10905 : node10722;
							assign node10722 = (inp[14]) ? node10814 : node10723;
								assign node10723 = (inp[0]) ? node10771 : node10724;
									assign node10724 = (inp[15]) ? node10748 : node10725;
										assign node10725 = (inp[11]) ? node10735 : node10726;
											assign node10726 = (inp[8]) ? node10728 : 16'b0000000111111111;
												assign node10728 = (inp[12]) ? 16'b0000000011111111 : node10729;
													assign node10729 = (inp[5]) ? node10731 : 16'b0000001111111111;
														assign node10731 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node10735 = (inp[5]) ? node10741 : node10736;
												assign node10736 = (inp[7]) ? 16'b0000000011111111 : node10737;
													assign node10737 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10741 = (inp[7]) ? node10743 : 16'b0000000111111111;
													assign node10743 = (inp[13]) ? 16'b0000000001111111 : node10744;
														assign node10744 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node10748 = (inp[13]) ? node10764 : node10749;
											assign node10749 = (inp[12]) ? node10755 : node10750;
												assign node10750 = (inp[8]) ? 16'b0000000011111111 : node10751;
													assign node10751 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10755 = (inp[7]) ? 16'b0000000001111111 : node10756;
													assign node10756 = (inp[8]) ? node10758 : 16'b0000000011111111;
														assign node10758 = (inp[11]) ? node10760 : 16'b0000000011111111;
															assign node10760 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10764 = (inp[11]) ? node10768 : node10765;
												assign node10765 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node10768 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node10771 = (inp[15]) ? node10803 : node10772;
										assign node10772 = (inp[12]) ? node10788 : node10773;
											assign node10773 = (inp[1]) ? node10779 : node10774;
												assign node10774 = (inp[7]) ? node10776 : 16'b0000000111111111;
													assign node10776 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000111111111;
												assign node10779 = (inp[11]) ? 16'b0000000001111111 : node10780;
													assign node10780 = (inp[5]) ? node10784 : node10781;
														assign node10781 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10784 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10788 = (inp[11]) ? node10800 : node10789;
												assign node10789 = (inp[1]) ? node10795 : node10790;
													assign node10790 = (inp[5]) ? 16'b0000000001111111 : node10791;
														assign node10791 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10795 = (inp[5]) ? node10797 : 16'b0000000001111111;
														assign node10797 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node10800 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node10803 = (inp[5]) ? node10805 : 16'b0000000000111111;
											assign node10805 = (inp[8]) ? node10807 : 16'b0000000000111111;
												assign node10807 = (inp[12]) ? 16'b0000000000011111 : node10808;
													assign node10808 = (inp[11]) ? node10810 : 16'b0000000000111111;
														assign node10810 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node10814 = (inp[5]) ? node10850 : node10815;
									assign node10815 = (inp[7]) ? node10833 : node10816;
										assign node10816 = (inp[12]) ? node10826 : node10817;
											assign node10817 = (inp[0]) ? node10821 : node10818;
												assign node10818 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10821 = (inp[13]) ? node10823 : 16'b0000000001111111;
													assign node10823 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10826 = (inp[0]) ? node10830 : node10827;
												assign node10827 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10830 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node10833 = (inp[15]) ? node10841 : node10834;
											assign node10834 = (inp[1]) ? node10838 : node10835;
												assign node10835 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node10838 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10841 = (inp[12]) ? node10845 : node10842;
												assign node10842 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10845 = (inp[11]) ? 16'b0000000000111111 : node10846;
													assign node10846 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node10850 = (inp[13]) ? node10882 : node10851;
										assign node10851 = (inp[7]) ? node10865 : node10852;
											assign node10852 = (inp[11]) ? node10860 : node10853;
												assign node10853 = (inp[1]) ? 16'b0000000001111111 : node10854;
													assign node10854 = (inp[15]) ? node10856 : 16'b0000000111111111;
														assign node10856 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10860 = (inp[8]) ? node10862 : 16'b0000000000111111;
													assign node10862 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node10865 = (inp[15]) ? node10871 : node10866;
												assign node10866 = (inp[12]) ? 16'b0000000000111111 : node10867;
													assign node10867 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10871 = (inp[1]) ? node10875 : node10872;
													assign node10872 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000000111111;
													assign node10875 = (inp[12]) ? node10877 : 16'b0000000000001111;
														assign node10877 = (inp[11]) ? 16'b0000000000011111 : node10878;
															assign node10878 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000011111;
										assign node10882 = (inp[0]) ? node10896 : node10883;
											assign node10883 = (inp[15]) ? node10885 : 16'b0000000000111111;
												assign node10885 = (inp[11]) ? node10893 : node10886;
													assign node10886 = (inp[8]) ? node10890 : node10887;
														assign node10887 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10890 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node10893 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node10896 = (inp[1]) ? node10900 : node10897;
												assign node10897 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10900 = (inp[12]) ? node10902 : 16'b0000000000111111;
													assign node10902 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000000111;
							assign node10905 = (inp[1]) ? node10997 : node10906;
								assign node10906 = (inp[0]) ? node10944 : node10907;
									assign node10907 = (inp[11]) ? node10929 : node10908;
										assign node10908 = (inp[14]) ? node10910 : 16'b0000000011111111;
											assign node10910 = (inp[12]) ? node10920 : node10911;
												assign node10911 = (inp[13]) ? node10915 : node10912;
													assign node10912 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10915 = (inp[7]) ? 16'b0000000001111111 : node10916;
														assign node10916 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10920 = (inp[15]) ? node10924 : node10921;
													assign node10921 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10924 = (inp[13]) ? node10926 : 16'b0000000000111111;
														assign node10926 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node10929 = (inp[13]) ? node10939 : node10930;
											assign node10930 = (inp[15]) ? 16'b0000000000111111 : node10931;
												assign node10931 = (inp[12]) ? node10933 : 16'b0000000011111111;
													assign node10933 = (inp[7]) ? node10935 : 16'b0000000001111111;
														assign node10935 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10939 = (inp[5]) ? node10941 : 16'b0000000000111111;
												assign node10941 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node10944 = (inp[12]) ? node10970 : node10945;
										assign node10945 = (inp[7]) ? node10959 : node10946;
											assign node10946 = (inp[14]) ? node10952 : node10947;
												assign node10947 = (inp[8]) ? 16'b0000000001111111 : node10948;
													assign node10948 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node10952 = (inp[8]) ? 16'b0000000000111111 : node10953;
													assign node10953 = (inp[15]) ? 16'b0000000001111111 : node10954;
														assign node10954 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10959 = (inp[15]) ? node10967 : node10960;
												assign node10960 = (inp[8]) ? node10962 : 16'b0000000001111111;
													assign node10962 = (inp[11]) ? 16'b0000000000111111 : node10963;
														assign node10963 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10967 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000001111;
										assign node10970 = (inp[8]) ? node10988 : node10971;
											assign node10971 = (inp[15]) ? node10981 : node10972;
												assign node10972 = (inp[14]) ? 16'b0000000000111111 : node10973;
													assign node10973 = (inp[13]) ? node10977 : node10974;
														assign node10974 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10977 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node10981 = (inp[11]) ? 16'b0000000000011111 : node10982;
													assign node10982 = (inp[5]) ? node10984 : 16'b0000000000111111;
														assign node10984 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node10988 = (inp[7]) ? 16'b0000000000011111 : node10989;
												assign node10989 = (inp[5]) ? node10991 : 16'b0000000000111111;
													assign node10991 = (inp[15]) ? 16'b0000000000011111 : node10992;
														assign node10992 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node10997 = (inp[15]) ? node11049 : node10998;
									assign node10998 = (inp[11]) ? node11014 : node10999;
										assign node10999 = (inp[5]) ? node11007 : node11000;
											assign node11000 = (inp[7]) ? node11004 : node11001;
												assign node11001 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node11004 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node11007 = (inp[8]) ? node11009 : 16'b0000000000111111;
												assign node11009 = (inp[7]) ? node11011 : 16'b0000000000111111;
													assign node11011 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node11014 = (inp[12]) ? node11034 : node11015;
											assign node11015 = (inp[13]) ? node11023 : node11016;
												assign node11016 = (inp[14]) ? node11018 : 16'b0000000001111111;
													assign node11018 = (inp[7]) ? 16'b0000000000111111 : node11019;
														assign node11019 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11023 = (inp[14]) ? node11031 : node11024;
													assign node11024 = (inp[0]) ? node11028 : node11025;
														assign node11025 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11028 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000011111;
													assign node11031 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node11034 = (inp[7]) ? node11044 : node11035;
												assign node11035 = (inp[13]) ? node11041 : node11036;
													assign node11036 = (inp[14]) ? 16'b0000000000011111 : node11037;
														assign node11037 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11041 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11044 = (inp[13]) ? node11046 : 16'b0000000000001111;
													assign node11046 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node11049 = (inp[13]) ? node11067 : node11050;
										assign node11050 = (inp[5]) ? node11058 : node11051;
											assign node11051 = (inp[12]) ? node11055 : node11052;
												assign node11052 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11055 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node11058 = (inp[12]) ? node11064 : node11059;
												assign node11059 = (inp[8]) ? 16'b0000000000011111 : node11060;
													assign node11060 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node11064 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node11067 = (inp[14]) ? node11073 : node11068;
											assign node11068 = (inp[0]) ? 16'b0000000000001111 : node11069;
												assign node11069 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node11073 = (inp[0]) ? node11077 : node11074;
												assign node11074 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node11077 = (inp[7]) ? node11079 : 16'b0000000000001111;
													assign node11079 = (inp[12]) ? 16'b0000000000000011 : 16'b0000000000001111;
						assign node11082 = (inp[12]) ? node11266 : node11083;
							assign node11083 = (inp[5]) ? node11181 : node11084;
								assign node11084 = (inp[8]) ? node11124 : node11085;
									assign node11085 = (inp[0]) ? node11101 : node11086;
										assign node11086 = (inp[11]) ? node11098 : node11087;
											assign node11087 = (inp[7]) ? node11091 : node11088;
												assign node11088 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node11091 = (inp[10]) ? 16'b0000000011111111 : node11092;
													assign node11092 = (inp[1]) ? node11094 : 16'b0000000111111111;
														assign node11094 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node11098 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node11101 = (inp[13]) ? node11107 : node11102;
											assign node11102 = (inp[1]) ? node11104 : 16'b0000000011111111;
												assign node11104 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node11107 = (inp[10]) ? node11113 : node11108;
												assign node11108 = (inp[15]) ? node11110 : 16'b0000000001111111;
													assign node11110 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11113 = (inp[1]) ? node11119 : node11114;
													assign node11114 = (inp[14]) ? node11116 : 16'b0000000000111111;
														assign node11116 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11119 = (inp[15]) ? 16'b0000000000001111 : node11120;
														assign node11120 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node11124 = (inp[13]) ? node11160 : node11125;
										assign node11125 = (inp[11]) ? node11145 : node11126;
											assign node11126 = (inp[7]) ? node11138 : node11127;
												assign node11127 = (inp[14]) ? node11133 : node11128;
													assign node11128 = (inp[0]) ? 16'b0000000011111111 : node11129;
														assign node11129 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11133 = (inp[15]) ? 16'b0000000000111111 : node11134;
														assign node11134 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11138 = (inp[0]) ? 16'b0000000000111111 : node11139;
													assign node11139 = (inp[1]) ? node11141 : 16'b0000000001111111;
														assign node11141 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node11145 = (inp[1]) ? node11157 : node11146;
												assign node11146 = (inp[10]) ? node11152 : node11147;
													assign node11147 = (inp[14]) ? 16'b0000000001111111 : node11148;
														assign node11148 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11152 = (inp[7]) ? 16'b0000000000111111 : node11153;
														assign node11153 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11157 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node11160 = (inp[15]) ? node11170 : node11161;
											assign node11161 = (inp[7]) ? node11167 : node11162;
												assign node11162 = (inp[14]) ? 16'b0000000000111111 : node11163;
													assign node11163 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11167 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node11170 = (inp[1]) ? node11176 : node11171;
												assign node11171 = (inp[11]) ? node11173 : 16'b0000000000111111;
													assign node11173 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11176 = (inp[7]) ? node11178 : 16'b0000000000011111;
													assign node11178 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node11181 = (inp[14]) ? node11223 : node11182;
									assign node11182 = (inp[10]) ? node11198 : node11183;
										assign node11183 = (inp[1]) ? node11191 : node11184;
											assign node11184 = (inp[11]) ? node11188 : node11185;
												assign node11185 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node11188 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node11191 = (inp[11]) ? 16'b0000000000111111 : node11192;
												assign node11192 = (inp[15]) ? node11194 : 16'b0000000001111111;
													assign node11194 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node11198 = (inp[8]) ? node11210 : node11199;
											assign node11199 = (inp[15]) ? node11207 : node11200;
												assign node11200 = (inp[13]) ? node11202 : 16'b0000000001111111;
													assign node11202 = (inp[1]) ? 16'b0000000001111111 : node11203;
														assign node11203 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11207 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node11210 = (inp[13]) ? node11214 : node11211;
												assign node11211 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11214 = (inp[11]) ? 16'b0000000000001111 : node11215;
													assign node11215 = (inp[1]) ? node11217 : 16'b0000000000011111;
														assign node11217 = (inp[15]) ? node11219 : 16'b0000000000011111;
															assign node11219 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node11223 = (inp[10]) ? node11243 : node11224;
										assign node11224 = (inp[15]) ? node11230 : node11225;
											assign node11225 = (inp[7]) ? node11227 : 16'b0000000001111111;
												assign node11227 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node11230 = (inp[13]) ? node11236 : node11231;
												assign node11231 = (inp[8]) ? node11233 : 16'b0000000000111111;
													assign node11233 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node11236 = (inp[1]) ? node11238 : 16'b0000000000011111;
													assign node11238 = (inp[0]) ? 16'b0000000000001111 : node11239;
														assign node11239 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node11243 = (inp[7]) ? node11251 : node11244;
											assign node11244 = (inp[15]) ? node11246 : 16'b0000000000011111;
												assign node11246 = (inp[13]) ? 16'b0000000000001111 : node11247;
													assign node11247 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node11251 = (inp[1]) ? node11261 : node11252;
												assign node11252 = (inp[15]) ? node11254 : 16'b0000000000011111;
													assign node11254 = (inp[0]) ? 16'b0000000000001111 : node11255;
														assign node11255 = (inp[8]) ? 16'b0000000000001111 : node11256;
															assign node11256 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node11261 = (inp[0]) ? node11263 : 16'b0000000000000111;
													assign node11263 = (inp[13]) ? 16'b0000000000000011 : 16'b0000000000001111;
							assign node11266 = (inp[8]) ? node11360 : node11267;
								assign node11267 = (inp[0]) ? node11309 : node11268;
									assign node11268 = (inp[11]) ? node11294 : node11269;
										assign node11269 = (inp[7]) ? node11283 : node11270;
											assign node11270 = (inp[1]) ? node11276 : node11271;
												assign node11271 = (inp[15]) ? node11273 : 16'b0000000111111111;
													assign node11273 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11276 = (inp[5]) ? 16'b0000000001111111 : node11277;
													assign node11277 = (inp[10]) ? 16'b0000000001111111 : node11278;
														assign node11278 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node11283 = (inp[14]) ? node11287 : node11284;
												assign node11284 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node11287 = (inp[13]) ? 16'b0000000000011111 : node11288;
													assign node11288 = (inp[1]) ? node11290 : 16'b0000000000111111;
														assign node11290 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node11294 = (inp[1]) ? node11302 : node11295;
											assign node11295 = (inp[14]) ? 16'b0000000000111111 : node11296;
												assign node11296 = (inp[5]) ? 16'b0000000000111111 : node11297;
													assign node11297 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node11302 = (inp[10]) ? 16'b0000000000000111 : node11303;
												assign node11303 = (inp[14]) ? 16'b0000000000011111 : node11304;
													assign node11304 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node11309 = (inp[13]) ? node11333 : node11310;
										assign node11310 = (inp[1]) ? node11324 : node11311;
											assign node11311 = (inp[5]) ? node11317 : node11312;
												assign node11312 = (inp[7]) ? node11314 : 16'b0000000001111111;
													assign node11314 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11317 = (inp[14]) ? 16'b0000000000000111 : node11318;
													assign node11318 = (inp[10]) ? 16'b0000000000011111 : node11319;
														assign node11319 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node11324 = (inp[15]) ? 16'b0000000000011111 : node11325;
												assign node11325 = (inp[5]) ? 16'b0000000000011111 : node11326;
													assign node11326 = (inp[7]) ? node11328 : 16'b0000000000111111;
														assign node11328 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000001111111;
										assign node11333 = (inp[1]) ? node11351 : node11334;
											assign node11334 = (inp[15]) ? node11340 : node11335;
												assign node11335 = (inp[11]) ? node11337 : 16'b0000000000011111;
													assign node11337 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11340 = (inp[7]) ? node11348 : node11341;
													assign node11341 = (inp[14]) ? node11343 : 16'b0000000000001111;
														assign node11343 = (inp[11]) ? 16'b0000000000011111 : node11344;
															assign node11344 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000011111;
													assign node11348 = (inp[10]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node11351 = (inp[10]) ? node11355 : node11352;
												assign node11352 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node11355 = (inp[7]) ? node11357 : 16'b0000000000001111;
													assign node11357 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000000111;
								assign node11360 = (inp[7]) ? node11414 : node11361;
									assign node11361 = (inp[14]) ? node11383 : node11362;
										assign node11362 = (inp[1]) ? node11370 : node11363;
											assign node11363 = (inp[13]) ? node11365 : 16'b0000000000111111;
												assign node11365 = (inp[5]) ? 16'b0000000000011111 : node11366;
													assign node11366 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node11370 = (inp[10]) ? node11376 : node11371;
												assign node11371 = (inp[11]) ? node11373 : 16'b0000000000111111;
													assign node11373 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11376 = (inp[15]) ? node11378 : 16'b0000000000011111;
													assign node11378 = (inp[13]) ? 16'b0000000000001111 : node11379;
														assign node11379 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node11383 = (inp[11]) ? node11399 : node11384;
											assign node11384 = (inp[13]) ? node11390 : node11385;
												assign node11385 = (inp[15]) ? node11387 : 16'b0000000000111111;
													assign node11387 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11390 = (inp[10]) ? 16'b0000000000001111 : node11391;
													assign node11391 = (inp[0]) ? node11395 : node11392;
														assign node11392 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11395 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node11399 = (inp[15]) ? node11405 : node11400;
												assign node11400 = (inp[0]) ? 16'b0000000000000111 : node11401;
													assign node11401 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11405 = (inp[1]) ? node11411 : node11406;
													assign node11406 = (inp[10]) ? node11408 : 16'b0000000000001111;
														assign node11408 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node11411 = (inp[0]) ? 16'b0000000000000011 : 16'b0000000000000111;
									assign node11414 = (inp[10]) ? node11450 : node11415;
										assign node11415 = (inp[5]) ? node11435 : node11416;
											assign node11416 = (inp[14]) ? node11428 : node11417;
												assign node11417 = (inp[1]) ? node11421 : node11418;
													assign node11418 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11421 = (inp[0]) ? node11425 : node11422;
														assign node11422 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node11425 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000001111;
												assign node11428 = (inp[11]) ? node11430 : 16'b0000000000011111;
													assign node11430 = (inp[1]) ? 16'b0000000000001111 : node11431;
														assign node11431 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node11435 = (inp[15]) ? node11447 : node11436;
												assign node11436 = (inp[14]) ? node11444 : node11437;
													assign node11437 = (inp[13]) ? node11441 : node11438;
														assign node11438 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node11441 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node11444 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node11447 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node11450 = (inp[13]) ? node11462 : node11451;
											assign node11451 = (inp[11]) ? node11457 : node11452;
												assign node11452 = (inp[15]) ? node11454 : 16'b0000000000111111;
													assign node11454 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000001111;
												assign node11457 = (inp[15]) ? 16'b0000000000001111 : node11458;
													assign node11458 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000001111;
											assign node11462 = (inp[14]) ? node11470 : node11463;
												assign node11463 = (inp[11]) ? 16'b0000000000000111 : node11464;
													assign node11464 = (inp[15]) ? node11466 : 16'b0000000000001111;
														assign node11466 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node11470 = (inp[11]) ? node11474 : node11471;
													assign node11471 = (inp[1]) ? 16'b0000000000000011 : 16'b0000000000000111;
													assign node11474 = (inp[1]) ? 16'b0000000000000000 : node11475;
														assign node11475 = (inp[0]) ? 16'b0000000000000001 : 16'b0000000000000011;

endmodule