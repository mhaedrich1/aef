module dtc_split05_bm25 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node5;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node11;
	wire [14-1:0] node12;
	wire [14-1:0] node13;
	wire [14-1:0] node17;
	wire [14-1:0] node20;
	wire [14-1:0] node21;
	wire [14-1:0] node24;
	wire [14-1:0] node27;
	wire [14-1:0] node28;
	wire [14-1:0] node29;
	wire [14-1:0] node30;
	wire [14-1:0] node35;
	wire [14-1:0] node36;
	wire [14-1:0] node39;
	wire [14-1:0] node40;
	wire [14-1:0] node44;
	wire [14-1:0] node45;
	wire [14-1:0] node46;
	wire [14-1:0] node47;
	wire [14-1:0] node48;
	wire [14-1:0] node52;
	wire [14-1:0] node54;
	wire [14-1:0] node57;
	wire [14-1:0] node60;
	wire [14-1:0] node61;
	wire [14-1:0] node62;
	wire [14-1:0] node63;
	wire [14-1:0] node67;
	wire [14-1:0] node68;
	wire [14-1:0] node69;
	wire [14-1:0] node74;
	wire [14-1:0] node76;
	wire [14-1:0] node79;
	wire [14-1:0] node80;
	wire [14-1:0] node81;
	wire [14-1:0] node82;
	wire [14-1:0] node84;
	wire [14-1:0] node85;
	wire [14-1:0] node87;
	wire [14-1:0] node88;
	wire [14-1:0] node93;
	wire [14-1:0] node94;
	wire [14-1:0] node96;
	wire [14-1:0] node100;
	wire [14-1:0] node101;
	wire [14-1:0] node102;
	wire [14-1:0] node103;
	wire [14-1:0] node107;
	wire [14-1:0] node110;
	wire [14-1:0] node111;
	wire [14-1:0] node112;
	wire [14-1:0] node116;
	wire [14-1:0] node119;
	wire [14-1:0] node120;
	wire [14-1:0] node121;
	wire [14-1:0] node122;
	wire [14-1:0] node125;
	wire [14-1:0] node126;
	wire [14-1:0] node129;
	wire [14-1:0] node132;
	wire [14-1:0] node135;
	wire [14-1:0] node137;
	wire [14-1:0] node138;
	wire [14-1:0] node140;
	wire [14-1:0] node141;
	wire [14-1:0] node142;
	wire [14-1:0] node147;
	wire [14-1:0] node148;
	wire [14-1:0] node152;
	wire [14-1:0] node153;
	wire [14-1:0] node154;
	wire [14-1:0] node155;
	wire [14-1:0] node156;
	wire [14-1:0] node159;
	wire [14-1:0] node160;
	wire [14-1:0] node161;
	wire [14-1:0] node165;
	wire [14-1:0] node168;
	wire [14-1:0] node169;
	wire [14-1:0] node170;
	wire [14-1:0] node171;
	wire [14-1:0] node174;
	wire [14-1:0] node177;
	wire [14-1:0] node178;
	wire [14-1:0] node180;
	wire [14-1:0] node183;
	wire [14-1:0] node184;
	wire [14-1:0] node188;
	wire [14-1:0] node191;
	wire [14-1:0] node192;
	wire [14-1:0] node193;
	wire [14-1:0] node194;
	wire [14-1:0] node195;
	wire [14-1:0] node198;
	wire [14-1:0] node201;
	wire [14-1:0] node203;
	wire [14-1:0] node206;
	wire [14-1:0] node209;
	wire [14-1:0] node210;
	wire [14-1:0] node211;
	wire [14-1:0] node215;
	wire [14-1:0] node216;
	wire [14-1:0] node219;
	wire [14-1:0] node221;
	wire [14-1:0] node224;
	wire [14-1:0] node225;
	wire [14-1:0] node226;
	wire [14-1:0] node227;
	wire [14-1:0] node228;
	wire [14-1:0] node230;
	wire [14-1:0] node233;
	wire [14-1:0] node235;
	wire [14-1:0] node238;
	wire [14-1:0] node240;
	wire [14-1:0] node243;
	wire [14-1:0] node244;
	wire [14-1:0] node245;
	wire [14-1:0] node247;
	wire [14-1:0] node251;
	wire [14-1:0] node252;
	wire [14-1:0] node254;
	wire [14-1:0] node256;
	wire [14-1:0] node260;
	wire [14-1:0] node261;
	wire [14-1:0] node262;
	wire [14-1:0] node263;
	wire [14-1:0] node264;
	wire [14-1:0] node267;
	wire [14-1:0] node269;
	wire [14-1:0] node272;
	wire [14-1:0] node273;
	wire [14-1:0] node274;
	wire [14-1:0] node279;
	wire [14-1:0] node281;
	wire [14-1:0] node282;
	wire [14-1:0] node286;
	wire [14-1:0] node287;
	wire [14-1:0] node289;
	wire [14-1:0] node291;
	wire [14-1:0] node294;
	wire [14-1:0] node295;
	wire [14-1:0] node298;
	wire [14-1:0] node299;
	wire [14-1:0] node300;
	wire [14-1:0] node302;
	wire [14-1:0] node307;
	wire [14-1:0] node308;
	wire [14-1:0] node309;
	wire [14-1:0] node310;
	wire [14-1:0] node311;
	wire [14-1:0] node312;
	wire [14-1:0] node313;
	wire [14-1:0] node317;
	wire [14-1:0] node318;
	wire [14-1:0] node319;
	wire [14-1:0] node323;
	wire [14-1:0] node326;
	wire [14-1:0] node327;
	wire [14-1:0] node328;
	wire [14-1:0] node329;
	wire [14-1:0] node333;
	wire [14-1:0] node334;
	wire [14-1:0] node338;
	wire [14-1:0] node339;
	wire [14-1:0] node340;
	wire [14-1:0] node343;
	wire [14-1:0] node345;
	wire [14-1:0] node348;
	wire [14-1:0] node351;
	wire [14-1:0] node352;
	wire [14-1:0] node353;
	wire [14-1:0] node355;
	wire [14-1:0] node358;
	wire [14-1:0] node359;
	wire [14-1:0] node361;
	wire [14-1:0] node364;
	wire [14-1:0] node367;
	wire [14-1:0] node368;
	wire [14-1:0] node370;
	wire [14-1:0] node372;
	wire [14-1:0] node375;
	wire [14-1:0] node376;
	wire [14-1:0] node379;
	wire [14-1:0] node382;
	wire [14-1:0] node383;
	wire [14-1:0] node384;
	wire [14-1:0] node385;
	wire [14-1:0] node386;
	wire [14-1:0] node390;
	wire [14-1:0] node391;
	wire [14-1:0] node392;
	wire [14-1:0] node396;
	wire [14-1:0] node398;
	wire [14-1:0] node401;
	wire [14-1:0] node402;
	wire [14-1:0] node403;
	wire [14-1:0] node404;
	wire [14-1:0] node408;
	wire [14-1:0] node411;
	wire [14-1:0] node412;
	wire [14-1:0] node413;
	wire [14-1:0] node417;
	wire [14-1:0] node420;
	wire [14-1:0] node421;
	wire [14-1:0] node422;
	wire [14-1:0] node423;
	wire [14-1:0] node424;
	wire [14-1:0] node428;
	wire [14-1:0] node429;
	wire [14-1:0] node433;
	wire [14-1:0] node436;
	wire [14-1:0] node437;
	wire [14-1:0] node438;
	wire [14-1:0] node442;
	wire [14-1:0] node444;
	wire [14-1:0] node447;
	wire [14-1:0] node448;
	wire [14-1:0] node449;
	wire [14-1:0] node450;
	wire [14-1:0] node451;
	wire [14-1:0] node452;
	wire [14-1:0] node455;
	wire [14-1:0] node458;
	wire [14-1:0] node460;
	wire [14-1:0] node461;
	wire [14-1:0] node463;
	wire [14-1:0] node467;
	wire [14-1:0] node468;
	wire [14-1:0] node469;
	wire [14-1:0] node470;
	wire [14-1:0] node473;
	wire [14-1:0] node477;
	wire [14-1:0] node478;
	wire [14-1:0] node480;
	wire [14-1:0] node484;
	wire [14-1:0] node485;
	wire [14-1:0] node486;
	wire [14-1:0] node487;
	wire [14-1:0] node490;
	wire [14-1:0] node493;
	wire [14-1:0] node495;
	wire [14-1:0] node498;
	wire [14-1:0] node499;
	wire [14-1:0] node501;
	wire [14-1:0] node503;
	wire [14-1:0] node504;
	wire [14-1:0] node508;
	wire [14-1:0] node510;
	wire [14-1:0] node513;
	wire [14-1:0] node514;
	wire [14-1:0] node515;
	wire [14-1:0] node516;
	wire [14-1:0] node517;
	wire [14-1:0] node519;
	wire [14-1:0] node523;
	wire [14-1:0] node524;
	wire [14-1:0] node527;
	wire [14-1:0] node528;
	wire [14-1:0] node532;
	wire [14-1:0] node533;
	wire [14-1:0] node534;
	wire [14-1:0] node536;
	wire [14-1:0] node540;
	wire [14-1:0] node541;
	wire [14-1:0] node545;
	wire [14-1:0] node546;
	wire [14-1:0] node547;
	wire [14-1:0] node549;
	wire [14-1:0] node550;
	wire [14-1:0] node554;
	wire [14-1:0] node555;
	wire [14-1:0] node556;
	wire [14-1:0] node559;
	wire [14-1:0] node560;
	wire [14-1:0] node562;
	wire [14-1:0] node567;
	wire [14-1:0] node568;
	wire [14-1:0] node569;
	wire [14-1:0] node573;
	wire [14-1:0] node574;
	wire [14-1:0] node577;
	wire [14-1:0] node578;
	wire [14-1:0] node582;
	wire [14-1:0] node583;
	wire [14-1:0] node584;
	wire [14-1:0] node585;
	wire [14-1:0] node586;
	wire [14-1:0] node587;
	wire [14-1:0] node588;
	wire [14-1:0] node589;
	wire [14-1:0] node592;
	wire [14-1:0] node593;
	wire [14-1:0] node595;
	wire [14-1:0] node599;
	wire [14-1:0] node600;
	wire [14-1:0] node603;
	wire [14-1:0] node605;
	wire [14-1:0] node608;
	wire [14-1:0] node609;
	wire [14-1:0] node611;
	wire [14-1:0] node614;
	wire [14-1:0] node615;
	wire [14-1:0] node616;
	wire [14-1:0] node617;
	wire [14-1:0] node619;
	wire [14-1:0] node623;
	wire [14-1:0] node627;
	wire [14-1:0] node628;
	wire [14-1:0] node629;
	wire [14-1:0] node631;
	wire [14-1:0] node634;
	wire [14-1:0] node635;
	wire [14-1:0] node638;
	wire [14-1:0] node641;
	wire [14-1:0] node642;
	wire [14-1:0] node643;
	wire [14-1:0] node646;
	wire [14-1:0] node649;
	wire [14-1:0] node651;
	wire [14-1:0] node652;
	wire [14-1:0] node655;
	wire [14-1:0] node657;
	wire [14-1:0] node660;
	wire [14-1:0] node661;
	wire [14-1:0] node662;
	wire [14-1:0] node663;
	wire [14-1:0] node666;
	wire [14-1:0] node667;
	wire [14-1:0] node669;
	wire [14-1:0] node671;
	wire [14-1:0] node674;
	wire [14-1:0] node677;
	wire [14-1:0] node678;
	wire [14-1:0] node680;
	wire [14-1:0] node681;
	wire [14-1:0] node685;
	wire [14-1:0] node686;
	wire [14-1:0] node687;
	wire [14-1:0] node690;
	wire [14-1:0] node691;
	wire [14-1:0] node696;
	wire [14-1:0] node697;
	wire [14-1:0] node698;
	wire [14-1:0] node699;
	wire [14-1:0] node700;
	wire [14-1:0] node704;
	wire [14-1:0] node707;
	wire [14-1:0] node708;
	wire [14-1:0] node709;
	wire [14-1:0] node711;
	wire [14-1:0] node716;
	wire [14-1:0] node717;
	wire [14-1:0] node719;
	wire [14-1:0] node720;
	wire [14-1:0] node724;
	wire [14-1:0] node726;
	wire [14-1:0] node728;
	wire [14-1:0] node731;
	wire [14-1:0] node732;
	wire [14-1:0] node733;
	wire [14-1:0] node734;
	wire [14-1:0] node735;
	wire [14-1:0] node736;
	wire [14-1:0] node741;
	wire [14-1:0] node742;
	wire [14-1:0] node744;
	wire [14-1:0] node747;
	wire [14-1:0] node748;
	wire [14-1:0] node752;
	wire [14-1:0] node753;
	wire [14-1:0] node754;
	wire [14-1:0] node755;
	wire [14-1:0] node757;
	wire [14-1:0] node760;
	wire [14-1:0] node761;
	wire [14-1:0] node765;
	wire [14-1:0] node766;
	wire [14-1:0] node768;
	wire [14-1:0] node771;
	wire [14-1:0] node774;
	wire [14-1:0] node775;
	wire [14-1:0] node776;
	wire [14-1:0] node777;
	wire [14-1:0] node780;
	wire [14-1:0] node783;
	wire [14-1:0] node784;
	wire [14-1:0] node787;
	wire [14-1:0] node790;
	wire [14-1:0] node791;
	wire [14-1:0] node792;
	wire [14-1:0] node796;
	wire [14-1:0] node798;
	wire [14-1:0] node801;
	wire [14-1:0] node802;
	wire [14-1:0] node803;
	wire [14-1:0] node804;
	wire [14-1:0] node805;
	wire [14-1:0] node809;
	wire [14-1:0] node810;
	wire [14-1:0] node812;
	wire [14-1:0] node813;
	wire [14-1:0] node815;
	wire [14-1:0] node819;
	wire [14-1:0] node820;
	wire [14-1:0] node824;
	wire [14-1:0] node825;
	wire [14-1:0] node826;
	wire [14-1:0] node827;
	wire [14-1:0] node828;
	wire [14-1:0] node833;
	wire [14-1:0] node836;
	wire [14-1:0] node839;
	wire [14-1:0] node840;
	wire [14-1:0] node841;
	wire [14-1:0] node843;
	wire [14-1:0] node846;
	wire [14-1:0] node847;
	wire [14-1:0] node850;
	wire [14-1:0] node851;
	wire [14-1:0] node852;
	wire [14-1:0] node857;
	wire [14-1:0] node858;
	wire [14-1:0] node859;
	wire [14-1:0] node863;
	wire [14-1:0] node864;
	wire [14-1:0] node865;
	wire [14-1:0] node869;
	wire [14-1:0] node871;
	wire [14-1:0] node874;
	wire [14-1:0] node875;
	wire [14-1:0] node876;
	wire [14-1:0] node877;
	wire [14-1:0] node878;
	wire [14-1:0] node879;
	wire [14-1:0] node880;
	wire [14-1:0] node883;
	wire [14-1:0] node886;
	wire [14-1:0] node888;
	wire [14-1:0] node889;
	wire [14-1:0] node893;
	wire [14-1:0] node894;
	wire [14-1:0] node896;
	wire [14-1:0] node899;
	wire [14-1:0] node900;
	wire [14-1:0] node904;
	wire [14-1:0] node905;
	wire [14-1:0] node906;
	wire [14-1:0] node907;
	wire [14-1:0] node910;
	wire [14-1:0] node913;
	wire [14-1:0] node916;
	wire [14-1:0] node917;
	wire [14-1:0] node920;
	wire [14-1:0] node922;
	wire [14-1:0] node924;
	wire [14-1:0] node927;
	wire [14-1:0] node928;
	wire [14-1:0] node929;
	wire [14-1:0] node931;
	wire [14-1:0] node932;
	wire [14-1:0] node933;
	wire [14-1:0] node934;
	wire [14-1:0] node938;
	wire [14-1:0] node941;
	wire [14-1:0] node944;
	wire [14-1:0] node945;
	wire [14-1:0] node946;
	wire [14-1:0] node949;
	wire [14-1:0] node950;
	wire [14-1:0] node953;
	wire [14-1:0] node954;
	wire [14-1:0] node958;
	wire [14-1:0] node960;
	wire [14-1:0] node961;
	wire [14-1:0] node965;
	wire [14-1:0] node966;
	wire [14-1:0] node967;
	wire [14-1:0] node968;
	wire [14-1:0] node969;
	wire [14-1:0] node972;
	wire [14-1:0] node974;
	wire [14-1:0] node977;
	wire [14-1:0] node979;
	wire [14-1:0] node980;
	wire [14-1:0] node984;
	wire [14-1:0] node986;
	wire [14-1:0] node988;
	wire [14-1:0] node990;
	wire [14-1:0] node993;
	wire [14-1:0] node994;
	wire [14-1:0] node995;
	wire [14-1:0] node997;
	wire [14-1:0] node1000;
	wire [14-1:0] node1001;
	wire [14-1:0] node1003;
	wire [14-1:0] node1007;
	wire [14-1:0] node1009;
	wire [14-1:0] node1010;
	wire [14-1:0] node1014;
	wire [14-1:0] node1015;
	wire [14-1:0] node1016;
	wire [14-1:0] node1017;
	wire [14-1:0] node1019;
	wire [14-1:0] node1020;
	wire [14-1:0] node1023;
	wire [14-1:0] node1026;
	wire [14-1:0] node1027;
	wire [14-1:0] node1028;
	wire [14-1:0] node1031;
	wire [14-1:0] node1032;
	wire [14-1:0] node1034;
	wire [14-1:0] node1037;
	wire [14-1:0] node1040;
	wire [14-1:0] node1043;
	wire [14-1:0] node1044;
	wire [14-1:0] node1045;
	wire [14-1:0] node1046;
	wire [14-1:0] node1050;
	wire [14-1:0] node1051;
	wire [14-1:0] node1052;
	wire [14-1:0] node1057;
	wire [14-1:0] node1058;
	wire [14-1:0] node1059;
	wire [14-1:0] node1062;
	wire [14-1:0] node1063;
	wire [14-1:0] node1067;
	wire [14-1:0] node1069;
	wire [14-1:0] node1071;
	wire [14-1:0] node1074;
	wire [14-1:0] node1075;
	wire [14-1:0] node1076;
	wire [14-1:0] node1077;
	wire [14-1:0] node1080;
	wire [14-1:0] node1082;
	wire [14-1:0] node1085;
	wire [14-1:0] node1086;
	wire [14-1:0] node1088;
	wire [14-1:0] node1090;
	wire [14-1:0] node1093;
	wire [14-1:0] node1094;
	wire [14-1:0] node1095;
	wire [14-1:0] node1099;
	wire [14-1:0] node1102;
	wire [14-1:0] node1103;
	wire [14-1:0] node1104;
	wire [14-1:0] node1106;
	wire [14-1:0] node1108;
	wire [14-1:0] node1111;
	wire [14-1:0] node1113;
	wire [14-1:0] node1116;
	wire [14-1:0] node1117;
	wire [14-1:0] node1119;
	wire [14-1:0] node1120;
	wire [14-1:0] node1122;
	wire [14-1:0] node1126;
	wire [14-1:0] node1127;
	wire [14-1:0] node1129;
	wire [14-1:0] node1132;
	wire [14-1:0] node1133;
	wire [14-1:0] node1135;
	wire [14-1:0] node1137;

	assign outp = (inp[4]) ? node582 : node1;
		assign node1 = (inp[1]) ? node307 : node2;
			assign node2 = (inp[0]) ? node152 : node3;
				assign node3 = (inp[7]) ? node79 : node4;
					assign node4 = (inp[3]) ? node44 : node5;
						assign node5 = (inp[13]) ? node27 : node6;
							assign node6 = (inp[12]) ? node20 : node7;
								assign node7 = (inp[5]) ? node11 : node8;
									assign node8 = (inp[2]) ? 14'b00011111111111 : 14'b00111111111111;
									assign node11 = (inp[6]) ? node17 : node12;
										assign node12 = (inp[10]) ? 14'b00011111111111 : node13;
											assign node13 = (inp[11]) ? 14'b00011111111111 : 14'b00111111111111;
										assign node17 = (inp[11]) ? 14'b00001111111111 : 14'b00011111111111;
								assign node20 = (inp[2]) ? node24 : node21;
									assign node21 = (inp[5]) ? 14'b00011111111111 : 14'b00001111111111;
									assign node24 = (inp[8]) ? 14'b00001111111111 : 14'b00000111111111;
							assign node27 = (inp[10]) ? node35 : node28;
								assign node28 = (inp[5]) ? 14'b00000111111111 : node29;
									assign node29 = (inp[6]) ? 14'b00011111111111 : node30;
										assign node30 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
								assign node35 = (inp[11]) ? node39 : node36;
									assign node36 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node39 = (inp[8]) ? 14'b00000011111111 : node40;
										assign node40 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
						assign node44 = (inp[6]) ? node60 : node45;
							assign node45 = (inp[5]) ? node57 : node46;
								assign node46 = (inp[13]) ? node52 : node47;
									assign node47 = (inp[11]) ? 14'b00001111111111 : node48;
										assign node48 = (inp[10]) ? 14'b00111111111111 : 14'b01111111111111;
									assign node52 = (inp[12]) ? node54 : 14'b00001111111111;
										assign node54 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
								assign node57 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
							assign node60 = (inp[2]) ? node74 : node61;
								assign node61 = (inp[9]) ? node67 : node62;
									assign node62 = (inp[8]) ? 14'b00000111111111 : node63;
										assign node63 = (inp[13]) ? 14'b00000011111111 : 14'b00001111111111;
									assign node67 = (inp[11]) ? 14'b00000000111111 : node68;
										assign node68 = (inp[13]) ? 14'b00000001111111 : node69;
											assign node69 = (inp[8]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node74 = (inp[13]) ? node76 : 14'b00000011111111;
									assign node76 = (inp[8]) ? 14'b00000011111111 : 14'b00000001111111;
					assign node79 = (inp[12]) ? node119 : node80;
						assign node80 = (inp[13]) ? node100 : node81;
							assign node81 = (inp[3]) ? node93 : node82;
								assign node82 = (inp[5]) ? node84 : 14'b00001111111111;
									assign node84 = (inp[11]) ? 14'b00000111111111 : node85;
										assign node85 = (inp[10]) ? node87 : 14'b00001111111111;
											assign node87 = (inp[6]) ? 14'b00000111111111 : node88;
												assign node88 = (inp[8]) ? 14'b00000111111111 : 14'b00001111111111;
								assign node93 = (inp[10]) ? 14'b00000011111111 : node94;
									assign node94 = (inp[5]) ? node96 : 14'b00000111111111;
										assign node96 = (inp[8]) ? 14'b00000001111111 : 14'b00000111111111;
							assign node100 = (inp[10]) ? node110 : node101;
								assign node101 = (inp[11]) ? node107 : node102;
									assign node102 = (inp[9]) ? 14'b00000111111111 : node103;
										assign node103 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
									assign node107 = (inp[8]) ? 14'b00000011111111 : 14'b00000001111111;
								assign node110 = (inp[3]) ? node116 : node111;
									assign node111 = (inp[2]) ? 14'b00000011111111 : node112;
										assign node112 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node116 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
						assign node119 = (inp[10]) ? node135 : node120;
							assign node120 = (inp[3]) ? node132 : node121;
								assign node121 = (inp[2]) ? node125 : node122;
									assign node122 = (inp[8]) ? 14'b00001111111111 : 14'b00000111111111;
									assign node125 = (inp[11]) ? node129 : node126;
										assign node126 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node129 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node132 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node135 = (inp[6]) ? node137 : 14'b00000011111111;
								assign node137 = (inp[3]) ? node147 : node138;
									assign node138 = (inp[8]) ? node140 : 14'b00000011111111;
										assign node140 = (inp[13]) ? 14'b00000001111111 : node141;
											assign node141 = (inp[9]) ? 14'b00000001111111 : node142;
												assign node142 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node147 = (inp[8]) ? 14'b00000000111111 : node148;
										assign node148 = (inp[9]) ? 14'b00000001111111 : 14'b00000000111111;
				assign node152 = (inp[12]) ? node224 : node153;
					assign node153 = (inp[5]) ? node191 : node154;
						assign node154 = (inp[11]) ? node168 : node155;
							assign node155 = (inp[2]) ? node159 : node156;
								assign node156 = (inp[7]) ? 14'b00001111111111 : 14'b00011111111111;
								assign node159 = (inp[9]) ? node165 : node160;
									assign node160 = (inp[7]) ? 14'b00000111111111 : node161;
										assign node161 = (inp[8]) ? 14'b00001111111111 : 14'b00011111111111;
									assign node165 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
							assign node168 = (inp[3]) ? node188 : node169;
								assign node169 = (inp[8]) ? node177 : node170;
									assign node170 = (inp[7]) ? node174 : node171;
										assign node171 = (inp[6]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node174 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node177 = (inp[2]) ? node183 : node178;
										assign node178 = (inp[9]) ? node180 : 14'b00000111111111;
											assign node180 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node183 = (inp[13]) ? 14'b00000011111111 : node184;
											assign node184 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node188 = (inp[8]) ? 14'b00000001111111 : 14'b00000011111111;
						assign node191 = (inp[8]) ? node209 : node192;
							assign node192 = (inp[6]) ? node206 : node193;
								assign node193 = (inp[7]) ? node201 : node194;
									assign node194 = (inp[9]) ? node198 : node195;
										assign node195 = (inp[3]) ? 14'b00000111111111 : 14'b00001111111111;
										assign node198 = (inp[13]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node201 = (inp[2]) ? node203 : 14'b00000011111111;
										assign node203 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node206 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node209 = (inp[7]) ? node215 : node210;
								assign node210 = (inp[9]) ? 14'b00000001111111 : node211;
									assign node211 = (inp[6]) ? 14'b00000011111111 : 14'b00001111111111;
								assign node215 = (inp[2]) ? node219 : node216;
									assign node216 = (inp[9]) ? 14'b00000000111111 : 14'b00000011111111;
									assign node219 = (inp[9]) ? node221 : 14'b00000000111111;
										assign node221 = (inp[3]) ? 14'b00000000001111 : 14'b00000000111111;
					assign node224 = (inp[10]) ? node260 : node225;
						assign node225 = (inp[2]) ? node243 : node226;
							assign node226 = (inp[11]) ? node238 : node227;
								assign node227 = (inp[3]) ? node233 : node228;
									assign node228 = (inp[5]) ? node230 : 14'b00011111111111;
										assign node230 = (inp[6]) ? 14'b00001111111111 : 14'b00000111111111;
									assign node233 = (inp[7]) ? node235 : 14'b00000011111111;
										assign node235 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node238 = (inp[9]) ? node240 : 14'b00000011111111;
									assign node240 = (inp[6]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node243 = (inp[6]) ? node251 : node244;
								assign node244 = (inp[11]) ? 14'b00000001111111 : node245;
									assign node245 = (inp[8]) ? node247 : 14'b00000111111111;
										assign node247 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node251 = (inp[7]) ? 14'b00000000001111 : node252;
									assign node252 = (inp[8]) ? node254 : 14'b00000000111111;
										assign node254 = (inp[9]) ? node256 : 14'b00000001111111;
											assign node256 = (inp[3]) ? 14'b00000000011111 : 14'b00000001111111;
						assign node260 = (inp[8]) ? node286 : node261;
							assign node261 = (inp[6]) ? node279 : node262;
								assign node262 = (inp[13]) ? node272 : node263;
									assign node263 = (inp[5]) ? node267 : node264;
										assign node264 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node267 = (inp[9]) ? node269 : 14'b00000011111111;
											assign node269 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node272 = (inp[5]) ? 14'b00000000011111 : node273;
										assign node273 = (inp[3]) ? 14'b00000001111111 : node274;
											assign node274 = (inp[11]) ? 14'b00000011111111 : 14'b00000001111111;
								assign node279 = (inp[5]) ? node281 : 14'b00000000111111;
									assign node281 = (inp[9]) ? 14'b00000000001111 : node282;
										assign node282 = (inp[2]) ? 14'b00000000111111 : 14'b00000000011111;
							assign node286 = (inp[3]) ? node294 : node287;
								assign node287 = (inp[13]) ? node289 : 14'b00000000111111;
									assign node289 = (inp[2]) ? node291 : 14'b00000000111111;
										assign node291 = (inp[7]) ? 14'b00000000000111 : 14'b00000000011111;
								assign node294 = (inp[7]) ? node298 : node295;
									assign node295 = (inp[9]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node298 = (inp[6]) ? 14'b00000000001111 : node299;
										assign node299 = (inp[9]) ? 14'b00000000001111 : node300;
											assign node300 = (inp[13]) ? node302 : 14'b00000000011111;
												assign node302 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
			assign node307 = (inp[3]) ? node447 : node308;
				assign node308 = (inp[6]) ? node382 : node309;
					assign node309 = (inp[8]) ? node351 : node310;
						assign node310 = (inp[13]) ? node326 : node311;
							assign node311 = (inp[11]) ? node317 : node312;
								assign node312 = (inp[7]) ? 14'b00001111111111 : node313;
									assign node313 = (inp[5]) ? 14'b00011111111111 : 14'b00111111111111;
								assign node317 = (inp[2]) ? node323 : node318;
									assign node318 = (inp[5]) ? 14'b00000111111111 : node319;
										assign node319 = (inp[12]) ? 14'b00011111111111 : 14'b00001111111111;
									assign node323 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
							assign node326 = (inp[9]) ? node338 : node327;
								assign node327 = (inp[10]) ? node333 : node328;
									assign node328 = (inp[11]) ? 14'b00000111111111 : node329;
										assign node329 = (inp[12]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node333 = (inp[7]) ? 14'b00000011111111 : node334;
										assign node334 = (inp[0]) ? 14'b00000011111111 : 14'b00001111111111;
								assign node338 = (inp[12]) ? node348 : node339;
									assign node339 = (inp[0]) ? node343 : node340;
										assign node340 = (inp[5]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node343 = (inp[11]) ? node345 : 14'b00000111111111;
											assign node345 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node348 = (inp[7]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node351 = (inp[9]) ? node367 : node352;
							assign node352 = (inp[13]) ? node358 : node353;
								assign node353 = (inp[10]) ? node355 : 14'b00000111111111;
									assign node355 = (inp[0]) ? 14'b00000001111111 : 14'b00000111111111;
								assign node358 = (inp[10]) ? node364 : node359;
									assign node359 = (inp[2]) ? node361 : 14'b00000111111111;
										assign node361 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node364 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node367 = (inp[2]) ? node375 : node368;
								assign node368 = (inp[11]) ? node370 : 14'b00000111111111;
									assign node370 = (inp[10]) ? node372 : 14'b00000001111111;
										assign node372 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node375 = (inp[13]) ? node379 : node376;
									assign node376 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node379 = (inp[12]) ? 14'b00000000001111 : 14'b00000000111111;
					assign node382 = (inp[7]) ? node420 : node383;
						assign node383 = (inp[2]) ? node401 : node384;
							assign node384 = (inp[0]) ? node390 : node385;
								assign node385 = (inp[11]) ? 14'b00001111111111 : node386;
									assign node386 = (inp[10]) ? 14'b00000111111111 : 14'b00000011111111;
								assign node390 = (inp[8]) ? node396 : node391;
									assign node391 = (inp[12]) ? 14'b00000000111111 : node392;
										assign node392 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node396 = (inp[13]) ? node398 : 14'b00000001111111;
										assign node398 = (inp[5]) ? 14'b00000001111111 : 14'b00000000111111;
							assign node401 = (inp[10]) ? node411 : node402;
								assign node402 = (inp[12]) ? node408 : node403;
									assign node403 = (inp[9]) ? 14'b00000001111111 : node404;
										assign node404 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node408 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node411 = (inp[11]) ? node417 : node412;
									assign node412 = (inp[12]) ? 14'b00000001111111 : node413;
										assign node413 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node417 = (inp[0]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node420 = (inp[8]) ? node436 : node421;
							assign node421 = (inp[0]) ? node433 : node422;
								assign node422 = (inp[10]) ? node428 : node423;
									assign node423 = (inp[5]) ? 14'b00000001111111 : node424;
										assign node424 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node428 = (inp[12]) ? 14'b00000001111111 : node429;
										assign node429 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node433 = (inp[2]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node436 = (inp[5]) ? node442 : node437;
								assign node437 = (inp[11]) ? 14'b00000000011111 : node438;
									assign node438 = (inp[9]) ? 14'b00000011111111 : 14'b00000001111111;
								assign node442 = (inp[12]) ? node444 : 14'b00000000111111;
									assign node444 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
				assign node447 = (inp[6]) ? node513 : node448;
					assign node448 = (inp[9]) ? node484 : node449;
						assign node449 = (inp[5]) ? node467 : node450;
							assign node450 = (inp[7]) ? node458 : node451;
								assign node451 = (inp[0]) ? node455 : node452;
									assign node452 = (inp[13]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node455 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node458 = (inp[2]) ? node460 : 14'b00000011111111;
									assign node460 = (inp[13]) ? 14'b00000001111111 : node461;
										assign node461 = (inp[8]) ? node463 : 14'b00000011111111;
											assign node463 = (inp[12]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node467 = (inp[11]) ? node477 : node468;
								assign node468 = (inp[13]) ? 14'b00000000111111 : node469;
									assign node469 = (inp[7]) ? node473 : node470;
										assign node470 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node473 = (inp[12]) ? 14'b00000011111111 : 14'b00000001111111;
								assign node477 = (inp[10]) ? 14'b00000000111111 : node478;
									assign node478 = (inp[0]) ? node480 : 14'b00000011111111;
										assign node480 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node484 = (inp[7]) ? node498 : node485;
							assign node485 = (inp[13]) ? node493 : node486;
								assign node486 = (inp[8]) ? node490 : node487;
									assign node487 = (inp[12]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node490 = (inp[12]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node493 = (inp[2]) ? node495 : 14'b00000001111111;
									assign node495 = (inp[10]) ? 14'b00000001111111 : 14'b00000000111111;
							assign node498 = (inp[5]) ? node508 : node499;
								assign node499 = (inp[0]) ? node501 : 14'b00000000111111;
									assign node501 = (inp[2]) ? node503 : 14'b00000000111111;
										assign node503 = (inp[12]) ? 14'b00000000011111 : node504;
											assign node504 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node508 = (inp[8]) ? node510 : 14'b00000000111111;
									assign node510 = (inp[11]) ? 14'b00000000011111 : 14'b00000000001111;
					assign node513 = (inp[12]) ? node545 : node514;
						assign node514 = (inp[0]) ? node532 : node515;
							assign node515 = (inp[8]) ? node523 : node516;
								assign node516 = (inp[11]) ? 14'b00000001111111 : node517;
									assign node517 = (inp[13]) ? node519 : 14'b00000011111111;
										assign node519 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node523 = (inp[2]) ? node527 : node524;
									assign node524 = (inp[13]) ? 14'b00000001111111 : 14'b00000000111111;
									assign node527 = (inp[10]) ? 14'b00000000011111 : node528;
										assign node528 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node532 = (inp[13]) ? node540 : node533;
								assign node533 = (inp[10]) ? 14'b00000000111111 : node534;
									assign node534 = (inp[9]) ? node536 : 14'b00000001111111;
										assign node536 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node540 = (inp[7]) ? 14'b00000000000111 : node541;
									assign node541 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
						assign node545 = (inp[7]) ? node567 : node546;
							assign node546 = (inp[2]) ? node554 : node547;
								assign node547 = (inp[11]) ? node549 : 14'b00000001111111;
									assign node549 = (inp[5]) ? 14'b00000000111111 : node550;
										assign node550 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node554 = (inp[13]) ? 14'b00000000001111 : node555;
									assign node555 = (inp[8]) ? node559 : node556;
										assign node556 = (inp[9]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node559 = (inp[5]) ? 14'b00000000011111 : node560;
											assign node560 = (inp[11]) ? node562 : 14'b00000000111111;
												assign node562 = (inp[9]) ? 14'b00000000111111 : 14'b00000000011111;
							assign node567 = (inp[10]) ? node573 : node568;
								assign node568 = (inp[2]) ? 14'b00000000011111 : node569;
									assign node569 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node573 = (inp[11]) ? node577 : node574;
									assign node574 = (inp[0]) ? 14'b00000000001111 : 14'b00000000011111;
									assign node577 = (inp[0]) ? 14'b00000000000011 : node578;
										assign node578 = (inp[9]) ? 14'b00000000000111 : 14'b00000000001111;
		assign node582 = (inp[12]) ? node874 : node583;
			assign node583 = (inp[6]) ? node731 : node584;
				assign node584 = (inp[8]) ? node660 : node585;
					assign node585 = (inp[13]) ? node627 : node586;
						assign node586 = (inp[5]) ? node608 : node587;
							assign node587 = (inp[1]) ? node599 : node588;
								assign node588 = (inp[9]) ? node592 : node589;
									assign node589 = (inp[3]) ? 14'b00001111111111 : 14'b00011111111111;
									assign node592 = (inp[7]) ? 14'b00000011111111 : node593;
										assign node593 = (inp[2]) ? node595 : 14'b00001111111111;
											assign node595 = (inp[10]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node599 = (inp[3]) ? node603 : node600;
									assign node600 = (inp[11]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node603 = (inp[7]) ? node605 : 14'b00000111111111;
										assign node605 = (inp[9]) ? 14'b00000001111111 : 14'b00000111111111;
							assign node608 = (inp[0]) ? node614 : node609;
								assign node609 = (inp[9]) ? node611 : 14'b00000111111111;
									assign node611 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node614 = (inp[11]) ? 14'b00000001111111 : node615;
									assign node615 = (inp[7]) ? node623 : node616;
										assign node616 = (inp[2]) ? 14'b00000011111111 : node617;
											assign node617 = (inp[3]) ? node619 : 14'b00000111111111;
												assign node619 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node623 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
						assign node627 = (inp[11]) ? node641 : node628;
							assign node628 = (inp[2]) ? node634 : node629;
								assign node629 = (inp[7]) ? node631 : 14'b00000111111111;
									assign node631 = (inp[9]) ? 14'b00001111111111 : 14'b00000111111111;
								assign node634 = (inp[1]) ? node638 : node635;
									assign node635 = (inp[9]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node638 = (inp[9]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node641 = (inp[5]) ? node649 : node642;
								assign node642 = (inp[10]) ? node646 : node643;
									assign node643 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node646 = (inp[9]) ? 14'b00000011111111 : 14'b00000001111111;
								assign node649 = (inp[7]) ? node651 : 14'b00000001111111;
									assign node651 = (inp[9]) ? node655 : node652;
										assign node652 = (inp[1]) ? 14'b00000000111111 : 14'b00000011111111;
										assign node655 = (inp[1]) ? node657 : 14'b00000000111111;
											assign node657 = (inp[10]) ? 14'b00000000011111 : 14'b00000000001111;
					assign node660 = (inp[13]) ? node696 : node661;
						assign node661 = (inp[2]) ? node677 : node662;
							assign node662 = (inp[5]) ? node666 : node663;
								assign node663 = (inp[7]) ? 14'b00000011111111 : 14'b00001111111111;
								assign node666 = (inp[9]) ? node674 : node667;
									assign node667 = (inp[0]) ? node669 : 14'b00000111111111;
										assign node669 = (inp[1]) ? node671 : 14'b00000011111111;
											assign node671 = (inp[3]) ? 14'b00000000111111 : 14'b00000011111111;
									assign node674 = (inp[10]) ? 14'b00000001111111 : 14'b00000000111111;
							assign node677 = (inp[10]) ? node685 : node678;
								assign node678 = (inp[7]) ? node680 : 14'b00000011111111;
									assign node680 = (inp[0]) ? 14'b00000001111111 : node681;
										assign node681 = (inp[1]) ? 14'b00000001111111 : 14'b00000111111111;
								assign node685 = (inp[0]) ? 14'b00000000111111 : node686;
									assign node686 = (inp[7]) ? node690 : node687;
										assign node687 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node690 = (inp[9]) ? 14'b00000000111111 : node691;
											assign node691 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
						assign node696 = (inp[11]) ? node716 : node697;
							assign node697 = (inp[3]) ? node707 : node698;
								assign node698 = (inp[10]) ? node704 : node699;
									assign node699 = (inp[9]) ? 14'b00000011111111 : node700;
										assign node700 = (inp[2]) ? 14'b00000111111111 : 14'b00000011111111;
									assign node704 = (inp[9]) ? 14'b00000000011111 : 14'b00000011111111;
								assign node707 = (inp[5]) ? 14'b00000000111111 : node708;
									assign node708 = (inp[0]) ? 14'b00000011111111 : node709;
										assign node709 = (inp[2]) ? node711 : 14'b00000001111111;
											assign node711 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node716 = (inp[7]) ? node724 : node717;
								assign node717 = (inp[10]) ? node719 : 14'b00000001111111;
									assign node719 = (inp[2]) ? 14'b00000000011111 : node720;
										assign node720 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node724 = (inp[9]) ? node726 : 14'b00000000111111;
									assign node726 = (inp[0]) ? node728 : 14'b00000000001111;
										assign node728 = (inp[2]) ? 14'b00000000001111 : 14'b00000000011111;
				assign node731 = (inp[13]) ? node801 : node732;
					assign node732 = (inp[8]) ? node752 : node733;
						assign node733 = (inp[3]) ? node741 : node734;
							assign node734 = (inp[5]) ? 14'b00000011111111 : node735;
								assign node735 = (inp[0]) ? 14'b00000011111111 : node736;
									assign node736 = (inp[1]) ? 14'b00000111111111 : 14'b00001111111111;
							assign node741 = (inp[7]) ? node747 : node742;
								assign node742 = (inp[2]) ? node744 : 14'b00000001111111;
									assign node744 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node747 = (inp[0]) ? 14'b00000000111111 : node748;
									assign node748 = (inp[9]) ? 14'b00000000011111 : 14'b00000111111111;
						assign node752 = (inp[7]) ? node774 : node753;
							assign node753 = (inp[2]) ? node765 : node754;
								assign node754 = (inp[3]) ? node760 : node755;
									assign node755 = (inp[9]) ? node757 : 14'b00000011111111;
										assign node757 = (inp[0]) ? 14'b00000011111111 : 14'b00000111111111;
									assign node760 = (inp[9]) ? 14'b00000001111111 : node761;
										assign node761 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node765 = (inp[1]) ? node771 : node766;
									assign node766 = (inp[5]) ? node768 : 14'b00000011111111;
										assign node768 = (inp[11]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node771 = (inp[10]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node774 = (inp[1]) ? node790 : node775;
								assign node775 = (inp[3]) ? node783 : node776;
									assign node776 = (inp[2]) ? node780 : node777;
										assign node777 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node780 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node783 = (inp[0]) ? node787 : node784;
										assign node784 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node787 = (inp[9]) ? 14'b00000000111111 : 14'b00000000011111;
								assign node790 = (inp[10]) ? node796 : node791;
									assign node791 = (inp[0]) ? 14'b00000000001111 : node792;
										assign node792 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node796 = (inp[9]) ? node798 : 14'b00000000011111;
										assign node798 = (inp[3]) ? 14'b00000000000111 : 14'b00000000001111;
					assign node801 = (inp[8]) ? node839 : node802;
						assign node802 = (inp[1]) ? node824 : node803;
							assign node803 = (inp[10]) ? node809 : node804;
								assign node804 = (inp[7]) ? 14'b00000001111111 : node805;
									assign node805 = (inp[11]) ? 14'b00000011111111 : 14'b00000111111111;
								assign node809 = (inp[7]) ? node819 : node810;
									assign node810 = (inp[0]) ? node812 : 14'b00000001111111;
										assign node812 = (inp[2]) ? 14'b00000000111111 : node813;
											assign node813 = (inp[9]) ? node815 : 14'b00000001111111;
												assign node815 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node819 = (inp[0]) ? 14'b00000000011111 : node820;
										assign node820 = (inp[9]) ? 14'b00000001111111 : 14'b00000000111111;
							assign node824 = (inp[3]) ? node836 : node825;
								assign node825 = (inp[9]) ? node833 : node826;
									assign node826 = (inp[11]) ? 14'b00000000111111 : node827;
										assign node827 = (inp[10]) ? 14'b00000000111111 : node828;
											assign node828 = (inp[2]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node833 = (inp[11]) ? 14'b00000000111111 : 14'b00000000011111;
								assign node836 = (inp[7]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node839 = (inp[9]) ? node857 : node840;
							assign node840 = (inp[0]) ? node846 : node841;
								assign node841 = (inp[2]) ? node843 : 14'b00000000111111;
									assign node843 = (inp[1]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node846 = (inp[3]) ? node850 : node847;
									assign node847 = (inp[10]) ? 14'b00000000111111 : 14'b00000000011111;
									assign node850 = (inp[2]) ? 14'b00000000000111 : node851;
										assign node851 = (inp[7]) ? 14'b00000000011111 : node852;
											assign node852 = (inp[11]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node857 = (inp[10]) ? node863 : node858;
								assign node858 = (inp[3]) ? 14'b00000000111111 : node859;
									assign node859 = (inp[2]) ? 14'b00000000001111 : 14'b00000000111111;
								assign node863 = (inp[1]) ? node869 : node864;
									assign node864 = (inp[7]) ? 14'b00000000001111 : node865;
										assign node865 = (inp[0]) ? 14'b00000000011111 : 14'b00000000001111;
									assign node869 = (inp[2]) ? node871 : 14'b00000000011111;
										assign node871 = (inp[11]) ? 14'b00000000000111 : 14'b00000000001111;
			assign node874 = (inp[11]) ? node1014 : node875;
				assign node875 = (inp[2]) ? node927 : node876;
					assign node876 = (inp[8]) ? node904 : node877;
						assign node877 = (inp[9]) ? node893 : node878;
							assign node878 = (inp[7]) ? node886 : node879;
								assign node879 = (inp[13]) ? node883 : node880;
									assign node880 = (inp[10]) ? 14'b00000111111111 : 14'b00001111111111;
									assign node883 = (inp[10]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node886 = (inp[6]) ? node888 : 14'b00000011111111;
									assign node888 = (inp[0]) ? 14'b00000001111111 : node889;
										assign node889 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
							assign node893 = (inp[5]) ? node899 : node894;
								assign node894 = (inp[13]) ? node896 : 14'b00000001111111;
									assign node896 = (inp[10]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node899 = (inp[6]) ? 14'b00000001111111 : node900;
									assign node900 = (inp[1]) ? 14'b00000011111111 : 14'b00000111111111;
						assign node904 = (inp[6]) ? node916 : node905;
							assign node905 = (inp[10]) ? node913 : node906;
								assign node906 = (inp[9]) ? node910 : node907;
									assign node907 = (inp[5]) ? 14'b00001111111111 : 14'b00000111111111;
									assign node910 = (inp[1]) ? 14'b00000011111111 : 14'b00000001111111;
								assign node913 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node916 = (inp[3]) ? node920 : node917;
								assign node917 = (inp[5]) ? 14'b00000000011111 : 14'b00000111111111;
								assign node920 = (inp[13]) ? node922 : 14'b00000000011111;
									assign node922 = (inp[7]) ? node924 : 14'b00000000111111;
										assign node924 = (inp[5]) ? 14'b00000000011111 : 14'b00000000111111;
					assign node927 = (inp[9]) ? node965 : node928;
						assign node928 = (inp[3]) ? node944 : node929;
							assign node929 = (inp[5]) ? node931 : 14'b00000001111111;
								assign node931 = (inp[6]) ? node941 : node932;
									assign node932 = (inp[0]) ? node938 : node933;
										assign node933 = (inp[1]) ? 14'b00000001111111 : node934;
											assign node934 = (inp[7]) ? 14'b00000011111111 : 14'b00000111111111;
										assign node938 = (inp[1]) ? 14'b00000000111111 : 14'b00000001111111;
									assign node941 = (inp[13]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node944 = (inp[1]) ? node958 : node945;
								assign node945 = (inp[0]) ? node949 : node946;
									assign node946 = (inp[7]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node949 = (inp[6]) ? node953 : node950;
										assign node950 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node953 = (inp[5]) ? 14'b00000000011111 : node954;
											assign node954 = (inp[8]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node958 = (inp[7]) ? node960 : 14'b00000000111111;
									assign node960 = (inp[0]) ? 14'b00000000011111 : node961;
										assign node961 = (inp[6]) ? 14'b00000000001111 : 14'b00000000011111;
						assign node965 = (inp[10]) ? node993 : node966;
							assign node966 = (inp[6]) ? node984 : node967;
								assign node967 = (inp[1]) ? node977 : node968;
									assign node968 = (inp[8]) ? node972 : node969;
										assign node969 = (inp[3]) ? 14'b00000001111111 : 14'b00000011111111;
										assign node972 = (inp[7]) ? node974 : 14'b00000001111111;
											assign node974 = (inp[3]) ? 14'b00000000111111 : 14'b00000000011111;
									assign node977 = (inp[13]) ? node979 : 14'b00000000111111;
										assign node979 = (inp[8]) ? 14'b00000000011111 : node980;
											assign node980 = (inp[3]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node984 = (inp[1]) ? node986 : 14'b00000000111111;
									assign node986 = (inp[13]) ? node988 : 14'b00000000011111;
										assign node988 = (inp[8]) ? node990 : 14'b00000000011111;
											assign node990 = (inp[3]) ? 14'b00000000001111 : 14'b00000000000111;
							assign node993 = (inp[7]) ? node1007 : node994;
								assign node994 = (inp[3]) ? node1000 : node995;
									assign node995 = (inp[5]) ? node997 : 14'b00000000111111;
										assign node997 = (inp[0]) ? 14'b00000000111111 : 14'b00000000011111;
									assign node1000 = (inp[8]) ? 14'b00000000001111 : node1001;
										assign node1001 = (inp[1]) ? node1003 : 14'b00000000011111;
											assign node1003 = (inp[13]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node1007 = (inp[8]) ? node1009 : 14'b00000000001111;
									assign node1009 = (inp[5]) ? 14'b00000000000111 : node1010;
										assign node1010 = (inp[13]) ? 14'b00000000000111 : 14'b00000000001111;
				assign node1014 = (inp[1]) ? node1074 : node1015;
					assign node1015 = (inp[9]) ? node1043 : node1016;
						assign node1016 = (inp[3]) ? node1026 : node1017;
							assign node1017 = (inp[0]) ? node1019 : 14'b00000111111111;
								assign node1019 = (inp[2]) ? node1023 : node1020;
									assign node1020 = (inp[5]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1023 = (inp[5]) ? 14'b00000000111111 : 14'b00000001111111;
							assign node1026 = (inp[8]) ? node1040 : node1027;
								assign node1027 = (inp[7]) ? node1031 : node1028;
									assign node1028 = (inp[13]) ? 14'b00000001111111 : 14'b00000011111111;
									assign node1031 = (inp[13]) ? node1037 : node1032;
										assign node1032 = (inp[5]) ? node1034 : 14'b00000011111111;
											assign node1034 = (inp[0]) ? 14'b00000000111111 : 14'b00000001111111;
										assign node1037 = (inp[0]) ? 14'b00000000001111 : 14'b00000000111111;
								assign node1040 = (inp[13]) ? 14'b00000000011111 : 14'b00000000001111;
						assign node1043 = (inp[5]) ? node1057 : node1044;
							assign node1044 = (inp[2]) ? node1050 : node1045;
								assign node1045 = (inp[13]) ? 14'b00000000011111 : node1046;
									assign node1046 = (inp[0]) ? 14'b00000001111111 : 14'b00000011111111;
								assign node1050 = (inp[8]) ? 14'b00000000011111 : node1051;
									assign node1051 = (inp[0]) ? 14'b00000000011111 : node1052;
										assign node1052 = (inp[7]) ? 14'b00000000011111 : 14'b00000000111111;
							assign node1057 = (inp[7]) ? node1067 : node1058;
								assign node1058 = (inp[6]) ? node1062 : node1059;
									assign node1059 = (inp[8]) ? 14'b00000000011111 : 14'b00000001111111;
									assign node1062 = (inp[13]) ? 14'b00000000000111 : node1063;
										assign node1063 = (inp[8]) ? 14'b00000000011111 : 14'b00000000001111;
								assign node1067 = (inp[8]) ? node1069 : 14'b00000000001111;
									assign node1069 = (inp[10]) ? node1071 : 14'b00000000001111;
										assign node1071 = (inp[13]) ? 14'b00000000000011 : 14'b00000000000111;
					assign node1074 = (inp[13]) ? node1102 : node1075;
						assign node1075 = (inp[5]) ? node1085 : node1076;
							assign node1076 = (inp[7]) ? node1080 : node1077;
								assign node1077 = (inp[8]) ? 14'b00000000111111 : 14'b00000001111111;
								assign node1080 = (inp[2]) ? node1082 : 14'b00000000011111;
									assign node1082 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node1085 = (inp[9]) ? node1093 : node1086;
								assign node1086 = (inp[8]) ? node1088 : 14'b00000000011111;
									assign node1088 = (inp[7]) ? node1090 : 14'b00000000011111;
										assign node1090 = (inp[2]) ? 14'b00000000011111 : 14'b00000000111111;
								assign node1093 = (inp[10]) ? node1099 : node1094;
									assign node1094 = (inp[0]) ? 14'b00000000000111 : node1095;
										assign node1095 = (inp[3]) ? 14'b00000000011111 : 14'b00000000111111;
									assign node1099 = (inp[3]) ? 14'b00000000000111 : 14'b00000000001111;
						assign node1102 = (inp[6]) ? node1116 : node1103;
							assign node1103 = (inp[2]) ? node1111 : node1104;
								assign node1104 = (inp[0]) ? node1106 : 14'b00000000111111;
									assign node1106 = (inp[3]) ? node1108 : 14'b00000000011111;
										assign node1108 = (inp[8]) ? 14'b00000000001111 : 14'b00000000011111;
								assign node1111 = (inp[3]) ? node1113 : 14'b00000000000111;
									assign node1113 = (inp[10]) ? 14'b00000000001111 : 14'b00000000011111;
							assign node1116 = (inp[10]) ? node1126 : node1117;
								assign node1117 = (inp[0]) ? node1119 : 14'b00000000011111;
									assign node1119 = (inp[7]) ? 14'b00000000000111 : node1120;
										assign node1120 = (inp[5]) ? node1122 : 14'b00000000001111;
											assign node1122 = (inp[9]) ? 14'b00000000001111 : 14'b00000000000111;
								assign node1126 = (inp[3]) ? node1132 : node1127;
									assign node1127 = (inp[7]) ? node1129 : 14'b00000000011111;
										assign node1129 = (inp[0]) ? 14'b00000000001111 : 14'b00000000000011;
									assign node1132 = (inp[7]) ? 14'b00000000000011 : node1133;
										assign node1133 = (inp[2]) ? node1135 : 14'b00000000001111;
											assign node1135 = (inp[0]) ? node1137 : 14'b00000000000111;
												assign node1137 = (inp[8]) ? 14'b00000000000011 : 14'b00000000000111;

endmodule