module dtc_split75_bm48 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node6;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node10;
	wire [14-1:0] node11;
	wire [14-1:0] node13;
	wire [14-1:0] node16;
	wire [14-1:0] node17;
	wire [14-1:0] node18;
	wire [14-1:0] node19;
	wire [14-1:0] node25;
	wire [14-1:0] node27;
	wire [14-1:0] node28;
	wire [14-1:0] node29;
	wire [14-1:0] node34;
	wire [14-1:0] node36;
	wire [14-1:0] node38;
	wire [14-1:0] node40;
	wire [14-1:0] node41;
	wire [14-1:0] node42;
	wire [14-1:0] node47;
	wire [14-1:0] node48;
	wire [14-1:0] node49;
	wire [14-1:0] node50;
	wire [14-1:0] node51;
	wire [14-1:0] node52;
	wire [14-1:0] node54;
	wire [14-1:0] node55;
	wire [14-1:0] node57;
	wire [14-1:0] node62;
	wire [14-1:0] node63;
	wire [14-1:0] node64;
	wire [14-1:0] node66;
	wire [14-1:0] node71;
	wire [14-1:0] node73;
	wire [14-1:0] node74;
	wire [14-1:0] node75;
	wire [14-1:0] node76;
	wire [14-1:0] node78;
	wire [14-1:0] node81;
	wire [14-1:0] node82;
	wire [14-1:0] node89;
	wire [14-1:0] node90;
	wire [14-1:0] node92;
	wire [14-1:0] node93;
	wire [14-1:0] node94;
	wire [14-1:0] node95;
	wire [14-1:0] node98;
	wire [14-1:0] node99;
	wire [14-1:0] node103;
	wire [14-1:0] node104;
	wire [14-1:0] node105;
	wire [14-1:0] node106;
	wire [14-1:0] node113;
	wire [14-1:0] node114;
	wire [14-1:0] node116;
	wire [14-1:0] node119;
	wire [14-1:0] node121;
	wire [14-1:0] node123;
	wire [14-1:0] node124;
	wire [14-1:0] node125;
	wire [14-1:0] node126;
	wire [14-1:0] node132;
	wire [14-1:0] node133;
	wire [14-1:0] node135;
	wire [14-1:0] node136;
	wire [14-1:0] node137;
	wire [14-1:0] node138;
	wire [14-1:0] node139;
	wire [14-1:0] node140;
	wire [14-1:0] node142;
	wire [14-1:0] node147;
	wire [14-1:0] node149;
	wire [14-1:0] node150;
	wire [14-1:0] node153;
	wire [14-1:0] node155;
	wire [14-1:0] node156;
	wire [14-1:0] node160;
	wire [14-1:0] node161;
	wire [14-1:0] node162;
	wire [14-1:0] node163;
	wire [14-1:0] node164;
	wire [14-1:0] node167;
	wire [14-1:0] node168;
	wire [14-1:0] node175;
	wire [14-1:0] node176;
	wire [14-1:0] node178;
	wire [14-1:0] node179;
	wire [14-1:0] node181;
	wire [14-1:0] node182;
	wire [14-1:0] node187;
	wire [14-1:0] node188;
	wire [14-1:0] node189;
	wire [14-1:0] node190;
	wire [14-1:0] node195;
	wire [14-1:0] node196;
	wire [14-1:0] node198;
	wire [14-1:0] node199;
	wire [14-1:0] node200;
	wire [14-1:0] node206;
	wire [14-1:0] node207;
	wire [14-1:0] node208;
	wire [14-1:0] node210;
	wire [14-1:0] node212;
	wire [14-1:0] node215;
	wire [14-1:0] node216;
	wire [14-1:0] node217;
	wire [14-1:0] node220;
	wire [14-1:0] node221;
	wire [14-1:0] node223;
	wire [14-1:0] node224;
	wire [14-1:0] node229;
	wire [14-1:0] node230;
	wire [14-1:0] node231;
	wire [14-1:0] node232;
	wire [14-1:0] node234;
	wire [14-1:0] node235;
	wire [14-1:0] node242;
	wire [14-1:0] node243;
	wire [14-1:0] node245;
	wire [14-1:0] node246;
	wire [14-1:0] node247;
	wire [14-1:0] node248;
	wire [14-1:0] node250;
	wire [14-1:0] node256;
	wire [14-1:0] node257;
	wire [14-1:0] node259;
	wire [14-1:0] node260;
	wire [14-1:0] node261;
	wire [14-1:0] node263;
	wire [14-1:0] node266;
	wire [14-1:0] node267;
	wire [14-1:0] node269;
	wire [14-1:0] node274;
	wire [14-1:0] node275;
	wire [14-1:0] node277;
	wire [14-1:0] node279;
	wire [14-1:0] node282;
	wire [14-1:0] node284;
	wire [14-1:0] node286;
	wire [14-1:0] node289;
	wire [14-1:0] node290;
	wire [14-1:0] node291;
	wire [14-1:0] node293;
	wire [14-1:0] node295;
	wire [14-1:0] node296;
	wire [14-1:0] node297;
	wire [14-1:0] node298;
	wire [14-1:0] node303;
	wire [14-1:0] node304;
	wire [14-1:0] node305;
	wire [14-1:0] node306;
	wire [14-1:0] node307;
	wire [14-1:0] node314;
	wire [14-1:0] node315;
	wire [14-1:0] node316;
	wire [14-1:0] node317;
	wire [14-1:0] node318;
	wire [14-1:0] node322;
	wire [14-1:0] node324;
	wire [14-1:0] node326;
	wire [14-1:0] node328;
	wire [14-1:0] node329;
	wire [14-1:0] node330;
	wire [14-1:0] node333;
	wire [14-1:0] node337;
	wire [14-1:0] node338;
	wire [14-1:0] node340;
	wire [14-1:0] node342;
	wire [14-1:0] node343;
	wire [14-1:0] node345;
	wire [14-1:0] node348;
	wire [14-1:0] node350;
	wire [14-1:0] node352;
	wire [14-1:0] node356;
	wire [14-1:0] node357;
	wire [14-1:0] node358;
	wire [14-1:0] node359;
	wire [14-1:0] node360;
	wire [14-1:0] node361;
	wire [14-1:0] node362;
	wire [14-1:0] node364;
	wire [14-1:0] node367;
	wire [14-1:0] node370;
	wire [14-1:0] node371;
	wire [14-1:0] node375;
	wire [14-1:0] node377;
	wire [14-1:0] node378;
	wire [14-1:0] node382;
	wire [14-1:0] node384;
	wire [14-1:0] node385;
	wire [14-1:0] node386;
	wire [14-1:0] node391;
	wire [14-1:0] node392;
	wire [14-1:0] node394;
	wire [14-1:0] node395;
	wire [14-1:0] node396;
	wire [14-1:0] node399;
	wire [14-1:0] node404;
	wire [14-1:0] node406;
	wire [14-1:0] node408;
	wire [14-1:0] node410;
	wire [14-1:0] node411;
	wire [14-1:0] node412;
	wire [14-1:0] node413;
	wire [14-1:0] node418;
	wire [14-1:0] node421;
	wire [14-1:0] node422;
	wire [14-1:0] node423;
	wire [14-1:0] node425;
	wire [14-1:0] node426;
	wire [14-1:0] node427;
	wire [14-1:0] node429;
	wire [14-1:0] node430;
	wire [14-1:0] node431;
	wire [14-1:0] node432;
	wire [14-1:0] node438;
	wire [14-1:0] node439;
	wire [14-1:0] node440;
	wire [14-1:0] node441;
	wire [14-1:0] node442;
	wire [14-1:0] node447;
	wire [14-1:0] node448;
	wire [14-1:0] node452;
	wire [14-1:0] node454;
	wire [14-1:0] node455;
	wire [14-1:0] node456;
	wire [14-1:0] node461;
	wire [14-1:0] node463;
	wire [14-1:0] node464;
	wire [14-1:0] node465;
	wire [14-1:0] node466;
	wire [14-1:0] node472;
	wire [14-1:0] node473;
	wire [14-1:0] node474;
	wire [14-1:0] node476;
	wire [14-1:0] node477;
	wire [14-1:0] node479;
	wire [14-1:0] node480;
	wire [14-1:0] node481;
	wire [14-1:0] node485;
	wire [14-1:0] node486;
	wire [14-1:0] node492;
	wire [14-1:0] node493;
	wire [14-1:0] node494;
	wire [14-1:0] node495;
	wire [14-1:0] node496;
	wire [14-1:0] node497;
	wire [14-1:0] node498;
	wire [14-1:0] node505;
	wire [14-1:0] node506;
	wire [14-1:0] node507;
	wire [14-1:0] node508;
	wire [14-1:0] node509;
	wire [14-1:0] node515;
	wire [14-1:0] node517;
	wire [14-1:0] node520;
	wire [14-1:0] node522;
	wire [14-1:0] node523;
	wire [14-1:0] node527;
	wire [14-1:0] node528;
	wire [14-1:0] node529;
	wire [14-1:0] node530;
	wire [14-1:0] node531;
	wire [14-1:0] node533;
	wire [14-1:0] node534;
	wire [14-1:0] node535;
	wire [14-1:0] node538;
	wire [14-1:0] node541;
	wire [14-1:0] node542;
	wire [14-1:0] node548;
	wire [14-1:0] node549;
	wire [14-1:0] node550;
	wire [14-1:0] node552;
	wire [14-1:0] node553;
	wire [14-1:0] node555;
	wire [14-1:0] node556;
	wire [14-1:0] node559;
	wire [14-1:0] node562;
	wire [14-1:0] node566;
	wire [14-1:0] node568;
	wire [14-1:0] node570;
	wire [14-1:0] node572;
	wire [14-1:0] node576;
	wire [14-1:0] node577;
	wire [14-1:0] node578;
	wire [14-1:0] node579;
	wire [14-1:0] node580;
	wire [14-1:0] node581;
	wire [14-1:0] node582;
	wire [14-1:0] node583;
	wire [14-1:0] node584;
	wire [14-1:0] node585;
	wire [14-1:0] node590;
	wire [14-1:0] node592;
	wire [14-1:0] node594;
	wire [14-1:0] node597;
	wire [14-1:0] node598;
	wire [14-1:0] node599;
	wire [14-1:0] node600;
	wire [14-1:0] node601;
	wire [14-1:0] node602;
	wire [14-1:0] node607;
	wire [14-1:0] node609;
	wire [14-1:0] node611;
	wire [14-1:0] node614;
	wire [14-1:0] node615;
	wire [14-1:0] node616;
	wire [14-1:0] node617;
	wire [14-1:0] node623;
	wire [14-1:0] node624;
	wire [14-1:0] node625;
	wire [14-1:0] node626;
	wire [14-1:0] node627;
	wire [14-1:0] node632;
	wire [14-1:0] node634;
	wire [14-1:0] node636;
	wire [14-1:0] node639;
	wire [14-1:0] node640;
	wire [14-1:0] node641;
	wire [14-1:0] node642;
	wire [14-1:0] node647;
	wire [14-1:0] node649;
	wire [14-1:0] node651;
	wire [14-1:0] node654;
	wire [14-1:0] node655;
	wire [14-1:0] node656;
	wire [14-1:0] node657;
	wire [14-1:0] node662;
	wire [14-1:0] node664;
	wire [14-1:0] node666;
	wire [14-1:0] node669;
	wire [14-1:0] node670;
	wire [14-1:0] node671;
	wire [14-1:0] node672;
	wire [14-1:0] node673;
	wire [14-1:0] node678;
	wire [14-1:0] node680;
	wire [14-1:0] node682;
	wire [14-1:0] node685;
	wire [14-1:0] node686;
	wire [14-1:0] node687;
	wire [14-1:0] node688;
	wire [14-1:0] node693;
	wire [14-1:0] node695;
	wire [14-1:0] node697;
	wire [14-1:0] node700;
	wire [14-1:0] node701;
	wire [14-1:0] node702;
	wire [14-1:0] node703;
	wire [14-1:0] node704;
	wire [14-1:0] node705;
	wire [14-1:0] node706;
	wire [14-1:0] node707;
	wire [14-1:0] node712;
	wire [14-1:0] node714;
	wire [14-1:0] node716;
	wire [14-1:0] node719;
	wire [14-1:0] node720;
	wire [14-1:0] node721;
	wire [14-1:0] node722;
	wire [14-1:0] node727;
	wire [14-1:0] node729;
	wire [14-1:0] node731;
	wire [14-1:0] node734;
	wire [14-1:0] node736;
	wire [14-1:0] node737;
	wire [14-1:0] node738;
	wire [14-1:0] node739;
	wire [14-1:0] node740;
	wire [14-1:0] node746;
	wire [14-1:0] node747;
	wire [14-1:0] node748;
	wire [14-1:0] node752;
	wire [14-1:0] node754;
	wire [14-1:0] node756;
	wire [14-1:0] node759;
	wire [14-1:0] node760;
	wire [14-1:0] node761;
	wire [14-1:0] node762;
	wire [14-1:0] node763;
	wire [14-1:0] node768;
	wire [14-1:0] node770;
	wire [14-1:0] node772;
	wire [14-1:0] node775;
	wire [14-1:0] node776;
	wire [14-1:0] node777;
	wire [14-1:0] node778;
	wire [14-1:0] node779;
	wire [14-1:0] node784;
	wire [14-1:0] node786;
	wire [14-1:0] node788;
	wire [14-1:0] node791;
	wire [14-1:0] node792;
	wire [14-1:0] node793;
	wire [14-1:0] node794;
	wire [14-1:0] node799;
	wire [14-1:0] node801;
	wire [14-1:0] node803;
	wire [14-1:0] node806;
	wire [14-1:0] node807;
	wire [14-1:0] node808;
	wire [14-1:0] node809;
	wire [14-1:0] node810;
	wire [14-1:0] node811;
	wire [14-1:0] node812;
	wire [14-1:0] node817;
	wire [14-1:0] node819;
	wire [14-1:0] node821;
	wire [14-1:0] node824;
	wire [14-1:0] node825;
	wire [14-1:0] node826;
	wire [14-1:0] node827;
	wire [14-1:0] node832;
	wire [14-1:0] node834;
	wire [14-1:0] node836;
	wire [14-1:0] node839;
	wire [14-1:0] node840;
	wire [14-1:0] node841;
	wire [14-1:0] node842;
	wire [14-1:0] node847;
	wire [14-1:0] node849;
	wire [14-1:0] node851;
	wire [14-1:0] node854;
	wire [14-1:0] node855;
	wire [14-1:0] node856;
	wire [14-1:0] node857;
	wire [14-1:0] node858;
	wire [14-1:0] node859;
	wire [14-1:0] node864;
	wire [14-1:0] node866;
	wire [14-1:0] node868;
	wire [14-1:0] node871;
	wire [14-1:0] node872;
	wire [14-1:0] node873;
	wire [14-1:0] node874;
	wire [14-1:0] node879;
	wire [14-1:0] node881;
	wire [14-1:0] node883;
	wire [14-1:0] node886;
	wire [14-1:0] node887;
	wire [14-1:0] node888;
	wire [14-1:0] node889;
	wire [14-1:0] node890;
	wire [14-1:0] node895;
	wire [14-1:0] node897;
	wire [14-1:0] node899;
	wire [14-1:0] node902;
	wire [14-1:0] node903;
	wire [14-1:0] node904;
	wire [14-1:0] node905;
	wire [14-1:0] node906;
	wire [14-1:0] node911;
	wire [14-1:0] node913;
	wire [14-1:0] node915;
	wire [14-1:0] node918;
	wire [14-1:0] node919;
	wire [14-1:0] node920;
	wire [14-1:0] node921;
	wire [14-1:0] node926;
	wire [14-1:0] node928;
	wire [14-1:0] node930;
	wire [14-1:0] node933;
	wire [14-1:0] node934;
	wire [14-1:0] node935;
	wire [14-1:0] node936;
	wire [14-1:0] node937;
	wire [14-1:0] node938;
	wire [14-1:0] node939;
	wire [14-1:0] node941;
	wire [14-1:0] node942;
	wire [14-1:0] node943;
	wire [14-1:0] node948;
	wire [14-1:0] node949;
	wire [14-1:0] node950;
	wire [14-1:0] node953;
	wire [14-1:0] node955;
	wire [14-1:0] node958;
	wire [14-1:0] node960;
	wire [14-1:0] node962;
	wire [14-1:0] node965;
	wire [14-1:0] node966;
	wire [14-1:0] node967;
	wire [14-1:0] node968;
	wire [14-1:0] node973;
	wire [14-1:0] node975;
	wire [14-1:0] node977;
	wire [14-1:0] node980;
	wire [14-1:0] node981;
	wire [14-1:0] node982;
	wire [14-1:0] node983;
	wire [14-1:0] node984;
	wire [14-1:0] node989;
	wire [14-1:0] node991;
	wire [14-1:0] node993;
	wire [14-1:0] node996;
	wire [14-1:0] node997;
	wire [14-1:0] node998;
	wire [14-1:0] node999;
	wire [14-1:0] node1000;
	wire [14-1:0] node1005;
	wire [14-1:0] node1007;
	wire [14-1:0] node1009;
	wire [14-1:0] node1012;
	wire [14-1:0] node1013;
	wire [14-1:0] node1014;
	wire [14-1:0] node1015;
	wire [14-1:0] node1020;
	wire [14-1:0] node1022;
	wire [14-1:0] node1024;
	wire [14-1:0] node1027;
	wire [14-1:0] node1028;
	wire [14-1:0] node1029;
	wire [14-1:0] node1030;
	wire [14-1:0] node1031;
	wire [14-1:0] node1036;
	wire [14-1:0] node1038;
	wire [14-1:0] node1040;
	wire [14-1:0] node1043;
	wire [14-1:0] node1044;
	wire [14-1:0] node1045;
	wire [14-1:0] node1046;
	wire [14-1:0] node1047;
	wire [14-1:0] node1052;
	wire [14-1:0] node1054;
	wire [14-1:0] node1056;
	wire [14-1:0] node1059;
	wire [14-1:0] node1060;
	wire [14-1:0] node1061;
	wire [14-1:0] node1062;
	wire [14-1:0] node1063;
	wire [14-1:0] node1068;
	wire [14-1:0] node1070;
	wire [14-1:0] node1072;
	wire [14-1:0] node1076;
	wire [14-1:0] node1077;
	wire [14-1:0] node1078;
	wire [14-1:0] node1079;
	wire [14-1:0] node1084;
	wire [14-1:0] node1086;
	wire [14-1:0] node1088;
	wire [14-1:0] node1091;
	wire [14-1:0] node1092;
	wire [14-1:0] node1093;
	wire [14-1:0] node1094;
	wire [14-1:0] node1098;
	wire [14-1:0] node1099;
	wire [14-1:0] node1101;
	wire [14-1:0] node1103;
	wire [14-1:0] node1104;
	wire [14-1:0] node1105;
	wire [14-1:0] node1106;
	wire [14-1:0] node1113;
	wire [14-1:0] node1114;
	wire [14-1:0] node1115;
	wire [14-1:0] node1116;
	wire [14-1:0] node1117;
	wire [14-1:0] node1118;
	wire [14-1:0] node1119;
	wire [14-1:0] node1120;
	wire [14-1:0] node1127;
	wire [14-1:0] node1130;
	wire [14-1:0] node1131;
	wire [14-1:0] node1135;
	wire [14-1:0] node1136;
	wire [14-1:0] node1137;
	wire [14-1:0] node1138;
	wire [14-1:0] node1139;
	wire [14-1:0] node1140;
	wire [14-1:0] node1141;
	wire [14-1:0] node1148;
	wire [14-1:0] node1151;
	wire [14-1:0] node1152;
	wire [14-1:0] node1156;
	wire [14-1:0] node1157;
	wire [14-1:0] node1158;
	wire [14-1:0] node1159;
	wire [14-1:0] node1161;
	wire [14-1:0] node1162;
	wire [14-1:0] node1163;
	wire [14-1:0] node1164;
	wire [14-1:0] node1165;
	wire [14-1:0] node1167;
	wire [14-1:0] node1168;
	wire [14-1:0] node1172;
	wire [14-1:0] node1173;
	wire [14-1:0] node1176;
	wire [14-1:0] node1179;
	wire [14-1:0] node1181;
	wire [14-1:0] node1183;
	wire [14-1:0] node1187;
	wire [14-1:0] node1189;
	wire [14-1:0] node1191;
	wire [14-1:0] node1193;
	wire [14-1:0] node1194;
	wire [14-1:0] node1198;
	wire [14-1:0] node1199;
	wire [14-1:0] node1200;
	wire [14-1:0] node1201;
	wire [14-1:0] node1202;
	wire [14-1:0] node1204;
	wire [14-1:0] node1205;
	wire [14-1:0] node1206;
	wire [14-1:0] node1211;
	wire [14-1:0] node1212;
	wire [14-1:0] node1213;
	wire [14-1:0] node1216;
	wire [14-1:0] node1219;
	wire [14-1:0] node1220;
	wire [14-1:0] node1223;
	wire [14-1:0] node1226;
	wire [14-1:0] node1227;
	wire [14-1:0] node1228;
	wire [14-1:0] node1229;
	wire [14-1:0] node1232;
	wire [14-1:0] node1234;
	wire [14-1:0] node1239;
	wire [14-1:0] node1240;
	wire [14-1:0] node1241;
	wire [14-1:0] node1242;
	wire [14-1:0] node1244;
	wire [14-1:0] node1250;
	wire [14-1:0] node1252;
	wire [14-1:0] node1254;
	wire [14-1:0] node1256;
	wire [14-1:0] node1257;
	wire [14-1:0] node1258;
	wire [14-1:0] node1259;
	wire [14-1:0] node1264;
	wire [14-1:0] node1266;
	wire [14-1:0] node1269;
	wire [14-1:0] node1270;
	wire [14-1:0] node1271;
	wire [14-1:0] node1272;
	wire [14-1:0] node1273;
	wire [14-1:0] node1275;
	wire [14-1:0] node1277;
	wire [14-1:0] node1278;
	wire [14-1:0] node1282;
	wire [14-1:0] node1283;
	wire [14-1:0] node1284;
	wire [14-1:0] node1285;
	wire [14-1:0] node1288;
	wire [14-1:0] node1291;
	wire [14-1:0] node1293;
	wire [14-1:0] node1297;
	wire [14-1:0] node1299;
	wire [14-1:0] node1300;
	wire [14-1:0] node1301;
	wire [14-1:0] node1302;
	wire [14-1:0] node1304;
	wire [14-1:0] node1307;
	wire [14-1:0] node1308;
	wire [14-1:0] node1312;
	wire [14-1:0] node1313;
	wire [14-1:0] node1315;
	wire [14-1:0] node1318;
	wire [14-1:0] node1321;
	wire [14-1:0] node1323;
	wire [14-1:0] node1325;
	wire [14-1:0] node1326;
	wire [14-1:0] node1330;
	wire [14-1:0] node1331;
	wire [14-1:0] node1332;
	wire [14-1:0] node1333;
	wire [14-1:0] node1334;
	wire [14-1:0] node1335;
	wire [14-1:0] node1336;
	wire [14-1:0] node1341;
	wire [14-1:0] node1343;
	wire [14-1:0] node1345;
	wire [14-1:0] node1349;
	wire [14-1:0] node1350;
	wire [14-1:0] node1351;
	wire [14-1:0] node1352;
	wire [14-1:0] node1353;
	wire [14-1:0] node1359;
	wire [14-1:0] node1361;
	wire [14-1:0] node1362;
	wire [14-1:0] node1364;
	wire [14-1:0] node1368;
	wire [14-1:0] node1369;
	wire [14-1:0] node1370;
	wire [14-1:0] node1372;
	wire [14-1:0] node1374;
	wire [14-1:0] node1375;
	wire [14-1:0] node1381;
	wire [14-1:0] node1382;
	wire [14-1:0] node1383;
	wire [14-1:0] node1384;
	wire [14-1:0] node1386;
	wire [14-1:0] node1387;
	wire [14-1:0] node1388;
	wire [14-1:0] node1389;
	wire [14-1:0] node1397;
	wire [14-1:0] node1398;
	wire [14-1:0] node1399;
	wire [14-1:0] node1400;
	wire [14-1:0] node1401;
	wire [14-1:0] node1402;
	wire [14-1:0] node1404;
	wire [14-1:0] node1411;
	wire [14-1:0] node1413;
	wire [14-1:0] node1415;
	wire [14-1:0] node1416;
	wire [14-1:0] node1417;
	wire [14-1:0] node1421;
	wire [14-1:0] node1422;
	wire [14-1:0] node1426;
	wire [14-1:0] node1427;
	wire [14-1:0] node1428;
	wire [14-1:0] node1429;
	wire [14-1:0] node1430;
	wire [14-1:0] node1431;
	wire [14-1:0] node1432;
	wire [14-1:0] node1434;
	wire [14-1:0] node1436;
	wire [14-1:0] node1440;
	wire [14-1:0] node1442;
	wire [14-1:0] node1443;
	wire [14-1:0] node1444;
	wire [14-1:0] node1445;
	wire [14-1:0] node1451;
	wire [14-1:0] node1452;
	wire [14-1:0] node1454;
	wire [14-1:0] node1456;
	wire [14-1:0] node1458;
	wire [14-1:0] node1459;
	wire [14-1:0] node1462;
	wire [14-1:0] node1466;
	wire [14-1:0] node1467;
	wire [14-1:0] node1468;
	wire [14-1:0] node1470;
	wire [14-1:0] node1471;
	wire [14-1:0] node1472;
	wire [14-1:0] node1478;
	wire [14-1:0] node1479;
	wire [14-1:0] node1480;
	wire [14-1:0] node1482;
	wire [14-1:0] node1483;
	wire [14-1:0] node1489;
	wire [14-1:0] node1490;
	wire [14-1:0] node1491;
	wire [14-1:0] node1492;
	wire [14-1:0] node1493;
	wire [14-1:0] node1494;
	wire [14-1:0] node1495;
	wire [14-1:0] node1497;
	wire [14-1:0] node1500;
	wire [14-1:0] node1503;
	wire [14-1:0] node1504;
	wire [14-1:0] node1505;
	wire [14-1:0] node1513;
	wire [14-1:0] node1514;
	wire [14-1:0] node1515;
	wire [14-1:0] node1516;
	wire [14-1:0] node1517;
	wire [14-1:0] node1518;
	wire [14-1:0] node1521;
	wire [14-1:0] node1524;
	wire [14-1:0] node1526;
	wire [14-1:0] node1531;
	wire [14-1:0] node1532;
	wire [14-1:0] node1534;
	wire [14-1:0] node1535;
	wire [14-1:0] node1536;
	wire [14-1:0] node1537;
	wire [14-1:0] node1542;
	wire [14-1:0] node1543;
	wire [14-1:0] node1544;
	wire [14-1:0] node1549;
	wire [14-1:0] node1550;
	wire [14-1:0] node1551;
	wire [14-1:0] node1555;
	wire [14-1:0] node1556;
	wire [14-1:0] node1559;
	wire [14-1:0] node1562;
	wire [14-1:0] node1563;
	wire [14-1:0] node1564;
	wire [14-1:0] node1565;
	wire [14-1:0] node1566;
	wire [14-1:0] node1567;
	wire [14-1:0] node1568;
	wire [14-1:0] node1572;
	wire [14-1:0] node1573;
	wire [14-1:0] node1575;
	wire [14-1:0] node1576;
	wire [14-1:0] node1581;
	wire [14-1:0] node1583;
	wire [14-1:0] node1584;
	wire [14-1:0] node1586;
	wire [14-1:0] node1587;
	wire [14-1:0] node1592;
	wire [14-1:0] node1594;
	wire [14-1:0] node1596;
	wire [14-1:0] node1597;
	wire [14-1:0] node1599;
	wire [14-1:0] node1601;
	wire [14-1:0] node1605;
	wire [14-1:0] node1606;
	wire [14-1:0] node1607;
	wire [14-1:0] node1608;
	wire [14-1:0] node1609;
	wire [14-1:0] node1610;
	wire [14-1:0] node1617;
	wire [14-1:0] node1619;
	wire [14-1:0] node1621;
	wire [14-1:0] node1622;
	wire [14-1:0] node1623;
	wire [14-1:0] node1624;
	wire [14-1:0] node1629;
	wire [14-1:0] node1632;
	wire [14-1:0] node1633;
	wire [14-1:0] node1634;
	wire [14-1:0] node1635;
	wire [14-1:0] node1636;
	wire [14-1:0] node1637;
	wire [14-1:0] node1638;
	wire [14-1:0] node1641;
	wire [14-1:0] node1645;
	wire [14-1:0] node1646;
	wire [14-1:0] node1647;
	wire [14-1:0] node1648;
	wire [14-1:0] node1654;
	wire [14-1:0] node1655;
	wire [14-1:0] node1657;
	wire [14-1:0] node1658;
	wire [14-1:0] node1659;
	wire [14-1:0] node1665;
	wire [14-1:0] node1666;
	wire [14-1:0] node1668;
	wire [14-1:0] node1670;

	assign outp = (inp[10]) ? node576 : node1;
		assign node1 = (inp[13]) ? node289 : node2;
			assign node2 = (inp[11]) ? node132 : node3;
				assign node3 = (inp[12]) ? node47 : node4;
					assign node4 = (inp[8]) ? node6 : 14'b00000100000011;
						assign node6 = (inp[1]) ? node8 : 14'b00000000000000;
							assign node8 = (inp[6]) ? node34 : node9;
								assign node9 = (inp[2]) ? node25 : node10;
									assign node10 = (inp[0]) ? node16 : node11;
										assign node11 = (inp[3]) ? node13 : 14'b00000000000000;
											assign node13 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
										assign node16 = (inp[5]) ? 14'b00000000000000 : node17;
											assign node17 = (inp[3]) ? 14'b00000000000000 : node18;
												assign node18 = (inp[9]) ? 14'b00000000000000 : node19;
													assign node19 = (inp[4]) ? 14'b00000000000000 : 14'b00100100001100;
									assign node25 = (inp[0]) ? node27 : 14'b00000000000000;
										assign node27 = (inp[4]) ? 14'b00000000000000 : node28;
											assign node28 = (inp[3]) ? 14'b00000000000000 : node29;
												assign node29 = (inp[9]) ? 14'b00000000000000 : 14'b10000000011010;
								assign node34 = (inp[3]) ? node36 : 14'b00000000000000;
									assign node36 = (inp[7]) ? node38 : 14'b00000000000000;
										assign node38 = (inp[9]) ? node40 : 14'b00000000000000;
											assign node40 = (inp[5]) ? 14'b00000000011100 : node41;
												assign node41 = (inp[0]) ? 14'b00000000000000 : node42;
													assign node42 = (inp[2]) ? 14'b00000000000000 : 14'b01000000010000;
					assign node47 = (inp[8]) ? node89 : node48;
						assign node48 = (inp[9]) ? 14'b00000000000000 : node49;
							assign node49 = (inp[7]) ? node71 : node50;
								assign node50 = (inp[3]) ? node62 : node51;
									assign node51 = (inp[4]) ? 14'b00000000000000 : node52;
										assign node52 = (inp[1]) ? node54 : 14'b00000000000000;
											assign node54 = (inp[6]) ? 14'b00000000000000 : node55;
												assign node55 = (inp[0]) ? node57 : 14'b00000000000000;
													assign node57 = (inp[5]) ? 14'b00000000000000 : 14'b00100000000011;
									assign node62 = (inp[0]) ? 14'b00000000000000 : node63;
										assign node63 = (inp[1]) ? 14'b00000000000000 : node64;
											assign node64 = (inp[6]) ? node66 : 14'b00000000000000;
												assign node66 = (inp[2]) ? 14'b00000000000000 : 14'b00100000000011;
								assign node71 = (inp[1]) ? node73 : 14'b00000000000000;
									assign node73 = (inp[3]) ? 14'b00000000000000 : node74;
										assign node74 = (inp[4]) ? 14'b00000000000000 : node75;
											assign node75 = (inp[0]) ? node81 : node76;
												assign node76 = (inp[5]) ? node78 : 14'b00000000000000;
													assign node78 = (inp[2]) ? 14'b00000000000000 : 14'b00000000000000;
												assign node81 = (inp[6]) ? 14'b00000000000000 : node82;
													assign node82 = (inp[5]) ? 14'b00000000000000 : 14'b00100000000011;
						assign node89 = (inp[6]) ? node113 : node90;
							assign node90 = (inp[1]) ? node92 : 14'b00000000000000;
								assign node92 = (inp[2]) ? 14'b00000000000000 : node93;
									assign node93 = (inp[0]) ? node103 : node94;
										assign node94 = (inp[3]) ? node98 : node95;
											assign node95 = (inp[9]) ? 14'b00000000000000 : 14'b00100000000011;
											assign node98 = (inp[7]) ? 14'b00000000000000 : node99;
												assign node99 = (inp[9]) ? 14'b00001000000101 : 14'b00001000000000;
										assign node103 = (inp[9]) ? 14'b00000000000000 : node104;
											assign node104 = (inp[3]) ? 14'b00000000000000 : node105;
												assign node105 = (inp[4]) ? 14'b00000000000000 : node106;
													assign node106 = (inp[5]) ? 14'b00000000000000 : 14'b00000000011100;
							assign node113 = (inp[1]) ? node119 : node114;
								assign node114 = (inp[9]) ? node116 : 14'b00000000000000;
									assign node116 = (inp[3]) ? 14'b11110111110010 : 14'b00000000000000;
								assign node119 = (inp[5]) ? node121 : 14'b00000000000000;
									assign node121 = (inp[7]) ? node123 : 14'b00000000000000;
										assign node123 = (inp[9]) ? 14'b00000000000000 : node124;
											assign node124 = (inp[3]) ? 14'b00000000000000 : node125;
												assign node125 = (inp[0]) ? 14'b00000000000000 : node126;
													assign node126 = (inp[2]) ? 14'b00000000000000 : 14'b10100100111111;
				assign node132 = (inp[12]) ? node206 : node133;
					assign node133 = (inp[1]) ? node135 : 14'b00000000000000;
						assign node135 = (inp[9]) ? node175 : node136;
							assign node136 = (inp[3]) ? node160 : node137;
								assign node137 = (inp[8]) ? node147 : node138;
									assign node138 = (inp[4]) ? 14'b00000000000000 : node139;
										assign node139 = (inp[6]) ? 14'b00000000000000 : node140;
											assign node140 = (inp[2]) ? node142 : 14'b00000000000000;
												assign node142 = (inp[0]) ? 14'b00100000000011 : 14'b00000000000000;
									assign node147 = (inp[6]) ? node149 : 14'b01001000000100;
										assign node149 = (inp[5]) ? node153 : node150;
											assign node150 = (inp[7]) ? 14'b00000000000000 : 14'b11000000000100;
											assign node153 = (inp[7]) ? node155 : 14'b00000000000000;
												assign node155 = (inp[2]) ? 14'b00000000000000 : node156;
													assign node156 = (inp[0]) ? 14'b00000000000000 : 14'b11000000000100;
								assign node160 = (inp[6]) ? 14'b00000000000000 : node161;
									assign node161 = (inp[2]) ? 14'b00000000000000 : node162;
										assign node162 = (inp[0]) ? 14'b00000000000000 : node163;
											assign node163 = (inp[7]) ? node167 : node164;
												assign node164 = (inp[8]) ? 14'b00000100000001 : 14'b00000000000000;
												assign node167 = (inp[8]) ? 14'b00000000000000 : node168;
													assign node168 = (inp[5]) ? 14'b10010000001101 : 14'b00000000000000;
							assign node175 = (inp[7]) ? node187 : node176;
								assign node176 = (inp[3]) ? node178 : 14'b00000000000000;
									assign node178 = (inp[0]) ? 14'b00000000000000 : node179;
										assign node179 = (inp[8]) ? node181 : 14'b00000000000000;
											assign node181 = (inp[6]) ? 14'b00000000000000 : node182;
												assign node182 = (inp[2]) ? 14'b00000000000000 : 14'b00000100000001;
								assign node187 = (inp[6]) ? node195 : node188;
									assign node188 = (inp[0]) ? 14'b00000000000000 : node189;
										assign node189 = (inp[2]) ? 14'b00000000000000 : node190;
											assign node190 = (inp[8]) ? 14'b00000000000000 : 14'b10010000001101;
									assign node195 = (inp[5]) ? 14'b00000000000000 : node196;
										assign node196 = (inp[3]) ? node198 : 14'b00000000000000;
											assign node198 = (inp[8]) ? 14'b01100000001010 : node199;
												assign node199 = (inp[0]) ? 14'b01001000000100 : node200;
													assign node200 = (inp[2]) ? 14'b01001000000100 : 14'b10100000101010;
					assign node206 = (inp[9]) ? node242 : node207;
						assign node207 = (inp[1]) ? node215 : node208;
							assign node208 = (inp[3]) ? node210 : 14'b00000000000000;
								assign node210 = (inp[6]) ? node212 : 14'b00000000000000;
									assign node212 = (inp[8]) ? 14'b00000000000000 : 14'b01100000001010;
							assign node215 = (inp[3]) ? node229 : node216;
								assign node216 = (inp[6]) ? node220 : node217;
									assign node217 = (inp[8]) ? 14'b00100100011111 : 14'b10000100011000;
									assign node220 = (inp[8]) ? 14'b01000100000100 : node221;
										assign node221 = (inp[5]) ? node223 : 14'b00000000000000;
											assign node223 = (inp[0]) ? 14'b00000000000000 : node224;
												assign node224 = (inp[2]) ? 14'b00000000000000 : 14'b10100000001000;
								assign node229 = (inp[2]) ? 14'b00000000000000 : node230;
									assign node230 = (inp[8]) ? 14'b00000000000000 : node231;
										assign node231 = (inp[0]) ? 14'b00000000000000 : node232;
											assign node232 = (inp[7]) ? node234 : 14'b00000000000000;
												assign node234 = (inp[6]) ? 14'b00000000000000 : node235;
													assign node235 = (inp[5]) ? 14'b01001000000100 : 14'b01001000000101;
						assign node242 = (inp[3]) ? node256 : node243;
							assign node243 = (inp[1]) ? node245 : 14'b00000000000000;
								assign node245 = (inp[8]) ? 14'b00000000000000 : node246;
									assign node246 = (inp[0]) ? 14'b00000000000000 : node247;
										assign node247 = (inp[2]) ? 14'b00000000000000 : node248;
											assign node248 = (inp[7]) ? node250 : 14'b00000000000000;
												assign node250 = (inp[6]) ? 14'b00000000000000 : 14'b01001000000100;
							assign node256 = (inp[6]) ? node274 : node257;
								assign node257 = (inp[1]) ? node259 : 14'b00000000000000;
									assign node259 = (inp[0]) ? 14'b00000000000000 : node260;
										assign node260 = (inp[8]) ? node266 : node261;
											assign node261 = (inp[7]) ? node263 : 14'b00000000000000;
												assign node263 = (inp[2]) ? 14'b00000000000000 : 14'b01001000000100;
											assign node266 = (inp[7]) ? 14'b00000000000000 : node267;
												assign node267 = (inp[5]) ? node269 : 14'b00000000000000;
													assign node269 = (inp[2]) ? 14'b00000000000000 : 14'b10000000101000;
								assign node274 = (inp[8]) ? node282 : node275;
									assign node275 = (inp[5]) ? node277 : 14'b00000000000000;
										assign node277 = (inp[1]) ? node279 : 14'b00000000000000;
											assign node279 = (inp[7]) ? 14'b00000000000000 : 14'b01001000001100;
									assign node282 = (inp[1]) ? node284 : 14'b10100010001100;
										assign node284 = (inp[5]) ? node286 : 14'b00000000000000;
											assign node286 = (inp[7]) ? 14'b10000000011010 : 14'b00000000000000;
			assign node289 = (inp[12]) ? node421 : node290;
				assign node290 = (inp[1]) ? node314 : node291;
					assign node291 = (inp[6]) ? node293 : 14'b00000000000000;
						assign node293 = (inp[3]) ? node295 : 14'b00000000000000;
							assign node295 = (inp[11]) ? node303 : node296;
								assign node296 = (inp[7]) ? 14'b00000000000000 : node297;
									assign node297 = (inp[8]) ? 14'b00000000000000 : node298;
										assign node298 = (inp[9]) ? 14'b00000000000000 : 14'b11000000000100;
								assign node303 = (inp[2]) ? 14'b00000000000000 : node304;
									assign node304 = (inp[7]) ? 14'b00000000000000 : node305;
										assign node305 = (inp[9]) ? 14'b00000000000000 : node306;
											assign node306 = (inp[0]) ? 14'b00000000000000 : node307;
												assign node307 = (inp[8]) ? 14'b00100000000011 : 14'b00000000000000;
					assign node314 = (inp[11]) ? node356 : node315;
						assign node315 = (inp[8]) ? node337 : node316;
							assign node316 = (inp[6]) ? node322 : node317;
								assign node317 = (inp[3]) ? 14'b00000000000000 : node318;
									assign node318 = (inp[9]) ? 14'b00000000000000 : 14'b11000000000100;
								assign node322 = (inp[7]) ? node324 : 14'b00000000000000;
									assign node324 = (inp[3]) ? node326 : 14'b00000000000000;
										assign node326 = (inp[9]) ? node328 : 14'b00000000000000;
											assign node328 = (inp[5]) ? 14'b00000000000000 : node329;
												assign node329 = (inp[0]) ? node333 : node330;
													assign node330 = (inp[2]) ? 14'b01100000000110 : 14'b00001000000101;
													assign node333 = (inp[2]) ? 14'b00000000000000 : 14'b01100000000110;
							assign node337 = (inp[0]) ? 14'b00000000000000 : node338;
								assign node338 = (inp[7]) ? node340 : 14'b00000000000000;
									assign node340 = (inp[3]) ? node342 : 14'b00000000000000;
										assign node342 = (inp[6]) ? node348 : node343;
											assign node343 = (inp[5]) ? node345 : 14'b00000000000000;
												assign node345 = (inp[9]) ? 14'b00000000000000 : 14'b10000000111000;
											assign node348 = (inp[9]) ? node350 : 14'b00000000000000;
												assign node350 = (inp[4]) ? node352 : 14'b00000000011100;
													assign node352 = (inp[5]) ? 14'b00000000000000 : 14'b00000000000000;
						assign node356 = (inp[6]) ? node404 : node357;
							assign node357 = (inp[9]) ? node391 : node358;
								assign node358 = (inp[8]) ? node382 : node359;
									assign node359 = (inp[4]) ? node375 : node360;
										assign node360 = (inp[3]) ? node370 : node361;
											assign node361 = (inp[2]) ? node367 : node362;
												assign node362 = (inp[7]) ? node364 : 14'b00000000000000;
													assign node364 = (inp[5]) ? 14'b00000000000000 : 14'b01001000000100;
												assign node367 = (inp[0]) ? 14'b10110101111111 : 14'b00000000000000;
											assign node370 = (inp[2]) ? 14'b00000000000000 : node371;
												assign node371 = (inp[0]) ? 14'b00000000000000 : 14'b10000100111010;
										assign node375 = (inp[3]) ? node377 : 14'b00000000000000;
											assign node377 = (inp[0]) ? 14'b00000000000000 : node378;
												assign node378 = (inp[2]) ? 14'b00000000000000 : 14'b10000100101010;
									assign node382 = (inp[3]) ? node384 : 14'b00000000011100;
										assign node384 = (inp[0]) ? 14'b00000000000000 : node385;
											assign node385 = (inp[2]) ? 14'b00000000000000 : node386;
												assign node386 = (inp[7]) ? 14'b00000000000000 : 14'b00000000011100;
								assign node391 = (inp[0]) ? 14'b00000000000000 : node392;
									assign node392 = (inp[3]) ? node394 : 14'b00000000000000;
										assign node394 = (inp[2]) ? 14'b00000000000000 : node395;
											assign node395 = (inp[8]) ? node399 : node396;
												assign node396 = (inp[4]) ? 14'b10000100101010 : 14'b10000100111010;
												assign node399 = (inp[7]) ? 14'b00000000000000 : 14'b00000000011100;
							assign node404 = (inp[7]) ? node406 : 14'b00000000000000;
								assign node406 = (inp[3]) ? node408 : 14'b00000000000000;
									assign node408 = (inp[9]) ? node410 : 14'b00000000000000;
										assign node410 = (inp[5]) ? node418 : node411;
											assign node411 = (inp[8]) ? 14'b10100010001100 : node412;
												assign node412 = (inp[2]) ? 14'b10000010001100 : node413;
													assign node413 = (inp[0]) ? 14'b10000010001100 : 14'b10000100101000;
											assign node418 = (inp[8]) ? 14'b00000000000000 : 14'b01001000000101;
				assign node421 = (inp[8]) ? node527 : node422;
					assign node422 = (inp[3]) ? node472 : node423;
						assign node423 = (inp[1]) ? node425 : 14'b00000000000000;
							assign node425 = (inp[2]) ? node461 : node426;
								assign node426 = (inp[7]) ? node438 : node427;
									assign node427 = (inp[11]) ? node429 : 14'b00000000000000;
										assign node429 = (inp[5]) ? 14'b00000000000000 : node430;
											assign node430 = (inp[9]) ? 14'b00000000000000 : node431;
												assign node431 = (inp[4]) ? 14'b00000000000000 : node432;
													assign node432 = (inp[6]) ? 14'b00000000000000 : 14'b01001000000101;
									assign node438 = (inp[6]) ? node452 : node439;
										assign node439 = (inp[9]) ? node447 : node440;
											assign node440 = (inp[5]) ? 14'b00000000000000 : node441;
												assign node441 = (inp[4]) ? 14'b00000000000000 : node442;
													assign node442 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001100;
											assign node447 = (inp[0]) ? 14'b00000000000000 : node448;
												assign node448 = (inp[11]) ? 14'b10100010001100 : 14'b11110111110010;
										assign node452 = (inp[5]) ? node454 : 14'b00000000000000;
											assign node454 = (inp[9]) ? 14'b00000000000000 : node455;
												assign node455 = (inp[0]) ? 14'b00000000000000 : node456;
													assign node456 = (inp[11]) ? 14'b00001000000001 : 14'b01001000000101;
								assign node461 = (inp[0]) ? node463 : 14'b00000000000000;
									assign node463 = (inp[4]) ? 14'b00000000000000 : node464;
										assign node464 = (inp[6]) ? 14'b00000000000000 : node465;
											assign node465 = (inp[11]) ? 14'b00000000000000 : node466;
												assign node466 = (inp[9]) ? 14'b00000000000000 : 14'b10000000101100;
						assign node472 = (inp[6]) ? node492 : node473;
							assign node473 = (inp[2]) ? 14'b00000000000000 : node474;
								assign node474 = (inp[1]) ? node476 : 14'b00000000000000;
									assign node476 = (inp[0]) ? 14'b00000000000000 : node477;
										assign node477 = (inp[7]) ? node479 : 14'b00000000000000;
											assign node479 = (inp[11]) ? node485 : node480;
												assign node480 = (inp[9]) ? 14'b11110111110010 : node481;
													assign node481 = (inp[4]) ? 14'b11110111110010 : 14'b00000000000000;
												assign node485 = (inp[9]) ? 14'b10100010001100 : node486;
													assign node486 = (inp[5]) ? 14'b10100010001100 : 14'b10010101111110;
							assign node492 = (inp[7]) ? node520 : node493;
								assign node493 = (inp[5]) ? node505 : node494;
									assign node494 = (inp[9]) ? 14'b00000000000000 : node495;
										assign node495 = (inp[1]) ? 14'b00000000000000 : node496;
											assign node496 = (inp[11]) ? 14'b00100100001101 : node497;
												assign node497 = (inp[2]) ? 14'b00000000000000 : node498;
													assign node498 = (inp[0]) ? 14'b00000000000000 : 14'b00000000011100;
									assign node505 = (inp[9]) ? node515 : node506;
										assign node506 = (inp[1]) ? 14'b00000000000000 : node507;
											assign node507 = (inp[11]) ? 14'b00100100001101 : node508;
												assign node508 = (inp[0]) ? 14'b00000000000000 : node509;
													assign node509 = (inp[2]) ? 14'b00000000000000 : 14'b00000000011100;
										assign node515 = (inp[1]) ? node517 : 14'b00000000000000;
											assign node517 = (inp[11]) ? 14'b00000000011100 : 14'b00000000011101;
								assign node520 = (inp[11]) ? node522 : 14'b00000000000000;
									assign node522 = (inp[1]) ? 14'b00000000000000 : node523;
										assign node523 = (inp[9]) ? 14'b00000000000000 : 14'b00100100001101;
					assign node527 = (inp[11]) ? 14'b01000000010100 : node528;
						assign node528 = (inp[6]) ? node548 : node529;
							assign node529 = (inp[0]) ? 14'b00000000000000 : node530;
								assign node530 = (inp[2]) ? 14'b00000000000000 : node531;
									assign node531 = (inp[1]) ? node533 : 14'b00000000000000;
										assign node533 = (inp[7]) ? node541 : node534;
											assign node534 = (inp[3]) ? node538 : node535;
												assign node535 = (inp[9]) ? 14'b00000000000000 : 14'b00000000011100;
												assign node538 = (inp[4]) ? 14'b10000100101010 : 14'b10000100111010;
											assign node541 = (inp[9]) ? 14'b00000000000000 : node542;
												assign node542 = (inp[3]) ? 14'b00000000000000 : 14'b00000000011100;
							assign node548 = (inp[3]) ? node566 : node549;
								assign node549 = (inp[9]) ? 14'b00000000000000 : node550;
									assign node550 = (inp[1]) ? node552 : 14'b00000000000000;
										assign node552 = (inp[5]) ? node562 : node553;
											assign node553 = (inp[7]) ? node555 : 14'b10010100011100;
												assign node555 = (inp[4]) ? node559 : node556;
													assign node556 = (inp[0]) ? 14'b00000000000000 : 14'b00000000000000;
													assign node559 = (inp[2]) ? 14'b10010010001100 : 14'b00000000000000;
											assign node562 = (inp[7]) ? 14'b11100100010100 : 14'b11100100000100;
								assign node566 = (inp[9]) ? node568 : 14'b00000000000000;
									assign node568 = (inp[1]) ? node570 : 14'b01001000000100;
										assign node570 = (inp[5]) ? node572 : 14'b00000000000000;
											assign node572 = (inp[7]) ? 14'b01001000001001 : 14'b00000000000000;
		assign node576 = (inp[1]) ? node1156 : node577;
			assign node577 = (inp[3]) ? node933 : node578;
				assign node578 = (inp[4]) ? node700 : node579;
					assign node579 = (inp[9]) ? node669 : node580;
						assign node580 = (inp[5]) ? node654 : node581;
							assign node581 = (inp[0]) ? node597 : node582;
								assign node582 = (inp[8]) ? node590 : node583;
									assign node583 = (inp[13]) ? 14'b00000000000000 : node584;
										assign node584 = (inp[12]) ? 14'b00000000000000 : node585;
											assign node585 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node590 = (inp[11]) ? node592 : 14'b00000000000000;
										assign node592 = (inp[13]) ? node594 : 14'b00000000000000;
											assign node594 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node597 = (inp[7]) ? node623 : node598;
									assign node598 = (inp[6]) ? node614 : node599;
										assign node599 = (inp[8]) ? node607 : node600;
											assign node600 = (inp[11]) ? 14'b00000000000000 : node601;
												assign node601 = (inp[13]) ? 14'b00000000000000 : node602;
													assign node602 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node607 = (inp[11]) ? node609 : 14'b00000000000000;
												assign node609 = (inp[12]) ? node611 : 14'b00000000000000;
													assign node611 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
										assign node614 = (inp[8]) ? 14'b00000000000000 : node615;
											assign node615 = (inp[12]) ? 14'b00000000000000 : node616;
												assign node616 = (inp[13]) ? 14'b00000000000000 : node617;
													assign node617 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node623 = (inp[6]) ? node639 : node624;
										assign node624 = (inp[2]) ? node632 : node625;
											assign node625 = (inp[8]) ? 14'b00000000000000 : node626;
												assign node626 = (inp[12]) ? 14'b00000000000000 : node627;
													assign node627 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node632 = (inp[12]) ? node634 : 14'b00000000000000;
												assign node634 = (inp[11]) ? node636 : 14'b00000000000000;
													assign node636 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
										assign node639 = (inp[12]) ? node647 : node640;
											assign node640 = (inp[13]) ? 14'b00000000000000 : node641;
												assign node641 = (inp[11]) ? 14'b00000000000000 : node642;
													assign node642 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node647 = (inp[11]) ? node649 : 14'b00000000000000;
												assign node649 = (inp[8]) ? node651 : 14'b00000000000000;
													assign node651 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node654 = (inp[13]) ? node662 : node655;
								assign node655 = (inp[11]) ? 14'b00000000000000 : node656;
									assign node656 = (inp[12]) ? 14'b00000000000000 : node657;
										assign node657 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node662 = (inp[8]) ? node664 : 14'b00000000000000;
									assign node664 = (inp[12]) ? node666 : 14'b00000000000000;
										assign node666 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
						assign node669 = (inp[6]) ? node685 : node670;
							assign node670 = (inp[8]) ? node678 : node671;
								assign node671 = (inp[12]) ? 14'b00000000000000 : node672;
									assign node672 = (inp[13]) ? 14'b00000000000000 : node673;
										assign node673 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node678 = (inp[12]) ? node680 : 14'b00000000000000;
									assign node680 = (inp[13]) ? node682 : 14'b00000000000000;
										assign node682 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node685 = (inp[12]) ? node693 : node686;
								assign node686 = (inp[13]) ? 14'b00000000000000 : node687;
									assign node687 = (inp[11]) ? 14'b00000000000000 : node688;
										assign node688 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node693 = (inp[8]) ? node695 : 14'b00000000000000;
									assign node695 = (inp[11]) ? node697 : 14'b00000000000000;
										assign node697 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
					assign node700 = (inp[2]) ? node806 : node701;
						assign node701 = (inp[5]) ? node759 : node702;
							assign node702 = (inp[7]) ? node734 : node703;
								assign node703 = (inp[0]) ? node719 : node704;
									assign node704 = (inp[11]) ? node712 : node705;
										assign node705 = (inp[8]) ? 14'b00000000000000 : node706;
											assign node706 = (inp[12]) ? 14'b00000000000000 : node707;
												assign node707 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node712 = (inp[8]) ? node714 : 14'b00000000000000;
											assign node714 = (inp[12]) ? node716 : 14'b00000000000000;
												assign node716 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node719 = (inp[13]) ? node727 : node720;
										assign node720 = (inp[12]) ? 14'b00000000000000 : node721;
											assign node721 = (inp[8]) ? 14'b00000000000000 : node722;
												assign node722 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node727 = (inp[12]) ? node729 : 14'b00000000000000;
											assign node729 = (inp[11]) ? node731 : 14'b00000000000000;
												assign node731 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node734 = (inp[6]) ? node736 : 14'b00000000000000;
									assign node736 = (inp[0]) ? node746 : node737;
										assign node737 = (inp[11]) ? 14'b00000000000000 : node738;
											assign node738 = (inp[13]) ? 14'b00000000000000 : node739;
												assign node739 = (inp[12]) ? 14'b00000000000000 : node740;
													assign node740 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node746 = (inp[12]) ? node752 : node747;
											assign node747 = (inp[11]) ? 14'b00000000000000 : node748;
												assign node748 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node752 = (inp[8]) ? node754 : 14'b00000000000000;
												assign node754 = (inp[13]) ? node756 : 14'b00000000000000;
													assign node756 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node759 = (inp[7]) ? node775 : node760;
								assign node760 = (inp[12]) ? node768 : node761;
									assign node761 = (inp[11]) ? 14'b00000000000000 : node762;
										assign node762 = (inp[8]) ? 14'b00000000000000 : node763;
											assign node763 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node768 = (inp[13]) ? node770 : 14'b00000000000000;
										assign node770 = (inp[11]) ? node772 : 14'b00000000000000;
											assign node772 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node775 = (inp[0]) ? node791 : node776;
									assign node776 = (inp[13]) ? node784 : node777;
										assign node777 = (inp[12]) ? 14'b00000000000000 : node778;
											assign node778 = (inp[8]) ? 14'b00000000000000 : node779;
												assign node779 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node784 = (inp[11]) ? node786 : 14'b00000000000000;
											assign node786 = (inp[12]) ? node788 : 14'b00000000000000;
												assign node788 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node791 = (inp[11]) ? node799 : node792;
										assign node792 = (inp[8]) ? 14'b00000000000000 : node793;
											assign node793 = (inp[13]) ? 14'b00000000000000 : node794;
												assign node794 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node799 = (inp[8]) ? node801 : 14'b00000000000000;
											assign node801 = (inp[13]) ? node803 : 14'b00000000000000;
												assign node803 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
						assign node806 = (inp[5]) ? node854 : node807;
							assign node807 = (inp[7]) ? node839 : node808;
								assign node808 = (inp[0]) ? node824 : node809;
									assign node809 = (inp[12]) ? node817 : node810;
										assign node810 = (inp[13]) ? 14'b00000000000000 : node811;
											assign node811 = (inp[8]) ? 14'b00000000000000 : node812;
												assign node812 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node817 = (inp[13]) ? node819 : 14'b00000000000000;
											assign node819 = (inp[8]) ? node821 : 14'b00000000000000;
												assign node821 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node824 = (inp[11]) ? node832 : node825;
										assign node825 = (inp[8]) ? 14'b00000000000000 : node826;
											assign node826 = (inp[13]) ? 14'b00000000000000 : node827;
												assign node827 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node832 = (inp[12]) ? node834 : 14'b00000000000000;
											assign node834 = (inp[13]) ? node836 : 14'b00000000000000;
												assign node836 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node839 = (inp[11]) ? node847 : node840;
									assign node840 = (inp[13]) ? 14'b00000000000000 : node841;
										assign node841 = (inp[12]) ? 14'b00000000000000 : node842;
											assign node842 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node847 = (inp[13]) ? node849 : 14'b00000000000000;
										assign node849 = (inp[12]) ? node851 : 14'b00000000000000;
											assign node851 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node854 = (inp[7]) ? node886 : node855;
								assign node855 = (inp[6]) ? node871 : node856;
									assign node856 = (inp[8]) ? node864 : node857;
										assign node857 = (inp[11]) ? 14'b00000000000000 : node858;
											assign node858 = (inp[13]) ? 14'b00000000000000 : node859;
												assign node859 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node864 = (inp[13]) ? node866 : 14'b00000000000000;
											assign node866 = (inp[12]) ? node868 : 14'b00000000000000;
												assign node868 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node871 = (inp[12]) ? node879 : node872;
										assign node872 = (inp[11]) ? 14'b00000000000000 : node873;
											assign node873 = (inp[8]) ? 14'b00000000000000 : node874;
												assign node874 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node879 = (inp[11]) ? node881 : 14'b00000000000000;
											assign node881 = (inp[13]) ? node883 : 14'b00000000000000;
												assign node883 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node886 = (inp[0]) ? node902 : node887;
									assign node887 = (inp[13]) ? node895 : node888;
										assign node888 = (inp[11]) ? 14'b00000000000000 : node889;
											assign node889 = (inp[12]) ? 14'b00000000000000 : node890;
												assign node890 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node895 = (inp[11]) ? node897 : 14'b00000000000000;
											assign node897 = (inp[8]) ? node899 : 14'b00000000000000;
												assign node899 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node902 = (inp[6]) ? node918 : node903;
										assign node903 = (inp[13]) ? node911 : node904;
											assign node904 = (inp[11]) ? 14'b00000000000000 : node905;
												assign node905 = (inp[8]) ? 14'b00000000000000 : node906;
													assign node906 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node911 = (inp[11]) ? node913 : 14'b00000000000000;
												assign node913 = (inp[12]) ? node915 : 14'b00000000000000;
													assign node915 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
										assign node918 = (inp[13]) ? node926 : node919;
											assign node919 = (inp[11]) ? 14'b00000000000000 : node920;
												assign node920 = (inp[8]) ? 14'b00000000000000 : node921;
													assign node921 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node926 = (inp[12]) ? node928 : 14'b00000000000000;
												assign node928 = (inp[8]) ? node930 : 14'b00000000000000;
													assign node930 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
				assign node933 = (inp[6]) ? node1091 : node934;
					assign node934 = (inp[4]) ? node1076 : node935;
						assign node935 = (inp[5]) ? node1027 : node936;
							assign node936 = (inp[9]) ? node980 : node937;
								assign node937 = (inp[7]) ? node965 : node938;
									assign node938 = (inp[0]) ? node948 : node939;
										assign node939 = (inp[2]) ? node941 : 14'b00000000000000;
											assign node941 = (inp[8]) ? 14'b00000000000000 : node942;
												assign node942 = (inp[13]) ? 14'b00000000000000 : node943;
													assign node943 = (inp[11]) ? 14'b00000000000000 : 14'b00000000000000;
										assign node948 = (inp[2]) ? node958 : node949;
											assign node949 = (inp[13]) ? node953 : node950;
												assign node950 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
												assign node953 = (inp[12]) ? node955 : 14'b00000000000000;
													assign node955 = (inp[11]) ? 14'b00000000000000 : 14'b00000000000000;
											assign node958 = (inp[13]) ? node960 : 14'b00000000000000;
												assign node960 = (inp[11]) ? node962 : 14'b00000000000000;
													assign node962 = (inp[8]) ? 14'b00000000000000 : 14'b00000000000000;
									assign node965 = (inp[12]) ? node973 : node966;
										assign node966 = (inp[8]) ? 14'b00000000000000 : node967;
											assign node967 = (inp[11]) ? 14'b00000000000000 : node968;
												assign node968 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node973 = (inp[8]) ? node975 : 14'b00000000000000;
											assign node975 = (inp[13]) ? node977 : 14'b00000000000000;
												assign node977 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node980 = (inp[2]) ? node996 : node981;
									assign node981 = (inp[13]) ? node989 : node982;
										assign node982 = (inp[11]) ? 14'b00000000000000 : node983;
											assign node983 = (inp[8]) ? 14'b00000000000000 : node984;
												assign node984 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node989 = (inp[12]) ? node991 : 14'b00000000000000;
											assign node991 = (inp[8]) ? node993 : 14'b00000000000000;
												assign node993 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node996 = (inp[7]) ? node1012 : node997;
										assign node997 = (inp[12]) ? node1005 : node998;
											assign node998 = (inp[8]) ? 14'b00000000000000 : node999;
												assign node999 = (inp[11]) ? 14'b00000000000000 : node1000;
													assign node1000 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node1005 = (inp[13]) ? node1007 : 14'b00000000000000;
												assign node1007 = (inp[8]) ? node1009 : 14'b00000000000000;
													assign node1009 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
										assign node1012 = (inp[12]) ? node1020 : node1013;
											assign node1013 = (inp[8]) ? 14'b00000000000000 : node1014;
												assign node1014 = (inp[11]) ? 14'b00000000000000 : node1015;
													assign node1015 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node1020 = (inp[11]) ? node1022 : 14'b00000000000000;
												assign node1022 = (inp[8]) ? node1024 : 14'b00000000000000;
													assign node1024 = (inp[0]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node1027 = (inp[7]) ? node1043 : node1028;
								assign node1028 = (inp[12]) ? node1036 : node1029;
									assign node1029 = (inp[8]) ? 14'b00000000000000 : node1030;
										assign node1030 = (inp[13]) ? 14'b00000000000000 : node1031;
											assign node1031 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node1036 = (inp[8]) ? node1038 : 14'b00000000000000;
										assign node1038 = (inp[13]) ? node1040 : 14'b00000000000000;
											assign node1040 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node1043 = (inp[0]) ? node1059 : node1044;
									assign node1044 = (inp[13]) ? node1052 : node1045;
										assign node1045 = (inp[11]) ? 14'b00000000000000 : node1046;
											assign node1046 = (inp[8]) ? 14'b00000000000000 : node1047;
												assign node1047 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node1052 = (inp[12]) ? node1054 : 14'b00000000000000;
											assign node1054 = (inp[8]) ? node1056 : 14'b00000000000000;
												assign node1056 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node1059 = (inp[9]) ? 14'b00000000000000 : node1060;
										assign node1060 = (inp[8]) ? node1068 : node1061;
											assign node1061 = (inp[11]) ? 14'b00000000000000 : node1062;
												assign node1062 = (inp[2]) ? 14'b00000000000000 : node1063;
													assign node1063 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node1068 = (inp[13]) ? node1070 : 14'b00000000000000;
												assign node1070 = (inp[12]) ? node1072 : 14'b00000000000000;
													assign node1072 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
						assign node1076 = (inp[13]) ? node1084 : node1077;
							assign node1077 = (inp[11]) ? 14'b00000000000000 : node1078;
								assign node1078 = (inp[8]) ? 14'b00000000000000 : node1079;
									assign node1079 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
							assign node1084 = (inp[8]) ? node1086 : 14'b00000000000000;
								assign node1086 = (inp[12]) ? node1088 : 14'b00000000000000;
									assign node1088 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
					assign node1091 = (inp[12]) ? node1113 : node1092;
						assign node1092 = (inp[13]) ? node1098 : node1093;
							assign node1093 = (inp[11]) ? 14'b00000000000000 : node1094;
								assign node1094 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
							assign node1098 = (inp[0]) ? 14'b00000000000000 : node1099;
								assign node1099 = (inp[8]) ? node1101 : 14'b00000000000000;
									assign node1101 = (inp[11]) ? node1103 : 14'b00000000000000;
										assign node1103 = (inp[9]) ? 14'b00000000000000 : node1104;
											assign node1104 = (inp[2]) ? 14'b00000000000000 : node1105;
												assign node1105 = (inp[7]) ? 14'b00000000000000 : node1106;
													assign node1106 = (inp[4]) ? 14'b10000100101010 : 14'b10000100111010;
						assign node1113 = (inp[13]) ? node1135 : node1114;
							assign node1114 = (inp[11]) ? node1130 : node1115;
								assign node1115 = (inp[9]) ? node1127 : node1116;
									assign node1116 = (inp[0]) ? 14'b00000000000000 : node1117;
										assign node1117 = (inp[7]) ? 14'b00000000000000 : node1118;
											assign node1118 = (inp[2]) ? 14'b00000000000000 : node1119;
												assign node1119 = (inp[8]) ? 14'b00000000000000 : node1120;
													assign node1120 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
									assign node1127 = (inp[8]) ? 14'b01100000001010 : 14'b00000000000000;
								assign node1130 = (inp[8]) ? 14'b00000000000000 : node1131;
									assign node1131 = (inp[9]) ? 14'b00000000000000 : 14'b01001000000101;
							assign node1135 = (inp[11]) ? node1151 : node1136;
								assign node1136 = (inp[9]) ? node1148 : node1137;
									assign node1137 = (inp[2]) ? 14'b00000000000000 : node1138;
										assign node1138 = (inp[7]) ? 14'b00000000000000 : node1139;
											assign node1139 = (inp[8]) ? 14'b00000000000000 : node1140;
												assign node1140 = (inp[0]) ? 14'b00000000000000 : node1141;
													assign node1141 = (inp[4]) ? 14'b10000000101000 : 14'b10000000111000;
									assign node1148 = (inp[8]) ? 14'b00100100001101 : 14'b00000000000000;
								assign node1151 = (inp[8]) ? 14'b10000100001000 : node1152;
									assign node1152 = (inp[9]) ? 14'b00000000000000 : 14'b10010101111110;
			assign node1156 = (inp[13]) ? node1426 : node1157;
				assign node1157 = (inp[12]) ? node1269 : node1158;
					assign node1158 = (inp[11]) ? node1198 : node1159;
						assign node1159 = (inp[8]) ? node1161 : 14'b10000100001000;
							assign node1161 = (inp[9]) ? node1187 : node1162;
								assign node1162 = (inp[6]) ? 14'b00000000000000 : node1163;
									assign node1163 = (inp[3]) ? node1179 : node1164;
										assign node1164 = (inp[2]) ? node1172 : node1165;
											assign node1165 = (inp[0]) ? node1167 : 14'b00100000000011;
												assign node1167 = (inp[7]) ? 14'b00100000000011 : node1168;
													assign node1168 = (inp[4]) ? 14'b00000000000000 : 14'b00000000000000;
											assign node1172 = (inp[0]) ? node1176 : node1173;
												assign node1173 = (inp[4]) ? 14'b00100000000011 : 14'b00000000000000;
												assign node1176 = (inp[4]) ? 14'b00000000000000 : 14'b00100000000011;
										assign node1179 = (inp[7]) ? node1181 : 14'b00000000000000;
											assign node1181 = (inp[5]) ? node1183 : 14'b00000000000000;
												assign node1183 = (inp[2]) ? 14'b00000000000000 : 14'b00000000011100;
								assign node1187 = (inp[3]) ? node1189 : 14'b00000000000000;
									assign node1189 = (inp[6]) ? node1191 : 14'b00000000000000;
										assign node1191 = (inp[7]) ? node1193 : 14'b00000000000000;
											assign node1193 = (inp[5]) ? 14'b10100000001000 : node1194;
												assign node1194 = (inp[0]) ? 14'b00000000000000 : 14'b00100000001010;
						assign node1198 = (inp[6]) ? node1250 : node1199;
							assign node1199 = (inp[9]) ? node1239 : node1200;
								assign node1200 = (inp[3]) ? node1226 : node1201;
									assign node1201 = (inp[8]) ? node1211 : node1202;
										assign node1202 = (inp[0]) ? node1204 : 14'b00000000000000;
											assign node1204 = (inp[4]) ? 14'b00000000000000 : node1205;
												assign node1205 = (inp[2]) ? 14'b01001000000101 : node1206;
													assign node1206 = (inp[7]) ? 14'b01100000001010 : 14'b00000000000000;
										assign node1211 = (inp[0]) ? node1219 : node1212;
											assign node1212 = (inp[4]) ? node1216 : node1213;
												assign node1213 = (inp[2]) ? 14'b00000000000000 : 14'b10000001001101;
												assign node1216 = (inp[2]) ? 14'b10000100001101 : 14'b10000010001101;
											assign node1219 = (inp[2]) ? node1223 : node1220;
												assign node1220 = (inp[4]) ? 14'b10000000011101 : 14'b00000000000000;
												assign node1223 = (inp[4]) ? 14'b00000000000000 : 14'b10010000001101;
									assign node1226 = (inp[2]) ? 14'b00000000000000 : node1227;
										assign node1227 = (inp[0]) ? 14'b00000000000000 : node1228;
											assign node1228 = (inp[7]) ? node1232 : node1229;
												assign node1229 = (inp[8]) ? 14'b00100000001010 : 14'b00100000000011;
												assign node1232 = (inp[5]) ? node1234 : 14'b00000000000000;
													assign node1234 = (inp[8]) ? 14'b00000000000000 : 14'b00100000000011;
								assign node1239 = (inp[2]) ? 14'b00000000000000 : node1240;
									assign node1240 = (inp[0]) ? 14'b00000000000000 : node1241;
										assign node1241 = (inp[7]) ? 14'b00000000000000 : node1242;
											assign node1242 = (inp[3]) ? node1244 : 14'b00000000000000;
												assign node1244 = (inp[8]) ? 14'b00100000001010 : 14'b00100000000011;
							assign node1250 = (inp[7]) ? node1252 : 14'b00000000000000;
								assign node1252 = (inp[3]) ? node1254 : 14'b00000000000000;
									assign node1254 = (inp[9]) ? node1256 : 14'b00000000000000;
										assign node1256 = (inp[5]) ? node1264 : node1257;
											assign node1257 = (inp[8]) ? 14'b01001000000100 : node1258;
												assign node1258 = (inp[0]) ? 14'b00000100001111 : node1259;
													assign node1259 = (inp[2]) ? 14'b00000100001111 : 14'b00100000000011;
											assign node1264 = (inp[0]) ? node1266 : 14'b00000000000000;
												assign node1266 = (inp[8]) ? 14'b00000000000000 : 14'b00100000000011;
					assign node1269 = (inp[2]) ? node1381 : node1270;
						assign node1270 = (inp[0]) ? node1330 : node1271;
							assign node1271 = (inp[6]) ? node1297 : node1272;
								assign node1272 = (inp[8]) ? node1282 : node1273;
									assign node1273 = (inp[11]) ? node1275 : 14'b00000000000000;
										assign node1275 = (inp[7]) ? node1277 : 14'b00000000000000;
											assign node1277 = (inp[3]) ? 14'b00100100001101 : node1278;
												assign node1278 = (inp[9]) ? 14'b00100100001101 : 14'b00000000000000;
									assign node1282 = (inp[11]) ? 14'b00000000000000 : node1283;
										assign node1283 = (inp[9]) ? node1291 : node1284;
											assign node1284 = (inp[3]) ? node1288 : node1285;
												assign node1285 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
												assign node1288 = (inp[7]) ? 14'b00000000000000 : 14'b00000000011100;
											assign node1291 = (inp[3]) ? node1293 : 14'b00000000000000;
												assign node1293 = (inp[7]) ? 14'b00000000000000 : 14'b00000000011100;
								assign node1297 = (inp[5]) ? node1299 : 14'b00000000000000;
									assign node1299 = (inp[8]) ? node1321 : node1300;
										assign node1300 = (inp[11]) ? node1312 : node1301;
											assign node1301 = (inp[7]) ? node1307 : node1302;
												assign node1302 = (inp[9]) ? node1304 : 14'b00000000000000;
													assign node1304 = (inp[3]) ? 14'b00001000001100 : 14'b00000000000000;
												assign node1307 = (inp[3]) ? 14'b00000000000000 : node1308;
													assign node1308 = (inp[9]) ? 14'b00000000000000 : 14'b00000100001101;
											assign node1312 = (inp[9]) ? node1318 : node1313;
												assign node1313 = (inp[7]) ? node1315 : 14'b00000000000000;
													assign node1315 = (inp[3]) ? 14'b00000000000000 : 14'b01100000000010;
												assign node1318 = (inp[7]) ? 14'b00000000000000 : 14'b00000100001111;
										assign node1321 = (inp[7]) ? node1323 : 14'b00000000000000;
											assign node1323 = (inp[3]) ? node1325 : 14'b00000000000000;
												assign node1325 = (inp[11]) ? 14'b00000000000000 : node1326;
													assign node1326 = (inp[9]) ? 14'b01100000000110 : 14'b00000000000000;
							assign node1330 = (inp[4]) ? node1368 : node1331;
								assign node1331 = (inp[8]) ? node1349 : node1332;
									assign node1332 = (inp[7]) ? 14'b00000000000000 : node1333;
										assign node1333 = (inp[3]) ? node1341 : node1334;
											assign node1334 = (inp[9]) ? 14'b00000000000000 : node1335;
												assign node1335 = (inp[6]) ? 14'b00000000000000 : node1336;
													assign node1336 = (inp[11]) ? 14'b00000000000000 : 14'b01001000000100;
											assign node1341 = (inp[6]) ? node1343 : 14'b00000000000000;
												assign node1343 = (inp[9]) ? node1345 : 14'b00000000000000;
													assign node1345 = (inp[11]) ? 14'b00000100001111 : 14'b00000000000000;
									assign node1349 = (inp[5]) ? node1359 : node1350;
										assign node1350 = (inp[3]) ? 14'b00000000000000 : node1351;
											assign node1351 = (inp[11]) ? 14'b00000000000000 : node1352;
												assign node1352 = (inp[9]) ? 14'b00000000000000 : node1353;
													assign node1353 = (inp[6]) ? 14'b00000000000000 : 14'b10000100011000;
										assign node1359 = (inp[3]) ? node1361 : 14'b00000000000000;
											assign node1361 = (inp[11]) ? 14'b00000000000000 : node1362;
												assign node1362 = (inp[6]) ? node1364 : 14'b00000000000000;
													assign node1364 = (inp[7]) ? 14'b00000000000000 : 14'b00000000000000;
								assign node1368 = (inp[8]) ? 14'b00000000000000 : node1369;
									assign node1369 = (inp[7]) ? 14'b00000000000000 : node1370;
										assign node1370 = (inp[9]) ? node1372 : 14'b00000000000000;
											assign node1372 = (inp[6]) ? node1374 : 14'b00000000000000;
												assign node1374 = (inp[11]) ? 14'b00000000000000 : node1375;
													assign node1375 = (inp[3]) ? 14'b00000000000000 : 14'b00000000000000;
						assign node1381 = (inp[5]) ? node1397 : node1382;
							assign node1382 = (inp[9]) ? 14'b00000000000000 : node1383;
								assign node1383 = (inp[3]) ? 14'b00000000000000 : node1384;
									assign node1384 = (inp[0]) ? node1386 : 14'b00000000000000;
										assign node1386 = (inp[6]) ? 14'b00000000000000 : node1387;
											assign node1387 = (inp[8]) ? 14'b00000000000000 : node1388;
												assign node1388 = (inp[4]) ? 14'b00000000000000 : node1389;
													assign node1389 = (inp[11]) ? 14'b00000000000000 : 14'b01001000000100;
							assign node1397 = (inp[9]) ? node1411 : node1398;
								assign node1398 = (inp[4]) ? 14'b00000000000000 : node1399;
									assign node1399 = (inp[6]) ? 14'b00000000000000 : node1400;
										assign node1400 = (inp[11]) ? 14'b00000000000000 : node1401;
											assign node1401 = (inp[3]) ? 14'b00000000000000 : node1402;
												assign node1402 = (inp[0]) ? node1404 : 14'b00000000000000;
													assign node1404 = (inp[8]) ? 14'b00000000000000 : 14'b01001000000100;
								assign node1411 = (inp[6]) ? node1413 : 14'b00000000000000;
									assign node1413 = (inp[3]) ? node1415 : 14'b00000000000000;
										assign node1415 = (inp[7]) ? node1421 : node1416;
											assign node1416 = (inp[8]) ? 14'b00000000000000 : node1417;
												assign node1417 = (inp[11]) ? 14'b00000100001111 : 14'b00001000001100;
											assign node1421 = (inp[11]) ? 14'b00000000000000 : node1422;
												assign node1422 = (inp[8]) ? 14'b01100000000110 : 14'b00000000000000;
				assign node1426 = (inp[8]) ? node1562 : node1427;
					assign node1427 = (inp[3]) ? node1489 : node1428;
						assign node1428 = (inp[9]) ? node1466 : node1429;
							assign node1429 = (inp[6]) ? node1451 : node1430;
								assign node1430 = (inp[12]) ? node1440 : node1431;
									assign node1431 = (inp[4]) ? 14'b00000000000000 : node1432;
										assign node1432 = (inp[11]) ? node1434 : 14'b00000000000000;
											assign node1434 = (inp[0]) ? node1436 : 14'b00000000000000;
												assign node1436 = (inp[2]) ? 14'b00000000011100 : 14'b00000000000000;
									assign node1440 = (inp[11]) ? node1442 : 14'b00000000011101;
										assign node1442 = (inp[4]) ? 14'b00000000000000 : node1443;
											assign node1443 = (inp[2]) ? 14'b00000000000000 : node1444;
												assign node1444 = (inp[5]) ? 14'b00000000000000 : node1445;
													assign node1445 = (inp[0]) ? 14'b10000000001111 : 14'b00000000000000;
								assign node1451 = (inp[2]) ? 14'b00000000000000 : node1452;
									assign node1452 = (inp[5]) ? node1454 : 14'b00000000000000;
										assign node1454 = (inp[7]) ? node1456 : 14'b00000000000000;
											assign node1456 = (inp[12]) ? node1458 : 14'b00000000000000;
												assign node1458 = (inp[11]) ? node1462 : node1459;
													assign node1459 = (inp[0]) ? 14'b00000000000000 : 14'b00000000011100;
													assign node1462 = (inp[0]) ? 14'b00000000000000 : 14'b01001000000101;
							assign node1466 = (inp[12]) ? node1478 : node1467;
								assign node1467 = (inp[2]) ? 14'b00000000000000 : node1468;
									assign node1468 = (inp[7]) ? node1470 : 14'b00000000000000;
										assign node1470 = (inp[11]) ? 14'b00000000000000 : node1471;
											assign node1471 = (inp[0]) ? 14'b00000000000000 : node1472;
												assign node1472 = (inp[6]) ? 14'b00000000000000 : 14'b00001000000100;
								assign node1478 = (inp[6]) ? 14'b00000000000000 : node1479;
									assign node1479 = (inp[0]) ? 14'b00000000000000 : node1480;
										assign node1480 = (inp[7]) ? node1482 : 14'b00000000000000;
											assign node1482 = (inp[11]) ? 14'b00000000000000 : node1483;
												assign node1483 = (inp[2]) ? 14'b00000000000000 : 14'b01100000001010;
						assign node1489 = (inp[9]) ? node1513 : node1490;
							assign node1490 = (inp[6]) ? 14'b00000000000000 : node1491;
								assign node1491 = (inp[0]) ? 14'b00000000000000 : node1492;
									assign node1492 = (inp[2]) ? 14'b00000000000000 : node1493;
										assign node1493 = (inp[11]) ? node1503 : node1494;
											assign node1494 = (inp[12]) ? node1500 : node1495;
												assign node1495 = (inp[5]) ? node1497 : 14'b00000000000000;
													assign node1497 = (inp[7]) ? 14'b00001000000100 : 14'b00000000000000;
												assign node1500 = (inp[7]) ? 14'b01100000001010 : 14'b00000000000000;
											assign node1503 = (inp[12]) ? 14'b00000000000000 : node1504;
												assign node1504 = (inp[5]) ? 14'b00100000000011 : node1505;
													assign node1505 = (inp[7]) ? 14'b00000000000000 : 14'b00100000000011;
							assign node1513 = (inp[6]) ? node1531 : node1514;
								assign node1514 = (inp[0]) ? 14'b00000000000000 : node1515;
									assign node1515 = (inp[2]) ? 14'b00000000000000 : node1516;
										assign node1516 = (inp[12]) ? node1524 : node1517;
											assign node1517 = (inp[11]) ? node1521 : node1518;
												assign node1518 = (inp[7]) ? 14'b00001000000100 : 14'b00000000000000;
												assign node1521 = (inp[7]) ? 14'b00000000000000 : 14'b00100000000011;
											assign node1524 = (inp[7]) ? node1526 : 14'b00000000000000;
												assign node1526 = (inp[11]) ? 14'b00000000000000 : 14'b01100000001010;
								assign node1531 = (inp[5]) ? node1549 : node1532;
									assign node1532 = (inp[7]) ? node1534 : 14'b00000000000000;
										assign node1534 = (inp[11]) ? node1542 : node1535;
											assign node1535 = (inp[0]) ? 14'b00000000000000 : node1536;
												assign node1536 = (inp[12]) ? 14'b00000000000000 : node1537;
													assign node1537 = (inp[2]) ? 14'b00000000000000 : 14'b00000000011101;
											assign node1542 = (inp[12]) ? 14'b00000000000000 : node1543;
												assign node1543 = (inp[0]) ? 14'b01000100000010 : node1544;
													assign node1544 = (inp[4]) ? 14'b01000100000010 : 14'b00001000001001;
									assign node1549 = (inp[11]) ? node1555 : node1550;
										assign node1550 = (inp[7]) ? 14'b00000000000000 : node1551;
											assign node1551 = (inp[12]) ? 14'b10100000001000 : 14'b00000000000000;
										assign node1555 = (inp[7]) ? node1559 : node1556;
											assign node1556 = (inp[12]) ? 14'b10100100001000 : 14'b00000000000000;
											assign node1559 = (inp[12]) ? 14'b00000000000000 : 14'b10100101111111;
					assign node1562 = (inp[11]) ? node1632 : node1563;
						assign node1563 = (inp[12]) ? node1605 : node1564;
							assign node1564 = (inp[2]) ? node1592 : node1565;
								assign node1565 = (inp[6]) ? node1581 : node1566;
									assign node1566 = (inp[7]) ? node1572 : node1567;
										assign node1567 = (inp[0]) ? 14'b00000000000000 : node1568;
											assign node1568 = (inp[3]) ? 14'b00001000001001 : 14'b00000000000000;
										assign node1572 = (inp[9]) ? 14'b00000000000000 : node1573;
											assign node1573 = (inp[0]) ? node1575 : 14'b00000000000000;
												assign node1575 = (inp[3]) ? 14'b00000000000000 : node1576;
													assign node1576 = (inp[4]) ? 14'b00000000000000 : 14'b10110111101111;
									assign node1581 = (inp[3]) ? node1583 : 14'b00000000000000;
										assign node1583 = (inp[5]) ? 14'b00000000000000 : node1584;
											assign node1584 = (inp[7]) ? node1586 : 14'b00000000000000;
												assign node1586 = (inp[0]) ? 14'b00000000000000 : node1587;
													assign node1587 = (inp[9]) ? 14'b10000100111000 : 14'b00000000000000;
								assign node1592 = (inp[7]) ? node1594 : 14'b00000000000000;
									assign node1594 = (inp[9]) ? node1596 : 14'b00000000000000;
										assign node1596 = (inp[0]) ? 14'b00000000000000 : node1597;
											assign node1597 = (inp[6]) ? node1599 : 14'b00000000000000;
												assign node1599 = (inp[3]) ? node1601 : 14'b00000000000000;
													assign node1601 = (inp[4]) ? 14'b00000000000000 : 14'b00000000000000;
							assign node1605 = (inp[3]) ? node1617 : node1606;
								assign node1606 = (inp[9]) ? 14'b00000000000000 : node1607;
									assign node1607 = (inp[6]) ? 14'b00000100001110 : node1608;
										assign node1608 = (inp[0]) ? 14'b00001000000100 : node1609;
											assign node1609 = (inp[2]) ? 14'b00001000000100 : node1610;
												assign node1610 = (inp[4]) ? 14'b10000000101000 : 14'b10000000111000;
								assign node1617 = (inp[5]) ? node1619 : 14'b00000000000000;
									assign node1619 = (inp[9]) ? node1621 : 14'b00000000000000;
										assign node1621 = (inp[6]) ? node1629 : node1622;
											assign node1622 = (inp[2]) ? 14'b00000000000000 : node1623;
												assign node1623 = (inp[0]) ? 14'b00000000000000 : node1624;
													assign node1624 = (inp[7]) ? 14'b00000000000000 : 14'b00000000011101;
											assign node1629 = (inp[7]) ? 14'b00000000011100 : 14'b00000000000000;
						assign node1632 = (inp[12]) ? 14'b10000100001000 : node1633;
							assign node1633 = (inp[6]) ? node1665 : node1634;
								assign node1634 = (inp[9]) ? node1654 : node1635;
									assign node1635 = (inp[3]) ? node1645 : node1636;
										assign node1636 = (inp[0]) ? 14'b10100100011000 : node1637;
											assign node1637 = (inp[4]) ? node1641 : node1638;
												assign node1638 = (inp[2]) ? 14'b00000000000000 : 14'b10000000001010;
												assign node1641 = (inp[2]) ? 14'b10100100011000 : 14'b10000000001010;
										assign node1645 = (inp[0]) ? 14'b00000000000000 : node1646;
											assign node1646 = (inp[2]) ? 14'b00000000000000 : node1647;
												assign node1647 = (inp[7]) ? 14'b00000000000000 : node1648;
													assign node1648 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
									assign node1654 = (inp[0]) ? 14'b00000000000000 : node1655;
										assign node1655 = (inp[3]) ? node1657 : 14'b00000000000000;
											assign node1657 = (inp[7]) ? 14'b00000000000000 : node1658;
												assign node1658 = (inp[2]) ? 14'b00000000000000 : node1659;
													assign node1659 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
								assign node1665 = (inp[5]) ? 14'b00000000000000 : node1666;
									assign node1666 = (inp[9]) ? node1668 : 14'b00000000000000;
										assign node1668 = (inp[7]) ? node1670 : 14'b00000000000000;
											assign node1670 = (inp[3]) ? 14'b00100100001101 : 14'b00000000000000;

endmodule