module dtc_split25_bm97 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node39;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node139;

	assign outp = (inp[3]) ? node28 : node1;
		assign node1 = (inp[9]) ? node3 : 3'b000;
			assign node3 = (inp[6]) ? node5 : 3'b000;
				assign node5 = (inp[7]) ? node7 : 3'b001;
					assign node7 = (inp[10]) ? node9 : 3'b000;
						assign node9 = (inp[4]) ? node19 : node10;
							assign node10 = (inp[11]) ? node12 : 3'b000;
								assign node12 = (inp[5]) ? node16 : node13;
									assign node13 = (inp[8]) ? 3'b100 : 3'b000;
									assign node16 = (inp[8]) ? 3'b101 : 3'b001;
							assign node19 = (inp[8]) ? node23 : node20;
								assign node20 = (inp[11]) ? 3'b000 : 3'b100;
								assign node23 = (inp[11]) ? node25 : 3'b100;
									assign node25 = (inp[2]) ? 3'b100 : 3'b110;
		assign node28 = (inp[9]) ? node44 : node29;
			assign node29 = (inp[7]) ? 3'b000 : node30;
				assign node30 = (inp[6]) ? 3'b000 : node31;
					assign node31 = (inp[4]) ? node33 : 3'b100;
						assign node33 = (inp[11]) ? node39 : node34;
							assign node34 = (inp[8]) ? 3'b100 : node35;
								assign node35 = (inp[2]) ? 3'b100 : 3'b000;
							assign node39 = (inp[8]) ? 3'b000 : 3'b100;
			assign node44 = (inp[4]) ? node98 : node45;
				assign node45 = (inp[10]) ? node79 : node46;
					assign node46 = (inp[2]) ? node72 : node47;
						assign node47 = (inp[1]) ? node63 : node48;
							assign node48 = (inp[11]) ? node56 : node49;
								assign node49 = (inp[6]) ? node53 : node50;
									assign node50 = (inp[7]) ? 3'b110 : 3'b000;
									assign node53 = (inp[7]) ? 3'b000 : 3'b110;
								assign node56 = (inp[7]) ? node60 : node57;
									assign node57 = (inp[6]) ? 3'b110 : 3'b000;
									assign node60 = (inp[6]) ? 3'b000 : 3'b110;
							assign node63 = (inp[11]) ? node65 : 3'b000;
								assign node65 = (inp[6]) ? node69 : node66;
									assign node66 = (inp[7]) ? 3'b110 : 3'b000;
									assign node69 = (inp[7]) ? 3'b000 : 3'b110;
						assign node72 = (inp[6]) ? node76 : node73;
							assign node73 = (inp[7]) ? 3'b110 : 3'b000;
							assign node76 = (inp[7]) ? 3'b000 : 3'b110;
					assign node79 = (inp[6]) ? node83 : node80;
						assign node80 = (inp[7]) ? 3'b110 : 3'b000;
						assign node83 = (inp[7]) ? node85 : 3'b110;
							assign node85 = (inp[5]) ? node91 : node86;
								assign node86 = (inp[2]) ? node88 : 3'b010;
									assign node88 = (inp[0]) ? 3'b000 : 3'b010;
								assign node91 = (inp[2]) ? node95 : node92;
									assign node92 = (inp[11]) ? 3'b100 : 3'b000;
									assign node95 = (inp[8]) ? 3'b010 : 3'b100;
				assign node98 = (inp[6]) ? node130 : node99;
					assign node99 = (inp[10]) ? node111 : node100;
						assign node100 = (inp[7]) ? 3'b001 : node101;
							assign node101 = (inp[11]) ? node103 : 3'b010;
								assign node103 = (inp[5]) ? node107 : node104;
									assign node104 = (inp[8]) ? 3'b010 : 3'b010;
									assign node107 = (inp[0]) ? 3'b110 : 3'b010;
						assign node111 = (inp[11]) ? node119 : node112;
							assign node112 = (inp[8]) ? 3'b001 : node113;
								assign node113 = (inp[7]) ? 3'b001 : node114;
									assign node114 = (inp[2]) ? 3'b001 : 3'b101;
							assign node119 = (inp[8]) ? node127 : node120;
								assign node120 = (inp[0]) ? node124 : node121;
									assign node121 = (inp[7]) ? 3'b001 : 3'b011;
									assign node124 = (inp[7]) ? 3'b001 : 3'b101;
								assign node127 = (inp[7]) ? 3'b110 : 3'b101;
					assign node130 = (inp[11]) ? node132 : 3'b000;
						assign node132 = (inp[8]) ? node138 : node133;
							assign node133 = (inp[10]) ? node135 : 3'b000;
								assign node135 = (inp[7]) ? 3'b000 : 3'b010;
							assign node138 = (inp[7]) ? 3'b000 : node139;
								assign node139 = (inp[10]) ? 3'b100 : 3'b000;

endmodule