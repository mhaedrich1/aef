module dtc_split66_bm14 (
	input  wire [13-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node7;
	wire [1-1:0] node9;
	wire [1-1:0] node11;
	wire [1-1:0] node13;
	wire [1-1:0] node15;
	wire [1-1:0] node18;
	wire [1-1:0] node19;
	wire [1-1:0] node21;
	wire [1-1:0] node23;
	wire [1-1:0] node25;
	wire [1-1:0] node27;
	wire [1-1:0] node30;
	wire [1-1:0] node31;
	wire [1-1:0] node33;
	wire [1-1:0] node34;
	wire [1-1:0] node36;
	wire [1-1:0] node39;
	wire [1-1:0] node40;
	wire [1-1:0] node43;
	wire [1-1:0] node46;
	wire [1-1:0] node47;
	wire [1-1:0] node49;
	wire [1-1:0] node50;
	wire [1-1:0] node53;
	wire [1-1:0] node56;
	wire [1-1:0] node57;
	wire [1-1:0] node59;
	wire [1-1:0] node62;
	wire [1-1:0] node63;
	wire [1-1:0] node67;
	wire [1-1:0] node68;
	wire [1-1:0] node69;
	wire [1-1:0] node71;
	wire [1-1:0] node73;
	wire [1-1:0] node75;
	wire [1-1:0] node77;
	wire [1-1:0] node80;
	wire [1-1:0] node81;
	wire [1-1:0] node83;
	wire [1-1:0] node85;
	wire [1-1:0] node87;
	wire [1-1:0] node90;
	wire [1-1:0] node91;
	wire [1-1:0] node92;
	wire [1-1:0] node94;
	wire [1-1:0] node97;
	wire [1-1:0] node98;
	wire [1-1:0] node101;
	wire [1-1:0] node104;
	wire [1-1:0] node105;
	wire [1-1:0] node107;
	wire [1-1:0] node110;
	wire [1-1:0] node111;
	wire [1-1:0] node115;
	wire [1-1:0] node116;
	wire [1-1:0] node117;
	wire [1-1:0] node119;
	wire [1-1:0] node120;
	wire [1-1:0] node122;
	wire [1-1:0] node125;
	wire [1-1:0] node126;
	wire [1-1:0] node129;
	wire [1-1:0] node132;
	wire [1-1:0] node133;
	wire [1-1:0] node135;
	wire [1-1:0] node136;
	wire [1-1:0] node139;
	wire [1-1:0] node142;
	wire [1-1:0] node143;
	wire [1-1:0] node145;
	wire [1-1:0] node148;
	wire [1-1:0] node149;
	wire [1-1:0] node153;
	wire [1-1:0] node154;
	wire [1-1:0] node155;
	wire [1-1:0] node157;
	wire [1-1:0] node159;
	wire [1-1:0] node162;
	wire [1-1:0] node163;
	wire [1-1:0] node165;
	wire [1-1:0] node168;
	wire [1-1:0] node169;
	wire [1-1:0] node173;
	wire [1-1:0] node174;
	wire [1-1:0] node175;
	wire [1-1:0] node177;
	wire [1-1:0] node180;
	wire [1-1:0] node181;
	wire [1-1:0] node185;
	wire [1-1:0] node186;
	wire [1-1:0] node187;
	wire [1-1:0] node192;
	wire [1-1:0] node193;
	wire [1-1:0] node194;
	wire [1-1:0] node195;
	wire [1-1:0] node197;
	wire [1-1:0] node199;
	wire [1-1:0] node201;
	wire [1-1:0] node203;
	wire [1-1:0] node206;
	wire [1-1:0] node207;
	wire [1-1:0] node209;
	wire [1-1:0] node211;
	wire [1-1:0] node213;
	wire [1-1:0] node216;
	wire [1-1:0] node217;
	wire [1-1:0] node219;
	wire [1-1:0] node221;
	wire [1-1:0] node224;
	wire [1-1:0] node225;
	wire [1-1:0] node226;
	wire [1-1:0] node229;
	wire [1-1:0] node232;
	wire [1-1:0] node233;
	wire [1-1:0] node237;
	wire [1-1:0] node238;
	wire [1-1:0] node239;
	wire [1-1:0] node241;
	wire [1-1:0] node243;
	wire [1-1:0] node245;
	wire [1-1:0] node248;
	wire [1-1:0] node249;
	wire [1-1:0] node251;
	wire [1-1:0] node253;
	wire [1-1:0] node256;
	wire [1-1:0] node257;
	wire [1-1:0] node259;
	wire [1-1:0] node262;
	wire [1-1:0] node263;
	wire [1-1:0] node267;
	wire [1-1:0] node268;
	wire [1-1:0] node269;
	wire [1-1:0] node271;
	wire [1-1:0] node272;
	wire [1-1:0] node275;
	wire [1-1:0] node278;
	wire [1-1:0] node279;
	wire [1-1:0] node281;
	wire [1-1:0] node284;
	wire [1-1:0] node285;
	wire [1-1:0] node289;
	wire [1-1:0] node290;
	wire [1-1:0] node291;
	wire [1-1:0] node293;
	wire [1-1:0] node296;
	wire [1-1:0] node297;
	wire [1-1:0] node301;
	wire [1-1:0] node302;
	wire [1-1:0] node303;
	wire [1-1:0] node308;
	wire [1-1:0] node309;
	wire [1-1:0] node310;
	wire [1-1:0] node311;
	wire [1-1:0] node313;
	wire [1-1:0] node315;
	wire [1-1:0] node317;
	wire [1-1:0] node320;
	wire [1-1:0] node321;
	wire [1-1:0] node323;
	wire [1-1:0] node325;
	wire [1-1:0] node328;
	wire [1-1:0] node329;
	wire [1-1:0] node331;
	wire [1-1:0] node334;
	wire [1-1:0] node335;
	wire [1-1:0] node339;
	wire [1-1:0] node340;
	wire [1-1:0] node341;
	wire [1-1:0] node343;
	wire [1-1:0] node345;
	wire [1-1:0] node348;
	wire [1-1:0] node349;
	wire [1-1:0] node350;
	wire [1-1:0] node353;
	wire [1-1:0] node356;
	wire [1-1:0] node357;
	wire [1-1:0] node361;
	wire [1-1:0] node362;
	wire [1-1:0] node363;
	wire [1-1:0] node365;
	wire [1-1:0] node368;
	wire [1-1:0] node369;
	wire [1-1:0] node373;
	wire [1-1:0] node374;
	wire [1-1:0] node375;
	wire [1-1:0] node380;
	wire [1-1:0] node381;
	wire [1-1:0] node382;
	wire [1-1:0] node383;
	wire [1-1:0] node385;
	wire [1-1:0] node387;
	wire [1-1:0] node390;
	wire [1-1:0] node391;
	wire [1-1:0] node393;
	wire [1-1:0] node396;
	wire [1-1:0] node397;
	wire [1-1:0] node401;
	wire [1-1:0] node402;
	wire [1-1:0] node403;
	wire [1-1:0] node405;
	wire [1-1:0] node408;
	wire [1-1:0] node409;
	wire [1-1:0] node413;
	wire [1-1:0] node414;
	wire [1-1:0] node415;
	wire [1-1:0] node420;
	wire [1-1:0] node421;
	wire [1-1:0] node422;
	wire [1-1:0] node423;
	wire [1-1:0] node425;
	wire [1-1:0] node428;
	wire [1-1:0] node429;
	wire [1-1:0] node433;
	wire [1-1:0] node434;
	wire [1-1:0] node435;
	wire [1-1:0] node440;
	wire [1-1:0] node441;
	wire [1-1:0] node442;
	wire [1-1:0] node443;
	wire [1-1:0] node449;
	wire [1-1:0] node450;
	wire [1-1:0] node451;
	wire [1-1:0] node452;
	wire [1-1:0] node453;
	wire [1-1:0] node455;
	wire [1-1:0] node457;
	wire [1-1:0] node459;
	wire [1-1:0] node460;
	wire [1-1:0] node463;
	wire [1-1:0] node466;
	wire [1-1:0] node467;
	wire [1-1:0] node469;
	wire [1-1:0] node471;
	wire [1-1:0] node473;
	wire [1-1:0] node476;
	wire [1-1:0] node477;
	wire [1-1:0] node479;
	wire [1-1:0] node481;
	wire [1-1:0] node484;
	wire [1-1:0] node485;
	wire [1-1:0] node487;
	wire [1-1:0] node490;
	wire [1-1:0] node491;
	wire [1-1:0] node495;
	wire [1-1:0] node496;
	wire [1-1:0] node497;
	wire [1-1:0] node499;
	wire [1-1:0] node501;
	wire [1-1:0] node503;
	wire [1-1:0] node506;
	wire [1-1:0] node507;
	wire [1-1:0] node509;
	wire [1-1:0] node511;
	wire [1-1:0] node514;
	wire [1-1:0] node515;
	wire [1-1:0] node517;
	wire [1-1:0] node520;
	wire [1-1:0] node521;
	wire [1-1:0] node525;
	wire [1-1:0] node526;
	wire [1-1:0] node527;
	wire [1-1:0] node529;
	wire [1-1:0] node531;
	wire [1-1:0] node534;
	wire [1-1:0] node535;
	wire [1-1:0] node537;
	wire [1-1:0] node540;
	wire [1-1:0] node541;
	wire [1-1:0] node545;
	wire [1-1:0] node546;
	wire [1-1:0] node547;
	wire [1-1:0] node549;
	wire [1-1:0] node552;
	wire [1-1:0] node553;
	wire [1-1:0] node557;
	wire [1-1:0] node558;
	wire [1-1:0] node559;
	wire [1-1:0] node564;
	wire [1-1:0] node565;
	wire [1-1:0] node566;
	wire [1-1:0] node567;
	wire [1-1:0] node569;
	wire [1-1:0] node571;
	wire [1-1:0] node573;
	wire [1-1:0] node576;
	wire [1-1:0] node577;
	wire [1-1:0] node579;
	wire [1-1:0] node581;
	wire [1-1:0] node584;
	wire [1-1:0] node585;
	wire [1-1:0] node587;
	wire [1-1:0] node590;
	wire [1-1:0] node591;
	wire [1-1:0] node595;
	wire [1-1:0] node596;
	wire [1-1:0] node597;
	wire [1-1:0] node599;
	wire [1-1:0] node601;
	wire [1-1:0] node604;
	wire [1-1:0] node605;
	wire [1-1:0] node607;
	wire [1-1:0] node610;
	wire [1-1:0] node611;
	wire [1-1:0] node615;
	wire [1-1:0] node616;
	wire [1-1:0] node617;
	wire [1-1:0] node619;
	wire [1-1:0] node622;
	wire [1-1:0] node623;
	wire [1-1:0] node627;
	wire [1-1:0] node628;
	wire [1-1:0] node632;
	wire [1-1:0] node633;
	wire [1-1:0] node634;
	wire [1-1:0] node635;
	wire [1-1:0] node637;
	wire [1-1:0] node638;
	wire [1-1:0] node641;
	wire [1-1:0] node644;
	wire [1-1:0] node645;
	wire [1-1:0] node647;
	wire [1-1:0] node650;
	wire [1-1:0] node651;
	wire [1-1:0] node655;
	wire [1-1:0] node656;
	wire [1-1:0] node657;
	wire [1-1:0] node659;
	wire [1-1:0] node662;
	wire [1-1:0] node663;
	wire [1-1:0] node667;
	wire [1-1:0] node668;
	wire [1-1:0] node669;
	wire [1-1:0] node674;
	wire [1-1:0] node675;
	wire [1-1:0] node676;
	wire [1-1:0] node677;
	wire [1-1:0] node679;
	wire [1-1:0] node682;
	wire [1-1:0] node683;
	wire [1-1:0] node687;
	wire [1-1:0] node688;
	wire [1-1:0] node689;
	wire [1-1:0] node692;
	wire [1-1:0] node696;
	wire [1-1:0] node697;
	wire [1-1:0] node698;
	wire [1-1:0] node699;
	wire [1-1:0] node705;
	wire [1-1:0] node706;
	wire [1-1:0] node707;
	wire [1-1:0] node708;
	wire [1-1:0] node709;
	wire [1-1:0] node711;
	wire [1-1:0] node713;
	wire [1-1:0] node715;
	wire [1-1:0] node718;
	wire [1-1:0] node719;
	wire [1-1:0] node721;
	wire [1-1:0] node723;
	wire [1-1:0] node726;
	wire [1-1:0] node727;
	wire [1-1:0] node729;
	wire [1-1:0] node732;
	wire [1-1:0] node733;
	wire [1-1:0] node737;
	wire [1-1:0] node738;
	wire [1-1:0] node739;
	wire [1-1:0] node741;
	wire [1-1:0] node743;
	wire [1-1:0] node746;
	wire [1-1:0] node747;
	wire [1-1:0] node749;
	wire [1-1:0] node752;
	wire [1-1:0] node753;
	wire [1-1:0] node757;
	wire [1-1:0] node758;
	wire [1-1:0] node759;
	wire [1-1:0] node761;
	wire [1-1:0] node764;
	wire [1-1:0] node765;
	wire [1-1:0] node769;
	wire [1-1:0] node770;
	wire [1-1:0] node771;
	wire [1-1:0] node776;
	wire [1-1:0] node777;
	wire [1-1:0] node778;
	wire [1-1:0] node779;
	wire [1-1:0] node781;
	wire [1-1:0] node783;
	wire [1-1:0] node786;
	wire [1-1:0] node787;
	wire [1-1:0] node789;
	wire [1-1:0] node792;
	wire [1-1:0] node793;
	wire [1-1:0] node797;
	wire [1-1:0] node798;
	wire [1-1:0] node799;
	wire [1-1:0] node801;
	wire [1-1:0] node804;
	wire [1-1:0] node805;
	wire [1-1:0] node809;
	wire [1-1:0] node810;
	wire [1-1:0] node811;
	wire [1-1:0] node816;
	wire [1-1:0] node817;
	wire [1-1:0] node818;
	wire [1-1:0] node819;
	wire [1-1:0] node821;
	wire [1-1:0] node824;
	wire [1-1:0] node825;
	wire [1-1:0] node829;
	wire [1-1:0] node830;
	wire [1-1:0] node831;
	wire [1-1:0] node836;
	wire [1-1:0] node837;
	wire [1-1:0] node838;
	wire [1-1:0] node839;
	wire [1-1:0] node845;
	wire [1-1:0] node846;
	wire [1-1:0] node847;
	wire [1-1:0] node848;
	wire [1-1:0] node849;
	wire [1-1:0] node851;
	wire [1-1:0] node853;
	wire [1-1:0] node856;
	wire [1-1:0] node857;
	wire [1-1:0] node859;
	wire [1-1:0] node862;
	wire [1-1:0] node863;
	wire [1-1:0] node867;
	wire [1-1:0] node868;
	wire [1-1:0] node869;
	wire [1-1:0] node871;
	wire [1-1:0] node874;
	wire [1-1:0] node875;
	wire [1-1:0] node879;
	wire [1-1:0] node880;
	wire [1-1:0] node881;
	wire [1-1:0] node884;
	wire [1-1:0] node888;
	wire [1-1:0] node889;
	wire [1-1:0] node890;
	wire [1-1:0] node891;
	wire [1-1:0] node893;
	wire [1-1:0] node896;
	wire [1-1:0] node897;
	wire [1-1:0] node901;
	wire [1-1:0] node902;
	wire [1-1:0] node903;
	wire [1-1:0] node906;
	wire [1-1:0] node910;
	wire [1-1:0] node911;
	wire [1-1:0] node912;
	wire [1-1:0] node913;
	wire [1-1:0] node919;
	wire [1-1:0] node920;
	wire [1-1:0] node921;
	wire [1-1:0] node922;
	wire [1-1:0] node923;
	wire [1-1:0] node925;
	wire [1-1:0] node928;
	wire [1-1:0] node929;
	wire [1-1:0] node933;
	wire [1-1:0] node934;
	wire [1-1:0] node935;
	wire [1-1:0] node940;
	wire [1-1:0] node941;
	wire [1-1:0] node942;
	wire [1-1:0] node943;
	wire [1-1:0] node949;
	wire [1-1:0] node950;
	wire [1-1:0] node951;
	wire [1-1:0] node952;
	wire [1-1:0] node953;
	wire [1-1:0] node960;
	wire [1-1:0] node961;
	wire [1-1:0] node962;
	wire [1-1:0] node963;
	wire [1-1:0] node964;
	wire [1-1:0] node965;
	wire [1-1:0] node967;
	wire [1-1:0] node969;
	wire [1-1:0] node971;
	wire [1-1:0] node973;
	wire [1-1:0] node976;
	wire [1-1:0] node977;
	wire [1-1:0] node979;
	wire [1-1:0] node981;
	wire [1-1:0] node983;
	wire [1-1:0] node986;
	wire [1-1:0] node987;
	wire [1-1:0] node989;
	wire [1-1:0] node991;
	wire [1-1:0] node994;
	wire [1-1:0] node995;
	wire [1-1:0] node997;
	wire [1-1:0] node1000;
	wire [1-1:0] node1001;
	wire [1-1:0] node1005;
	wire [1-1:0] node1006;
	wire [1-1:0] node1007;
	wire [1-1:0] node1009;
	wire [1-1:0] node1011;
	wire [1-1:0] node1013;
	wire [1-1:0] node1016;
	wire [1-1:0] node1017;
	wire [1-1:0] node1019;
	wire [1-1:0] node1021;
	wire [1-1:0] node1024;
	wire [1-1:0] node1025;
	wire [1-1:0] node1027;
	wire [1-1:0] node1030;
	wire [1-1:0] node1031;
	wire [1-1:0] node1035;
	wire [1-1:0] node1036;
	wire [1-1:0] node1037;
	wire [1-1:0] node1039;
	wire [1-1:0] node1041;
	wire [1-1:0] node1044;
	wire [1-1:0] node1045;
	wire [1-1:0] node1047;
	wire [1-1:0] node1050;
	wire [1-1:0] node1051;
	wire [1-1:0] node1055;
	wire [1-1:0] node1056;
	wire [1-1:0] node1057;
	wire [1-1:0] node1059;
	wire [1-1:0] node1062;
	wire [1-1:0] node1063;
	wire [1-1:0] node1067;
	wire [1-1:0] node1068;
	wire [1-1:0] node1069;
	wire [1-1:0] node1074;
	wire [1-1:0] node1075;
	wire [1-1:0] node1076;
	wire [1-1:0] node1077;
	wire [1-1:0] node1079;
	wire [1-1:0] node1081;
	wire [1-1:0] node1083;
	wire [1-1:0] node1086;
	wire [1-1:0] node1087;
	wire [1-1:0] node1088;
	wire [1-1:0] node1090;
	wire [1-1:0] node1093;
	wire [1-1:0] node1094;
	wire [1-1:0] node1097;
	wire [1-1:0] node1100;
	wire [1-1:0] node1101;
	wire [1-1:0] node1103;
	wire [1-1:0] node1106;
	wire [1-1:0] node1107;
	wire [1-1:0] node1111;
	wire [1-1:0] node1112;
	wire [1-1:0] node1113;
	wire [1-1:0] node1115;
	wire [1-1:0] node1116;
	wire [1-1:0] node1119;
	wire [1-1:0] node1122;
	wire [1-1:0] node1123;
	wire [1-1:0] node1124;
	wire [1-1:0] node1127;
	wire [1-1:0] node1130;
	wire [1-1:0] node1131;
	wire [1-1:0] node1135;
	wire [1-1:0] node1136;
	wire [1-1:0] node1137;
	wire [1-1:0] node1139;
	wire [1-1:0] node1142;
	wire [1-1:0] node1143;
	wire [1-1:0] node1147;
	wire [1-1:0] node1148;
	wire [1-1:0] node1149;
	wire [1-1:0] node1154;
	wire [1-1:0] node1155;
	wire [1-1:0] node1156;
	wire [1-1:0] node1157;
	wire [1-1:0] node1159;
	wire [1-1:0] node1161;
	wire [1-1:0] node1164;
	wire [1-1:0] node1165;
	wire [1-1:0] node1167;
	wire [1-1:0] node1170;
	wire [1-1:0] node1171;
	wire [1-1:0] node1175;
	wire [1-1:0] node1176;
	wire [1-1:0] node1177;
	wire [1-1:0] node1179;
	wire [1-1:0] node1182;
	wire [1-1:0] node1183;
	wire [1-1:0] node1187;
	wire [1-1:0] node1188;
	wire [1-1:0] node1189;
	wire [1-1:0] node1194;
	wire [1-1:0] node1195;
	wire [1-1:0] node1196;
	wire [1-1:0] node1197;
	wire [1-1:0] node1199;
	wire [1-1:0] node1202;
	wire [1-1:0] node1203;
	wire [1-1:0] node1207;
	wire [1-1:0] node1208;
	wire [1-1:0] node1209;
	wire [1-1:0] node1214;
	wire [1-1:0] node1215;
	wire [1-1:0] node1216;
	wire [1-1:0] node1217;
	wire [1-1:0] node1223;
	wire [1-1:0] node1224;
	wire [1-1:0] node1225;
	wire [1-1:0] node1226;
	wire [1-1:0] node1227;
	wire [1-1:0] node1229;
	wire [1-1:0] node1231;
	wire [1-1:0] node1233;
	wire [1-1:0] node1236;
	wire [1-1:0] node1237;
	wire [1-1:0] node1239;
	wire [1-1:0] node1241;
	wire [1-1:0] node1244;
	wire [1-1:0] node1245;
	wire [1-1:0] node1247;
	wire [1-1:0] node1250;
	wire [1-1:0] node1251;
	wire [1-1:0] node1255;
	wire [1-1:0] node1256;
	wire [1-1:0] node1257;
	wire [1-1:0] node1259;
	wire [1-1:0] node1261;
	wire [1-1:0] node1264;
	wire [1-1:0] node1265;
	wire [1-1:0] node1267;
	wire [1-1:0] node1270;
	wire [1-1:0] node1271;
	wire [1-1:0] node1275;
	wire [1-1:0] node1276;
	wire [1-1:0] node1277;
	wire [1-1:0] node1279;
	wire [1-1:0] node1282;
	wire [1-1:0] node1283;
	wire [1-1:0] node1287;
	wire [1-1:0] node1288;
	wire [1-1:0] node1289;
	wire [1-1:0] node1294;
	wire [1-1:0] node1295;
	wire [1-1:0] node1296;
	wire [1-1:0] node1297;
	wire [1-1:0] node1299;
	wire [1-1:0] node1301;
	wire [1-1:0] node1304;
	wire [1-1:0] node1305;
	wire [1-1:0] node1306;
	wire [1-1:0] node1309;
	wire [1-1:0] node1312;
	wire [1-1:0] node1313;
	wire [1-1:0] node1316;
	wire [1-1:0] node1319;
	wire [1-1:0] node1320;
	wire [1-1:0] node1321;
	wire [1-1:0] node1323;
	wire [1-1:0] node1326;
	wire [1-1:0] node1327;
	wire [1-1:0] node1330;
	wire [1-1:0] node1333;
	wire [1-1:0] node1334;
	wire [1-1:0] node1335;
	wire [1-1:0] node1340;
	wire [1-1:0] node1341;
	wire [1-1:0] node1342;
	wire [1-1:0] node1343;
	wire [1-1:0] node1345;
	wire [1-1:0] node1348;
	wire [1-1:0] node1349;
	wire [1-1:0] node1353;
	wire [1-1:0] node1354;
	wire [1-1:0] node1355;
	wire [1-1:0] node1360;
	wire [1-1:0] node1361;
	wire [1-1:0] node1362;
	wire [1-1:0] node1363;
	wire [1-1:0] node1369;
	wire [1-1:0] node1370;
	wire [1-1:0] node1371;
	wire [1-1:0] node1372;
	wire [1-1:0] node1373;
	wire [1-1:0] node1375;
	wire [1-1:0] node1376;
	wire [1-1:0] node1379;
	wire [1-1:0] node1382;
	wire [1-1:0] node1383;
	wire [1-1:0] node1385;
	wire [1-1:0] node1388;
	wire [1-1:0] node1389;
	wire [1-1:0] node1393;
	wire [1-1:0] node1394;
	wire [1-1:0] node1395;
	wire [1-1:0] node1397;
	wire [1-1:0] node1400;
	wire [1-1:0] node1401;
	wire [1-1:0] node1405;
	wire [1-1:0] node1406;
	wire [1-1:0] node1407;
	wire [1-1:0] node1412;
	wire [1-1:0] node1413;
	wire [1-1:0] node1414;
	wire [1-1:0] node1415;
	wire [1-1:0] node1417;
	wire [1-1:0] node1420;
	wire [1-1:0] node1421;
	wire [1-1:0] node1425;
	wire [1-1:0] node1426;
	wire [1-1:0] node1427;
	wire [1-1:0] node1432;
	wire [1-1:0] node1433;
	wire [1-1:0] node1434;
	wire [1-1:0] node1435;
	wire [1-1:0] node1441;
	wire [1-1:0] node1442;
	wire [1-1:0] node1443;
	wire [1-1:0] node1444;
	wire [1-1:0] node1445;
	wire [1-1:0] node1447;
	wire [1-1:0] node1450;
	wire [1-1:0] node1451;
	wire [1-1:0] node1455;
	wire [1-1:0] node1456;
	wire [1-1:0] node1457;
	wire [1-1:0] node1462;
	wire [1-1:0] node1463;
	wire [1-1:0] node1464;
	wire [1-1:0] node1465;
	wire [1-1:0] node1471;
	wire [1-1:0] node1472;
	wire [1-1:0] node1473;
	wire [1-1:0] node1474;
	wire [1-1:0] node1480;
	wire [1-1:0] node1481;
	wire [1-1:0] node1482;
	wire [1-1:0] node1483;
	wire [1-1:0] node1484;
	wire [1-1:0] node1485;
	wire [1-1:0] node1487;
	wire [1-1:0] node1489;
	wire [1-1:0] node1491;
	wire [1-1:0] node1494;
	wire [1-1:0] node1495;
	wire [1-1:0] node1497;
	wire [1-1:0] node1499;
	wire [1-1:0] node1502;
	wire [1-1:0] node1503;
	wire [1-1:0] node1505;
	wire [1-1:0] node1508;
	wire [1-1:0] node1509;
	wire [1-1:0] node1513;
	wire [1-1:0] node1514;
	wire [1-1:0] node1515;
	wire [1-1:0] node1517;
	wire [1-1:0] node1519;
	wire [1-1:0] node1522;
	wire [1-1:0] node1523;
	wire [1-1:0] node1525;
	wire [1-1:0] node1528;
	wire [1-1:0] node1529;
	wire [1-1:0] node1532;
	wire [1-1:0] node1535;
	wire [1-1:0] node1536;
	wire [1-1:0] node1537;
	wire [1-1:0] node1539;
	wire [1-1:0] node1542;
	wire [1-1:0] node1543;
	wire [1-1:0] node1547;
	wire [1-1:0] node1548;
	wire [1-1:0] node1549;
	wire [1-1:0] node1554;
	wire [1-1:0] node1555;
	wire [1-1:0] node1556;
	wire [1-1:0] node1557;
	wire [1-1:0] node1559;
	wire [1-1:0] node1560;
	wire [1-1:0] node1564;
	wire [1-1:0] node1565;
	wire [1-1:0] node1567;
	wire [1-1:0] node1570;
	wire [1-1:0] node1571;
	wire [1-1:0] node1575;
	wire [1-1:0] node1576;
	wire [1-1:0] node1577;
	wire [1-1:0] node1579;
	wire [1-1:0] node1582;
	wire [1-1:0] node1583;
	wire [1-1:0] node1587;
	wire [1-1:0] node1588;
	wire [1-1:0] node1589;
	wire [1-1:0] node1594;
	wire [1-1:0] node1595;
	wire [1-1:0] node1596;
	wire [1-1:0] node1597;
	wire [1-1:0] node1599;
	wire [1-1:0] node1602;
	wire [1-1:0] node1603;
	wire [1-1:0] node1607;
	wire [1-1:0] node1608;
	wire [1-1:0] node1609;
	wire [1-1:0] node1612;
	wire [1-1:0] node1616;
	wire [1-1:0] node1617;
	wire [1-1:0] node1618;
	wire [1-1:0] node1619;
	wire [1-1:0] node1625;
	wire [1-1:0] node1626;
	wire [1-1:0] node1627;
	wire [1-1:0] node1628;
	wire [1-1:0] node1629;
	wire [1-1:0] node1631;
	wire [1-1:0] node1633;
	wire [1-1:0] node1636;
	wire [1-1:0] node1637;
	wire [1-1:0] node1639;
	wire [1-1:0] node1642;
	wire [1-1:0] node1643;
	wire [1-1:0] node1647;
	wire [1-1:0] node1648;
	wire [1-1:0] node1649;
	wire [1-1:0] node1651;
	wire [1-1:0] node1654;
	wire [1-1:0] node1655;
	wire [1-1:0] node1658;
	wire [1-1:0] node1661;
	wire [1-1:0] node1662;
	wire [1-1:0] node1663;
	wire [1-1:0] node1668;
	wire [1-1:0] node1669;
	wire [1-1:0] node1670;
	wire [1-1:0] node1671;
	wire [1-1:0] node1673;
	wire [1-1:0] node1676;
	wire [1-1:0] node1677;
	wire [1-1:0] node1681;
	wire [1-1:0] node1682;
	wire [1-1:0] node1683;
	wire [1-1:0] node1688;
	wire [1-1:0] node1689;
	wire [1-1:0] node1690;
	wire [1-1:0] node1691;
	wire [1-1:0] node1697;
	wire [1-1:0] node1698;
	wire [1-1:0] node1699;
	wire [1-1:0] node1700;
	wire [1-1:0] node1701;
	wire [1-1:0] node1703;
	wire [1-1:0] node1706;
	wire [1-1:0] node1707;
	wire [1-1:0] node1710;
	wire [1-1:0] node1713;
	wire [1-1:0] node1714;
	wire [1-1:0] node1715;
	wire [1-1:0] node1720;
	wire [1-1:0] node1721;
	wire [1-1:0] node1722;
	wire [1-1:0] node1723;
	wire [1-1:0] node1729;
	wire [1-1:0] node1730;
	wire [1-1:0] node1731;
	wire [1-1:0] node1732;
	wire [1-1:0] node1733;
	wire [1-1:0] node1740;
	wire [1-1:0] node1741;
	wire [1-1:0] node1742;
	wire [1-1:0] node1743;
	wire [1-1:0] node1744;
	wire [1-1:0] node1745;
	wire [1-1:0] node1747;
	wire [1-1:0] node1749;
	wire [1-1:0] node1752;
	wire [1-1:0] node1753;
	wire [1-1:0] node1754;
	wire [1-1:0] node1757;
	wire [1-1:0] node1760;
	wire [1-1:0] node1761;
	wire [1-1:0] node1765;
	wire [1-1:0] node1766;
	wire [1-1:0] node1767;
	wire [1-1:0] node1769;
	wire [1-1:0] node1772;
	wire [1-1:0] node1773;
	wire [1-1:0] node1777;
	wire [1-1:0] node1778;
	wire [1-1:0] node1779;
	wire [1-1:0] node1784;
	wire [1-1:0] node1785;
	wire [1-1:0] node1786;
	wire [1-1:0] node1787;
	wire [1-1:0] node1789;
	wire [1-1:0] node1792;
	wire [1-1:0] node1793;
	wire [1-1:0] node1797;
	wire [1-1:0] node1798;
	wire [1-1:0] node1799;
	wire [1-1:0] node1802;
	wire [1-1:0] node1806;
	wire [1-1:0] node1807;
	wire [1-1:0] node1808;
	wire [1-1:0] node1809;
	wire [1-1:0] node1815;
	wire [1-1:0] node1816;
	wire [1-1:0] node1817;
	wire [1-1:0] node1818;
	wire [1-1:0] node1819;
	wire [1-1:0] node1821;
	wire [1-1:0] node1824;
	wire [1-1:0] node1825;
	wire [1-1:0] node1829;
	wire [1-1:0] node1830;
	wire [1-1:0] node1831;
	wire [1-1:0] node1834;
	wire [1-1:0] node1838;
	wire [1-1:0] node1839;
	wire [1-1:0] node1840;
	wire [1-1:0] node1841;
	wire [1-1:0] node1844;
	wire [1-1:0] node1849;
	wire [1-1:0] node1850;
	wire [1-1:0] node1851;
	wire [1-1:0] node1852;
	wire [1-1:0] node1853;
	wire [1-1:0] node1860;
	wire [1-1:0] node1861;
	wire [1-1:0] node1862;
	wire [1-1:0] node1863;
	wire [1-1:0] node1864;
	wire [1-1:0] node1865;
	wire [1-1:0] node1867;
	wire [1-1:0] node1870;
	wire [1-1:0] node1871;
	wire [1-1:0] node1875;
	wire [1-1:0] node1876;
	wire [1-1:0] node1877;
	wire [1-1:0] node1882;
	wire [1-1:0] node1883;
	wire [1-1:0] node1884;
	wire [1-1:0] node1885;
	wire [1-1:0] node1888;
	wire [1-1:0] node1893;
	wire [1-1:0] node1894;
	wire [1-1:0] node1895;
	wire [1-1:0] node1896;
	wire [1-1:0] node1897;
	wire [1-1:0] node1904;
	wire [1-1:0] node1905;
	wire [1-1:0] node1906;
	wire [1-1:0] node1907;
	wire [1-1:0] node1908;
	wire [1-1:0] node1909;

	assign outp = (inp[11]) ? node960 : node1;
		assign node1 = (inp[2]) ? node449 : node2;
			assign node2 = (inp[0]) ? node192 : node3;
				assign node3 = (inp[4]) ? node67 : node4;
					assign node4 = (inp[5]) ? node18 : node5;
						assign node5 = (inp[3]) ? node7 : 1'b1;
							assign node7 = (inp[1]) ? node9 : 1'b1;
								assign node9 = (inp[7]) ? node11 : 1'b1;
									assign node11 = (inp[6]) ? node13 : 1'b1;
										assign node13 = (inp[9]) ? node15 : 1'b1;
											assign node15 = (inp[12]) ? 1'b0 : 1'b1;
						assign node18 = (inp[12]) ? node30 : node19;
							assign node19 = (inp[10]) ? node21 : 1'b1;
								assign node21 = (inp[7]) ? node23 : 1'b1;
									assign node23 = (inp[8]) ? node25 : 1'b1;
										assign node25 = (inp[6]) ? node27 : 1'b1;
											assign node27 = (inp[1]) ? 1'b0 : 1'b1;
							assign node30 = (inp[10]) ? node46 : node31;
								assign node31 = (inp[1]) ? node33 : 1'b1;
									assign node33 = (inp[3]) ? node39 : node34;
										assign node34 = (inp[9]) ? node36 : 1'b1;
											assign node36 = (inp[6]) ? 1'b1 : 1'b1;
										assign node39 = (inp[9]) ? node43 : node40;
											assign node40 = (inp[7]) ? 1'b1 : 1'b1;
											assign node43 = (inp[6]) ? 1'b0 : 1'b0;
								assign node46 = (inp[9]) ? node56 : node47;
									assign node47 = (inp[1]) ? node49 : 1'b1;
										assign node49 = (inp[3]) ? node53 : node50;
											assign node50 = (inp[6]) ? 1'b1 : 1'b1;
											assign node53 = (inp[7]) ? 1'b0 : 1'b0;
									assign node56 = (inp[7]) ? node62 : node57;
										assign node57 = (inp[8]) ? node59 : 1'b1;
											assign node59 = (inp[6]) ? 1'b0 : 1'b1;
										assign node62 = (inp[1]) ? 1'b0 : node63;
											assign node63 = (inp[8]) ? 1'b0 : 1'b1;
					assign node67 = (inp[3]) ? node115 : node68;
						assign node68 = (inp[7]) ? node80 : node69;
							assign node69 = (inp[5]) ? node71 : 1'b1;
								assign node71 = (inp[8]) ? node73 : 1'b1;
									assign node73 = (inp[10]) ? node75 : 1'b1;
										assign node75 = (inp[9]) ? node77 : 1'b1;
											assign node77 = (inp[1]) ? 1'b0 : 1'b1;
							assign node80 = (inp[9]) ? node90 : node81;
								assign node81 = (inp[6]) ? node83 : 1'b1;
									assign node83 = (inp[5]) ? node85 : 1'b1;
										assign node85 = (inp[12]) ? node87 : 1'b1;
											assign node87 = (inp[8]) ? 1'b0 : 1'b1;
								assign node90 = (inp[1]) ? node104 : node91;
									assign node91 = (inp[8]) ? node97 : node92;
										assign node92 = (inp[10]) ? node94 : 1'b1;
											assign node94 = (inp[6]) ? 1'b1 : 1'b1;
										assign node97 = (inp[12]) ? node101 : node98;
											assign node98 = (inp[10]) ? 1'b1 : 1'b1;
											assign node101 = (inp[6]) ? 1'b0 : 1'b1;
									assign node104 = (inp[8]) ? node110 : node105;
										assign node105 = (inp[10]) ? node107 : 1'b1;
											assign node107 = (inp[6]) ? 1'b0 : 1'b0;
										assign node110 = (inp[5]) ? 1'b0 : node111;
											assign node111 = (inp[6]) ? 1'b1 : 1'b0;
						assign node115 = (inp[9]) ? node153 : node116;
							assign node116 = (inp[7]) ? node132 : node117;
								assign node117 = (inp[5]) ? node119 : 1'b1;
									assign node119 = (inp[10]) ? node125 : node120;
										assign node120 = (inp[6]) ? node122 : 1'b1;
											assign node122 = (inp[1]) ? 1'b1 : 1'b1;
										assign node125 = (inp[1]) ? node129 : node126;
											assign node126 = (inp[12]) ? 1'b1 : 1'b1;
											assign node129 = (inp[6]) ? 1'b0 : 1'b1;
								assign node132 = (inp[12]) ? node142 : node133;
									assign node133 = (inp[10]) ? node135 : 1'b1;
										assign node135 = (inp[6]) ? node139 : node136;
											assign node136 = (inp[1]) ? 1'b1 : 1'b1;
											assign node139 = (inp[5]) ? 1'b0 : 1'b1;
									assign node142 = (inp[6]) ? node148 : node143;
										assign node143 = (inp[10]) ? node145 : 1'b1;
											assign node145 = (inp[8]) ? 1'b0 : 1'b1;
										assign node148 = (inp[5]) ? 1'b0 : node149;
											assign node149 = (inp[8]) ? 1'b0 : 1'b1;
							assign node153 = (inp[10]) ? node173 : node154;
								assign node154 = (inp[1]) ? node162 : node155;
									assign node155 = (inp[12]) ? node157 : 1'b1;
										assign node157 = (inp[6]) ? node159 : 1'b1;
											assign node159 = (inp[7]) ? 1'b0 : 1'b1;
									assign node162 = (inp[8]) ? node168 : node163;
										assign node163 = (inp[7]) ? node165 : 1'b1;
											assign node165 = (inp[5]) ? 1'b0 : 1'b1;
										assign node168 = (inp[5]) ? 1'b0 : node169;
											assign node169 = (inp[6]) ? 1'b0 : 1'b1;
								assign node173 = (inp[6]) ? node185 : node174;
									assign node174 = (inp[8]) ? node180 : node175;
										assign node175 = (inp[7]) ? node177 : 1'b1;
											assign node177 = (inp[12]) ? 1'b0 : 1'b1;
										assign node180 = (inp[5]) ? 1'b0 : node181;
											assign node181 = (inp[1]) ? 1'b0 : 1'b1;
									assign node185 = (inp[12]) ? 1'b0 : node186;
										assign node186 = (inp[8]) ? 1'b0 : node187;
											assign node187 = (inp[5]) ? 1'b0 : 1'b1;
				assign node192 = (inp[7]) ? node308 : node193;
					assign node193 = (inp[10]) ? node237 : node194;
						assign node194 = (inp[1]) ? node206 : node195;
							assign node195 = (inp[8]) ? node197 : 1'b1;
								assign node197 = (inp[4]) ? node199 : 1'b1;
									assign node199 = (inp[12]) ? node201 : 1'b1;
										assign node201 = (inp[5]) ? node203 : 1'b1;
											assign node203 = (inp[3]) ? 1'b0 : 1'b1;
							assign node206 = (inp[4]) ? node216 : node207;
								assign node207 = (inp[3]) ? node209 : 1'b1;
									assign node209 = (inp[12]) ? node211 : 1'b1;
										assign node211 = (inp[5]) ? node213 : 1'b1;
											assign node213 = (inp[6]) ? 1'b0 : 1'b0;
								assign node216 = (inp[6]) ? node224 : node217;
									assign node217 = (inp[12]) ? node219 : 1'b1;
										assign node219 = (inp[3]) ? node221 : 1'b1;
											assign node221 = (inp[5]) ? 1'b0 : 1'b1;
									assign node224 = (inp[8]) ? node232 : node225;
										assign node225 = (inp[12]) ? node229 : node226;
											assign node226 = (inp[9]) ? 1'b1 : 1'b1;
											assign node229 = (inp[3]) ? 1'b0 : 1'b1;
										assign node232 = (inp[5]) ? 1'b0 : node233;
											assign node233 = (inp[3]) ? 1'b0 : 1'b1;
						assign node237 = (inp[9]) ? node267 : node238;
							assign node238 = (inp[1]) ? node248 : node239;
								assign node239 = (inp[6]) ? node241 : 1'b1;
									assign node241 = (inp[8]) ? node243 : 1'b1;
										assign node243 = (inp[4]) ? node245 : 1'b1;
											assign node245 = (inp[5]) ? 1'b0 : 1'b1;
								assign node248 = (inp[6]) ? node256 : node249;
									assign node249 = (inp[5]) ? node251 : 1'b1;
										assign node251 = (inp[3]) ? node253 : 1'b1;
											assign node253 = (inp[4]) ? 1'b0 : 1'b1;
									assign node256 = (inp[8]) ? node262 : node257;
										assign node257 = (inp[3]) ? node259 : 1'b1;
											assign node259 = (inp[5]) ? 1'b0 : 1'b1;
										assign node262 = (inp[12]) ? 1'b0 : node263;
											assign node263 = (inp[3]) ? 1'b0 : 1'b1;
							assign node267 = (inp[8]) ? node289 : node268;
								assign node268 = (inp[5]) ? node278 : node269;
									assign node269 = (inp[12]) ? node271 : 1'b1;
										assign node271 = (inp[3]) ? node275 : node272;
											assign node272 = (inp[1]) ? 1'b1 : 1'b1;
											assign node275 = (inp[1]) ? 1'b0 : 1'b0;
									assign node278 = (inp[1]) ? node284 : node279;
										assign node279 = (inp[3]) ? node281 : 1'b1;
											assign node281 = (inp[12]) ? 1'b0 : 1'b1;
										assign node284 = (inp[6]) ? 1'b0 : node285;
											assign node285 = (inp[4]) ? 1'b0 : 1'b1;
								assign node289 = (inp[6]) ? node301 : node290;
									assign node290 = (inp[12]) ? node296 : node291;
										assign node291 = (inp[1]) ? node293 : 1'b1;
											assign node293 = (inp[5]) ? 1'b0 : 1'b1;
										assign node296 = (inp[5]) ? 1'b0 : node297;
											assign node297 = (inp[1]) ? 1'b0 : 1'b1;
									assign node301 = (inp[5]) ? 1'b0 : node302;
										assign node302 = (inp[12]) ? 1'b0 : node303;
											assign node303 = (inp[3]) ? 1'b0 : 1'b1;
					assign node308 = (inp[5]) ? node380 : node309;
						assign node309 = (inp[6]) ? node339 : node310;
							assign node310 = (inp[9]) ? node320 : node311;
								assign node311 = (inp[3]) ? node313 : 1'b1;
									assign node313 = (inp[10]) ? node315 : 1'b1;
										assign node315 = (inp[12]) ? node317 : 1'b1;
											assign node317 = (inp[4]) ? 1'b0 : 1'b1;
								assign node320 = (inp[1]) ? node328 : node321;
									assign node321 = (inp[12]) ? node323 : 1'b1;
										assign node323 = (inp[8]) ? node325 : 1'b1;
											assign node325 = (inp[4]) ? 1'b0 : 1'b1;
									assign node328 = (inp[10]) ? node334 : node329;
										assign node329 = (inp[3]) ? node331 : 1'b1;
											assign node331 = (inp[12]) ? 1'b0 : 1'b1;
										assign node334 = (inp[3]) ? 1'b0 : node335;
											assign node335 = (inp[4]) ? 1'b0 : 1'b1;
							assign node339 = (inp[8]) ? node361 : node340;
								assign node340 = (inp[12]) ? node348 : node341;
									assign node341 = (inp[3]) ? node343 : 1'b1;
										assign node343 = (inp[10]) ? node345 : 1'b1;
											assign node345 = (inp[9]) ? 1'b0 : 1'b1;
									assign node348 = (inp[9]) ? node356 : node349;
										assign node349 = (inp[4]) ? node353 : node350;
											assign node350 = (inp[1]) ? 1'b1 : 1'b1;
											assign node353 = (inp[1]) ? 1'b0 : 1'b1;
										assign node356 = (inp[3]) ? 1'b0 : node357;
											assign node357 = (inp[10]) ? 1'b0 : 1'b1;
								assign node361 = (inp[4]) ? node373 : node362;
									assign node362 = (inp[9]) ? node368 : node363;
										assign node363 = (inp[3]) ? node365 : 1'b1;
											assign node365 = (inp[10]) ? 1'b0 : 1'b1;
										assign node368 = (inp[1]) ? 1'b0 : node369;
											assign node369 = (inp[12]) ? 1'b0 : 1'b1;
									assign node373 = (inp[9]) ? 1'b0 : node374;
										assign node374 = (inp[1]) ? 1'b0 : node375;
											assign node375 = (inp[3]) ? 1'b0 : 1'b1;
						assign node380 = (inp[1]) ? node420 : node381;
							assign node381 = (inp[4]) ? node401 : node382;
								assign node382 = (inp[3]) ? node390 : node383;
									assign node383 = (inp[8]) ? node385 : 1'b1;
										assign node385 = (inp[12]) ? node387 : 1'b1;
											assign node387 = (inp[9]) ? 1'b0 : 1'b1;
									assign node390 = (inp[9]) ? node396 : node391;
										assign node391 = (inp[6]) ? node393 : 1'b1;
											assign node393 = (inp[12]) ? 1'b0 : 1'b1;
										assign node396 = (inp[8]) ? 1'b0 : node397;
											assign node397 = (inp[6]) ? 1'b0 : 1'b1;
								assign node401 = (inp[12]) ? node413 : node402;
									assign node402 = (inp[8]) ? node408 : node403;
										assign node403 = (inp[9]) ? node405 : 1'b1;
											assign node405 = (inp[6]) ? 1'b0 : 1'b1;
										assign node408 = (inp[3]) ? 1'b0 : node409;
											assign node409 = (inp[6]) ? 1'b0 : 1'b1;
									assign node413 = (inp[8]) ? 1'b0 : node414;
										assign node414 = (inp[6]) ? 1'b0 : node415;
											assign node415 = (inp[3]) ? 1'b0 : 1'b1;
							assign node420 = (inp[12]) ? node440 : node421;
								assign node421 = (inp[8]) ? node433 : node422;
									assign node422 = (inp[9]) ? node428 : node423;
										assign node423 = (inp[4]) ? node425 : 1'b1;
											assign node425 = (inp[6]) ? 1'b0 : 1'b1;
										assign node428 = (inp[10]) ? 1'b0 : node429;
											assign node429 = (inp[3]) ? 1'b0 : 1'b1;
									assign node433 = (inp[6]) ? 1'b0 : node434;
										assign node434 = (inp[4]) ? 1'b0 : node435;
											assign node435 = (inp[9]) ? 1'b0 : 1'b1;
								assign node440 = (inp[9]) ? 1'b0 : node441;
									assign node441 = (inp[6]) ? 1'b0 : node442;
										assign node442 = (inp[3]) ? 1'b0 : node443;
											assign node443 = (inp[4]) ? 1'b0 : 1'b1;
			assign node449 = (inp[10]) ? node705 : node450;
				assign node450 = (inp[5]) ? node564 : node451;
					assign node451 = (inp[1]) ? node495 : node452;
						assign node452 = (inp[12]) ? node466 : node453;
							assign node453 = (inp[0]) ? node455 : 1'b1;
								assign node455 = (inp[9]) ? node457 : 1'b1;
									assign node457 = (inp[6]) ? node459 : 1'b1;
										assign node459 = (inp[7]) ? node463 : node460;
											assign node460 = (inp[8]) ? 1'b0 : 1'b1;
											assign node463 = (inp[4]) ? 1'b0 : 1'b1;
							assign node466 = (inp[7]) ? node476 : node467;
								assign node467 = (inp[6]) ? node469 : 1'b1;
									assign node469 = (inp[9]) ? node471 : 1'b1;
										assign node471 = (inp[3]) ? node473 : 1'b1;
											assign node473 = (inp[0]) ? 1'b0 : 1'b1;
								assign node476 = (inp[4]) ? node484 : node477;
									assign node477 = (inp[8]) ? node479 : 1'b1;
										assign node479 = (inp[6]) ? node481 : 1'b1;
											assign node481 = (inp[9]) ? 1'b0 : 1'b1;
									assign node484 = (inp[3]) ? node490 : node485;
										assign node485 = (inp[9]) ? node487 : 1'b1;
											assign node487 = (inp[0]) ? 1'b0 : 1'b1;
										assign node490 = (inp[0]) ? 1'b0 : node491;
											assign node491 = (inp[6]) ? 1'b0 : 1'b1;
						assign node495 = (inp[8]) ? node525 : node496;
							assign node496 = (inp[9]) ? node506 : node497;
								assign node497 = (inp[3]) ? node499 : 1'b1;
									assign node499 = (inp[7]) ? node501 : 1'b1;
										assign node501 = (inp[12]) ? node503 : 1'b1;
											assign node503 = (inp[6]) ? 1'b0 : 1'b1;
								assign node506 = (inp[0]) ? node514 : node507;
									assign node507 = (inp[3]) ? node509 : 1'b1;
										assign node509 = (inp[12]) ? node511 : 1'b1;
											assign node511 = (inp[4]) ? 1'b0 : 1'b1;
									assign node514 = (inp[6]) ? node520 : node515;
										assign node515 = (inp[7]) ? node517 : 1'b1;
											assign node517 = (inp[4]) ? 1'b0 : 1'b1;
										assign node520 = (inp[3]) ? 1'b0 : node521;
											assign node521 = (inp[7]) ? 1'b0 : 1'b1;
							assign node525 = (inp[6]) ? node545 : node526;
								assign node526 = (inp[0]) ? node534 : node527;
									assign node527 = (inp[9]) ? node529 : 1'b1;
										assign node529 = (inp[7]) ? node531 : 1'b1;
											assign node531 = (inp[4]) ? 1'b0 : 1'b1;
									assign node534 = (inp[3]) ? node540 : node535;
										assign node535 = (inp[4]) ? node537 : 1'b1;
											assign node537 = (inp[12]) ? 1'b0 : 1'b1;
										assign node540 = (inp[9]) ? 1'b0 : node541;
											assign node541 = (inp[4]) ? 1'b0 : 1'b1;
								assign node545 = (inp[7]) ? node557 : node546;
									assign node546 = (inp[4]) ? node552 : node547;
										assign node547 = (inp[12]) ? node549 : 1'b1;
											assign node549 = (inp[3]) ? 1'b0 : 1'b1;
										assign node552 = (inp[3]) ? 1'b0 : node553;
											assign node553 = (inp[0]) ? 1'b0 : 1'b1;
									assign node557 = (inp[12]) ? 1'b0 : node558;
										assign node558 = (inp[4]) ? 1'b0 : node559;
											assign node559 = (inp[3]) ? 1'b0 : 1'b1;
					assign node564 = (inp[3]) ? node632 : node565;
						assign node565 = (inp[4]) ? node595 : node566;
							assign node566 = (inp[7]) ? node576 : node567;
								assign node567 = (inp[9]) ? node569 : 1'b1;
									assign node569 = (inp[1]) ? node571 : 1'b1;
										assign node571 = (inp[6]) ? node573 : 1'b1;
											assign node573 = (inp[12]) ? 1'b0 : 1'b1;
								assign node576 = (inp[9]) ? node584 : node577;
									assign node577 = (inp[1]) ? node579 : 1'b1;
										assign node579 = (inp[8]) ? node581 : 1'b1;
											assign node581 = (inp[12]) ? 1'b0 : 1'b1;
									assign node584 = (inp[12]) ? node590 : node585;
										assign node585 = (inp[6]) ? node587 : 1'b1;
											assign node587 = (inp[8]) ? 1'b0 : 1'b1;
										assign node590 = (inp[8]) ? 1'b0 : node591;
											assign node591 = (inp[0]) ? 1'b0 : 1'b1;
							assign node595 = (inp[9]) ? node615 : node596;
								assign node596 = (inp[1]) ? node604 : node597;
									assign node597 = (inp[6]) ? node599 : 1'b1;
										assign node599 = (inp[8]) ? node601 : 1'b1;
											assign node601 = (inp[12]) ? 1'b0 : 1'b1;
									assign node604 = (inp[12]) ? node610 : node605;
										assign node605 = (inp[7]) ? node607 : 1'b1;
											assign node607 = (inp[8]) ? 1'b0 : 1'b1;
										assign node610 = (inp[0]) ? 1'b0 : node611;
											assign node611 = (inp[7]) ? 1'b0 : 1'b1;
								assign node615 = (inp[0]) ? node627 : node616;
									assign node616 = (inp[7]) ? node622 : node617;
										assign node617 = (inp[8]) ? node619 : 1'b1;
											assign node619 = (inp[12]) ? 1'b0 : 1'b1;
										assign node622 = (inp[6]) ? 1'b0 : node623;
											assign node623 = (inp[8]) ? 1'b0 : 1'b1;
									assign node627 = (inp[1]) ? 1'b0 : node628;
										assign node628 = (inp[6]) ? 1'b0 : 1'b1;
						assign node632 = (inp[12]) ? node674 : node633;
							assign node633 = (inp[6]) ? node655 : node634;
								assign node634 = (inp[0]) ? node644 : node635;
									assign node635 = (inp[7]) ? node637 : 1'b1;
										assign node637 = (inp[4]) ? node641 : node638;
											assign node638 = (inp[8]) ? 1'b1 : 1'b1;
											assign node641 = (inp[8]) ? 1'b0 : 1'b1;
									assign node644 = (inp[1]) ? node650 : node645;
										assign node645 = (inp[8]) ? node647 : 1'b1;
											assign node647 = (inp[9]) ? 1'b0 : 1'b1;
										assign node650 = (inp[9]) ? 1'b0 : node651;
											assign node651 = (inp[4]) ? 1'b0 : 1'b1;
								assign node655 = (inp[1]) ? node667 : node656;
									assign node656 = (inp[0]) ? node662 : node657;
										assign node657 = (inp[4]) ? node659 : 1'b1;
											assign node659 = (inp[7]) ? 1'b0 : 1'b1;
										assign node662 = (inp[7]) ? 1'b0 : node663;
											assign node663 = (inp[4]) ? 1'b0 : 1'b1;
									assign node667 = (inp[8]) ? 1'b0 : node668;
										assign node668 = (inp[7]) ? 1'b0 : node669;
											assign node669 = (inp[0]) ? 1'b0 : 1'b1;
							assign node674 = (inp[7]) ? node696 : node675;
								assign node675 = (inp[4]) ? node687 : node676;
									assign node676 = (inp[6]) ? node682 : node677;
										assign node677 = (inp[0]) ? node679 : 1'b1;
											assign node679 = (inp[8]) ? 1'b0 : 1'b1;
										assign node682 = (inp[9]) ? 1'b0 : node683;
											assign node683 = (inp[0]) ? 1'b0 : 1'b1;
									assign node687 = (inp[9]) ? 1'b0 : node688;
										assign node688 = (inp[6]) ? node692 : node689;
											assign node689 = (inp[1]) ? 1'b0 : 1'b1;
											assign node692 = (inp[0]) ? 1'b0 : 1'b0;
								assign node696 = (inp[1]) ? 1'b0 : node697;
									assign node697 = (inp[8]) ? 1'b0 : node698;
										assign node698 = (inp[6]) ? 1'b0 : node699;
											assign node699 = (inp[0]) ? 1'b0 : 1'b1;
				assign node705 = (inp[0]) ? node845 : node706;
					assign node706 = (inp[12]) ? node776 : node707;
						assign node707 = (inp[9]) ? node737 : node708;
							assign node708 = (inp[1]) ? node718 : node709;
								assign node709 = (inp[8]) ? node711 : 1'b1;
									assign node711 = (inp[7]) ? node713 : 1'b1;
										assign node713 = (inp[6]) ? node715 : 1'b1;
											assign node715 = (inp[3]) ? 1'b0 : 1'b1;
								assign node718 = (inp[6]) ? node726 : node719;
									assign node719 = (inp[7]) ? node721 : 1'b1;
										assign node721 = (inp[3]) ? node723 : 1'b1;
											assign node723 = (inp[4]) ? 1'b0 : 1'b1;
									assign node726 = (inp[4]) ? node732 : node727;
										assign node727 = (inp[7]) ? node729 : 1'b1;
											assign node729 = (inp[5]) ? 1'b0 : 1'b1;
										assign node732 = (inp[5]) ? 1'b0 : node733;
											assign node733 = (inp[7]) ? 1'b0 : 1'b1;
							assign node737 = (inp[3]) ? node757 : node738;
								assign node738 = (inp[7]) ? node746 : node739;
									assign node739 = (inp[4]) ? node741 : 1'b1;
										assign node741 = (inp[1]) ? node743 : 1'b1;
											assign node743 = (inp[6]) ? 1'b0 : 1'b1;
									assign node746 = (inp[5]) ? node752 : node747;
										assign node747 = (inp[4]) ? node749 : 1'b1;
											assign node749 = (inp[8]) ? 1'b0 : 1'b1;
										assign node752 = (inp[6]) ? 1'b0 : node753;
											assign node753 = (inp[4]) ? 1'b0 : 1'b1;
								assign node757 = (inp[5]) ? node769 : node758;
									assign node758 = (inp[1]) ? node764 : node759;
										assign node759 = (inp[6]) ? node761 : 1'b1;
											assign node761 = (inp[7]) ? 1'b0 : 1'b1;
										assign node764 = (inp[6]) ? 1'b0 : node765;
											assign node765 = (inp[7]) ? 1'b0 : 1'b1;
									assign node769 = (inp[8]) ? 1'b0 : node770;
										assign node770 = (inp[4]) ? 1'b0 : node771;
											assign node771 = (inp[7]) ? 1'b0 : 1'b1;
						assign node776 = (inp[4]) ? node816 : node777;
							assign node777 = (inp[3]) ? node797 : node778;
								assign node778 = (inp[8]) ? node786 : node779;
									assign node779 = (inp[7]) ? node781 : 1'b1;
										assign node781 = (inp[1]) ? node783 : 1'b1;
											assign node783 = (inp[9]) ? 1'b0 : 1'b1;
									assign node786 = (inp[5]) ? node792 : node787;
										assign node787 = (inp[9]) ? node789 : 1'b1;
											assign node789 = (inp[6]) ? 1'b0 : 1'b1;
										assign node792 = (inp[1]) ? 1'b0 : node793;
											assign node793 = (inp[9]) ? 1'b0 : 1'b1;
								assign node797 = (inp[5]) ? node809 : node798;
									assign node798 = (inp[9]) ? node804 : node799;
										assign node799 = (inp[1]) ? node801 : 1'b1;
											assign node801 = (inp[8]) ? 1'b0 : 1'b1;
										assign node804 = (inp[6]) ? 1'b0 : node805;
											assign node805 = (inp[7]) ? 1'b0 : 1'b1;
									assign node809 = (inp[9]) ? 1'b0 : node810;
										assign node810 = (inp[6]) ? 1'b0 : node811;
											assign node811 = (inp[7]) ? 1'b0 : 1'b1;
							assign node816 = (inp[5]) ? node836 : node817;
								assign node817 = (inp[7]) ? node829 : node818;
									assign node818 = (inp[3]) ? node824 : node819;
										assign node819 = (inp[9]) ? node821 : 1'b1;
											assign node821 = (inp[6]) ? 1'b0 : 1'b1;
										assign node824 = (inp[1]) ? 1'b0 : node825;
											assign node825 = (inp[6]) ? 1'b0 : 1'b1;
									assign node829 = (inp[9]) ? 1'b0 : node830;
										assign node830 = (inp[1]) ? 1'b0 : node831;
											assign node831 = (inp[3]) ? 1'b0 : 1'b1;
								assign node836 = (inp[6]) ? 1'b0 : node837;
									assign node837 = (inp[9]) ? 1'b0 : node838;
										assign node838 = (inp[3]) ? 1'b0 : node839;
											assign node839 = (inp[8]) ? 1'b0 : 1'b1;
					assign node845 = (inp[6]) ? node919 : node846;
						assign node846 = (inp[4]) ? node888 : node847;
							assign node847 = (inp[9]) ? node867 : node848;
								assign node848 = (inp[8]) ? node856 : node849;
									assign node849 = (inp[1]) ? node851 : 1'b1;
										assign node851 = (inp[12]) ? node853 : 1'b1;
											assign node853 = (inp[3]) ? 1'b0 : 1'b1;
									assign node856 = (inp[7]) ? node862 : node857;
										assign node857 = (inp[1]) ? node859 : 1'b1;
											assign node859 = (inp[5]) ? 1'b0 : 1'b1;
										assign node862 = (inp[3]) ? 1'b0 : node863;
											assign node863 = (inp[5]) ? 1'b0 : 1'b1;
								assign node867 = (inp[1]) ? node879 : node868;
									assign node868 = (inp[3]) ? node874 : node869;
										assign node869 = (inp[7]) ? node871 : 1'b1;
											assign node871 = (inp[12]) ? 1'b0 : 1'b1;
										assign node874 = (inp[7]) ? 1'b0 : node875;
											assign node875 = (inp[8]) ? 1'b0 : 1'b1;
									assign node879 = (inp[12]) ? 1'b0 : node880;
										assign node880 = (inp[7]) ? node884 : node881;
											assign node881 = (inp[5]) ? 1'b0 : 1'b1;
											assign node884 = (inp[5]) ? 1'b0 : 1'b0;
							assign node888 = (inp[8]) ? node910 : node889;
								assign node889 = (inp[7]) ? node901 : node890;
									assign node890 = (inp[5]) ? node896 : node891;
										assign node891 = (inp[1]) ? node893 : 1'b1;
											assign node893 = (inp[9]) ? 1'b0 : 1'b1;
										assign node896 = (inp[3]) ? 1'b0 : node897;
											assign node897 = (inp[9]) ? 1'b0 : 1'b1;
									assign node901 = (inp[5]) ? 1'b0 : node902;
										assign node902 = (inp[1]) ? node906 : node903;
											assign node903 = (inp[9]) ? 1'b0 : 1'b1;
											assign node906 = (inp[12]) ? 1'b0 : 1'b0;
								assign node910 = (inp[7]) ? 1'b0 : node911;
									assign node911 = (inp[5]) ? 1'b0 : node912;
										assign node912 = (inp[1]) ? 1'b0 : node913;
											assign node913 = (inp[3]) ? 1'b0 : 1'b1;
						assign node919 = (inp[12]) ? node949 : node920;
							assign node920 = (inp[1]) ? node940 : node921;
								assign node921 = (inp[9]) ? node933 : node922;
									assign node922 = (inp[7]) ? node928 : node923;
										assign node923 = (inp[8]) ? node925 : 1'b1;
											assign node925 = (inp[5]) ? 1'b0 : 1'b1;
										assign node928 = (inp[4]) ? 1'b0 : node929;
											assign node929 = (inp[5]) ? 1'b0 : 1'b1;
									assign node933 = (inp[4]) ? 1'b0 : node934;
										assign node934 = (inp[3]) ? 1'b0 : node935;
											assign node935 = (inp[8]) ? 1'b0 : 1'b1;
								assign node940 = (inp[8]) ? 1'b0 : node941;
									assign node941 = (inp[3]) ? 1'b0 : node942;
										assign node942 = (inp[7]) ? 1'b0 : node943;
											assign node943 = (inp[5]) ? 1'b0 : 1'b1;
							assign node949 = (inp[5]) ? 1'b0 : node950;
								assign node950 = (inp[4]) ? 1'b0 : node951;
									assign node951 = (inp[3]) ? 1'b0 : node952;
										assign node952 = (inp[1]) ? 1'b0 : node953;
											assign node953 = (inp[8]) ? 1'b0 : 1'b1;
		assign node960 = (inp[12]) ? node1480 : node961;
			assign node961 = (inp[8]) ? node1223 : node962;
				assign node962 = (inp[10]) ? node1074 : node963;
					assign node963 = (inp[4]) ? node1005 : node964;
						assign node964 = (inp[9]) ? node976 : node965;
							assign node965 = (inp[7]) ? node967 : 1'b1;
								assign node967 = (inp[1]) ? node969 : 1'b1;
									assign node969 = (inp[0]) ? node971 : 1'b1;
										assign node971 = (inp[5]) ? node973 : 1'b1;
											assign node973 = (inp[2]) ? 1'b0 : 1'b1;
							assign node976 = (inp[6]) ? node986 : node977;
								assign node977 = (inp[1]) ? node979 : 1'b1;
									assign node979 = (inp[3]) ? node981 : 1'b1;
										assign node981 = (inp[5]) ? node983 : 1'b1;
											assign node983 = (inp[0]) ? 1'b0 : 1'b1;
								assign node986 = (inp[2]) ? node994 : node987;
									assign node987 = (inp[1]) ? node989 : 1'b1;
										assign node989 = (inp[5]) ? node991 : 1'b1;
											assign node991 = (inp[0]) ? 1'b0 : 1'b1;
									assign node994 = (inp[0]) ? node1000 : node995;
										assign node995 = (inp[3]) ? node997 : 1'b1;
											assign node997 = (inp[5]) ? 1'b0 : 1'b1;
										assign node1000 = (inp[7]) ? 1'b0 : node1001;
											assign node1001 = (inp[1]) ? 1'b0 : 1'b1;
						assign node1005 = (inp[1]) ? node1035 : node1006;
							assign node1006 = (inp[7]) ? node1016 : node1007;
								assign node1007 = (inp[0]) ? node1009 : 1'b1;
									assign node1009 = (inp[2]) ? node1011 : 1'b1;
										assign node1011 = (inp[5]) ? node1013 : 1'b1;
											assign node1013 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1016 = (inp[6]) ? node1024 : node1017;
									assign node1017 = (inp[2]) ? node1019 : 1'b1;
										assign node1019 = (inp[3]) ? node1021 : 1'b1;
											assign node1021 = (inp[0]) ? 1'b0 : 1'b0;
									assign node1024 = (inp[0]) ? node1030 : node1025;
										assign node1025 = (inp[2]) ? node1027 : 1'b1;
											assign node1027 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1030 = (inp[2]) ? 1'b0 : node1031;
											assign node1031 = (inp[9]) ? 1'b0 : 1'b1;
							assign node1035 = (inp[9]) ? node1055 : node1036;
								assign node1036 = (inp[3]) ? node1044 : node1037;
									assign node1037 = (inp[5]) ? node1039 : 1'b1;
										assign node1039 = (inp[6]) ? node1041 : 1'b1;
											assign node1041 = (inp[0]) ? 1'b0 : 1'b1;
									assign node1044 = (inp[6]) ? node1050 : node1045;
										assign node1045 = (inp[7]) ? node1047 : 1'b1;
											assign node1047 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1050 = (inp[2]) ? 1'b0 : node1051;
											assign node1051 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1055 = (inp[2]) ? node1067 : node1056;
									assign node1056 = (inp[5]) ? node1062 : node1057;
										assign node1057 = (inp[7]) ? node1059 : 1'b1;
											assign node1059 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1062 = (inp[6]) ? 1'b0 : node1063;
											assign node1063 = (inp[0]) ? 1'b0 : 1'b1;
									assign node1067 = (inp[0]) ? 1'b0 : node1068;
										assign node1068 = (inp[5]) ? 1'b0 : node1069;
											assign node1069 = (inp[6]) ? 1'b0 : 1'b1;
					assign node1074 = (inp[3]) ? node1154 : node1075;
						assign node1075 = (inp[0]) ? node1111 : node1076;
							assign node1076 = (inp[4]) ? node1086 : node1077;
								assign node1077 = (inp[5]) ? node1079 : 1'b1;
									assign node1079 = (inp[2]) ? node1081 : 1'b1;
										assign node1081 = (inp[1]) ? node1083 : 1'b1;
											assign node1083 = (inp[6]) ? 1'b0 : 1'b1;
								assign node1086 = (inp[1]) ? node1100 : node1087;
									assign node1087 = (inp[2]) ? node1093 : node1088;
										assign node1088 = (inp[7]) ? node1090 : 1'b1;
											assign node1090 = (inp[6]) ? 1'b1 : 1'b1;
										assign node1093 = (inp[6]) ? node1097 : node1094;
											assign node1094 = (inp[5]) ? 1'b1 : 1'b1;
											assign node1097 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1100 = (inp[7]) ? node1106 : node1101;
										assign node1101 = (inp[5]) ? node1103 : 1'b1;
											assign node1103 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1106 = (inp[6]) ? 1'b0 : node1107;
											assign node1107 = (inp[5]) ? 1'b0 : 1'b1;
							assign node1111 = (inp[5]) ? node1135 : node1112;
								assign node1112 = (inp[9]) ? node1122 : node1113;
									assign node1113 = (inp[6]) ? node1115 : 1'b1;
										assign node1115 = (inp[1]) ? node1119 : node1116;
											assign node1116 = (inp[7]) ? 1'b1 : 1'b1;
											assign node1119 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1122 = (inp[7]) ? node1130 : node1123;
										assign node1123 = (inp[2]) ? node1127 : node1124;
											assign node1124 = (inp[1]) ? 1'b1 : 1'b1;
											assign node1127 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1130 = (inp[4]) ? 1'b0 : node1131;
											assign node1131 = (inp[1]) ? 1'b0 : 1'b0;
								assign node1135 = (inp[2]) ? node1147 : node1136;
									assign node1136 = (inp[1]) ? node1142 : node1137;
										assign node1137 = (inp[4]) ? node1139 : 1'b1;
											assign node1139 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1142 = (inp[6]) ? 1'b0 : node1143;
											assign node1143 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1147 = (inp[7]) ? 1'b0 : node1148;
										assign node1148 = (inp[9]) ? 1'b0 : node1149;
											assign node1149 = (inp[4]) ? 1'b0 : 1'b1;
						assign node1154 = (inp[2]) ? node1194 : node1155;
							assign node1155 = (inp[9]) ? node1175 : node1156;
								assign node1156 = (inp[7]) ? node1164 : node1157;
									assign node1157 = (inp[4]) ? node1159 : 1'b1;
										assign node1159 = (inp[0]) ? node1161 : 1'b1;
											assign node1161 = (inp[5]) ? 1'b0 : 1'b0;
									assign node1164 = (inp[1]) ? node1170 : node1165;
										assign node1165 = (inp[4]) ? node1167 : 1'b1;
											assign node1167 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1170 = (inp[6]) ? 1'b0 : node1171;
											assign node1171 = (inp[0]) ? 1'b0 : 1'b1;
								assign node1175 = (inp[0]) ? node1187 : node1176;
									assign node1176 = (inp[4]) ? node1182 : node1177;
										assign node1177 = (inp[5]) ? node1179 : 1'b1;
											assign node1179 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1182 = (inp[1]) ? 1'b0 : node1183;
											assign node1183 = (inp[6]) ? 1'b0 : 1'b1;
									assign node1187 = (inp[7]) ? 1'b0 : node1188;
										assign node1188 = (inp[1]) ? 1'b0 : node1189;
											assign node1189 = (inp[6]) ? 1'b0 : 1'b1;
							assign node1194 = (inp[9]) ? node1214 : node1195;
								assign node1195 = (inp[6]) ? node1207 : node1196;
									assign node1196 = (inp[4]) ? node1202 : node1197;
										assign node1197 = (inp[5]) ? node1199 : 1'b1;
											assign node1199 = (inp[1]) ? 1'b0 : 1'b1;
										assign node1202 = (inp[7]) ? 1'b0 : node1203;
											assign node1203 = (inp[1]) ? 1'b0 : 1'b1;
									assign node1207 = (inp[7]) ? 1'b0 : node1208;
										assign node1208 = (inp[5]) ? 1'b0 : node1209;
											assign node1209 = (inp[1]) ? 1'b0 : 1'b1;
								assign node1214 = (inp[4]) ? 1'b0 : node1215;
									assign node1215 = (inp[6]) ? 1'b0 : node1216;
										assign node1216 = (inp[1]) ? 1'b0 : node1217;
											assign node1217 = (inp[0]) ? 1'b0 : 1'b1;
				assign node1223 = (inp[5]) ? node1369 : node1224;
					assign node1224 = (inp[3]) ? node1294 : node1225;
						assign node1225 = (inp[0]) ? node1255 : node1226;
							assign node1226 = (inp[1]) ? node1236 : node1227;
								assign node1227 = (inp[4]) ? node1229 : 1'b1;
									assign node1229 = (inp[10]) ? node1231 : 1'b1;
										assign node1231 = (inp[9]) ? node1233 : 1'b1;
											assign node1233 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1236 = (inp[9]) ? node1244 : node1237;
									assign node1237 = (inp[7]) ? node1239 : 1'b1;
										assign node1239 = (inp[2]) ? node1241 : 1'b1;
											assign node1241 = (inp[4]) ? 1'b0 : 1'b1;
									assign node1244 = (inp[6]) ? node1250 : node1245;
										assign node1245 = (inp[4]) ? node1247 : 1'b1;
											assign node1247 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1250 = (inp[2]) ? 1'b0 : node1251;
											assign node1251 = (inp[10]) ? 1'b0 : 1'b1;
							assign node1255 = (inp[4]) ? node1275 : node1256;
								assign node1256 = (inp[2]) ? node1264 : node1257;
									assign node1257 = (inp[6]) ? node1259 : 1'b1;
										assign node1259 = (inp[1]) ? node1261 : 1'b1;
											assign node1261 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1264 = (inp[9]) ? node1270 : node1265;
										assign node1265 = (inp[1]) ? node1267 : 1'b1;
											assign node1267 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1270 = (inp[1]) ? 1'b0 : node1271;
											assign node1271 = (inp[6]) ? 1'b0 : 1'b1;
								assign node1275 = (inp[1]) ? node1287 : node1276;
									assign node1276 = (inp[10]) ? node1282 : node1277;
										assign node1277 = (inp[6]) ? node1279 : 1'b1;
											assign node1279 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1282 = (inp[7]) ? 1'b0 : node1283;
											assign node1283 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1287 = (inp[6]) ? 1'b0 : node1288;
										assign node1288 = (inp[9]) ? 1'b0 : node1289;
											assign node1289 = (inp[2]) ? 1'b0 : 1'b1;
						assign node1294 = (inp[1]) ? node1340 : node1295;
							assign node1295 = (inp[4]) ? node1319 : node1296;
								assign node1296 = (inp[7]) ? node1304 : node1297;
									assign node1297 = (inp[6]) ? node1299 : 1'b1;
										assign node1299 = (inp[9]) ? node1301 : 1'b1;
											assign node1301 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1304 = (inp[6]) ? node1312 : node1305;
										assign node1305 = (inp[9]) ? node1309 : node1306;
											assign node1306 = (inp[2]) ? 1'b1 : 1'b1;
											assign node1309 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1312 = (inp[0]) ? node1316 : node1313;
											assign node1313 = (inp[9]) ? 1'b0 : 1'b1;
											assign node1316 = (inp[2]) ? 1'b0 : 1'b0;
								assign node1319 = (inp[2]) ? node1333 : node1320;
									assign node1320 = (inp[9]) ? node1326 : node1321;
										assign node1321 = (inp[7]) ? node1323 : 1'b1;
											assign node1323 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1326 = (inp[0]) ? node1330 : node1327;
											assign node1327 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1330 = (inp[7]) ? 1'b0 : 1'b0;
									assign node1333 = (inp[10]) ? 1'b0 : node1334;
										assign node1334 = (inp[0]) ? 1'b0 : node1335;
											assign node1335 = (inp[6]) ? 1'b0 : 1'b1;
							assign node1340 = (inp[2]) ? node1360 : node1341;
								assign node1341 = (inp[6]) ? node1353 : node1342;
									assign node1342 = (inp[4]) ? node1348 : node1343;
										assign node1343 = (inp[10]) ? node1345 : 1'b1;
											assign node1345 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1348 = (inp[0]) ? 1'b0 : node1349;
											assign node1349 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1353 = (inp[7]) ? 1'b0 : node1354;
										assign node1354 = (inp[0]) ? 1'b0 : node1355;
											assign node1355 = (inp[4]) ? 1'b0 : 1'b1;
								assign node1360 = (inp[0]) ? 1'b0 : node1361;
									assign node1361 = (inp[10]) ? 1'b0 : node1362;
										assign node1362 = (inp[4]) ? 1'b0 : node1363;
											assign node1363 = (inp[9]) ? 1'b0 : 1'b1;
					assign node1369 = (inp[7]) ? node1441 : node1370;
						assign node1370 = (inp[2]) ? node1412 : node1371;
							assign node1371 = (inp[4]) ? node1393 : node1372;
								assign node1372 = (inp[9]) ? node1382 : node1373;
									assign node1373 = (inp[10]) ? node1375 : 1'b1;
										assign node1375 = (inp[6]) ? node1379 : node1376;
											assign node1376 = (inp[0]) ? 1'b1 : 1'b1;
											assign node1379 = (inp[1]) ? 1'b0 : 1'b1;
									assign node1382 = (inp[6]) ? node1388 : node1383;
										assign node1383 = (inp[3]) ? node1385 : 1'b1;
											assign node1385 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1388 = (inp[0]) ? 1'b0 : node1389;
											assign node1389 = (inp[1]) ? 1'b0 : 1'b1;
								assign node1393 = (inp[1]) ? node1405 : node1394;
									assign node1394 = (inp[10]) ? node1400 : node1395;
										assign node1395 = (inp[3]) ? node1397 : 1'b1;
											assign node1397 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1400 = (inp[6]) ? 1'b0 : node1401;
											assign node1401 = (inp[0]) ? 1'b0 : 1'b1;
									assign node1405 = (inp[10]) ? 1'b0 : node1406;
										assign node1406 = (inp[9]) ? 1'b0 : node1407;
											assign node1407 = (inp[0]) ? 1'b0 : 1'b1;
							assign node1412 = (inp[9]) ? node1432 : node1413;
								assign node1413 = (inp[3]) ? node1425 : node1414;
									assign node1414 = (inp[1]) ? node1420 : node1415;
										assign node1415 = (inp[10]) ? node1417 : 1'b1;
											assign node1417 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1420 = (inp[10]) ? 1'b0 : node1421;
											assign node1421 = (inp[4]) ? 1'b0 : 1'b1;
									assign node1425 = (inp[6]) ? 1'b0 : node1426;
										assign node1426 = (inp[1]) ? 1'b0 : node1427;
											assign node1427 = (inp[0]) ? 1'b0 : 1'b1;
								assign node1432 = (inp[0]) ? 1'b0 : node1433;
									assign node1433 = (inp[10]) ? 1'b0 : node1434;
										assign node1434 = (inp[6]) ? 1'b0 : node1435;
											assign node1435 = (inp[1]) ? 1'b0 : 1'b1;
						assign node1441 = (inp[0]) ? node1471 : node1442;
							assign node1442 = (inp[4]) ? node1462 : node1443;
								assign node1443 = (inp[9]) ? node1455 : node1444;
									assign node1444 = (inp[10]) ? node1450 : node1445;
										assign node1445 = (inp[6]) ? node1447 : 1'b1;
											assign node1447 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1450 = (inp[1]) ? 1'b0 : node1451;
											assign node1451 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1455 = (inp[3]) ? 1'b0 : node1456;
										assign node1456 = (inp[6]) ? 1'b0 : node1457;
											assign node1457 = (inp[1]) ? 1'b0 : 1'b1;
								assign node1462 = (inp[2]) ? 1'b0 : node1463;
									assign node1463 = (inp[6]) ? 1'b0 : node1464;
										assign node1464 = (inp[10]) ? 1'b0 : node1465;
											assign node1465 = (inp[9]) ? 1'b0 : 1'b1;
							assign node1471 = (inp[3]) ? 1'b0 : node1472;
								assign node1472 = (inp[2]) ? 1'b0 : node1473;
									assign node1473 = (inp[6]) ? 1'b0 : node1474;
										assign node1474 = (inp[4]) ? 1'b0 : 1'b1;
			assign node1480 = (inp[10]) ? node1740 : node1481;
				assign node1481 = (inp[1]) ? node1625 : node1482;
					assign node1482 = (inp[3]) ? node1554 : node1483;
						assign node1483 = (inp[5]) ? node1513 : node1484;
							assign node1484 = (inp[2]) ? node1494 : node1485;
								assign node1485 = (inp[9]) ? node1487 : 1'b1;
									assign node1487 = (inp[8]) ? node1489 : 1'b1;
										assign node1489 = (inp[6]) ? node1491 : 1'b1;
											assign node1491 = (inp[4]) ? 1'b0 : 1'b0;
								assign node1494 = (inp[7]) ? node1502 : node1495;
									assign node1495 = (inp[8]) ? node1497 : 1'b1;
										assign node1497 = (inp[6]) ? node1499 : 1'b1;
											assign node1499 = (inp[0]) ? 1'b0 : 1'b1;
									assign node1502 = (inp[8]) ? node1508 : node1503;
										assign node1503 = (inp[9]) ? node1505 : 1'b1;
											assign node1505 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1508 = (inp[0]) ? 1'b0 : node1509;
											assign node1509 = (inp[6]) ? 1'b0 : 1'b0;
							assign node1513 = (inp[4]) ? node1535 : node1514;
								assign node1514 = (inp[8]) ? node1522 : node1515;
									assign node1515 = (inp[9]) ? node1517 : 1'b1;
										assign node1517 = (inp[7]) ? node1519 : 1'b1;
											assign node1519 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1522 = (inp[7]) ? node1528 : node1523;
										assign node1523 = (inp[6]) ? node1525 : 1'b1;
											assign node1525 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1528 = (inp[2]) ? node1532 : node1529;
											assign node1529 = (inp[0]) ? 1'b0 : 1'b1;
											assign node1532 = (inp[6]) ? 1'b0 : 1'b0;
								assign node1535 = (inp[8]) ? node1547 : node1536;
									assign node1536 = (inp[9]) ? node1542 : node1537;
										assign node1537 = (inp[6]) ? node1539 : 1'b1;
											assign node1539 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1542 = (inp[7]) ? 1'b0 : node1543;
											assign node1543 = (inp[6]) ? 1'b0 : 1'b1;
									assign node1547 = (inp[2]) ? 1'b0 : node1548;
										assign node1548 = (inp[9]) ? 1'b0 : node1549;
											assign node1549 = (inp[6]) ? 1'b0 : 1'b1;
						assign node1554 = (inp[4]) ? node1594 : node1555;
							assign node1555 = (inp[9]) ? node1575 : node1556;
								assign node1556 = (inp[7]) ? node1564 : node1557;
									assign node1557 = (inp[0]) ? node1559 : 1'b1;
										assign node1559 = (inp[6]) ? 1'b0 : node1560;
											assign node1560 = (inp[2]) ? 1'b1 : 1'b1;
									assign node1564 = (inp[5]) ? node1570 : node1565;
										assign node1565 = (inp[6]) ? node1567 : 1'b1;
											assign node1567 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1570 = (inp[2]) ? 1'b0 : node1571;
											assign node1571 = (inp[0]) ? 1'b0 : 1'b1;
								assign node1575 = (inp[8]) ? node1587 : node1576;
									assign node1576 = (inp[2]) ? node1582 : node1577;
										assign node1577 = (inp[0]) ? node1579 : 1'b1;
											assign node1579 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1582 = (inp[0]) ? 1'b0 : node1583;
											assign node1583 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1587 = (inp[7]) ? 1'b0 : node1588;
										assign node1588 = (inp[2]) ? 1'b0 : node1589;
											assign node1589 = (inp[0]) ? 1'b0 : 1'b1;
							assign node1594 = (inp[7]) ? node1616 : node1595;
								assign node1595 = (inp[0]) ? node1607 : node1596;
									assign node1596 = (inp[9]) ? node1602 : node1597;
										assign node1597 = (inp[2]) ? node1599 : 1'b1;
											assign node1599 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1602 = (inp[5]) ? 1'b0 : node1603;
											assign node1603 = (inp[8]) ? 1'b0 : 1'b1;
									assign node1607 = (inp[6]) ? 1'b0 : node1608;
										assign node1608 = (inp[5]) ? node1612 : node1609;
											assign node1609 = (inp[8]) ? 1'b0 : 1'b1;
											assign node1612 = (inp[8]) ? 1'b0 : 1'b0;
								assign node1616 = (inp[5]) ? 1'b0 : node1617;
									assign node1617 = (inp[6]) ? 1'b0 : node1618;
										assign node1618 = (inp[9]) ? 1'b0 : node1619;
											assign node1619 = (inp[8]) ? 1'b0 : 1'b1;
					assign node1625 = (inp[6]) ? node1697 : node1626;
						assign node1626 = (inp[7]) ? node1668 : node1627;
							assign node1627 = (inp[9]) ? node1647 : node1628;
								assign node1628 = (inp[4]) ? node1636 : node1629;
									assign node1629 = (inp[8]) ? node1631 : 1'b1;
										assign node1631 = (inp[5]) ? node1633 : 1'b1;
											assign node1633 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1636 = (inp[5]) ? node1642 : node1637;
										assign node1637 = (inp[2]) ? node1639 : 1'b1;
											assign node1639 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1642 = (inp[2]) ? 1'b0 : node1643;
											assign node1643 = (inp[3]) ? 1'b0 : 1'b1;
								assign node1647 = (inp[3]) ? node1661 : node1648;
									assign node1648 = (inp[4]) ? node1654 : node1649;
										assign node1649 = (inp[5]) ? node1651 : 1'b1;
											assign node1651 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1654 = (inp[2]) ? node1658 : node1655;
											assign node1655 = (inp[0]) ? 1'b0 : 1'b1;
											assign node1658 = (inp[0]) ? 1'b0 : 1'b0;
									assign node1661 = (inp[5]) ? 1'b0 : node1662;
										assign node1662 = (inp[2]) ? 1'b0 : node1663;
											assign node1663 = (inp[0]) ? 1'b0 : 1'b1;
							assign node1668 = (inp[8]) ? node1688 : node1669;
								assign node1669 = (inp[0]) ? node1681 : node1670;
									assign node1670 = (inp[2]) ? node1676 : node1671;
										assign node1671 = (inp[3]) ? node1673 : 1'b1;
											assign node1673 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1676 = (inp[4]) ? 1'b0 : node1677;
											assign node1677 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1681 = (inp[3]) ? 1'b0 : node1682;
										assign node1682 = (inp[5]) ? 1'b0 : node1683;
											assign node1683 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1688 = (inp[9]) ? 1'b0 : node1689;
									assign node1689 = (inp[3]) ? 1'b0 : node1690;
										assign node1690 = (inp[5]) ? 1'b0 : node1691;
											assign node1691 = (inp[2]) ? 1'b0 : 1'b1;
						assign node1697 = (inp[4]) ? node1729 : node1698;
							assign node1698 = (inp[0]) ? node1720 : node1699;
								assign node1699 = (inp[9]) ? node1713 : node1700;
									assign node1700 = (inp[8]) ? node1706 : node1701;
										assign node1701 = (inp[2]) ? node1703 : 1'b1;
											assign node1703 = (inp[5]) ? 1'b0 : 1'b1;
										assign node1706 = (inp[7]) ? node1710 : node1707;
											assign node1707 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1710 = (inp[5]) ? 1'b0 : 1'b0;
									assign node1713 = (inp[7]) ? 1'b0 : node1714;
										assign node1714 = (inp[3]) ? 1'b0 : node1715;
											assign node1715 = (inp[5]) ? 1'b0 : 1'b1;
								assign node1720 = (inp[7]) ? 1'b0 : node1721;
									assign node1721 = (inp[5]) ? 1'b0 : node1722;
										assign node1722 = (inp[3]) ? 1'b0 : node1723;
											assign node1723 = (inp[8]) ? 1'b0 : 1'b1;
							assign node1729 = (inp[3]) ? 1'b0 : node1730;
								assign node1730 = (inp[0]) ? 1'b0 : node1731;
									assign node1731 = (inp[9]) ? 1'b0 : node1732;
										assign node1732 = (inp[8]) ? 1'b0 : node1733;
											assign node1733 = (inp[7]) ? 1'b0 : 1'b1;
				assign node1740 = (inp[6]) ? node1860 : node1741;
					assign node1741 = (inp[5]) ? node1815 : node1742;
						assign node1742 = (inp[9]) ? node1784 : node1743;
							assign node1743 = (inp[2]) ? node1765 : node1744;
								assign node1744 = (inp[0]) ? node1752 : node1745;
									assign node1745 = (inp[1]) ? node1747 : 1'b1;
										assign node1747 = (inp[8]) ? node1749 : 1'b1;
											assign node1749 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1752 = (inp[8]) ? node1760 : node1753;
										assign node1753 = (inp[7]) ? node1757 : node1754;
											assign node1754 = (inp[4]) ? 1'b1 : 1'b1;
											assign node1757 = (inp[1]) ? 1'b0 : 1'b1;
										assign node1760 = (inp[7]) ? 1'b0 : node1761;
											assign node1761 = (inp[3]) ? 1'b0 : 1'b1;
								assign node1765 = (inp[4]) ? node1777 : node1766;
									assign node1766 = (inp[7]) ? node1772 : node1767;
										assign node1767 = (inp[3]) ? node1769 : 1'b1;
											assign node1769 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1772 = (inp[8]) ? 1'b0 : node1773;
											assign node1773 = (inp[0]) ? 1'b0 : 1'b1;
									assign node1777 = (inp[3]) ? 1'b0 : node1778;
										assign node1778 = (inp[7]) ? 1'b0 : node1779;
											assign node1779 = (inp[8]) ? 1'b0 : 1'b1;
							assign node1784 = (inp[3]) ? node1806 : node1785;
								assign node1785 = (inp[1]) ? node1797 : node1786;
									assign node1786 = (inp[7]) ? node1792 : node1787;
										assign node1787 = (inp[8]) ? node1789 : 1'b1;
											assign node1789 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1792 = (inp[4]) ? 1'b0 : node1793;
											assign node1793 = (inp[0]) ? 1'b0 : 1'b1;
									assign node1797 = (inp[4]) ? 1'b0 : node1798;
										assign node1798 = (inp[7]) ? node1802 : node1799;
											assign node1799 = (inp[8]) ? 1'b0 : 1'b1;
											assign node1802 = (inp[0]) ? 1'b0 : 1'b0;
								assign node1806 = (inp[0]) ? 1'b0 : node1807;
									assign node1807 = (inp[7]) ? 1'b0 : node1808;
										assign node1808 = (inp[1]) ? 1'b0 : node1809;
											assign node1809 = (inp[8]) ? 1'b0 : 1'b1;
						assign node1815 = (inp[3]) ? node1849 : node1816;
							assign node1816 = (inp[7]) ? node1838 : node1817;
								assign node1817 = (inp[4]) ? node1829 : node1818;
									assign node1818 = (inp[1]) ? node1824 : node1819;
										assign node1819 = (inp[8]) ? node1821 : 1'b1;
											assign node1821 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1824 = (inp[9]) ? 1'b0 : node1825;
											assign node1825 = (inp[8]) ? 1'b0 : 1'b1;
									assign node1829 = (inp[8]) ? 1'b0 : node1830;
										assign node1830 = (inp[1]) ? node1834 : node1831;
											assign node1831 = (inp[9]) ? 1'b0 : 1'b1;
											assign node1834 = (inp[9]) ? 1'b0 : 1'b0;
								assign node1838 = (inp[0]) ? 1'b0 : node1839;
									assign node1839 = (inp[8]) ? 1'b0 : node1840;
										assign node1840 = (inp[4]) ? node1844 : node1841;
											assign node1841 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1844 = (inp[1]) ? 1'b0 : 1'b0;
							assign node1849 = (inp[1]) ? 1'b0 : node1850;
								assign node1850 = (inp[4]) ? 1'b0 : node1851;
									assign node1851 = (inp[9]) ? 1'b0 : node1852;
										assign node1852 = (inp[2]) ? 1'b0 : node1853;
											assign node1853 = (inp[0]) ? 1'b0 : 1'b1;
					assign node1860 = (inp[8]) ? node1904 : node1861;
						assign node1861 = (inp[9]) ? node1893 : node1862;
							assign node1862 = (inp[5]) ? node1882 : node1863;
								assign node1863 = (inp[4]) ? node1875 : node1864;
									assign node1864 = (inp[2]) ? node1870 : node1865;
										assign node1865 = (inp[3]) ? node1867 : 1'b1;
											assign node1867 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1870 = (inp[1]) ? 1'b0 : node1871;
											assign node1871 = (inp[0]) ? 1'b0 : 1'b1;
									assign node1875 = (inp[1]) ? 1'b0 : node1876;
										assign node1876 = (inp[0]) ? 1'b0 : node1877;
											assign node1877 = (inp[3]) ? 1'b0 : 1'b1;
								assign node1882 = (inp[0]) ? 1'b0 : node1883;
									assign node1883 = (inp[1]) ? 1'b0 : node1884;
										assign node1884 = (inp[4]) ? node1888 : node1885;
											assign node1885 = (inp[2]) ? 1'b0 : 1'b1;
											assign node1888 = (inp[7]) ? 1'b0 : 1'b0;
							assign node1893 = (inp[2]) ? 1'b0 : node1894;
								assign node1894 = (inp[1]) ? 1'b0 : node1895;
									assign node1895 = (inp[3]) ? 1'b0 : node1896;
										assign node1896 = (inp[7]) ? 1'b0 : node1897;
											assign node1897 = (inp[4]) ? 1'b0 : 1'b1;
						assign node1904 = (inp[3]) ? 1'b0 : node1905;
							assign node1905 = (inp[5]) ? 1'b0 : node1906;
								assign node1906 = (inp[4]) ? 1'b0 : node1907;
									assign node1907 = (inp[1]) ? 1'b0 : node1908;
										assign node1908 = (inp[7]) ? 1'b0 : node1909;
											assign node1909 = (inp[2]) ? 1'b0 : 1'b1;

endmodule