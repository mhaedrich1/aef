module dtc_split05_bm14 (
	input  wire [13-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node5;
	wire [1-1:0] node7;
	wire [1-1:0] node8;
	wire [1-1:0] node10;
	wire [1-1:0] node13;
	wire [1-1:0] node16;
	wire [1-1:0] node17;
	wire [1-1:0] node19;
	wire [1-1:0] node21;
	wire [1-1:0] node22;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node29;
	wire [1-1:0] node30;
	wire [1-1:0] node32;
	wire [1-1:0] node36;
	wire [1-1:0] node37;
	wire [1-1:0] node41;
	wire [1-1:0] node42;
	wire [1-1:0] node43;
	wire [1-1:0] node45;
	wire [1-1:0] node48;
	wire [1-1:0] node49;
	wire [1-1:0] node51;
	wire [1-1:0] node55;
	wire [1-1:0] node56;
	wire [1-1:0] node57;
	wire [1-1:0] node59;
	wire [1-1:0] node62;
	wire [1-1:0] node63;
	wire [1-1:0] node66;
	wire [1-1:0] node67;
	wire [1-1:0] node71;
	wire [1-1:0] node72;
	wire [1-1:0] node73;
	wire [1-1:0] node75;
	wire [1-1:0] node78;
	wire [1-1:0] node79;
	wire [1-1:0] node84;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node87;
	wire [1-1:0] node89;
	wire [1-1:0] node91;
	wire [1-1:0] node92;
	wire [1-1:0] node94;
	wire [1-1:0] node98;
	wire [1-1:0] node99;
	wire [1-1:0] node101;
	wire [1-1:0] node102;
	wire [1-1:0] node105;
	wire [1-1:0] node106;
	wire [1-1:0] node110;
	wire [1-1:0] node111;
	wire [1-1:0] node114;
	wire [1-1:0] node115;
	wire [1-1:0] node116;
	wire [1-1:0] node121;
	wire [1-1:0] node122;
	wire [1-1:0] node124;
	wire [1-1:0] node126;
	wire [1-1:0] node127;
	wire [1-1:0] node131;
	wire [1-1:0] node132;
	wire [1-1:0] node133;
	wire [1-1:0] node136;
	wire [1-1:0] node137;
	wire [1-1:0] node142;
	wire [1-1:0] node143;
	wire [1-1:0] node144;
	wire [1-1:0] node145;
	wire [1-1:0] node147;
	wire [1-1:0] node148;
	wire [1-1:0] node152;
	wire [1-1:0] node153;
	wire [1-1:0] node154;
	wire [1-1:0] node155;
	wire [1-1:0] node157;
	wire [1-1:0] node163;
	wire [1-1:0] node164;
	wire [1-1:0] node165;
	wire [1-1:0] node166;
	wire [1-1:0] node168;
	wire [1-1:0] node174;
	wire [1-1:0] node175;
	wire [1-1:0] node176;
	wire [1-1:0] node177;
	wire [1-1:0] node178;
	wire [1-1:0] node181;
	wire [1-1:0] node182;
	wire [1-1:0] node186;
	wire [1-1:0] node187;

	assign outp = (inp[0]) ? node84 : node1;
		assign node1 = (inp[11]) ? node41 : node2;
			assign node2 = (inp[12]) ? node16 : node3;
				assign node3 = (inp[8]) ? node5 : 1'b1;
					assign node5 = (inp[10]) ? node7 : 1'b1;
						assign node7 = (inp[6]) ? node13 : node8;
							assign node8 = (inp[7]) ? node10 : 1'b1;
								assign node10 = (inp[1]) ? 1'b0 : 1'b1;
							assign node13 = (inp[2]) ? 1'b0 : 1'b1;
				assign node16 = (inp[8]) ? node26 : node17;
					assign node17 = (inp[9]) ? node19 : 1'b1;
						assign node19 = (inp[10]) ? node21 : 1'b1;
							assign node21 = (inp[7]) ? 1'b0 : node22;
								assign node22 = (inp[4]) ? 1'b0 : 1'b1;
					assign node26 = (inp[6]) ? node36 : node27;
						assign node27 = (inp[5]) ? node29 : 1'b1;
							assign node29 = (inp[9]) ? 1'b0 : node30;
								assign node30 = (inp[7]) ? node32 : 1'b1;
									assign node32 = (inp[10]) ? 1'b0 : 1'b1;
						assign node36 = (inp[1]) ? 1'b0 : node37;
							assign node37 = (inp[10]) ? 1'b0 : 1'b1;
			assign node41 = (inp[10]) ? node55 : node42;
				assign node42 = (inp[1]) ? node48 : node43;
					assign node43 = (inp[5]) ? node45 : 1'b1;
						assign node45 = (inp[4]) ? 1'b0 : 1'b1;
					assign node48 = (inp[12]) ? 1'b0 : node49;
						assign node49 = (inp[7]) ? node51 : 1'b1;
							assign node51 = (inp[9]) ? 1'b0 : 1'b1;
				assign node55 = (inp[2]) ? node71 : node56;
					assign node56 = (inp[5]) ? node62 : node57;
						assign node57 = (inp[9]) ? node59 : 1'b1;
							assign node59 = (inp[8]) ? 1'b0 : 1'b1;
						assign node62 = (inp[8]) ? node66 : node63;
							assign node63 = (inp[3]) ? 1'b0 : 1'b1;
							assign node66 = (inp[1]) ? 1'b0 : node67;
								assign node67 = (inp[4]) ? 1'b0 : 1'b1;
					assign node71 = (inp[5]) ? 1'b0 : node72;
						assign node72 = (inp[9]) ? node78 : node73;
							assign node73 = (inp[4]) ? node75 : 1'b1;
								assign node75 = (inp[8]) ? 1'b0 : 1'b1;
							assign node78 = (inp[7]) ? 1'b0 : node79;
								assign node79 = (inp[8]) ? 1'b0 : 1'b1;
		assign node84 = (inp[1]) ? node142 : node85;
			assign node85 = (inp[10]) ? node121 : node86;
				assign node86 = (inp[11]) ? node98 : node87;
					assign node87 = (inp[9]) ? node89 : 1'b1;
						assign node89 = (inp[5]) ? node91 : 1'b1;
							assign node91 = (inp[3]) ? 1'b0 : node92;
								assign node92 = (inp[12]) ? node94 : 1'b1;
									assign node94 = (inp[8]) ? 1'b0 : 1'b1;
					assign node98 = (inp[9]) ? node110 : node99;
						assign node99 = (inp[4]) ? node101 : 1'b1;
							assign node101 = (inp[5]) ? node105 : node102;
								assign node102 = (inp[2]) ? 1'b0 : 1'b1;
								assign node105 = (inp[7]) ? 1'b0 : node106;
									assign node106 = (inp[8]) ? 1'b0 : 1'b1;
						assign node110 = (inp[3]) ? node114 : node111;
							assign node111 = (inp[8]) ? 1'b0 : 1'b1;
							assign node114 = (inp[5]) ? 1'b0 : node115;
								assign node115 = (inp[2]) ? 1'b0 : node116;
									assign node116 = (inp[6]) ? 1'b0 : 1'b1;
				assign node121 = (inp[7]) ? node131 : node122;
					assign node122 = (inp[12]) ? node124 : 1'b1;
						assign node124 = (inp[8]) ? node126 : 1'b1;
							assign node126 = (inp[9]) ? 1'b0 : node127;
								assign node127 = (inp[2]) ? 1'b0 : 1'b1;
					assign node131 = (inp[9]) ? 1'b0 : node132;
						assign node132 = (inp[3]) ? node136 : node133;
							assign node133 = (inp[8]) ? 1'b0 : 1'b1;
							assign node136 = (inp[5]) ? 1'b0 : node137;
								assign node137 = (inp[6]) ? 1'b0 : 1'b1;
			assign node142 = (inp[3]) ? node174 : node143;
				assign node143 = (inp[9]) ? node163 : node144;
					assign node144 = (inp[11]) ? node152 : node145;
						assign node145 = (inp[4]) ? node147 : 1'b1;
							assign node147 = (inp[12]) ? 1'b0 : node148;
								assign node148 = (inp[2]) ? 1'b0 : 1'b1;
						assign node152 = (inp[2]) ? 1'b0 : node153;
							assign node153 = (inp[6]) ? 1'b0 : node154;
								assign node154 = (inp[8]) ? 1'b0 : node155;
									assign node155 = (inp[7]) ? node157 : 1'b1;
										assign node157 = (inp[4]) ? 1'b0 : 1'b1;
					assign node163 = (inp[12]) ? 1'b0 : node164;
						assign node164 = (inp[10]) ? 1'b0 : node165;
							assign node165 = (inp[6]) ? 1'b0 : node166;
								assign node166 = (inp[2]) ? node168 : 1'b1;
									assign node168 = (inp[8]) ? 1'b0 : 1'b1;
				assign node174 = (inp[2]) ? 1'b0 : node175;
					assign node175 = (inp[10]) ? 1'b0 : node176;
						assign node176 = (inp[12]) ? node186 : node177;
							assign node177 = (inp[8]) ? node181 : node178;
								assign node178 = (inp[6]) ? 1'b0 : 1'b1;
								assign node181 = (inp[4]) ? 1'b0 : node182;
									assign node182 = (inp[5]) ? 1'b0 : 1'b1;
							assign node186 = (inp[7]) ? 1'b0 : node187;
								assign node187 = (inp[5]) ? 1'b0 : 1'b1;

endmodule