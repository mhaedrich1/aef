module dtc_split05_bm62 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node13;
	wire [4-1:0] node17;
	wire [4-1:0] node18;
	wire [4-1:0] node20;
	wire [4-1:0] node23;
	wire [4-1:0] node24;
	wire [4-1:0] node28;
	wire [4-1:0] node29;
	wire [4-1:0] node30;
	wire [4-1:0] node31;
	wire [4-1:0] node34;
	wire [4-1:0] node38;
	wire [4-1:0] node39;
	wire [4-1:0] node40;
	wire [4-1:0] node43;
	wire [4-1:0] node46;
	wire [4-1:0] node47;
	wire [4-1:0] node50;
	wire [4-1:0] node53;
	wire [4-1:0] node54;
	wire [4-1:0] node55;
	wire [4-1:0] node57;
	wire [4-1:0] node58;
	wire [4-1:0] node62;
	wire [4-1:0] node63;
	wire [4-1:0] node64;
	wire [4-1:0] node68;
	wire [4-1:0] node69;
	wire [4-1:0] node72;
	wire [4-1:0] node75;
	wire [4-1:0] node76;
	wire [4-1:0] node77;
	wire [4-1:0] node79;
	wire [4-1:0] node82;
	wire [4-1:0] node83;
	wire [4-1:0] node86;
	wire [4-1:0] node89;
	wire [4-1:0] node90;
	wire [4-1:0] node91;
	wire [4-1:0] node95;
	wire [4-1:0] node97;
	wire [4-1:0] node100;
	wire [4-1:0] node101;
	wire [4-1:0] node102;
	wire [4-1:0] node103;
	wire [4-1:0] node104;
	wire [4-1:0] node105;
	wire [4-1:0] node108;
	wire [4-1:0] node111;
	wire [4-1:0] node112;
	wire [4-1:0] node115;
	wire [4-1:0] node118;
	wire [4-1:0] node119;
	wire [4-1:0] node122;
	wire [4-1:0] node123;
	wire [4-1:0] node126;
	wire [4-1:0] node129;
	wire [4-1:0] node130;
	wire [4-1:0] node131;
	wire [4-1:0] node132;
	wire [4-1:0] node135;
	wire [4-1:0] node138;
	wire [4-1:0] node139;
	wire [4-1:0] node142;
	wire [4-1:0] node145;
	wire [4-1:0] node146;
	wire [4-1:0] node147;
	wire [4-1:0] node150;
	wire [4-1:0] node153;
	wire [4-1:0] node154;
	wire [4-1:0] node157;
	wire [4-1:0] node160;
	wire [4-1:0] node161;
	wire [4-1:0] node162;
	wire [4-1:0] node163;
	wire [4-1:0] node164;
	wire [4-1:0] node167;
	wire [4-1:0] node170;
	wire [4-1:0] node172;
	wire [4-1:0] node175;
	wire [4-1:0] node176;
	wire [4-1:0] node179;
	wire [4-1:0] node180;
	wire [4-1:0] node183;
	wire [4-1:0] node186;
	wire [4-1:0] node187;
	wire [4-1:0] node188;
	wire [4-1:0] node189;
	wire [4-1:0] node192;
	wire [4-1:0] node195;
	wire [4-1:0] node196;
	wire [4-1:0] node199;
	wire [4-1:0] node202;
	wire [4-1:0] node204;
	wire [4-1:0] node205;
	wire [4-1:0] node209;
	wire [4-1:0] node210;
	wire [4-1:0] node211;
	wire [4-1:0] node212;
	wire [4-1:0] node213;
	wire [4-1:0] node214;
	wire [4-1:0] node216;
	wire [4-1:0] node219;
	wire [4-1:0] node220;
	wire [4-1:0] node223;
	wire [4-1:0] node226;
	wire [4-1:0] node227;
	wire [4-1:0] node228;
	wire [4-1:0] node231;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node238;
	wire [4-1:0] node241;
	wire [4-1:0] node242;
	wire [4-1:0] node243;
	wire [4-1:0] node244;
	wire [4-1:0] node248;
	wire [4-1:0] node249;
	wire [4-1:0] node253;
	wire [4-1:0] node254;
	wire [4-1:0] node256;
	wire [4-1:0] node259;
	wire [4-1:0] node260;
	wire [4-1:0] node263;
	wire [4-1:0] node266;
	wire [4-1:0] node267;
	wire [4-1:0] node268;
	wire [4-1:0] node269;
	wire [4-1:0] node271;
	wire [4-1:0] node274;
	wire [4-1:0] node275;
	wire [4-1:0] node278;
	wire [4-1:0] node281;
	wire [4-1:0] node282;
	wire [4-1:0] node283;
	wire [4-1:0] node287;
	wire [4-1:0] node289;
	wire [4-1:0] node292;
	wire [4-1:0] node293;
	wire [4-1:0] node294;
	wire [4-1:0] node295;
	wire [4-1:0] node298;
	wire [4-1:0] node301;
	wire [4-1:0] node302;
	wire [4-1:0] node305;
	wire [4-1:0] node308;
	wire [4-1:0] node309;
	wire [4-1:0] node312;
	wire [4-1:0] node313;
	wire [4-1:0] node316;
	wire [4-1:0] node319;
	wire [4-1:0] node320;
	wire [4-1:0] node321;
	wire [4-1:0] node322;
	wire [4-1:0] node323;
	wire [4-1:0] node325;
	wire [4-1:0] node328;
	wire [4-1:0] node329;
	wire [4-1:0] node333;
	wire [4-1:0] node334;
	wire [4-1:0] node337;
	wire [4-1:0] node338;
	wire [4-1:0] node341;
	wire [4-1:0] node344;
	wire [4-1:0] node345;
	wire [4-1:0] node346;
	wire [4-1:0] node347;
	wire [4-1:0] node351;
	wire [4-1:0] node352;
	wire [4-1:0] node356;
	wire [4-1:0] node357;
	wire [4-1:0] node358;
	wire [4-1:0] node361;
	wire [4-1:0] node365;
	wire [4-1:0] node366;
	wire [4-1:0] node367;
	wire [4-1:0] node368;
	wire [4-1:0] node369;
	wire [4-1:0] node373;
	wire [4-1:0] node374;
	wire [4-1:0] node378;
	wire [4-1:0] node379;
	wire [4-1:0] node380;
	wire [4-1:0] node384;
	wire [4-1:0] node385;
	wire [4-1:0] node388;
	wire [4-1:0] node391;
	wire [4-1:0] node392;
	wire [4-1:0] node393;
	wire [4-1:0] node394;
	wire [4-1:0] node398;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node404;
	wire [4-1:0] node407;
	wire [4-1:0] node408;
	wire [4-1:0] node411;
	wire [4-1:0] node414;
	wire [4-1:0] node415;
	wire [4-1:0] node416;
	wire [4-1:0] node417;
	wire [4-1:0] node418;
	wire [4-1:0] node419;
	wire [4-1:0] node420;
	wire [4-1:0] node421;
	wire [4-1:0] node424;
	wire [4-1:0] node427;
	wire [4-1:0] node429;
	wire [4-1:0] node432;
	wire [4-1:0] node433;
	wire [4-1:0] node435;
	wire [4-1:0] node438;
	wire [4-1:0] node439;
	wire [4-1:0] node442;
	wire [4-1:0] node445;
	wire [4-1:0] node446;
	wire [4-1:0] node447;
	wire [4-1:0] node448;
	wire [4-1:0] node451;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node459;
	wire [4-1:0] node460;
	wire [4-1:0] node462;
	wire [4-1:0] node465;
	wire [4-1:0] node466;
	wire [4-1:0] node469;
	wire [4-1:0] node472;
	wire [4-1:0] node473;
	wire [4-1:0] node474;
	wire [4-1:0] node476;
	wire [4-1:0] node477;
	wire [4-1:0] node480;
	wire [4-1:0] node483;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node490;
	wire [4-1:0] node491;
	wire [4-1:0] node492;
	wire [4-1:0] node493;
	wire [4-1:0] node496;
	wire [4-1:0] node499;
	wire [4-1:0] node501;
	wire [4-1:0] node504;
	wire [4-1:0] node505;
	wire [4-1:0] node506;
	wire [4-1:0] node509;
	wire [4-1:0] node512;
	wire [4-1:0] node513;
	wire [4-1:0] node517;
	wire [4-1:0] node518;
	wire [4-1:0] node519;
	wire [4-1:0] node520;
	wire [4-1:0] node521;
	wire [4-1:0] node522;
	wire [4-1:0] node526;
	wire [4-1:0] node527;
	wire [4-1:0] node530;
	wire [4-1:0] node533;
	wire [4-1:0] node534;
	wire [4-1:0] node535;
	wire [4-1:0] node539;
	wire [4-1:0] node540;
	wire [4-1:0] node543;
	wire [4-1:0] node546;
	wire [4-1:0] node547;
	wire [4-1:0] node548;
	wire [4-1:0] node549;
	wire [4-1:0] node553;
	wire [4-1:0] node554;
	wire [4-1:0] node557;
	wire [4-1:0] node560;
	wire [4-1:0] node561;
	wire [4-1:0] node562;
	wire [4-1:0] node565;
	wire [4-1:0] node568;
	wire [4-1:0] node569;
	wire [4-1:0] node573;
	wire [4-1:0] node574;
	wire [4-1:0] node575;
	wire [4-1:0] node576;
	wire [4-1:0] node580;
	wire [4-1:0] node581;
	wire [4-1:0] node582;
	wire [4-1:0] node586;
	wire [4-1:0] node587;
	wire [4-1:0] node591;
	wire [4-1:0] node592;
	wire [4-1:0] node593;
	wire [4-1:0] node594;
	wire [4-1:0] node597;
	wire [4-1:0] node600;
	wire [4-1:0] node601;
	wire [4-1:0] node604;
	wire [4-1:0] node607;
	wire [4-1:0] node608;
	wire [4-1:0] node610;
	wire [4-1:0] node613;
	wire [4-1:0] node615;
	wire [4-1:0] node618;
	wire [4-1:0] node619;
	wire [4-1:0] node620;
	wire [4-1:0] node621;
	wire [4-1:0] node622;
	wire [4-1:0] node623;
	wire [4-1:0] node624;
	wire [4-1:0] node627;
	wire [4-1:0] node630;
	wire [4-1:0] node631;
	wire [4-1:0] node635;
	wire [4-1:0] node636;
	wire [4-1:0] node637;
	wire [4-1:0] node640;
	wire [4-1:0] node644;
	wire [4-1:0] node645;
	wire [4-1:0] node646;
	wire [4-1:0] node647;
	wire [4-1:0] node650;
	wire [4-1:0] node653;
	wire [4-1:0] node654;
	wire [4-1:0] node657;
	wire [4-1:0] node660;
	wire [4-1:0] node661;
	wire [4-1:0] node663;
	wire [4-1:0] node666;
	wire [4-1:0] node668;
	wire [4-1:0] node671;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node674;
	wire [4-1:0] node677;
	wire [4-1:0] node678;
	wire [4-1:0] node682;
	wire [4-1:0] node683;
	wire [4-1:0] node684;
	wire [4-1:0] node688;
	wire [4-1:0] node689;
	wire [4-1:0] node692;
	wire [4-1:0] node695;
	wire [4-1:0] node696;
	wire [4-1:0] node698;
	wire [4-1:0] node699;
	wire [4-1:0] node702;
	wire [4-1:0] node705;
	wire [4-1:0] node706;
	wire [4-1:0] node707;
	wire [4-1:0] node710;
	wire [4-1:0] node713;
	wire [4-1:0] node714;
	wire [4-1:0] node717;
	wire [4-1:0] node720;
	wire [4-1:0] node721;
	wire [4-1:0] node722;
	wire [4-1:0] node723;
	wire [4-1:0] node724;
	wire [4-1:0] node726;
	wire [4-1:0] node729;
	wire [4-1:0] node730;
	wire [4-1:0] node733;
	wire [4-1:0] node736;
	wire [4-1:0] node737;
	wire [4-1:0] node739;
	wire [4-1:0] node742;
	wire [4-1:0] node743;
	wire [4-1:0] node747;
	wire [4-1:0] node748;
	wire [4-1:0] node750;
	wire [4-1:0] node751;
	wire [4-1:0] node754;
	wire [4-1:0] node757;
	wire [4-1:0] node758;
	wire [4-1:0] node759;
	wire [4-1:0] node762;
	wire [4-1:0] node765;
	wire [4-1:0] node767;
	wire [4-1:0] node770;
	wire [4-1:0] node771;
	wire [4-1:0] node772;
	wire [4-1:0] node773;
	wire [4-1:0] node774;
	wire [4-1:0] node777;
	wire [4-1:0] node780;
	wire [4-1:0] node782;
	wire [4-1:0] node785;
	wire [4-1:0] node786;
	wire [4-1:0] node787;
	wire [4-1:0] node791;
	wire [4-1:0] node792;
	wire [4-1:0] node795;
	wire [4-1:0] node798;
	wire [4-1:0] node799;
	wire [4-1:0] node800;
	wire [4-1:0] node802;
	wire [4-1:0] node805;
	wire [4-1:0] node806;
	wire [4-1:0] node810;
	wire [4-1:0] node811;
	wire [4-1:0] node813;
	wire [4-1:0] node816;
	wire [4-1:0] node817;
	wire [4-1:0] node821;
	wire [4-1:0] node822;
	wire [4-1:0] node823;
	wire [4-1:0] node824;
	wire [4-1:0] node825;
	wire [4-1:0] node826;
	wire [4-1:0] node827;
	wire [4-1:0] node828;
	wire [4-1:0] node829;
	wire [4-1:0] node832;
	wire [4-1:0] node835;
	wire [4-1:0] node836;
	wire [4-1:0] node839;
	wire [4-1:0] node842;
	wire [4-1:0] node843;
	wire [4-1:0] node844;
	wire [4-1:0] node847;
	wire [4-1:0] node850;
	wire [4-1:0] node853;
	wire [4-1:0] node854;
	wire [4-1:0] node855;
	wire [4-1:0] node856;
	wire [4-1:0] node859;
	wire [4-1:0] node862;
	wire [4-1:0] node863;
	wire [4-1:0] node866;
	wire [4-1:0] node869;
	wire [4-1:0] node870;
	wire [4-1:0] node872;
	wire [4-1:0] node875;
	wire [4-1:0] node876;
	wire [4-1:0] node880;
	wire [4-1:0] node881;
	wire [4-1:0] node882;
	wire [4-1:0] node883;
	wire [4-1:0] node884;
	wire [4-1:0] node887;
	wire [4-1:0] node890;
	wire [4-1:0] node892;
	wire [4-1:0] node895;
	wire [4-1:0] node896;
	wire [4-1:0] node897;
	wire [4-1:0] node900;
	wire [4-1:0] node903;
	wire [4-1:0] node904;
	wire [4-1:0] node907;
	wire [4-1:0] node910;
	wire [4-1:0] node911;
	wire [4-1:0] node912;
	wire [4-1:0] node913;
	wire [4-1:0] node917;
	wire [4-1:0] node918;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node924;
	wire [4-1:0] node927;
	wire [4-1:0] node930;
	wire [4-1:0] node931;
	wire [4-1:0] node934;
	wire [4-1:0] node937;
	wire [4-1:0] node938;
	wire [4-1:0] node939;
	wire [4-1:0] node940;
	wire [4-1:0] node941;
	wire [4-1:0] node942;
	wire [4-1:0] node945;
	wire [4-1:0] node948;
	wire [4-1:0] node949;
	wire [4-1:0] node952;
	wire [4-1:0] node955;
	wire [4-1:0] node956;
	wire [4-1:0] node957;
	wire [4-1:0] node961;
	wire [4-1:0] node962;
	wire [4-1:0] node966;
	wire [4-1:0] node967;
	wire [4-1:0] node968;
	wire [4-1:0] node969;
	wire [4-1:0] node973;
	wire [4-1:0] node975;
	wire [4-1:0] node979;
	wire [4-1:0] node980;
	wire [4-1:0] node981;
	wire [4-1:0] node982;
	wire [4-1:0] node984;
	wire [4-1:0] node987;
	wire [4-1:0] node988;
	wire [4-1:0] node992;
	wire [4-1:0] node993;
	wire [4-1:0] node995;
	wire [4-1:0] node998;
	wire [4-1:0] node999;
	wire [4-1:0] node1003;
	wire [4-1:0] node1004;
	wire [4-1:0] node1005;
	wire [4-1:0] node1006;
	wire [4-1:0] node1010;
	wire [4-1:0] node1011;
	wire [4-1:0] node1014;
	wire [4-1:0] node1017;
	wire [4-1:0] node1018;
	wire [4-1:0] node1019;
	wire [4-1:0] node1022;
	wire [4-1:0] node1025;
	wire [4-1:0] node1026;
	wire [4-1:0] node1030;
	wire [4-1:0] node1031;
	wire [4-1:0] node1032;
	wire [4-1:0] node1033;
	wire [4-1:0] node1034;
	wire [4-1:0] node1035;
	wire [4-1:0] node1038;
	wire [4-1:0] node1041;
	wire [4-1:0] node1042;
	wire [4-1:0] node1043;
	wire [4-1:0] node1046;
	wire [4-1:0] node1049;
	wire [4-1:0] node1052;
	wire [4-1:0] node1053;
	wire [4-1:0] node1054;
	wire [4-1:0] node1055;
	wire [4-1:0] node1059;
	wire [4-1:0] node1060;
	wire [4-1:0] node1063;
	wire [4-1:0] node1066;
	wire [4-1:0] node1067;
	wire [4-1:0] node1068;
	wire [4-1:0] node1071;
	wire [4-1:0] node1074;
	wire [4-1:0] node1075;
	wire [4-1:0] node1078;
	wire [4-1:0] node1081;
	wire [4-1:0] node1082;
	wire [4-1:0] node1083;
	wire [4-1:0] node1084;
	wire [4-1:0] node1085;
	wire [4-1:0] node1088;
	wire [4-1:0] node1091;
	wire [4-1:0] node1092;
	wire [4-1:0] node1096;
	wire [4-1:0] node1097;
	wire [4-1:0] node1100;
	wire [4-1:0] node1101;
	wire [4-1:0] node1105;
	wire [4-1:0] node1106;
	wire [4-1:0] node1107;
	wire [4-1:0] node1108;
	wire [4-1:0] node1112;
	wire [4-1:0] node1114;
	wire [4-1:0] node1117;
	wire [4-1:0] node1118;
	wire [4-1:0] node1120;
	wire [4-1:0] node1123;
	wire [4-1:0] node1124;
	wire [4-1:0] node1127;
	wire [4-1:0] node1130;
	wire [4-1:0] node1131;
	wire [4-1:0] node1132;
	wire [4-1:0] node1133;
	wire [4-1:0] node1134;
	wire [4-1:0] node1135;
	wire [4-1:0] node1138;
	wire [4-1:0] node1141;
	wire [4-1:0] node1143;
	wire [4-1:0] node1146;
	wire [4-1:0] node1147;
	wire [4-1:0] node1148;
	wire [4-1:0] node1152;
	wire [4-1:0] node1153;
	wire [4-1:0] node1157;
	wire [4-1:0] node1158;
	wire [4-1:0] node1159;
	wire [4-1:0] node1161;
	wire [4-1:0] node1164;
	wire [4-1:0] node1165;
	wire [4-1:0] node1168;
	wire [4-1:0] node1171;
	wire [4-1:0] node1172;
	wire [4-1:0] node1174;
	wire [4-1:0] node1177;
	wire [4-1:0] node1178;
	wire [4-1:0] node1182;
	wire [4-1:0] node1183;
	wire [4-1:0] node1184;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1189;
	wire [4-1:0] node1192;
	wire [4-1:0] node1195;
	wire [4-1:0] node1196;
	wire [4-1:0] node1197;
	wire [4-1:0] node1200;
	wire [4-1:0] node1203;
	wire [4-1:0] node1205;
	wire [4-1:0] node1208;
	wire [4-1:0] node1209;
	wire [4-1:0] node1210;
	wire [4-1:0] node1211;
	wire [4-1:0] node1215;
	wire [4-1:0] node1216;
	wire [4-1:0] node1219;
	wire [4-1:0] node1222;
	wire [4-1:0] node1223;
	wire [4-1:0] node1224;
	wire [4-1:0] node1227;
	wire [4-1:0] node1230;
	wire [4-1:0] node1231;
	wire [4-1:0] node1235;
	wire [4-1:0] node1236;
	wire [4-1:0] node1237;
	wire [4-1:0] node1238;
	wire [4-1:0] node1239;
	wire [4-1:0] node1240;
	wire [4-1:0] node1241;
	wire [4-1:0] node1242;
	wire [4-1:0] node1246;
	wire [4-1:0] node1249;
	wire [4-1:0] node1250;
	wire [4-1:0] node1251;
	wire [4-1:0] node1255;
	wire [4-1:0] node1258;
	wire [4-1:0] node1259;
	wire [4-1:0] node1260;
	wire [4-1:0] node1262;
	wire [4-1:0] node1265;
	wire [4-1:0] node1267;
	wire [4-1:0] node1270;
	wire [4-1:0] node1271;
	wire [4-1:0] node1272;
	wire [4-1:0] node1275;
	wire [4-1:0] node1278;
	wire [4-1:0] node1279;
	wire [4-1:0] node1282;
	wire [4-1:0] node1285;
	wire [4-1:0] node1286;
	wire [4-1:0] node1287;
	wire [4-1:0] node1288;
	wire [4-1:0] node1289;
	wire [4-1:0] node1292;
	wire [4-1:0] node1295;
	wire [4-1:0] node1297;
	wire [4-1:0] node1300;
	wire [4-1:0] node1301;
	wire [4-1:0] node1303;
	wire [4-1:0] node1306;
	wire [4-1:0] node1307;
	wire [4-1:0] node1311;
	wire [4-1:0] node1312;
	wire [4-1:0] node1313;
	wire [4-1:0] node1314;
	wire [4-1:0] node1317;
	wire [4-1:0] node1320;
	wire [4-1:0] node1321;
	wire [4-1:0] node1324;
	wire [4-1:0] node1327;
	wire [4-1:0] node1328;
	wire [4-1:0] node1329;
	wire [4-1:0] node1333;
	wire [4-1:0] node1334;
	wire [4-1:0] node1337;
	wire [4-1:0] node1340;
	wire [4-1:0] node1341;
	wire [4-1:0] node1342;
	wire [4-1:0] node1343;
	wire [4-1:0] node1344;
	wire [4-1:0] node1345;
	wire [4-1:0] node1349;
	wire [4-1:0] node1350;
	wire [4-1:0] node1353;
	wire [4-1:0] node1356;
	wire [4-1:0] node1357;
	wire [4-1:0] node1358;
	wire [4-1:0] node1361;
	wire [4-1:0] node1364;
	wire [4-1:0] node1365;
	wire [4-1:0] node1368;
	wire [4-1:0] node1371;
	wire [4-1:0] node1372;
	wire [4-1:0] node1373;
	wire [4-1:0] node1374;
	wire [4-1:0] node1377;
	wire [4-1:0] node1380;
	wire [4-1:0] node1381;
	wire [4-1:0] node1384;
	wire [4-1:0] node1387;
	wire [4-1:0] node1388;
	wire [4-1:0] node1389;
	wire [4-1:0] node1392;
	wire [4-1:0] node1395;
	wire [4-1:0] node1397;
	wire [4-1:0] node1400;
	wire [4-1:0] node1401;
	wire [4-1:0] node1402;
	wire [4-1:0] node1403;
	wire [4-1:0] node1404;
	wire [4-1:0] node1408;
	wire [4-1:0] node1409;
	wire [4-1:0] node1413;
	wire [4-1:0] node1414;
	wire [4-1:0] node1417;
	wire [4-1:0] node1418;
	wire [4-1:0] node1421;
	wire [4-1:0] node1424;
	wire [4-1:0] node1425;
	wire [4-1:0] node1426;
	wire [4-1:0] node1427;
	wire [4-1:0] node1430;
	wire [4-1:0] node1433;
	wire [4-1:0] node1435;
	wire [4-1:0] node1438;
	wire [4-1:0] node1439;
	wire [4-1:0] node1440;
	wire [4-1:0] node1444;
	wire [4-1:0] node1446;
	wire [4-1:0] node1449;
	wire [4-1:0] node1450;
	wire [4-1:0] node1451;
	wire [4-1:0] node1452;
	wire [4-1:0] node1453;
	wire [4-1:0] node1454;
	wire [4-1:0] node1455;
	wire [4-1:0] node1459;
	wire [4-1:0] node1461;
	wire [4-1:0] node1464;
	wire [4-1:0] node1465;
	wire [4-1:0] node1466;
	wire [4-1:0] node1469;
	wire [4-1:0] node1472;
	wire [4-1:0] node1474;
	wire [4-1:0] node1477;
	wire [4-1:0] node1478;
	wire [4-1:0] node1479;
	wire [4-1:0] node1480;
	wire [4-1:0] node1484;
	wire [4-1:0] node1485;
	wire [4-1:0] node1488;
	wire [4-1:0] node1491;
	wire [4-1:0] node1492;
	wire [4-1:0] node1493;
	wire [4-1:0] node1496;
	wire [4-1:0] node1499;
	wire [4-1:0] node1500;
	wire [4-1:0] node1503;
	wire [4-1:0] node1506;
	wire [4-1:0] node1507;
	wire [4-1:0] node1508;
	wire [4-1:0] node1509;
	wire [4-1:0] node1513;
	wire [4-1:0] node1514;
	wire [4-1:0] node1515;
	wire [4-1:0] node1518;
	wire [4-1:0] node1521;
	wire [4-1:0] node1522;
	wire [4-1:0] node1526;
	wire [4-1:0] node1527;
	wire [4-1:0] node1528;
	wire [4-1:0] node1529;
	wire [4-1:0] node1532;
	wire [4-1:0] node1535;
	wire [4-1:0] node1536;
	wire [4-1:0] node1540;
	wire [4-1:0] node1541;
	wire [4-1:0] node1542;
	wire [4-1:0] node1546;
	wire [4-1:0] node1547;
	wire [4-1:0] node1550;
	wire [4-1:0] node1553;
	wire [4-1:0] node1554;
	wire [4-1:0] node1555;
	wire [4-1:0] node1556;
	wire [4-1:0] node1557;
	wire [4-1:0] node1558;
	wire [4-1:0] node1561;
	wire [4-1:0] node1564;
	wire [4-1:0] node1567;
	wire [4-1:0] node1568;
	wire [4-1:0] node1569;
	wire [4-1:0] node1572;
	wire [4-1:0] node1575;
	wire [4-1:0] node1577;
	wire [4-1:0] node1580;
	wire [4-1:0] node1581;
	wire [4-1:0] node1582;
	wire [4-1:0] node1584;
	wire [4-1:0] node1587;
	wire [4-1:0] node1588;
	wire [4-1:0] node1591;
	wire [4-1:0] node1594;
	wire [4-1:0] node1595;
	wire [4-1:0] node1596;
	wire [4-1:0] node1599;
	wire [4-1:0] node1602;
	wire [4-1:0] node1604;
	wire [4-1:0] node1607;
	wire [4-1:0] node1608;
	wire [4-1:0] node1609;
	wire [4-1:0] node1610;
	wire [4-1:0] node1611;
	wire [4-1:0] node1615;
	wire [4-1:0] node1616;
	wire [4-1:0] node1620;
	wire [4-1:0] node1621;
	wire [4-1:0] node1622;
	wire [4-1:0] node1625;
	wire [4-1:0] node1628;
	wire [4-1:0] node1629;
	wire [4-1:0] node1632;
	wire [4-1:0] node1635;
	wire [4-1:0] node1636;
	wire [4-1:0] node1637;
	wire [4-1:0] node1638;
	wire [4-1:0] node1642;
	wire [4-1:0] node1645;
	wire [4-1:0] node1646;
	wire [4-1:0] node1647;
	wire [4-1:0] node1650;
	wire [4-1:0] node1653;
	wire [4-1:0] node1654;
	wire [4-1:0] node1657;
	wire [4-1:0] node1660;
	wire [4-1:0] node1661;
	wire [4-1:0] node1662;
	wire [4-1:0] node1663;
	wire [4-1:0] node1664;
	wire [4-1:0] node1665;
	wire [4-1:0] node1666;
	wire [4-1:0] node1667;
	wire [4-1:0] node1668;
	wire [4-1:0] node1669;
	wire [4-1:0] node1672;
	wire [4-1:0] node1675;
	wire [4-1:0] node1676;
	wire [4-1:0] node1679;
	wire [4-1:0] node1682;
	wire [4-1:0] node1683;
	wire [4-1:0] node1684;
	wire [4-1:0] node1687;
	wire [4-1:0] node1690;
	wire [4-1:0] node1691;
	wire [4-1:0] node1694;
	wire [4-1:0] node1697;
	wire [4-1:0] node1698;
	wire [4-1:0] node1699;
	wire [4-1:0] node1701;
	wire [4-1:0] node1704;
	wire [4-1:0] node1705;
	wire [4-1:0] node1708;
	wire [4-1:0] node1711;
	wire [4-1:0] node1712;
	wire [4-1:0] node1713;
	wire [4-1:0] node1716;
	wire [4-1:0] node1719;
	wire [4-1:0] node1720;
	wire [4-1:0] node1724;
	wire [4-1:0] node1725;
	wire [4-1:0] node1726;
	wire [4-1:0] node1727;
	wire [4-1:0] node1728;
	wire [4-1:0] node1732;
	wire [4-1:0] node1734;
	wire [4-1:0] node1737;
	wire [4-1:0] node1738;
	wire [4-1:0] node1739;
	wire [4-1:0] node1742;
	wire [4-1:0] node1745;
	wire [4-1:0] node1746;
	wire [4-1:0] node1750;
	wire [4-1:0] node1751;
	wire [4-1:0] node1752;
	wire [4-1:0] node1753;
	wire [4-1:0] node1757;
	wire [4-1:0] node1759;
	wire [4-1:0] node1762;
	wire [4-1:0] node1763;
	wire [4-1:0] node1764;
	wire [4-1:0] node1767;
	wire [4-1:0] node1770;
	wire [4-1:0] node1771;
	wire [4-1:0] node1775;
	wire [4-1:0] node1776;
	wire [4-1:0] node1777;
	wire [4-1:0] node1778;
	wire [4-1:0] node1779;
	wire [4-1:0] node1782;
	wire [4-1:0] node1783;
	wire [4-1:0] node1786;
	wire [4-1:0] node1789;
	wire [4-1:0] node1790;
	wire [4-1:0] node1791;
	wire [4-1:0] node1795;
	wire [4-1:0] node1798;
	wire [4-1:0] node1799;
	wire [4-1:0] node1800;
	wire [4-1:0] node1801;
	wire [4-1:0] node1804;
	wire [4-1:0] node1807;
	wire [4-1:0] node1808;
	wire [4-1:0] node1812;
	wire [4-1:0] node1813;
	wire [4-1:0] node1814;
	wire [4-1:0] node1817;
	wire [4-1:0] node1820;
	wire [4-1:0] node1821;
	wire [4-1:0] node1824;
	wire [4-1:0] node1827;
	wire [4-1:0] node1828;
	wire [4-1:0] node1829;
	wire [4-1:0] node1830;
	wire [4-1:0] node1831;
	wire [4-1:0] node1834;
	wire [4-1:0] node1837;
	wire [4-1:0] node1838;
	wire [4-1:0] node1841;
	wire [4-1:0] node1844;
	wire [4-1:0] node1845;
	wire [4-1:0] node1847;
	wire [4-1:0] node1850;
	wire [4-1:0] node1851;
	wire [4-1:0] node1854;
	wire [4-1:0] node1857;
	wire [4-1:0] node1858;
	wire [4-1:0] node1859;
	wire [4-1:0] node1862;
	wire [4-1:0] node1865;
	wire [4-1:0] node1867;
	wire [4-1:0] node1868;
	wire [4-1:0] node1871;
	wire [4-1:0] node1874;
	wire [4-1:0] node1875;
	wire [4-1:0] node1876;
	wire [4-1:0] node1877;
	wire [4-1:0] node1878;
	wire [4-1:0] node1879;
	wire [4-1:0] node1882;
	wire [4-1:0] node1883;
	wire [4-1:0] node1886;
	wire [4-1:0] node1889;
	wire [4-1:0] node1890;
	wire [4-1:0] node1892;
	wire [4-1:0] node1895;
	wire [4-1:0] node1897;
	wire [4-1:0] node1900;
	wire [4-1:0] node1901;
	wire [4-1:0] node1903;
	wire [4-1:0] node1904;
	wire [4-1:0] node1907;
	wire [4-1:0] node1910;
	wire [4-1:0] node1912;
	wire [4-1:0] node1913;
	wire [4-1:0] node1917;
	wire [4-1:0] node1918;
	wire [4-1:0] node1919;
	wire [4-1:0] node1920;
	wire [4-1:0] node1921;
	wire [4-1:0] node1924;
	wire [4-1:0] node1928;
	wire [4-1:0] node1929;
	wire [4-1:0] node1931;
	wire [4-1:0] node1934;
	wire [4-1:0] node1935;
	wire [4-1:0] node1938;
	wire [4-1:0] node1941;
	wire [4-1:0] node1942;
	wire [4-1:0] node1943;
	wire [4-1:0] node1944;
	wire [4-1:0] node1947;
	wire [4-1:0] node1950;
	wire [4-1:0] node1952;
	wire [4-1:0] node1955;
	wire [4-1:0] node1956;
	wire [4-1:0] node1957;
	wire [4-1:0] node1960;
	wire [4-1:0] node1963;
	wire [4-1:0] node1964;
	wire [4-1:0] node1968;
	wire [4-1:0] node1969;
	wire [4-1:0] node1970;
	wire [4-1:0] node1971;
	wire [4-1:0] node1972;
	wire [4-1:0] node1973;
	wire [4-1:0] node1977;
	wire [4-1:0] node1978;
	wire [4-1:0] node1981;
	wire [4-1:0] node1984;
	wire [4-1:0] node1985;
	wire [4-1:0] node1987;
	wire [4-1:0] node1990;
	wire [4-1:0] node1992;
	wire [4-1:0] node1995;
	wire [4-1:0] node1996;
	wire [4-1:0] node1997;
	wire [4-1:0] node1999;
	wire [4-1:0] node2002;
	wire [4-1:0] node2004;
	wire [4-1:0] node2007;
	wire [4-1:0] node2008;
	wire [4-1:0] node2011;
	wire [4-1:0] node2012;
	wire [4-1:0] node2015;
	wire [4-1:0] node2018;
	wire [4-1:0] node2019;
	wire [4-1:0] node2020;
	wire [4-1:0] node2021;
	wire [4-1:0] node2023;
	wire [4-1:0] node2026;
	wire [4-1:0] node2028;
	wire [4-1:0] node2031;
	wire [4-1:0] node2032;
	wire [4-1:0] node2033;
	wire [4-1:0] node2037;
	wire [4-1:0] node2038;
	wire [4-1:0] node2042;
	wire [4-1:0] node2043;
	wire [4-1:0] node2044;
	wire [4-1:0] node2046;
	wire [4-1:0] node2049;
	wire [4-1:0] node2050;
	wire [4-1:0] node2053;
	wire [4-1:0] node2056;
	wire [4-1:0] node2057;
	wire [4-1:0] node2058;
	wire [4-1:0] node2061;
	wire [4-1:0] node2064;
	wire [4-1:0] node2065;
	wire [4-1:0] node2068;
	wire [4-1:0] node2071;
	wire [4-1:0] node2072;
	wire [4-1:0] node2073;
	wire [4-1:0] node2074;
	wire [4-1:0] node2075;
	wire [4-1:0] node2076;
	wire [4-1:0] node2077;
	wire [4-1:0] node2078;
	wire [4-1:0] node2081;
	wire [4-1:0] node2084;
	wire [4-1:0] node2085;
	wire [4-1:0] node2089;
	wire [4-1:0] node2090;
	wire [4-1:0] node2091;
	wire [4-1:0] node2094;
	wire [4-1:0] node2097;
	wire [4-1:0] node2098;
	wire [4-1:0] node2102;
	wire [4-1:0] node2103;
	wire [4-1:0] node2104;
	wire [4-1:0] node2105;
	wire [4-1:0] node2108;
	wire [4-1:0] node2111;
	wire [4-1:0] node2112;
	wire [4-1:0] node2116;
	wire [4-1:0] node2117;
	wire [4-1:0] node2119;
	wire [4-1:0] node2122;
	wire [4-1:0] node2123;
	wire [4-1:0] node2126;
	wire [4-1:0] node2129;
	wire [4-1:0] node2130;
	wire [4-1:0] node2131;
	wire [4-1:0] node2132;
	wire [4-1:0] node2133;
	wire [4-1:0] node2136;
	wire [4-1:0] node2139;
	wire [4-1:0] node2140;
	wire [4-1:0] node2143;
	wire [4-1:0] node2146;
	wire [4-1:0] node2147;
	wire [4-1:0] node2148;
	wire [4-1:0] node2151;
	wire [4-1:0] node2154;
	wire [4-1:0] node2155;
	wire [4-1:0] node2158;
	wire [4-1:0] node2161;
	wire [4-1:0] node2162;
	wire [4-1:0] node2163;
	wire [4-1:0] node2165;
	wire [4-1:0] node2169;
	wire [4-1:0] node2170;
	wire [4-1:0] node2171;
	wire [4-1:0] node2174;
	wire [4-1:0] node2177;
	wire [4-1:0] node2178;
	wire [4-1:0] node2181;
	wire [4-1:0] node2184;
	wire [4-1:0] node2185;
	wire [4-1:0] node2186;
	wire [4-1:0] node2187;
	wire [4-1:0] node2188;
	wire [4-1:0] node2189;
	wire [4-1:0] node2192;
	wire [4-1:0] node2195;
	wire [4-1:0] node2197;
	wire [4-1:0] node2200;
	wire [4-1:0] node2201;
	wire [4-1:0] node2202;
	wire [4-1:0] node2206;
	wire [4-1:0] node2209;
	wire [4-1:0] node2210;
	wire [4-1:0] node2211;
	wire [4-1:0] node2212;
	wire [4-1:0] node2215;
	wire [4-1:0] node2218;
	wire [4-1:0] node2219;
	wire [4-1:0] node2222;
	wire [4-1:0] node2225;
	wire [4-1:0] node2226;
	wire [4-1:0] node2228;
	wire [4-1:0] node2231;
	wire [4-1:0] node2232;
	wire [4-1:0] node2235;
	wire [4-1:0] node2238;
	wire [4-1:0] node2239;
	wire [4-1:0] node2240;
	wire [4-1:0] node2241;
	wire [4-1:0] node2242;
	wire [4-1:0] node2245;
	wire [4-1:0] node2248;
	wire [4-1:0] node2250;
	wire [4-1:0] node2253;
	wire [4-1:0] node2254;
	wire [4-1:0] node2255;
	wire [4-1:0] node2258;
	wire [4-1:0] node2261;
	wire [4-1:0] node2262;
	wire [4-1:0] node2265;
	wire [4-1:0] node2268;
	wire [4-1:0] node2269;
	wire [4-1:0] node2270;
	wire [4-1:0] node2271;
	wire [4-1:0] node2274;
	wire [4-1:0] node2277;
	wire [4-1:0] node2278;
	wire [4-1:0] node2282;
	wire [4-1:0] node2283;
	wire [4-1:0] node2284;
	wire [4-1:0] node2287;
	wire [4-1:0] node2290;
	wire [4-1:0] node2291;
	wire [4-1:0] node2294;
	wire [4-1:0] node2297;
	wire [4-1:0] node2298;
	wire [4-1:0] node2299;
	wire [4-1:0] node2300;
	wire [4-1:0] node2301;
	wire [4-1:0] node2302;
	wire [4-1:0] node2304;
	wire [4-1:0] node2307;
	wire [4-1:0] node2308;
	wire [4-1:0] node2312;
	wire [4-1:0] node2313;
	wire [4-1:0] node2314;
	wire [4-1:0] node2317;
	wire [4-1:0] node2320;
	wire [4-1:0] node2321;
	wire [4-1:0] node2325;
	wire [4-1:0] node2326;
	wire [4-1:0] node2327;
	wire [4-1:0] node2329;
	wire [4-1:0] node2332;
	wire [4-1:0] node2333;
	wire [4-1:0] node2336;
	wire [4-1:0] node2339;
	wire [4-1:0] node2340;
	wire [4-1:0] node2341;
	wire [4-1:0] node2344;
	wire [4-1:0] node2347;
	wire [4-1:0] node2350;
	wire [4-1:0] node2351;
	wire [4-1:0] node2352;
	wire [4-1:0] node2354;
	wire [4-1:0] node2355;
	wire [4-1:0] node2359;
	wire [4-1:0] node2360;
	wire [4-1:0] node2362;
	wire [4-1:0] node2365;
	wire [4-1:0] node2366;
	wire [4-1:0] node2369;
	wire [4-1:0] node2372;
	wire [4-1:0] node2373;
	wire [4-1:0] node2374;
	wire [4-1:0] node2376;
	wire [4-1:0] node2379;
	wire [4-1:0] node2380;
	wire [4-1:0] node2384;
	wire [4-1:0] node2385;
	wire [4-1:0] node2386;
	wire [4-1:0] node2390;
	wire [4-1:0] node2392;
	wire [4-1:0] node2395;
	wire [4-1:0] node2396;
	wire [4-1:0] node2397;
	wire [4-1:0] node2398;
	wire [4-1:0] node2399;
	wire [4-1:0] node2400;
	wire [4-1:0] node2404;
	wire [4-1:0] node2405;
	wire [4-1:0] node2408;
	wire [4-1:0] node2411;
	wire [4-1:0] node2412;
	wire [4-1:0] node2413;
	wire [4-1:0] node2416;
	wire [4-1:0] node2419;
	wire [4-1:0] node2420;
	wire [4-1:0] node2424;
	wire [4-1:0] node2425;
	wire [4-1:0] node2426;
	wire [4-1:0] node2427;
	wire [4-1:0] node2430;
	wire [4-1:0] node2433;
	wire [4-1:0] node2434;
	wire [4-1:0] node2438;
	wire [4-1:0] node2439;
	wire [4-1:0] node2440;
	wire [4-1:0] node2444;
	wire [4-1:0] node2445;
	wire [4-1:0] node2448;
	wire [4-1:0] node2451;
	wire [4-1:0] node2452;
	wire [4-1:0] node2453;
	wire [4-1:0] node2454;
	wire [4-1:0] node2456;
	wire [4-1:0] node2459;
	wire [4-1:0] node2461;
	wire [4-1:0] node2464;
	wire [4-1:0] node2465;
	wire [4-1:0] node2466;
	wire [4-1:0] node2470;
	wire [4-1:0] node2471;
	wire [4-1:0] node2475;
	wire [4-1:0] node2476;
	wire [4-1:0] node2477;
	wire [4-1:0] node2478;
	wire [4-1:0] node2481;
	wire [4-1:0] node2484;
	wire [4-1:0] node2485;
	wire [4-1:0] node2488;
	wire [4-1:0] node2491;
	wire [4-1:0] node2492;
	wire [4-1:0] node2493;
	wire [4-1:0] node2496;
	wire [4-1:0] node2499;
	wire [4-1:0] node2500;
	wire [4-1:0] node2503;
	wire [4-1:0] node2506;
	wire [4-1:0] node2507;
	wire [4-1:0] node2508;
	wire [4-1:0] node2509;
	wire [4-1:0] node2510;
	wire [4-1:0] node2511;
	wire [4-1:0] node2512;
	wire [4-1:0] node2513;
	wire [4-1:0] node2516;
	wire [4-1:0] node2517;
	wire [4-1:0] node2521;
	wire [4-1:0] node2522;
	wire [4-1:0] node2524;
	wire [4-1:0] node2527;
	wire [4-1:0] node2528;
	wire [4-1:0] node2532;
	wire [4-1:0] node2533;
	wire [4-1:0] node2534;
	wire [4-1:0] node2535;
	wire [4-1:0] node2538;
	wire [4-1:0] node2541;
	wire [4-1:0] node2544;
	wire [4-1:0] node2545;
	wire [4-1:0] node2548;
	wire [4-1:0] node2549;
	wire [4-1:0] node2553;
	wire [4-1:0] node2554;
	wire [4-1:0] node2555;
	wire [4-1:0] node2556;
	wire [4-1:0] node2557;
	wire [4-1:0] node2561;
	wire [4-1:0] node2562;
	wire [4-1:0] node2566;
	wire [4-1:0] node2567;
	wire [4-1:0] node2570;
	wire [4-1:0] node2571;
	wire [4-1:0] node2575;
	wire [4-1:0] node2576;
	wire [4-1:0] node2577;
	wire [4-1:0] node2578;
	wire [4-1:0] node2581;
	wire [4-1:0] node2584;
	wire [4-1:0] node2585;
	wire [4-1:0] node2588;
	wire [4-1:0] node2591;
	wire [4-1:0] node2592;
	wire [4-1:0] node2593;
	wire [4-1:0] node2596;
	wire [4-1:0] node2599;
	wire [4-1:0] node2600;
	wire [4-1:0] node2604;
	wire [4-1:0] node2605;
	wire [4-1:0] node2606;
	wire [4-1:0] node2607;
	wire [4-1:0] node2608;
	wire [4-1:0] node2609;
	wire [4-1:0] node2612;
	wire [4-1:0] node2615;
	wire [4-1:0] node2617;
	wire [4-1:0] node2620;
	wire [4-1:0] node2621;
	wire [4-1:0] node2623;
	wire [4-1:0] node2626;
	wire [4-1:0] node2629;
	wire [4-1:0] node2630;
	wire [4-1:0] node2631;
	wire [4-1:0] node2632;
	wire [4-1:0] node2636;
	wire [4-1:0] node2639;
	wire [4-1:0] node2640;
	wire [4-1:0] node2642;
	wire [4-1:0] node2645;
	wire [4-1:0] node2647;
	wire [4-1:0] node2650;
	wire [4-1:0] node2651;
	wire [4-1:0] node2652;
	wire [4-1:0] node2653;
	wire [4-1:0] node2655;
	wire [4-1:0] node2658;
	wire [4-1:0] node2659;
	wire [4-1:0] node2663;
	wire [4-1:0] node2664;
	wire [4-1:0] node2665;
	wire [4-1:0] node2669;
	wire [4-1:0] node2671;
	wire [4-1:0] node2674;
	wire [4-1:0] node2675;
	wire [4-1:0] node2676;
	wire [4-1:0] node2679;
	wire [4-1:0] node2682;
	wire [4-1:0] node2683;
	wire [4-1:0] node2684;
	wire [4-1:0] node2687;
	wire [4-1:0] node2690;
	wire [4-1:0] node2691;
	wire [4-1:0] node2695;
	wire [4-1:0] node2696;
	wire [4-1:0] node2697;
	wire [4-1:0] node2698;
	wire [4-1:0] node2699;
	wire [4-1:0] node2700;
	wire [4-1:0] node2702;
	wire [4-1:0] node2705;
	wire [4-1:0] node2706;
	wire [4-1:0] node2709;
	wire [4-1:0] node2712;
	wire [4-1:0] node2713;
	wire [4-1:0] node2714;
	wire [4-1:0] node2717;
	wire [4-1:0] node2720;
	wire [4-1:0] node2721;
	wire [4-1:0] node2725;
	wire [4-1:0] node2726;
	wire [4-1:0] node2727;
	wire [4-1:0] node2728;
	wire [4-1:0] node2731;
	wire [4-1:0] node2734;
	wire [4-1:0] node2735;
	wire [4-1:0] node2738;
	wire [4-1:0] node2741;
	wire [4-1:0] node2742;
	wire [4-1:0] node2743;
	wire [4-1:0] node2747;
	wire [4-1:0] node2749;
	wire [4-1:0] node2752;
	wire [4-1:0] node2753;
	wire [4-1:0] node2754;
	wire [4-1:0] node2755;
	wire [4-1:0] node2756;
	wire [4-1:0] node2760;
	wire [4-1:0] node2761;
	wire [4-1:0] node2765;
	wire [4-1:0] node2766;
	wire [4-1:0] node2769;
	wire [4-1:0] node2770;
	wire [4-1:0] node2774;
	wire [4-1:0] node2775;
	wire [4-1:0] node2776;
	wire [4-1:0] node2779;
	wire [4-1:0] node2780;
	wire [4-1:0] node2783;
	wire [4-1:0] node2786;
	wire [4-1:0] node2787;
	wire [4-1:0] node2789;
	wire [4-1:0] node2792;
	wire [4-1:0] node2793;
	wire [4-1:0] node2796;
	wire [4-1:0] node2799;
	wire [4-1:0] node2800;
	wire [4-1:0] node2801;
	wire [4-1:0] node2802;
	wire [4-1:0] node2803;
	wire [4-1:0] node2805;
	wire [4-1:0] node2808;
	wire [4-1:0] node2809;
	wire [4-1:0] node2812;
	wire [4-1:0] node2815;
	wire [4-1:0] node2816;
	wire [4-1:0] node2819;
	wire [4-1:0] node2821;
	wire [4-1:0] node2824;
	wire [4-1:0] node2825;
	wire [4-1:0] node2826;
	wire [4-1:0] node2827;
	wire [4-1:0] node2830;
	wire [4-1:0] node2833;
	wire [4-1:0] node2835;
	wire [4-1:0] node2838;
	wire [4-1:0] node2839;
	wire [4-1:0] node2840;
	wire [4-1:0] node2844;
	wire [4-1:0] node2847;
	wire [4-1:0] node2848;
	wire [4-1:0] node2849;
	wire [4-1:0] node2850;
	wire [4-1:0] node2851;
	wire [4-1:0] node2854;
	wire [4-1:0] node2857;
	wire [4-1:0] node2859;
	wire [4-1:0] node2862;
	wire [4-1:0] node2863;
	wire [4-1:0] node2864;
	wire [4-1:0] node2867;
	wire [4-1:0] node2870;
	wire [4-1:0] node2871;
	wire [4-1:0] node2875;
	wire [4-1:0] node2876;
	wire [4-1:0] node2877;
	wire [4-1:0] node2878;
	wire [4-1:0] node2881;
	wire [4-1:0] node2884;
	wire [4-1:0] node2887;
	wire [4-1:0] node2888;
	wire [4-1:0] node2889;
	wire [4-1:0] node2892;
	wire [4-1:0] node2895;
	wire [4-1:0] node2896;
	wire [4-1:0] node2900;
	wire [4-1:0] node2901;
	wire [4-1:0] node2902;
	wire [4-1:0] node2903;
	wire [4-1:0] node2904;
	wire [4-1:0] node2905;
	wire [4-1:0] node2906;
	wire [4-1:0] node2908;
	wire [4-1:0] node2911;
	wire [4-1:0] node2913;
	wire [4-1:0] node2916;
	wire [4-1:0] node2917;
	wire [4-1:0] node2920;
	wire [4-1:0] node2922;
	wire [4-1:0] node2925;
	wire [4-1:0] node2926;
	wire [4-1:0] node2927;
	wire [4-1:0] node2928;
	wire [4-1:0] node2931;
	wire [4-1:0] node2934;
	wire [4-1:0] node2937;
	wire [4-1:0] node2938;
	wire [4-1:0] node2939;
	wire [4-1:0] node2942;
	wire [4-1:0] node2945;
	wire [4-1:0] node2946;
	wire [4-1:0] node2949;
	wire [4-1:0] node2952;
	wire [4-1:0] node2953;
	wire [4-1:0] node2954;
	wire [4-1:0] node2955;
	wire [4-1:0] node2956;
	wire [4-1:0] node2959;
	wire [4-1:0] node2962;
	wire [4-1:0] node2963;
	wire [4-1:0] node2967;
	wire [4-1:0] node2968;
	wire [4-1:0] node2971;
	wire [4-1:0] node2973;
	wire [4-1:0] node2976;
	wire [4-1:0] node2977;
	wire [4-1:0] node2978;
	wire [4-1:0] node2979;
	wire [4-1:0] node2983;
	wire [4-1:0] node2984;
	wire [4-1:0] node2988;
	wire [4-1:0] node2989;
	wire [4-1:0] node2990;
	wire [4-1:0] node2994;
	wire [4-1:0] node2995;
	wire [4-1:0] node2998;
	wire [4-1:0] node3001;
	wire [4-1:0] node3002;
	wire [4-1:0] node3003;
	wire [4-1:0] node3004;
	wire [4-1:0] node3005;
	wire [4-1:0] node3007;
	wire [4-1:0] node3010;
	wire [4-1:0] node3011;
	wire [4-1:0] node3014;
	wire [4-1:0] node3017;
	wire [4-1:0] node3018;
	wire [4-1:0] node3019;
	wire [4-1:0] node3022;
	wire [4-1:0] node3026;
	wire [4-1:0] node3027;
	wire [4-1:0] node3028;
	wire [4-1:0] node3029;
	wire [4-1:0] node3032;
	wire [4-1:0] node3035;
	wire [4-1:0] node3036;
	wire [4-1:0] node3039;
	wire [4-1:0] node3042;
	wire [4-1:0] node3043;
	wire [4-1:0] node3044;
	wire [4-1:0] node3048;
	wire [4-1:0] node3049;
	wire [4-1:0] node3052;
	wire [4-1:0] node3055;
	wire [4-1:0] node3056;
	wire [4-1:0] node3057;
	wire [4-1:0] node3058;
	wire [4-1:0] node3061;
	wire [4-1:0] node3062;
	wire [4-1:0] node3065;
	wire [4-1:0] node3068;
	wire [4-1:0] node3069;
	wire [4-1:0] node3071;
	wire [4-1:0] node3075;
	wire [4-1:0] node3076;
	wire [4-1:0] node3077;
	wire [4-1:0] node3078;
	wire [4-1:0] node3081;
	wire [4-1:0] node3084;
	wire [4-1:0] node3085;
	wire [4-1:0] node3088;
	wire [4-1:0] node3091;
	wire [4-1:0] node3092;
	wire [4-1:0] node3093;
	wire [4-1:0] node3097;
	wire [4-1:0] node3098;
	wire [4-1:0] node3102;
	wire [4-1:0] node3103;
	wire [4-1:0] node3104;
	wire [4-1:0] node3105;
	wire [4-1:0] node3106;
	wire [4-1:0] node3107;
	wire [4-1:0] node3110;
	wire [4-1:0] node3112;
	wire [4-1:0] node3115;
	wire [4-1:0] node3116;
	wire [4-1:0] node3119;
	wire [4-1:0] node3120;
	wire [4-1:0] node3123;
	wire [4-1:0] node3126;
	wire [4-1:0] node3127;
	wire [4-1:0] node3128;
	wire [4-1:0] node3131;
	wire [4-1:0] node3132;
	wire [4-1:0] node3135;
	wire [4-1:0] node3138;
	wire [4-1:0] node3139;
	wire [4-1:0] node3140;
	wire [4-1:0] node3144;
	wire [4-1:0] node3145;
	wire [4-1:0] node3149;
	wire [4-1:0] node3150;
	wire [4-1:0] node3151;
	wire [4-1:0] node3152;
	wire [4-1:0] node3153;
	wire [4-1:0] node3157;
	wire [4-1:0] node3158;
	wire [4-1:0] node3161;
	wire [4-1:0] node3164;
	wire [4-1:0] node3165;
	wire [4-1:0] node3166;
	wire [4-1:0] node3170;
	wire [4-1:0] node3173;
	wire [4-1:0] node3174;
	wire [4-1:0] node3175;
	wire [4-1:0] node3176;
	wire [4-1:0] node3179;
	wire [4-1:0] node3183;
	wire [4-1:0] node3184;
	wire [4-1:0] node3185;
	wire [4-1:0] node3189;
	wire [4-1:0] node3190;
	wire [4-1:0] node3194;
	wire [4-1:0] node3195;
	wire [4-1:0] node3196;
	wire [4-1:0] node3197;
	wire [4-1:0] node3198;
	wire [4-1:0] node3200;
	wire [4-1:0] node3203;
	wire [4-1:0] node3204;
	wire [4-1:0] node3207;
	wire [4-1:0] node3210;
	wire [4-1:0] node3211;
	wire [4-1:0] node3212;
	wire [4-1:0] node3215;
	wire [4-1:0] node3218;
	wire [4-1:0] node3219;
	wire [4-1:0] node3223;
	wire [4-1:0] node3224;
	wire [4-1:0] node3225;
	wire [4-1:0] node3227;
	wire [4-1:0] node3230;
	wire [4-1:0] node3232;
	wire [4-1:0] node3235;
	wire [4-1:0] node3236;
	wire [4-1:0] node3237;
	wire [4-1:0] node3241;
	wire [4-1:0] node3243;
	wire [4-1:0] node3246;
	wire [4-1:0] node3247;
	wire [4-1:0] node3248;
	wire [4-1:0] node3249;
	wire [4-1:0] node3250;
	wire [4-1:0] node3254;
	wire [4-1:0] node3255;
	wire [4-1:0] node3258;
	wire [4-1:0] node3261;
	wire [4-1:0] node3262;
	wire [4-1:0] node3263;
	wire [4-1:0] node3267;
	wire [4-1:0] node3268;
	wire [4-1:0] node3271;
	wire [4-1:0] node3274;
	wire [4-1:0] node3275;
	wire [4-1:0] node3276;
	wire [4-1:0] node3277;
	wire [4-1:0] node3280;
	wire [4-1:0] node3283;
	wire [4-1:0] node3285;
	wire [4-1:0] node3288;
	wire [4-1:0] node3289;
	wire [4-1:0] node3292;
	wire [4-1:0] node3293;
	wire [4-1:0] node3296;

	assign outp = (inp[0]) ? node1660 : node1;
		assign node1 = (inp[10]) ? node821 : node2;
			assign node2 = (inp[15]) ? node414 : node3;
				assign node3 = (inp[3]) ? node209 : node4;
					assign node4 = (inp[5]) ? node100 : node5;
						assign node5 = (inp[4]) ? node53 : node6;
							assign node6 = (inp[9]) ? node28 : node7;
								assign node7 = (inp[12]) ? node17 : node8;
									assign node8 = (inp[11]) ? 4'b1110 : node9;
										assign node9 = (inp[14]) ? node13 : node10;
											assign node10 = (inp[6]) ? 4'b1111 : 4'b1110;
											assign node13 = (inp[6]) ? 4'b1111 : 4'b0111;
									assign node17 = (inp[8]) ? node23 : node18;
										assign node18 = (inp[1]) ? node20 : 4'b0110;
											assign node20 = (inp[11]) ? 4'b0010 : 4'b1010;
										assign node23 = (inp[6]) ? 4'b1011 : node24;
											assign node24 = (inp[7]) ? 4'b0110 : 4'b1111;
								assign node28 = (inp[12]) ? node38 : node29;
									assign node29 = (inp[11]) ? 4'b0010 : node30;
										assign node30 = (inp[8]) ? node34 : node31;
											assign node31 = (inp[7]) ? 4'b0010 : 4'b1010;
											assign node34 = (inp[1]) ? 4'b1011 : 4'b0011;
									assign node38 = (inp[11]) ? node46 : node39;
										assign node39 = (inp[2]) ? node43 : node40;
											assign node40 = (inp[6]) ? 4'b0010 : 4'b1010;
											assign node43 = (inp[6]) ? 4'b1110 : 4'b0010;
										assign node46 = (inp[6]) ? node50 : node47;
											assign node47 = (inp[13]) ? 4'b1111 : 4'b1110;
											assign node50 = (inp[7]) ? 4'b0110 : 4'b1110;
							assign node53 = (inp[9]) ? node75 : node54;
								assign node54 = (inp[7]) ? node62 : node55;
									assign node55 = (inp[12]) ? node57 : 4'b1010;
										assign node57 = (inp[14]) ? 4'b1111 : node58;
											assign node58 = (inp[1]) ? 4'b1111 : 4'b0111;
									assign node62 = (inp[8]) ? node68 : node63;
										assign node63 = (inp[6]) ? 4'b0011 : node64;
											assign node64 = (inp[12]) ? 4'b0011 : 4'b1011;
										assign node68 = (inp[11]) ? node72 : node69;
											assign node69 = (inp[13]) ? 4'b0010 : 4'b0010;
											assign node72 = (inp[6]) ? 4'b0010 : 4'b1010;
								assign node75 = (inp[7]) ? node89 : node76;
									assign node76 = (inp[6]) ? node82 : node77;
										assign node77 = (inp[14]) ? node79 : 4'b1110;
											assign node79 = (inp[11]) ? 4'b1111 : 4'b0111;
										assign node82 = (inp[13]) ? node86 : node83;
											assign node83 = (inp[2]) ? 4'b0011 : 4'b0110;
											assign node86 = (inp[2]) ? 4'b0110 : 4'b0111;
									assign node89 = (inp[8]) ? node95 : node90;
										assign node90 = (inp[6]) ? 4'b1010 : node91;
											assign node91 = (inp[11]) ? 4'b0110 : 4'b1110;
										assign node95 = (inp[14]) ? node97 : 4'b0111;
											assign node97 = (inp[2]) ? 4'b0110 : 4'b0110;
						assign node100 = (inp[9]) ? node160 : node101;
							assign node101 = (inp[4]) ? node129 : node102;
								assign node102 = (inp[12]) ? node118 : node103;
									assign node103 = (inp[11]) ? node111 : node104;
										assign node104 = (inp[7]) ? node108 : node105;
											assign node105 = (inp[1]) ? 4'b1110 : 4'b1110;
											assign node108 = (inp[8]) ? 4'b1110 : 4'b1111;
										assign node111 = (inp[1]) ? node115 : node112;
											assign node112 = (inp[2]) ? 4'b0110 : 4'b1111;
											assign node115 = (inp[7]) ? 4'b0111 : 4'b0110;
									assign node118 = (inp[13]) ? node122 : node119;
										assign node119 = (inp[14]) ? 4'b0110 : 4'b0111;
										assign node122 = (inp[11]) ? node126 : node123;
											assign node123 = (inp[6]) ? 4'b1010 : 4'b0111;
											assign node126 = (inp[7]) ? 4'b0011 : 4'b1011;
								assign node129 = (inp[12]) ? node145 : node130;
									assign node130 = (inp[13]) ? node138 : node131;
										assign node131 = (inp[2]) ? node135 : node132;
											assign node132 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node135 = (inp[14]) ? 4'b1011 : 4'b1010;
										assign node138 = (inp[8]) ? node142 : node139;
											assign node139 = (inp[1]) ? 4'b0010 : 4'b1010;
											assign node142 = (inp[11]) ? 4'b0010 : 4'b0011;
									assign node145 = (inp[6]) ? node153 : node146;
										assign node146 = (inp[13]) ? node150 : node147;
											assign node147 = (inp[11]) ? 4'b0010 : 4'b1010;
											assign node150 = (inp[2]) ? 4'b0011 : 4'b1101;
										assign node153 = (inp[13]) ? node157 : node154;
											assign node154 = (inp[14]) ? 4'b0011 : 4'b0101;
											assign node157 = (inp[1]) ? 4'b1101 : 4'b1100;
							assign node160 = (inp[4]) ? node186 : node161;
								assign node161 = (inp[6]) ? node175 : node162;
									assign node162 = (inp[13]) ? node170 : node163;
										assign node163 = (inp[12]) ? node167 : node164;
											assign node164 = (inp[1]) ? 4'b1011 : 4'b1010;
											assign node167 = (inp[11]) ? 4'b0011 : 4'b1010;
										assign node170 = (inp[12]) ? node172 : 4'b0011;
											assign node172 = (inp[14]) ? 4'b1100 : 4'b0010;
									assign node175 = (inp[12]) ? node179 : node176;
										assign node176 = (inp[11]) ? 4'b0010 : 4'b0011;
										assign node179 = (inp[1]) ? node183 : node180;
											assign node180 = (inp[13]) ? 4'b1100 : 4'b0010;
											assign node183 = (inp[11]) ? 4'b0101 : 4'b1101;
								assign node186 = (inp[12]) ? node202 : node187;
									assign node187 = (inp[2]) ? node195 : node188;
										assign node188 = (inp[1]) ? node192 : node189;
											assign node189 = (inp[14]) ? 4'b0100 : 4'b1100;
											assign node192 = (inp[7]) ? 4'b0101 : 4'b0100;
										assign node195 = (inp[7]) ? node199 : node196;
											assign node196 = (inp[1]) ? 4'b1101 : 4'b0101;
											assign node199 = (inp[1]) ? 4'b1100 : 4'b1101;
									assign node202 = (inp[7]) ? node204 : 4'b0100;
										assign node204 = (inp[1]) ? 4'b1001 : node205;
											assign node205 = (inp[11]) ? 4'b0101 : 4'b1000;
					assign node209 = (inp[5]) ? node319 : node210;
						assign node210 = (inp[12]) ? node266 : node211;
							assign node211 = (inp[1]) ? node241 : node212;
								assign node212 = (inp[8]) ? node226 : node213;
									assign node213 = (inp[7]) ? node219 : node214;
										assign node214 = (inp[13]) ? node216 : 4'b1110;
											assign node216 = (inp[9]) ? 4'b0010 : 4'b0110;
										assign node219 = (inp[4]) ? node223 : node220;
											assign node220 = (inp[6]) ? 4'b0011 : 4'b1011;
											assign node223 = (inp[9]) ? 4'b1101 : 4'b1010;
									assign node226 = (inp[11]) ? node234 : node227;
										assign node227 = (inp[2]) ? node231 : node228;
											assign node228 = (inp[4]) ? 4'b0011 : 4'b1010;
											assign node231 = (inp[9]) ? 4'b1010 : 4'b1010;
										assign node234 = (inp[14]) ? node238 : node235;
											assign node235 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node238 = (inp[13]) ? 4'b1011 : 4'b0011;
								assign node241 = (inp[2]) ? node253 : node242;
									assign node242 = (inp[6]) ? node248 : node243;
										assign node243 = (inp[11]) ? 4'b1011 : node244;
											assign node244 = (inp[14]) ? 4'b0011 : 4'b0111;
										assign node248 = (inp[9]) ? 4'b0101 : node249;
											assign node249 = (inp[8]) ? 4'b1111 : 4'b0111;
									assign node253 = (inp[8]) ? node259 : node254;
										assign node254 = (inp[7]) ? node256 : 4'b0010;
											assign node256 = (inp[13]) ? 4'b0011 : 4'b1111;
										assign node259 = (inp[7]) ? node263 : node260;
											assign node260 = (inp[11]) ? 4'b1101 : 4'b0011;
											assign node263 = (inp[14]) ? 4'b0010 : 4'b0010;
							assign node266 = (inp[4]) ? node292 : node267;
								assign node267 = (inp[9]) ? node281 : node268;
									assign node268 = (inp[13]) ? node274 : node269;
										assign node269 = (inp[11]) ? node271 : 4'b1110;
											assign node271 = (inp[6]) ? 4'b1010 : 4'b1011;
										assign node274 = (inp[1]) ? node278 : node275;
											assign node275 = (inp[8]) ? 4'b0011 : 4'b0110;
											assign node278 = (inp[7]) ? 4'b1011 : 4'b1010;
									assign node281 = (inp[11]) ? node287 : node282;
										assign node282 = (inp[7]) ? 4'b0010 : node283;
											assign node283 = (inp[8]) ? 4'b0010 : 4'b1011;
										assign node287 = (inp[7]) ? node289 : 4'b1100;
											assign node289 = (inp[8]) ? 4'b1100 : 4'b0101;
								assign node292 = (inp[9]) ? node308 : node293;
									assign node293 = (inp[11]) ? node301 : node294;
										assign node294 = (inp[6]) ? node298 : node295;
											assign node295 = (inp[14]) ? 4'b0011 : 4'b0010;
											assign node298 = (inp[7]) ? 4'b1100 : 4'b0010;
										assign node301 = (inp[1]) ? node305 : node302;
											assign node302 = (inp[13]) ? 4'b1100 : 4'b0010;
											assign node305 = (inp[14]) ? 4'b1100 : 4'b0100;
									assign node308 = (inp[6]) ? node312 : node309;
										assign node309 = (inp[2]) ? 4'b0100 : 4'b1100;
										assign node312 = (inp[7]) ? node316 : node313;
											assign node313 = (inp[2]) ? 4'b1001 : 4'b0101;
											assign node316 = (inp[11]) ? 4'b0000 : 4'b1001;
						assign node319 = (inp[9]) ? node365 : node320;
							assign node320 = (inp[4]) ? node344 : node321;
								assign node321 = (inp[12]) ? node333 : node322;
									assign node322 = (inp[7]) ? node328 : node323;
										assign node323 = (inp[8]) ? node325 : 4'b0100;
											assign node325 = (inp[14]) ? 4'b1101 : 4'b0101;
										assign node328 = (inp[8]) ? 4'b0100 : node329;
											assign node329 = (inp[11]) ? 4'b0101 : 4'b1101;
									assign node333 = (inp[6]) ? node337 : node334;
										assign node334 = (inp[7]) ? 4'b0100 : 4'b1100;
										assign node337 = (inp[1]) ? node341 : node338;
											assign node338 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node341 = (inp[13]) ? 4'b0001 : 4'b0000;
								assign node344 = (inp[12]) ? node356 : node345;
									assign node345 = (inp[6]) ? node351 : node346;
										assign node346 = (inp[7]) ? 4'b1001 : node347;
											assign node347 = (inp[2]) ? 4'b1000 : 4'b0000;
										assign node351 = (inp[13]) ? 4'b0000 : node352;
											assign node352 = (inp[8]) ? 4'b0001 : 4'b0001;
									assign node356 = (inp[1]) ? 4'b1100 : node357;
										assign node357 = (inp[11]) ? node361 : node358;
											assign node358 = (inp[6]) ? 4'b1100 : 4'b0000;
											assign node361 = (inp[6]) ? 4'b0101 : 4'b0001;
							assign node365 = (inp[4]) ? node391 : node366;
								assign node366 = (inp[12]) ? node378 : node367;
									assign node367 = (inp[6]) ? node373 : node368;
										assign node368 = (inp[8]) ? 4'b0001 : node369;
											assign node369 = (inp[14]) ? 4'b1000 : 4'b1001;
										assign node373 = (inp[2]) ? 4'b0000 : node374;
											assign node374 = (inp[11]) ? 4'b1000 : 4'b0000;
									assign node378 = (inp[6]) ? node384 : node379;
										assign node379 = (inp[14]) ? 4'b1001 : node380;
											assign node380 = (inp[2]) ? 4'b0000 : 4'b0000;
										assign node384 = (inp[13]) ? node388 : node385;
											assign node385 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node388 = (inp[14]) ? 4'b0101 : 4'b1101;
								assign node391 = (inp[14]) ? node401 : node392;
									assign node392 = (inp[6]) ? node398 : node393;
										assign node393 = (inp[11]) ? 4'b1001 : node394;
											assign node394 = (inp[1]) ? 4'b1100 : 4'b1100;
										assign node398 = (inp[12]) ? 4'b1001 : 4'b1101;
									assign node401 = (inp[6]) ? node407 : node402;
										assign node402 = (inp[2]) ? node404 : 4'b1101;
											assign node404 = (inp[11]) ? 4'b0101 : 4'b0101;
										assign node407 = (inp[7]) ? node411 : node408;
											assign node408 = (inp[11]) ? 4'b1100 : 4'b0100;
											assign node411 = (inp[8]) ? 4'b0000 : 4'b0001;
				assign node414 = (inp[3]) ? node618 : node415;
					assign node415 = (inp[5]) ? node517 : node416;
						assign node416 = (inp[8]) ? node472 : node417;
							assign node417 = (inp[7]) ? node445 : node418;
								assign node418 = (inp[2]) ? node432 : node419;
									assign node419 = (inp[14]) ? node427 : node420;
										assign node420 = (inp[9]) ? node424 : node421;
											assign node421 = (inp[6]) ? 4'b1101 : 4'b1001;
											assign node424 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node427 = (inp[12]) ? node429 : 4'b1000;
											assign node429 = (inp[6]) ? 4'b0100 : 4'b1000;
									assign node432 = (inp[1]) ? node438 : node433;
										assign node433 = (inp[14]) ? node435 : 4'b0100;
											assign node435 = (inp[11]) ? 4'b0100 : 4'b0000;
										assign node438 = (inp[13]) ? node442 : node439;
											assign node439 = (inp[14]) ? 4'b1100 : 4'b0000;
											assign node442 = (inp[4]) ? 4'b1000 : 4'b0000;
								assign node445 = (inp[14]) ? node459 : node446;
									assign node446 = (inp[2]) ? node454 : node447;
										assign node447 = (inp[1]) ? node451 : node448;
											assign node448 = (inp[6]) ? 4'b1000 : 4'b1000;
											assign node451 = (inp[6]) ? 4'b1000 : 4'b1100;
										assign node454 = (inp[6]) ? 4'b0001 : node455;
											assign node455 = (inp[12]) ? 4'b0101 : 4'b0001;
									assign node459 = (inp[1]) ? node465 : node460;
										assign node460 = (inp[11]) ? node462 : 4'b0001;
											assign node462 = (inp[4]) ? 4'b1001 : 4'b0001;
										assign node465 = (inp[9]) ? node469 : node466;
											assign node466 = (inp[4]) ? 4'b1001 : 4'b0101;
											assign node469 = (inp[4]) ? 4'b1101 : 4'b0001;
							assign node472 = (inp[7]) ? node490 : node473;
								assign node473 = (inp[2]) ? node483 : node474;
									assign node474 = (inp[14]) ? node476 : 4'b0000;
										assign node476 = (inp[11]) ? node480 : node477;
											assign node477 = (inp[1]) ? 4'b1001 : 4'b0001;
											assign node480 = (inp[6]) ? 4'b0101 : 4'b1101;
									assign node483 = (inp[6]) ? 4'b0101 : node484;
										assign node484 = (inp[12]) ? 4'b1101 : node485;
											assign node485 = (inp[1]) ? 4'b1001 : 4'b1101;
								assign node490 = (inp[14]) ? node504 : node491;
									assign node491 = (inp[2]) ? node499 : node492;
										assign node492 = (inp[12]) ? node496 : node493;
											assign node493 = (inp[6]) ? 4'b0101 : 4'b1101;
											assign node496 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node499 = (inp[11]) ? node501 : 4'b1100;
											assign node501 = (inp[13]) ? 4'b0100 : 4'b0000;
									assign node504 = (inp[4]) ? node512 : node505;
										assign node505 = (inp[6]) ? node509 : node506;
											assign node506 = (inp[9]) ? 4'b0000 : 4'b0100;
											assign node509 = (inp[1]) ? 4'b1100 : 4'b1000;
										assign node512 = (inp[11]) ? 4'b0100 : node513;
											assign node513 = (inp[1]) ? 4'b0100 : 4'b1100;
						assign node517 = (inp[9]) ? node573 : node518;
							assign node518 = (inp[4]) ? node546 : node519;
								assign node519 = (inp[12]) ? node533 : node520;
									assign node520 = (inp[11]) ? node526 : node521;
										assign node521 = (inp[14]) ? 4'b1100 : node522;
											assign node522 = (inp[13]) ? 4'b1100 : 4'b0101;
										assign node526 = (inp[13]) ? node530 : node527;
											assign node527 = (inp[6]) ? 4'b0101 : 4'b0100;
											assign node530 = (inp[6]) ? 4'b0101 : 4'b1100;
									assign node533 = (inp[14]) ? node539 : node534;
										assign node534 = (inp[8]) ? 4'b1100 : node535;
											assign node535 = (inp[6]) ? 4'b0100 : 4'b0100;
										assign node539 = (inp[2]) ? node543 : node540;
											assign node540 = (inp[11]) ? 4'b1000 : 4'b1000;
											assign node543 = (inp[1]) ? 4'b1000 : 4'b0100;
								assign node546 = (inp[12]) ? node560 : node547;
									assign node547 = (inp[11]) ? node553 : node548;
										assign node548 = (inp[14]) ? 4'b1001 : node549;
											assign node549 = (inp[7]) ? 4'b0001 : 4'b0001;
										assign node553 = (inp[1]) ? node557 : node554;
											assign node554 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node557 = (inp[6]) ? 4'b0000 : 4'b1000;
									assign node560 = (inp[1]) ? node568 : node561;
										assign node561 = (inp[7]) ? node565 : node562;
											assign node562 = (inp[6]) ? 4'b0000 : 4'b1000;
											assign node565 = (inp[8]) ? 4'b0001 : 4'b1111;
										assign node568 = (inp[8]) ? 4'b0111 : node569;
											assign node569 = (inp[2]) ? 4'b1111 : 4'b1110;
							assign node573 = (inp[4]) ? node591 : node574;
								assign node574 = (inp[12]) ? node580 : node575;
									assign node575 = (inp[2]) ? 4'b1001 : node576;
										assign node576 = (inp[13]) ? 4'b1000 : 4'b0000;
									assign node580 = (inp[14]) ? node586 : node581;
										assign node581 = (inp[6]) ? 4'b1111 : node582;
											assign node582 = (inp[2]) ? 4'b1111 : 4'b1001;
										assign node586 = (inp[6]) ? 4'b0111 : node587;
											assign node587 = (inp[7]) ? 4'b1110 : 4'b1111;
								assign node591 = (inp[1]) ? node607 : node592;
									assign node592 = (inp[12]) ? node600 : node593;
										assign node593 = (inp[11]) ? node597 : node594;
											assign node594 = (inp[6]) ? 4'b0110 : 4'b0111;
											assign node597 = (inp[14]) ? 4'b1110 : 4'b1111;
										assign node600 = (inp[6]) ? node604 : node601;
											assign node601 = (inp[11]) ? 4'b0110 : 4'b1111;
											assign node604 = (inp[11]) ? 4'b1010 : 4'b0011;
									assign node607 = (inp[14]) ? node613 : node608;
										assign node608 = (inp[11]) ? node610 : 4'b0110;
											assign node610 = (inp[13]) ? 4'b0010 : 4'b0011;
										assign node613 = (inp[11]) ? node615 : 4'b0111;
											assign node615 = (inp[13]) ? 4'b0011 : 4'b0111;
					assign node618 = (inp[5]) ? node720 : node619;
						assign node619 = (inp[9]) ? node671 : node620;
							assign node620 = (inp[4]) ? node644 : node621;
								assign node621 = (inp[7]) ? node635 : node622;
									assign node622 = (inp[8]) ? node630 : node623;
										assign node623 = (inp[11]) ? node627 : node624;
											assign node624 = (inp[13]) ? 4'b0100 : 4'b1100;
											assign node627 = (inp[1]) ? 4'b1100 : 4'b0100;
										assign node630 = (inp[11]) ? 4'b0100 : node631;
											assign node631 = (inp[14]) ? 4'b1101 : 4'b1000;
									assign node635 = (inp[2]) ? 4'b0101 : node636;
										assign node636 = (inp[1]) ? node640 : node637;
											assign node637 = (inp[12]) ? 4'b1000 : 4'b1101;
											assign node640 = (inp[8]) ? 4'b0101 : 4'b0100;
								assign node644 = (inp[1]) ? node660 : node645;
									assign node645 = (inp[7]) ? node653 : node646;
										assign node646 = (inp[2]) ? node650 : node647;
											assign node647 = (inp[14]) ? 4'b1001 : 4'b1000;
											assign node650 = (inp[8]) ? 4'b0111 : 4'b0000;
										assign node653 = (inp[14]) ? node657 : node654;
											assign node654 = (inp[11]) ? 4'b1001 : 4'b0001;
											assign node657 = (inp[13]) ? 4'b0001 : 4'b0000;
									assign node660 = (inp[6]) ? node666 : node661;
										assign node661 = (inp[2]) ? node663 : 4'b0000;
											assign node663 = (inp[8]) ? 4'b1000 : 4'b1000;
										assign node666 = (inp[12]) ? node668 : 4'b0000;
											assign node668 = (inp[11]) ? 4'b0110 : 4'b1110;
							assign node671 = (inp[4]) ? node695 : node672;
								assign node672 = (inp[12]) ? node682 : node673;
									assign node673 = (inp[1]) ? node677 : node674;
										assign node674 = (inp[7]) ? 4'b1000 : 4'b0001;
										assign node677 = (inp[7]) ? 4'b0001 : node678;
											assign node678 = (inp[11]) ? 4'b0000 : 4'b1001;
									assign node682 = (inp[6]) ? node688 : node683;
										assign node683 = (inp[7]) ? 4'b1111 : node684;
											assign node684 = (inp[11]) ? 4'b0001 : 4'b1000;
										assign node688 = (inp[1]) ? node692 : node689;
											assign node689 = (inp[13]) ? 4'b0111 : 4'b1110;
											assign node692 = (inp[2]) ? 4'b0111 : 4'b1111;
								assign node695 = (inp[12]) ? node705 : node696;
									assign node696 = (inp[6]) ? node698 : 4'b1111;
										assign node698 = (inp[8]) ? node702 : node699;
											assign node699 = (inp[14]) ? 4'b0111 : 4'b0110;
											assign node702 = (inp[2]) ? 4'b0111 : 4'b0111;
									assign node705 = (inp[6]) ? node713 : node706;
										assign node706 = (inp[11]) ? node710 : node707;
											assign node707 = (inp[1]) ? 4'b0110 : 4'b1111;
											assign node710 = (inp[13]) ? 4'b1010 : 4'b0110;
										assign node713 = (inp[8]) ? node717 : node714;
											assign node714 = (inp[14]) ? 4'b0010 : 4'b1010;
											assign node717 = (inp[1]) ? 4'b0011 : 4'b0110;
						assign node720 = (inp[14]) ? node770 : node721;
							assign node721 = (inp[12]) ? node747 : node722;
								assign node722 = (inp[7]) ? node736 : node723;
									assign node723 = (inp[13]) ? node729 : node724;
										assign node724 = (inp[2]) ? node726 : 4'b1010;
											assign node726 = (inp[8]) ? 4'b0011 : 4'b0010;
										assign node729 = (inp[8]) ? node733 : node730;
											assign node730 = (inp[2]) ? 4'b1010 : 4'b0111;
											assign node733 = (inp[2]) ? 4'b1011 : 4'b1010;
									assign node736 = (inp[6]) ? node742 : node737;
										assign node737 = (inp[2]) ? node739 : 4'b1011;
											assign node739 = (inp[8]) ? 4'b0110 : 4'b0011;
										assign node742 = (inp[9]) ? 4'b0110 : node743;
											assign node743 = (inp[13]) ? 4'b0011 : 4'b0111;
								assign node747 = (inp[13]) ? node757 : node748;
									assign node748 = (inp[8]) ? node750 : 4'b0111;
										assign node750 = (inp[1]) ? node754 : node751;
											assign node751 = (inp[9]) ? 4'b0011 : 4'b0110;
											assign node754 = (inp[6]) ? 4'b0110 : 4'b0110;
									assign node757 = (inp[4]) ? node765 : node758;
										assign node758 = (inp[8]) ? node762 : node759;
											assign node759 = (inp[6]) ? 4'b1111 : 4'b1010;
											assign node762 = (inp[9]) ? 4'b0110 : 4'b0110;
										assign node765 = (inp[2]) ? node767 : 4'b1010;
											assign node767 = (inp[7]) ? 4'b0010 : 4'b0110;
							assign node770 = (inp[1]) ? node798 : node771;
								assign node771 = (inp[11]) ? node785 : node772;
									assign node772 = (inp[9]) ? node780 : node773;
										assign node773 = (inp[8]) ? node777 : node774;
											assign node774 = (inp[13]) ? 4'b1010 : 4'b1111;
											assign node777 = (inp[12]) ? 4'b0110 : 4'b0110;
										assign node780 = (inp[8]) ? node782 : 4'b1110;
											assign node782 = (inp[7]) ? 4'b1110 : 4'b1111;
									assign node785 = (inp[6]) ? node791 : node786;
										assign node786 = (inp[13]) ? 4'b1011 : node787;
											assign node787 = (inp[2]) ? 4'b0110 : 4'b0011;
										assign node791 = (inp[7]) ? node795 : node792;
											assign node792 = (inp[8]) ? 4'b0011 : 4'b1010;
											assign node795 = (inp[8]) ? 4'b1110 : 4'b1111;
								assign node798 = (inp[7]) ? node810 : node799;
									assign node799 = (inp[8]) ? node805 : node800;
										assign node800 = (inp[4]) ? node802 : 4'b0010;
											assign node802 = (inp[11]) ? 4'b0010 : 4'b0110;
										assign node805 = (inp[6]) ? 4'b1011 : node806;
											assign node806 = (inp[11]) ? 4'b1011 : 4'b0111;
									assign node810 = (inp[8]) ? node816 : node811;
										assign node811 = (inp[2]) ? node813 : 4'b1111;
											assign node813 = (inp[11]) ? 4'b0011 : 4'b1011;
										assign node816 = (inp[12]) ? 4'b0010 : node817;
											assign node817 = (inp[4]) ? 4'b1010 : 4'b1110;
			assign node821 = (inp[15]) ? node1235 : node822;
				assign node822 = (inp[3]) ? node1030 : node823;
					assign node823 = (inp[5]) ? node937 : node824;
						assign node824 = (inp[2]) ? node880 : node825;
							assign node825 = (inp[13]) ? node853 : node826;
								assign node826 = (inp[11]) ? node842 : node827;
									assign node827 = (inp[12]) ? node835 : node828;
										assign node828 = (inp[9]) ? node832 : node829;
											assign node829 = (inp[6]) ? 4'b1111 : 4'b1110;
											assign node832 = (inp[7]) ? 4'b0111 : 4'b0110;
										assign node835 = (inp[4]) ? node839 : node836;
											assign node836 = (inp[14]) ? 4'b0010 : 4'b0011;
											assign node839 = (inp[7]) ? 4'b0011 : 4'b1111;
									assign node842 = (inp[8]) ? node850 : node843;
										assign node843 = (inp[1]) ? node847 : node844;
											assign node844 = (inp[6]) ? 4'b1111 : 4'b0111;
											assign node847 = (inp[7]) ? 4'b0111 : 4'b0111;
										assign node850 = (inp[4]) ? 4'b0110 : 4'b0111;
								assign node853 = (inp[14]) ? node869 : node854;
									assign node854 = (inp[11]) ? node862 : node855;
										assign node855 = (inp[6]) ? node859 : node856;
											assign node856 = (inp[12]) ? 4'b0111 : 4'b0110;
											assign node859 = (inp[8]) ? 4'b1011 : 4'b1110;
										assign node862 = (inp[12]) ? node866 : node863;
											assign node863 = (inp[9]) ? 4'b0011 : 4'b0011;
											assign node866 = (inp[7]) ? 4'b1010 : 4'b0010;
									assign node869 = (inp[4]) ? node875 : node870;
										assign node870 = (inp[9]) ? node872 : 4'b0010;
											assign node872 = (inp[1]) ? 4'b1110 : 4'b0110;
										assign node875 = (inp[9]) ? 4'b1010 : node876;
											assign node876 = (inp[1]) ? 4'b1110 : 4'b1111;
							assign node880 = (inp[1]) ? node910 : node881;
								assign node881 = (inp[13]) ? node895 : node882;
									assign node882 = (inp[7]) ? node890 : node883;
										assign node883 = (inp[8]) ? node887 : node884;
											assign node884 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node887 = (inp[9]) ? 4'b1111 : 4'b0111;
										assign node890 = (inp[4]) ? node892 : 4'b1011;
											assign node892 = (inp[14]) ? 4'b1111 : 4'b1110;
									assign node895 = (inp[12]) ? node903 : node896;
										assign node896 = (inp[7]) ? node900 : node897;
											assign node897 = (inp[8]) ? 4'b0111 : 4'b0010;
											assign node900 = (inp[8]) ? 4'b1010 : 4'b0011;
										assign node903 = (inp[7]) ? node907 : node904;
											assign node904 = (inp[9]) ? 4'b1011 : 4'b0111;
											assign node907 = (inp[8]) ? 4'b0110 : 4'b1111;
								assign node910 = (inp[8]) ? node922 : node911;
									assign node911 = (inp[7]) ? node917 : node912;
										assign node912 = (inp[14]) ? 4'b0010 : node913;
											assign node913 = (inp[6]) ? 4'b1110 : 4'b0010;
										assign node917 = (inp[6]) ? 4'b0011 : node918;
											assign node918 = (inp[13]) ? 4'b0011 : 4'b1011;
									assign node922 = (inp[7]) ? node930 : node923;
										assign node923 = (inp[14]) ? node927 : node924;
											assign node924 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node927 = (inp[4]) ? 4'b1011 : 4'b0111;
										assign node930 = (inp[14]) ? node934 : node931;
											assign node931 = (inp[4]) ? 4'b0010 : 4'b1010;
											assign node934 = (inp[12]) ? 4'b0110 : 4'b1110;
						assign node937 = (inp[4]) ? node979 : node938;
							assign node938 = (inp[9]) ? node966 : node939;
								assign node939 = (inp[12]) ? node955 : node940;
									assign node940 = (inp[6]) ? node948 : node941;
										assign node941 = (inp[2]) ? node945 : node942;
											assign node942 = (inp[14]) ? 4'b1110 : 4'b0110;
											assign node945 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node948 = (inp[7]) ? node952 : node949;
											assign node949 = (inp[8]) ? 4'b1010 : 4'b0110;
											assign node952 = (inp[11]) ? 4'b0010 : 4'b1011;
									assign node955 = (inp[7]) ? node961 : node956;
										assign node956 = (inp[8]) ? 4'b1011 : node957;
											assign node957 = (inp[13]) ? 4'b1011 : 4'b0010;
										assign node961 = (inp[8]) ? 4'b0010 : node962;
											assign node962 = (inp[13]) ? 4'b1011 : 4'b0011;
								assign node966 = (inp[11]) ? 4'b1101 : node967;
									assign node967 = (inp[12]) ? node973 : node968;
										assign node968 = (inp[2]) ? 4'b0010 : node969;
											assign node969 = (inp[13]) ? 4'b1101 : 4'b1011;
										assign node973 = (inp[2]) ? node975 : 4'b1100;
											assign node975 = (inp[7]) ? 4'b0100 : 4'b0100;
							assign node979 = (inp[9]) ? node1003 : node980;
								assign node980 = (inp[12]) ? node992 : node981;
									assign node981 = (inp[11]) ? node987 : node982;
										assign node982 = (inp[1]) ? node984 : 4'b1010;
											assign node984 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node987 = (inp[7]) ? 4'b1100 : node988;
											assign node988 = (inp[13]) ? 4'b0100 : 4'b0010;
									assign node992 = (inp[14]) ? node998 : node993;
										assign node993 = (inp[2]) ? node995 : 4'b0100;
											assign node995 = (inp[8]) ? 4'b1100 : 4'b0100;
										assign node998 = (inp[6]) ? 4'b1100 : node999;
											assign node999 = (inp[8]) ? 4'b0101 : 4'b1100;
								assign node1003 = (inp[1]) ? node1017 : node1004;
									assign node1004 = (inp[12]) ? node1010 : node1005;
										assign node1005 = (inp[8]) ? 4'b1100 : node1006;
											assign node1006 = (inp[13]) ? 4'b0001 : 4'b0101;
										assign node1010 = (inp[6]) ? node1014 : node1011;
											assign node1011 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node1014 = (inp[13]) ? 4'b1001 : 4'b0001;
									assign node1017 = (inp[14]) ? node1025 : node1018;
										assign node1018 = (inp[8]) ? node1022 : node1019;
											assign node1019 = (inp[12]) ? 4'b0001 : 4'b1100;
											assign node1022 = (inp[2]) ? 4'b0001 : 4'b1000;
										assign node1025 = (inp[7]) ? 4'b1001 : node1026;
											assign node1026 = (inp[8]) ? 4'b1001 : 4'b1000;
					assign node1030 = (inp[5]) ? node1130 : node1031;
						assign node1031 = (inp[9]) ? node1081 : node1032;
							assign node1032 = (inp[4]) ? node1052 : node1033;
								assign node1033 = (inp[1]) ? node1041 : node1034;
									assign node1034 = (inp[12]) ? node1038 : node1035;
										assign node1035 = (inp[6]) ? 4'b0110 : 4'b1110;
										assign node1038 = (inp[7]) ? 4'b0011 : 4'b0010;
									assign node1041 = (inp[7]) ? node1049 : node1042;
										assign node1042 = (inp[13]) ? node1046 : node1043;
											assign node1043 = (inp[8]) ? 4'b1011 : 4'b0010;
											assign node1046 = (inp[11]) ? 4'b1011 : 4'b1010;
										assign node1049 = (inp[8]) ? 4'b0010 : 4'b0011;
								assign node1052 = (inp[6]) ? node1066 : node1053;
									assign node1053 = (inp[12]) ? node1059 : node1054;
										assign node1054 = (inp[7]) ? 4'b0010 : node1055;
											assign node1055 = (inp[13]) ? 4'b1100 : 4'b1010;
										assign node1059 = (inp[8]) ? node1063 : node1060;
											assign node1060 = (inp[7]) ? 4'b1101 : 4'b1100;
											assign node1063 = (inp[2]) ? 4'b1100 : 4'b0100;
									assign node1066 = (inp[13]) ? node1074 : node1067;
										assign node1067 = (inp[8]) ? node1071 : node1068;
											assign node1068 = (inp[7]) ? 4'b1101 : 4'b0100;
											assign node1071 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node1074 = (inp[7]) ? node1078 : node1075;
											assign node1075 = (inp[1]) ? 4'b1101 : 4'b1100;
											assign node1078 = (inp[11]) ? 4'b0100 : 4'b1100;
							assign node1081 = (inp[4]) ? node1105 : node1082;
								assign node1082 = (inp[14]) ? node1096 : node1083;
									assign node1083 = (inp[11]) ? node1091 : node1084;
										assign node1084 = (inp[12]) ? node1088 : node1085;
											assign node1085 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node1088 = (inp[13]) ? 4'b0101 : 4'b0100;
										assign node1091 = (inp[12]) ? 4'b0100 : node1092;
											assign node1092 = (inp[2]) ? 4'b1100 : 4'b0100;
									assign node1096 = (inp[1]) ? node1100 : node1097;
										assign node1097 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node1100 = (inp[12]) ? 4'b0100 : node1101;
											assign node1101 = (inp[7]) ? 4'b1101 : 4'b0100;
								assign node1105 = (inp[12]) ? node1117 : node1106;
									assign node1106 = (inp[11]) ? node1112 : node1107;
										assign node1107 = (inp[7]) ? 4'b0101 : node1108;
											assign node1108 = (inp[2]) ? 4'b1100 : 4'b0100;
										assign node1112 = (inp[2]) ? node1114 : 4'b0100;
											assign node1114 = (inp[6]) ? 4'b0001 : 4'b1000;
									assign node1117 = (inp[11]) ? node1123 : node1118;
										assign node1118 = (inp[6]) ? node1120 : 4'b0001;
											assign node1120 = (inp[13]) ? 4'b1001 : 4'b0000;
										assign node1123 = (inp[8]) ? node1127 : node1124;
											assign node1124 = (inp[1]) ? 4'b0000 : 4'b0000;
											assign node1127 = (inp[13]) ? 4'b0001 : 4'b1000;
						assign node1130 = (inp[4]) ? node1182 : node1131;
							assign node1131 = (inp[9]) ? node1157 : node1132;
								assign node1132 = (inp[12]) ? node1146 : node1133;
									assign node1133 = (inp[2]) ? node1141 : node1134;
										assign node1134 = (inp[14]) ? node1138 : node1135;
											assign node1135 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node1138 = (inp[7]) ? 4'b1001 : 4'b1000;
										assign node1141 = (inp[13]) ? node1143 : 4'b0000;
											assign node1143 = (inp[11]) ? 4'b0001 : 4'b0101;
									assign node1146 = (inp[13]) ? node1152 : node1147;
										assign node1147 = (inp[11]) ? 4'b0000 : node1148;
											assign node1148 = (inp[14]) ? 4'b0001 : 4'b1001;
										assign node1152 = (inp[14]) ? 4'b1001 : node1153;
											assign node1153 = (inp[7]) ? 4'b1001 : 4'b0001;
								assign node1157 = (inp[12]) ? node1171 : node1158;
									assign node1158 = (inp[8]) ? node1164 : node1159;
										assign node1159 = (inp[14]) ? node1161 : 4'b0001;
											assign node1161 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node1164 = (inp[1]) ? node1168 : node1165;
											assign node1165 = (inp[6]) ? 4'b1101 : 4'b0000;
											assign node1168 = (inp[2]) ? 4'b1100 : 4'b1101;
									assign node1171 = (inp[13]) ? node1177 : node1172;
										assign node1172 = (inp[8]) ? node1174 : 4'b0101;
											assign node1174 = (inp[11]) ? 4'b0100 : 4'b1100;
										assign node1177 = (inp[1]) ? 4'b1100 : node1178;
											assign node1178 = (inp[6]) ? 4'b0100 : 4'b0101;
							assign node1182 = (inp[9]) ? node1208 : node1183;
								assign node1183 = (inp[6]) ? node1195 : node1184;
									assign node1184 = (inp[12]) ? node1192 : node1185;
										assign node1185 = (inp[8]) ? node1189 : node1186;
											assign node1186 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node1189 = (inp[1]) ? 4'b0000 : 4'b1100;
										assign node1192 = (inp[8]) ? 4'b0101 : 4'b0100;
									assign node1195 = (inp[8]) ? node1203 : node1196;
										assign node1196 = (inp[7]) ? node1200 : node1197;
											assign node1197 = (inp[13]) ? 4'b0100 : 4'b0000;
											assign node1200 = (inp[12]) ? 4'b1101 : 4'b0101;
										assign node1203 = (inp[7]) ? node1205 : 4'b0101;
											assign node1205 = (inp[11]) ? 4'b0100 : 4'b1100;
								assign node1208 = (inp[12]) ? node1222 : node1209;
									assign node1209 = (inp[13]) ? node1215 : node1210;
										assign node1210 = (inp[11]) ? 4'b0100 : node1211;
											assign node1211 = (inp[6]) ? 4'b0100 : 4'b0101;
										assign node1215 = (inp[8]) ? node1219 : node1216;
											assign node1216 = (inp[2]) ? 4'b0100 : 4'b0000;
											assign node1219 = (inp[6]) ? 4'b0000 : 4'b1001;
									assign node1222 = (inp[6]) ? node1230 : node1223;
										assign node1223 = (inp[2]) ? node1227 : node1224;
											assign node1224 = (inp[14]) ? 4'b1001 : 4'b1000;
											assign node1227 = (inp[13]) ? 4'b1000 : 4'b0000;
										assign node1230 = (inp[13]) ? 4'b0001 : node1231;
											assign node1231 = (inp[14]) ? 4'b1000 : 4'b1001;
				assign node1235 = (inp[5]) ? node1449 : node1236;
					assign node1236 = (inp[3]) ? node1340 : node1237;
						assign node1237 = (inp[7]) ? node1285 : node1238;
							assign node1238 = (inp[8]) ? node1258 : node1239;
								assign node1239 = (inp[2]) ? node1249 : node1240;
									assign node1240 = (inp[14]) ? node1246 : node1241;
										assign node1241 = (inp[1]) ? 4'b0001 : node1242;
											assign node1242 = (inp[9]) ? 4'b0101 : 4'b1001;
										assign node1246 = (inp[1]) ? 4'b1100 : 4'b1000;
									assign node1249 = (inp[4]) ? node1255 : node1250;
										assign node1250 = (inp[6]) ? 4'b0000 : node1251;
											assign node1251 = (inp[11]) ? 4'b1000 : 4'b1100;
										assign node1255 = (inp[14]) ? 4'b1100 : 4'b0100;
								assign node1258 = (inp[2]) ? node1270 : node1259;
									assign node1259 = (inp[14]) ? node1265 : node1260;
										assign node1260 = (inp[11]) ? node1262 : 4'b1100;
											assign node1262 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node1265 = (inp[13]) ? node1267 : 4'b1101;
											assign node1267 = (inp[9]) ? 4'b0001 : 4'b1101;
									assign node1270 = (inp[1]) ? node1278 : node1271;
										assign node1271 = (inp[13]) ? node1275 : node1272;
											assign node1272 = (inp[6]) ? 4'b1001 : 4'b1101;
											assign node1275 = (inp[14]) ? 4'b1101 : 4'b0101;
										assign node1278 = (inp[9]) ? node1282 : node1279;
											assign node1279 = (inp[4]) ? 4'b1101 : 4'b0001;
											assign node1282 = (inp[11]) ? 4'b0101 : 4'b0001;
							assign node1285 = (inp[8]) ? node1311 : node1286;
								assign node1286 = (inp[14]) ? node1300 : node1287;
									assign node1287 = (inp[2]) ? node1295 : node1288;
										assign node1288 = (inp[6]) ? node1292 : node1289;
											assign node1289 = (inp[11]) ? 4'b0000 : 4'b1000;
											assign node1292 = (inp[1]) ? 4'b0100 : 4'b0000;
										assign node1295 = (inp[12]) ? node1297 : 4'b0001;
											assign node1297 = (inp[6]) ? 4'b1001 : 4'b0101;
									assign node1300 = (inp[9]) ? node1306 : node1301;
										assign node1301 = (inp[4]) ? node1303 : 4'b1001;
											assign node1303 = (inp[12]) ? 4'b1101 : 4'b0101;
										assign node1306 = (inp[2]) ? 4'b0101 : node1307;
											assign node1307 = (inp[1]) ? 4'b0001 : 4'b0001;
								assign node1311 = (inp[2]) ? node1327 : node1312;
									assign node1312 = (inp[14]) ? node1320 : node1313;
										assign node1313 = (inp[4]) ? node1317 : node1314;
											assign node1314 = (inp[6]) ? 4'b1101 : 4'b0101;
											assign node1317 = (inp[6]) ? 4'b0001 : 4'b0101;
										assign node1320 = (inp[13]) ? node1324 : node1321;
											assign node1321 = (inp[11]) ? 4'b0000 : 4'b0100;
											assign node1324 = (inp[6]) ? 4'b0100 : 4'b0100;
									assign node1327 = (inp[1]) ? node1333 : node1328;
										assign node1328 = (inp[14]) ? 4'b0100 : node1329;
											assign node1329 = (inp[9]) ? 4'b0000 : 4'b0100;
										assign node1333 = (inp[13]) ? node1337 : node1334;
											assign node1334 = (inp[11]) ? 4'b1000 : 4'b1100;
											assign node1337 = (inp[14]) ? 4'b0100 : 4'b0000;
						assign node1340 = (inp[9]) ? node1400 : node1341;
							assign node1341 = (inp[4]) ? node1371 : node1342;
								assign node1342 = (inp[12]) ? node1356 : node1343;
									assign node1343 = (inp[11]) ? node1349 : node1344;
										assign node1344 = (inp[8]) ? 4'b0101 : node1345;
											assign node1345 = (inp[6]) ? 4'b0100 : 4'b1100;
										assign node1349 = (inp[1]) ? node1353 : node1350;
											assign node1350 = (inp[2]) ? 4'b1000 : 4'b0100;
											assign node1353 = (inp[14]) ? 4'b1001 : 4'b0001;
									assign node1356 = (inp[14]) ? node1364 : node1357;
										assign node1357 = (inp[8]) ? node1361 : node1358;
											assign node1358 = (inp[1]) ? 4'b0000 : 4'b0000;
											assign node1361 = (inp[13]) ? 4'b1000 : 4'b1001;
										assign node1364 = (inp[11]) ? node1368 : node1365;
											assign node1365 = (inp[7]) ? 4'b1001 : 4'b0000;
											assign node1368 = (inp[8]) ? 4'b0000 : 4'b0001;
								assign node1371 = (inp[12]) ? node1387 : node1372;
									assign node1372 = (inp[7]) ? node1380 : node1373;
										assign node1373 = (inp[11]) ? node1377 : node1374;
											assign node1374 = (inp[1]) ? 4'b0000 : 4'b1000;
											assign node1377 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node1380 = (inp[1]) ? node1384 : node1381;
											assign node1381 = (inp[13]) ? 4'b0111 : 4'b0001;
											assign node1384 = (inp[8]) ? 4'b1110 : 4'b1111;
									assign node1387 = (inp[1]) ? node1395 : node1388;
										assign node1388 = (inp[6]) ? node1392 : node1389;
											assign node1389 = (inp[8]) ? 4'b0111 : 4'b0110;
											assign node1392 = (inp[11]) ? 4'b1111 : 4'b0110;
										assign node1395 = (inp[8]) ? node1397 : 4'b1111;
											assign node1397 = (inp[2]) ? 4'b1111 : 4'b0110;
							assign node1400 = (inp[4]) ? node1424 : node1401;
								assign node1401 = (inp[2]) ? node1413 : node1402;
									assign node1402 = (inp[8]) ? node1408 : node1403;
										assign node1403 = (inp[12]) ? 4'b0110 : node1404;
											assign node1404 = (inp[6]) ? 4'b1111 : 4'b1110;
										assign node1408 = (inp[14]) ? 4'b0111 : node1409;
											assign node1409 = (inp[6]) ? 4'b0111 : 4'b1111;
									assign node1413 = (inp[12]) ? node1417 : node1414;
										assign node1414 = (inp[11]) ? 4'b1110 : 4'b0000;
										assign node1417 = (inp[7]) ? node1421 : node1418;
											assign node1418 = (inp[8]) ? 4'b1111 : 4'b1110;
											assign node1421 = (inp[8]) ? 4'b0110 : 4'b0111;
								assign node1424 = (inp[6]) ? node1438 : node1425;
									assign node1425 = (inp[12]) ? node1433 : node1426;
										assign node1426 = (inp[11]) ? node1430 : node1427;
											assign node1427 = (inp[7]) ? 4'b0110 : 4'b1111;
											assign node1430 = (inp[14]) ? 4'b1010 : 4'b0110;
										assign node1433 = (inp[1]) ? node1435 : 4'b0010;
											assign node1435 = (inp[7]) ? 4'b1010 : 4'b0010;
									assign node1438 = (inp[8]) ? node1444 : node1439;
										assign node1439 = (inp[1]) ? 4'b1010 : node1440;
											assign node1440 = (inp[7]) ? 4'b1011 : 4'b1010;
										assign node1444 = (inp[13]) ? node1446 : 4'b0010;
											assign node1446 = (inp[7]) ? 4'b1010 : 4'b1011;
					assign node1449 = (inp[3]) ? node1553 : node1450;
						assign node1450 = (inp[9]) ? node1506 : node1451;
							assign node1451 = (inp[4]) ? node1477 : node1452;
								assign node1452 = (inp[12]) ? node1464 : node1453;
									assign node1453 = (inp[2]) ? node1459 : node1454;
										assign node1454 = (inp[6]) ? 4'b0001 : node1455;
											assign node1455 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node1459 = (inp[1]) ? node1461 : 4'b1100;
											assign node1461 = (inp[6]) ? 4'b0000 : 4'b1000;
									assign node1464 = (inp[8]) ? node1472 : node1465;
										assign node1465 = (inp[7]) ? node1469 : node1466;
											assign node1466 = (inp[13]) ? 4'b1000 : 4'b0000;
											assign node1469 = (inp[11]) ? 4'b0001 : 4'b1001;
										assign node1472 = (inp[13]) ? node1474 : 4'b0001;
											assign node1474 = (inp[11]) ? 4'b0001 : 4'b1000;
								assign node1477 = (inp[6]) ? node1491 : node1478;
									assign node1478 = (inp[8]) ? node1484 : node1479;
										assign node1479 = (inp[14]) ? 4'b0000 : node1480;
											assign node1480 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node1484 = (inp[11]) ? node1488 : node1485;
											assign node1485 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node1488 = (inp[1]) ? 4'b1110 : 4'b0111;
									assign node1491 = (inp[8]) ? node1499 : node1492;
										assign node1492 = (inp[12]) ? node1496 : node1493;
											assign node1493 = (inp[13]) ? 4'b0110 : 4'b0000;
											assign node1496 = (inp[7]) ? 4'b1110 : 4'b1110;
										assign node1499 = (inp[7]) ? node1503 : node1500;
											assign node1500 = (inp[2]) ? 4'b1111 : 4'b0110;
											assign node1503 = (inp[14]) ? 4'b1110 : 4'b1111;
							assign node1506 = (inp[4]) ? node1526 : node1507;
								assign node1507 = (inp[11]) ? node1513 : node1508;
									assign node1508 = (inp[12]) ? 4'b0110 : node1509;
										assign node1509 = (inp[1]) ? 4'b0001 : 4'b1000;
									assign node1513 = (inp[6]) ? node1521 : node1514;
										assign node1514 = (inp[12]) ? node1518 : node1515;
											assign node1515 = (inp[13]) ? 4'b1110 : 4'b1111;
											assign node1518 = (inp[7]) ? 4'b0110 : 4'b1111;
										assign node1521 = (inp[12]) ? 4'b1111 : node1522;
											assign node1522 = (inp[8]) ? 4'b0110 : 4'b0111;
								assign node1526 = (inp[6]) ? node1540 : node1527;
									assign node1527 = (inp[12]) ? node1535 : node1528;
										assign node1528 = (inp[14]) ? node1532 : node1529;
											assign node1529 = (inp[11]) ? 4'b1011 : 4'b1110;
											assign node1532 = (inp[1]) ? 4'b0111 : 4'b0110;
										assign node1535 = (inp[2]) ? 4'b1010 : node1536;
											assign node1536 = (inp[13]) ? 4'b0010 : 4'b0011;
									assign node1540 = (inp[11]) ? node1546 : node1541;
										assign node1541 = (inp[12]) ? 4'b0011 : node1542;
											assign node1542 = (inp[2]) ? 4'b1011 : 4'b1010;
										assign node1546 = (inp[13]) ? node1550 : node1547;
											assign node1547 = (inp[8]) ? 4'b0010 : 4'b1010;
											assign node1550 = (inp[14]) ? 4'b0010 : 4'b0011;
						assign node1553 = (inp[7]) ? node1607 : node1554;
							assign node1554 = (inp[6]) ? node1580 : node1555;
								assign node1555 = (inp[11]) ? node1567 : node1556;
									assign node1556 = (inp[8]) ? node1564 : node1557;
										assign node1557 = (inp[9]) ? node1561 : node1558;
											assign node1558 = (inp[13]) ? 4'b1010 : 4'b1110;
											assign node1561 = (inp[12]) ? 4'b0110 : 4'b1110;
										assign node1564 = (inp[2]) ? 4'b0111 : 4'b1110;
									assign node1567 = (inp[1]) ? node1575 : node1568;
										assign node1568 = (inp[13]) ? node1572 : node1569;
											assign node1569 = (inp[8]) ? 4'b0111 : 4'b0010;
											assign node1572 = (inp[12]) ? 4'b0111 : 4'b0110;
										assign node1575 = (inp[13]) ? node1577 : 4'b0011;
											assign node1577 = (inp[2]) ? 4'b1011 : 4'b1010;
								assign node1580 = (inp[4]) ? node1594 : node1581;
									assign node1581 = (inp[8]) ? node1587 : node1582;
										assign node1582 = (inp[12]) ? node1584 : 4'b0110;
											assign node1584 = (inp[13]) ? 4'b0110 : 4'b1110;
										assign node1587 = (inp[2]) ? node1591 : node1588;
											assign node1588 = (inp[14]) ? 4'b1011 : 4'b0010;
											assign node1591 = (inp[9]) ? 4'b0111 : 4'b0111;
									assign node1594 = (inp[2]) ? node1602 : node1595;
										assign node1595 = (inp[1]) ? node1599 : node1596;
											assign node1596 = (inp[11]) ? 4'b1111 : 4'b0111;
											assign node1599 = (inp[8]) ? 4'b0111 : 4'b0011;
										assign node1602 = (inp[9]) ? node1604 : 4'b1111;
											assign node1604 = (inp[14]) ? 4'b1011 : 4'b1010;
							assign node1607 = (inp[8]) ? node1635 : node1608;
								assign node1608 = (inp[2]) ? node1620 : node1609;
									assign node1609 = (inp[14]) ? node1615 : node1610;
										assign node1610 = (inp[1]) ? 4'b0010 : node1611;
											assign node1611 = (inp[12]) ? 4'b1110 : 4'b0010;
										assign node1615 = (inp[6]) ? 4'b1111 : node1616;
											assign node1616 = (inp[4]) ? 4'b0011 : 4'b0111;
									assign node1620 = (inp[6]) ? node1628 : node1621;
										assign node1621 = (inp[11]) ? node1625 : node1622;
											assign node1622 = (inp[1]) ? 4'b0011 : 4'b0111;
											assign node1625 = (inp[4]) ? 4'b0011 : 4'b1011;
										assign node1628 = (inp[1]) ? node1632 : node1629;
											assign node1629 = (inp[9]) ? 4'b1111 : 4'b0111;
											assign node1632 = (inp[13]) ? 4'b0011 : 4'b0111;
								assign node1635 = (inp[14]) ? node1645 : node1636;
									assign node1636 = (inp[2]) ? node1642 : node1637;
										assign node1637 = (inp[1]) ? 4'b0111 : node1638;
											assign node1638 = (inp[13]) ? 4'b1011 : 4'b0011;
										assign node1642 = (inp[4]) ? 4'b1010 : 4'b0010;
									assign node1645 = (inp[4]) ? node1653 : node1646;
										assign node1646 = (inp[2]) ? node1650 : node1647;
											assign node1647 = (inp[12]) ? 4'b1110 : 4'b1010;
											assign node1650 = (inp[9]) ? 4'b0110 : 4'b0010;
										assign node1653 = (inp[9]) ? node1657 : node1654;
											assign node1654 = (inp[12]) ? 4'b0110 : 4'b0010;
											assign node1657 = (inp[12]) ? 4'b0010 : 4'b0010;
		assign node1660 = (inp[7]) ? node2506 : node1661;
			assign node1661 = (inp[8]) ? node2071 : node1662;
				assign node1662 = (inp[2]) ? node1874 : node1663;
					assign node1663 = (inp[14]) ? node1775 : node1664;
						assign node1664 = (inp[3]) ? node1724 : node1665;
							assign node1665 = (inp[15]) ? node1697 : node1666;
								assign node1666 = (inp[9]) ? node1682 : node1667;
									assign node1667 = (inp[13]) ? node1675 : node1668;
										assign node1668 = (inp[6]) ? node1672 : node1669;
											assign node1669 = (inp[10]) ? 4'b0101 : 4'b0001;
											assign node1672 = (inp[11]) ? 4'b1001 : 4'b0001;
										assign node1675 = (inp[11]) ? node1679 : node1676;
											assign node1676 = (inp[1]) ? 4'b1101 : 4'b1001;
											assign node1679 = (inp[6]) ? 4'b0001 : 4'b1001;
									assign node1682 = (inp[5]) ? node1690 : node1683;
										assign node1683 = (inp[11]) ? node1687 : node1684;
											assign node1684 = (inp[6]) ? 4'b0101 : 4'b1001;
											assign node1687 = (inp[12]) ? 4'b0001 : 4'b0101;
										assign node1690 = (inp[11]) ? node1694 : node1691;
											assign node1691 = (inp[13]) ? 4'b0011 : 4'b0001;
											assign node1694 = (inp[12]) ? 4'b0111 : 4'b0001;
								assign node1697 = (inp[5]) ? node1711 : node1698;
									assign node1698 = (inp[4]) ? node1704 : node1699;
										assign node1699 = (inp[13]) ? node1701 : 4'b0111;
											assign node1701 = (inp[10]) ? 4'b0011 : 4'b0111;
										assign node1704 = (inp[11]) ? node1708 : node1705;
											assign node1705 = (inp[9]) ? 4'b0111 : 4'b0011;
											assign node1708 = (inp[12]) ? 4'b1011 : 4'b1111;
									assign node1711 = (inp[1]) ? node1719 : node1712;
										assign node1712 = (inp[10]) ? node1716 : node1713;
											assign node1713 = (inp[4]) ? 4'b0101 : 4'b0011;
											assign node1716 = (inp[6]) ? 4'b1101 : 4'b0111;
										assign node1719 = (inp[11]) ? 4'b1111 : node1720;
											assign node1720 = (inp[13]) ? 4'b1011 : 4'b0011;
							assign node1724 = (inp[15]) ? node1750 : node1725;
								assign node1725 = (inp[5]) ? node1737 : node1726;
									assign node1726 = (inp[6]) ? node1732 : node1727;
										assign node1727 = (inp[4]) ? 4'b0001 : node1728;
											assign node1728 = (inp[13]) ? 4'b1001 : 4'b1101;
										assign node1732 = (inp[11]) ? node1734 : 4'b0101;
											assign node1734 = (inp[1]) ? 4'b0111 : 4'b1111;
									assign node1737 = (inp[6]) ? node1745 : node1738;
										assign node1738 = (inp[13]) ? node1742 : node1739;
											assign node1739 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node1742 = (inp[1]) ? 4'b1111 : 4'b0111;
										assign node1745 = (inp[12]) ? 4'b0011 : node1746;
											assign node1746 = (inp[1]) ? 4'b1011 : 4'b1111;
								assign node1750 = (inp[5]) ? node1762 : node1751;
									assign node1751 = (inp[12]) ? node1757 : node1752;
										assign node1752 = (inp[4]) ? 4'b0011 : node1753;
											assign node1753 = (inp[9]) ? 4'b1011 : 4'b1111;
										assign node1757 = (inp[11]) ? node1759 : 4'b0101;
											assign node1759 = (inp[4]) ? 4'b1001 : 4'b0011;
									assign node1762 = (inp[10]) ? node1770 : node1763;
										assign node1763 = (inp[4]) ? node1767 : node1764;
											assign node1764 = (inp[11]) ? 4'b1001 : 4'b0101;
											assign node1767 = (inp[12]) ? 4'b0101 : 4'b1101;
										assign node1770 = (inp[6]) ? 4'b0001 : node1771;
											assign node1771 = (inp[12]) ? 4'b0101 : 4'b1101;
						assign node1775 = (inp[6]) ? node1827 : node1776;
							assign node1776 = (inp[13]) ? node1798 : node1777;
								assign node1777 = (inp[11]) ? node1789 : node1778;
									assign node1778 = (inp[5]) ? node1782 : node1779;
										assign node1779 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node1782 = (inp[15]) ? node1786 : node1783;
											assign node1783 = (inp[3]) ? 4'b1010 : 4'b1110;
											assign node1786 = (inp[1]) ? 4'b1100 : 4'b1100;
									assign node1789 = (inp[15]) ? node1795 : node1790;
										assign node1790 = (inp[10]) ? 4'b0100 : node1791;
											assign node1791 = (inp[5]) ? 4'b0100 : 4'b0000;
										assign node1795 = (inp[9]) ? 4'b0000 : 4'b0010;
								assign node1798 = (inp[12]) ? node1812 : node1799;
									assign node1799 = (inp[15]) ? node1807 : node1800;
										assign node1800 = (inp[3]) ? node1804 : node1801;
											assign node1801 = (inp[4]) ? 4'b1000 : 4'b0000;
											assign node1804 = (inp[5]) ? 4'b0010 : 4'b0000;
										assign node1807 = (inp[4]) ? 4'b0100 : node1808;
											assign node1808 = (inp[3]) ? 4'b1100 : 4'b1010;
									assign node1812 = (inp[5]) ? node1820 : node1813;
										assign node1813 = (inp[10]) ? node1817 : node1814;
											assign node1814 = (inp[9]) ? 4'b1110 : 4'b0100;
											assign node1817 = (inp[3]) ? 4'b0100 : 4'b0010;
										assign node1820 = (inp[4]) ? node1824 : node1821;
											assign node1821 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node1824 = (inp[11]) ? 4'b1000 : 4'b0100;
							assign node1827 = (inp[11]) ? node1857 : node1828;
								assign node1828 = (inp[13]) ? node1844 : node1829;
									assign node1829 = (inp[3]) ? node1837 : node1830;
										assign node1830 = (inp[9]) ? node1834 : node1831;
											assign node1831 = (inp[15]) ? 4'b0110 : 4'b0100;
											assign node1834 = (inp[12]) ? 4'b0110 : 4'b0010;
										assign node1837 = (inp[15]) ? node1841 : node1838;
											assign node1838 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node1841 = (inp[9]) ? 4'b0000 : 4'b0100;
									assign node1844 = (inp[1]) ? node1850 : node1845;
										assign node1845 = (inp[3]) ? node1847 : 4'b0000;
											assign node1847 = (inp[5]) ? 4'b0110 : 4'b0010;
										assign node1850 = (inp[3]) ? node1854 : node1851;
											assign node1851 = (inp[12]) ? 4'b1110 : 4'b1010;
											assign node1854 = (inp[12]) ? 4'b1000 : 4'b1010;
								assign node1857 = (inp[13]) ? node1865 : node1858;
									assign node1858 = (inp[3]) ? node1862 : node1859;
										assign node1859 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node1862 = (inp[15]) ? 4'b1100 : 4'b1010;
									assign node1865 = (inp[1]) ? node1867 : 4'b1100;
										assign node1867 = (inp[12]) ? node1871 : node1868;
											assign node1868 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node1871 = (inp[4]) ? 4'b0100 : 4'b0000;
					assign node1874 = (inp[1]) ? node1968 : node1875;
						assign node1875 = (inp[3]) ? node1917 : node1876;
							assign node1876 = (inp[15]) ? node1900 : node1877;
								assign node1877 = (inp[6]) ? node1889 : node1878;
									assign node1878 = (inp[11]) ? node1882 : node1879;
										assign node1879 = (inp[14]) ? 4'b1100 : 4'b1000;
										assign node1882 = (inp[13]) ? node1886 : node1883;
											assign node1883 = (inp[14]) ? 4'b0000 : 4'b0100;
											assign node1886 = (inp[5]) ? 4'b0110 : 4'b0100;
									assign node1889 = (inp[5]) ? node1895 : node1890;
										assign node1890 = (inp[12]) ? node1892 : 4'b0100;
											assign node1892 = (inp[4]) ? 4'b0000 : 4'b0000;
										assign node1895 = (inp[12]) ? node1897 : 4'b0000;
											assign node1897 = (inp[4]) ? 4'b0010 : 4'b0000;
								assign node1900 = (inp[6]) ? node1910 : node1901;
									assign node1901 = (inp[11]) ? node1903 : 4'b1110;
										assign node1903 = (inp[9]) ? node1907 : node1904;
											assign node1904 = (inp[14]) ? 4'b0010 : 4'b0010;
											assign node1907 = (inp[13]) ? 4'b0100 : 4'b0000;
									assign node1910 = (inp[11]) ? node1912 : 4'b0010;
										assign node1912 = (inp[10]) ? 4'b1010 : node1913;
											assign node1913 = (inp[4]) ? 4'b1100 : 4'b1010;
							assign node1917 = (inp[15]) ? node1941 : node1918;
								assign node1918 = (inp[4]) ? node1928 : node1919;
									assign node1919 = (inp[5]) ? 4'b1010 : node1920;
										assign node1920 = (inp[9]) ? node1924 : node1921;
											assign node1921 = (inp[12]) ? 4'b0000 : 4'b0100;
											assign node1924 = (inp[13]) ? 4'b0000 : 4'b0000;
									assign node1928 = (inp[14]) ? node1934 : node1929;
										assign node1929 = (inp[9]) ? node1931 : 4'b0010;
											assign node1931 = (inp[11]) ? 4'b0110 : 4'b0110;
										assign node1934 = (inp[6]) ? node1938 : node1935;
											assign node1935 = (inp[5]) ? 4'b1110 : 4'b0000;
											assign node1938 = (inp[10]) ? 4'b1110 : 4'b1010;
								assign node1941 = (inp[5]) ? node1955 : node1942;
									assign node1942 = (inp[4]) ? node1950 : node1943;
										assign node1943 = (inp[13]) ? node1947 : node1944;
											assign node1944 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node1947 = (inp[6]) ? 4'b1100 : 4'b1110;
										assign node1950 = (inp[6]) ? node1952 : 4'b1100;
											assign node1952 = (inp[12]) ? 4'b0000 : 4'b0100;
									assign node1955 = (inp[4]) ? node1963 : node1956;
										assign node1956 = (inp[10]) ? node1960 : node1957;
											assign node1957 = (inp[11]) ? 4'b1100 : 4'b1000;
											assign node1960 = (inp[14]) ? 4'b0100 : 4'b0000;
										assign node1963 = (inp[13]) ? 4'b0000 : node1964;
											assign node1964 = (inp[10]) ? 4'b0100 : 4'b0100;
						assign node1968 = (inp[15]) ? node2018 : node1969;
							assign node1969 = (inp[3]) ? node1995 : node1970;
								assign node1970 = (inp[11]) ? node1984 : node1971;
									assign node1971 = (inp[13]) ? node1977 : node1972;
										assign node1972 = (inp[6]) ? 4'b0000 : node1973;
											assign node1973 = (inp[10]) ? 4'b1000 : 4'b1000;
										assign node1977 = (inp[5]) ? node1981 : node1978;
											assign node1978 = (inp[10]) ? 4'b0100 : 4'b0000;
											assign node1981 = (inp[10]) ? 4'b1110 : 4'b1100;
									assign node1984 = (inp[13]) ? node1990 : node1985;
										assign node1985 = (inp[9]) ? node1987 : 4'b0100;
											assign node1987 = (inp[14]) ? 4'b1100 : 4'b1110;
										assign node1990 = (inp[6]) ? node1992 : 4'b1100;
											assign node1992 = (inp[5]) ? 4'b0000 : 4'b0100;
								assign node1995 = (inp[5]) ? node2007 : node1996;
									assign node1996 = (inp[4]) ? node2002 : node1997;
										assign node1997 = (inp[6]) ? node1999 : 4'b0100;
											assign node1999 = (inp[14]) ? 4'b0100 : 4'b0000;
										assign node2002 = (inp[12]) ? node2004 : 4'b1110;
											assign node2004 = (inp[6]) ? 4'b0010 : 4'b1010;
									assign node2007 = (inp[9]) ? node2011 : node2008;
										assign node2008 = (inp[4]) ? 4'b1110 : 4'b1010;
										assign node2011 = (inp[11]) ? node2015 : node2012;
											assign node2012 = (inp[14]) ? 4'b0110 : 4'b1010;
											assign node2015 = (inp[4]) ? 4'b0010 : 4'b0010;
							assign node2018 = (inp[3]) ? node2042 : node2019;
								assign node2019 = (inp[12]) ? node2031 : node2020;
									assign node2020 = (inp[6]) ? node2026 : node2021;
										assign node2021 = (inp[11]) ? node2023 : 4'b0010;
											assign node2023 = (inp[13]) ? 4'b1010 : 4'b0010;
										assign node2026 = (inp[10]) ? node2028 : 4'b1010;
											assign node2028 = (inp[4]) ? 4'b1000 : 4'b1010;
									assign node2031 = (inp[11]) ? node2037 : node2032;
										assign node2032 = (inp[13]) ? 4'b1110 : node2033;
											assign node2033 = (inp[14]) ? 4'b1010 : 4'b1010;
										assign node2037 = (inp[6]) ? 4'b0000 : node2038;
											assign node2038 = (inp[9]) ? 4'b1110 : 4'b1100;
								assign node2042 = (inp[5]) ? node2056 : node2043;
									assign node2043 = (inp[9]) ? node2049 : node2044;
										assign node2044 = (inp[12]) ? node2046 : 4'b1010;
											assign node2046 = (inp[6]) ? 4'b1100 : 4'b0010;
										assign node2049 = (inp[13]) ? node2053 : node2050;
											assign node2050 = (inp[10]) ? 4'b0100 : 4'b1010;
											assign node2053 = (inp[4]) ? 4'b1000 : 4'b1100;
									assign node2056 = (inp[6]) ? node2064 : node2057;
										assign node2057 = (inp[14]) ? node2061 : node2058;
											assign node2058 = (inp[10]) ? 4'b1000 : 4'b1100;
											assign node2061 = (inp[10]) ? 4'b0000 : 4'b1000;
										assign node2064 = (inp[13]) ? node2068 : node2065;
											assign node2065 = (inp[11]) ? 4'b1100 : 4'b0000;
											assign node2068 = (inp[4]) ? 4'b0000 : 4'b0000;
				assign node2071 = (inp[14]) ? node2297 : node2072;
					assign node2072 = (inp[2]) ? node2184 : node2073;
						assign node2073 = (inp[12]) ? node2129 : node2074;
							assign node2074 = (inp[11]) ? node2102 : node2075;
								assign node2075 = (inp[6]) ? node2089 : node2076;
									assign node2076 = (inp[1]) ? node2084 : node2077;
										assign node2077 = (inp[13]) ? node2081 : node2078;
											assign node2078 = (inp[4]) ? 4'b1110 : 4'b1100;
											assign node2081 = (inp[5]) ? 4'b1000 : 4'b1000;
										assign node2084 = (inp[13]) ? 4'b0000 : node2085;
											assign node2085 = (inp[5]) ? 4'b1100 : 4'b1000;
									assign node2089 = (inp[1]) ? node2097 : node2090;
										assign node2090 = (inp[9]) ? node2094 : node2091;
											assign node2091 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node2094 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node2097 = (inp[15]) ? 4'b1010 : node2098;
											assign node2098 = (inp[13]) ? 4'b1100 : 4'b0000;
								assign node2102 = (inp[6]) ? node2116 : node2103;
									assign node2103 = (inp[1]) ? node2111 : node2104;
										assign node2104 = (inp[10]) ? node2108 : node2105;
											assign node2105 = (inp[9]) ? 4'b0000 : 4'b0010;
											assign node2108 = (inp[9]) ? 4'b0110 : 4'b0000;
										assign node2111 = (inp[13]) ? 4'b1110 : node2112;
											assign node2112 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node2116 = (inp[1]) ? node2122 : node2117;
										assign node2117 = (inp[5]) ? node2119 : 4'b1110;
											assign node2119 = (inp[15]) ? 4'b1100 : 4'b1000;
										assign node2122 = (inp[9]) ? node2126 : node2123;
											assign node2123 = (inp[5]) ? 4'b0000 : 4'b0100;
											assign node2126 = (inp[13]) ? 4'b0010 : 4'b1010;
							assign node2129 = (inp[10]) ? node2161 : node2130;
								assign node2130 = (inp[6]) ? node2146 : node2131;
									assign node2131 = (inp[4]) ? node2139 : node2132;
										assign node2132 = (inp[11]) ? node2136 : node2133;
											assign node2133 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node2136 = (inp[13]) ? 4'b1100 : 4'b0100;
										assign node2139 = (inp[9]) ? node2143 : node2140;
											assign node2140 = (inp[11]) ? 4'b0010 : 4'b0000;
											assign node2143 = (inp[1]) ? 4'b1010 : 4'b0110;
									assign node2146 = (inp[11]) ? node2154 : node2147;
										assign node2147 = (inp[3]) ? node2151 : node2148;
											assign node2148 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node2151 = (inp[5]) ? 4'b0110 : 4'b0100;
										assign node2154 = (inp[1]) ? node2158 : node2155;
											assign node2155 = (inp[13]) ? 4'b1110 : 4'b1000;
											assign node2158 = (inp[3]) ? 4'b1110 : 4'b0110;
								assign node2161 = (inp[15]) ? node2169 : node2162;
									assign node2162 = (inp[9]) ? 4'b1010 : node2163;
										assign node2163 = (inp[3]) ? node2165 : 4'b1000;
											assign node2165 = (inp[4]) ? 4'b0110 : 4'b0010;
									assign node2169 = (inp[5]) ? node2177 : node2170;
										assign node2170 = (inp[13]) ? node2174 : node2171;
											assign node2171 = (inp[11]) ? 4'b0010 : 4'b0010;
											assign node2174 = (inp[3]) ? 4'b0000 : 4'b1110;
										assign node2177 = (inp[13]) ? node2181 : node2178;
											assign node2178 = (inp[11]) ? 4'b0000 : 4'b0000;
											assign node2181 = (inp[6]) ? 4'b0100 : 4'b0000;
						assign node2184 = (inp[11]) ? node2238 : node2185;
							assign node2185 = (inp[6]) ? node2209 : node2186;
								assign node2186 = (inp[13]) ? node2200 : node2187;
									assign node2187 = (inp[1]) ? node2195 : node2188;
										assign node2188 = (inp[10]) ? node2192 : node2189;
											assign node2189 = (inp[5]) ? 4'b1101 : 4'b1001;
											assign node2192 = (inp[15]) ? 4'b1011 : 4'b1001;
										assign node2195 = (inp[10]) ? node2197 : 4'b0101;
											assign node2197 = (inp[9]) ? 4'b0001 : 4'b0011;
									assign node2200 = (inp[4]) ? node2206 : node2201;
										assign node2201 = (inp[1]) ? 4'b0101 : node2202;
											assign node2202 = (inp[5]) ? 4'b0001 : 4'b0101;
										assign node2206 = (inp[3]) ? 4'b0101 : 4'b0111;
								assign node2209 = (inp[1]) ? node2225 : node2210;
									assign node2210 = (inp[13]) ? node2218 : node2211;
										assign node2211 = (inp[5]) ? node2215 : node2212;
											assign node2212 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node2215 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node2218 = (inp[5]) ? node2222 : node2219;
											assign node2219 = (inp[15]) ? 4'b1001 : 4'b1001;
											assign node2222 = (inp[9]) ? 4'b1111 : 4'b1011;
									assign node2225 = (inp[15]) ? node2231 : node2226;
										assign node2226 = (inp[10]) ? node2228 : 4'b1111;
											assign node2228 = (inp[4]) ? 4'b1011 : 4'b1001;
										assign node2231 = (inp[3]) ? node2235 : node2232;
											assign node2232 = (inp[10]) ? 4'b1101 : 4'b1011;
											assign node2235 = (inp[4]) ? 4'b1101 : 4'b1001;
							assign node2238 = (inp[6]) ? node2268 : node2239;
								assign node2239 = (inp[13]) ? node2253 : node2240;
									assign node2240 = (inp[1]) ? node2248 : node2241;
										assign node2241 = (inp[5]) ? node2245 : node2242;
											assign node2242 = (inp[10]) ? 4'b0011 : 4'b0111;
											assign node2245 = (inp[9]) ? 4'b0001 : 4'b0101;
										assign node2248 = (inp[15]) ? node2250 : 4'b1111;
											assign node2250 = (inp[4]) ? 4'b1011 : 4'b1001;
									assign node2253 = (inp[12]) ? node2261 : node2254;
										assign node2254 = (inp[3]) ? node2258 : node2255;
											assign node2255 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node2258 = (inp[15]) ? 4'b1001 : 4'b1001;
										assign node2261 = (inp[1]) ? node2265 : node2262;
											assign node2262 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node2265 = (inp[5]) ? 4'b1001 : 4'b1101;
								assign node2268 = (inp[1]) ? node2282 : node2269;
									assign node2269 = (inp[13]) ? node2277 : node2270;
										assign node2270 = (inp[15]) ? node2274 : node2271;
											assign node2271 = (inp[10]) ? 4'b1001 : 4'b1001;
											assign node2274 = (inp[10]) ? 4'b1101 : 4'b1011;
										assign node2277 = (inp[9]) ? 4'b0001 : node2278;
											assign node2278 = (inp[5]) ? 4'b0001 : 4'b0101;
									assign node2282 = (inp[4]) ? node2290 : node2283;
										assign node2283 = (inp[15]) ? node2287 : node2284;
											assign node2284 = (inp[3]) ? 4'b0101 : 4'b0001;
											assign node2287 = (inp[5]) ? 4'b0001 : 4'b0011;
										assign node2290 = (inp[13]) ? node2294 : node2291;
											assign node2291 = (inp[12]) ? 4'b0001 : 4'b0001;
											assign node2294 = (inp[15]) ? 4'b0001 : 4'b0011;
					assign node2297 = (inp[11]) ? node2395 : node2298;
						assign node2298 = (inp[6]) ? node2350 : node2299;
							assign node2299 = (inp[13]) ? node2325 : node2300;
								assign node2300 = (inp[1]) ? node2312 : node2301;
									assign node2301 = (inp[2]) ? node2307 : node2302;
										assign node2302 = (inp[15]) ? node2304 : 4'b1101;
											assign node2304 = (inp[9]) ? 4'b1011 : 4'b1111;
										assign node2307 = (inp[3]) ? 4'b1001 : node2308;
											assign node2308 = (inp[4]) ? 4'b1001 : 4'b1101;
									assign node2312 = (inp[9]) ? node2320 : node2313;
										assign node2313 = (inp[4]) ? node2317 : node2314;
											assign node2314 = (inp[3]) ? 4'b0101 : 4'b0101;
											assign node2317 = (inp[3]) ? 4'b0011 : 4'b0001;
										assign node2320 = (inp[10]) ? 4'b0111 : node2321;
											assign node2321 = (inp[2]) ? 4'b0111 : 4'b0101;
								assign node2325 = (inp[4]) ? node2339 : node2326;
									assign node2326 = (inp[10]) ? node2332 : node2327;
										assign node2327 = (inp[9]) ? node2329 : 4'b0111;
											assign node2329 = (inp[5]) ? 4'b0011 : 4'b0001;
										assign node2332 = (inp[3]) ? node2336 : node2333;
											assign node2333 = (inp[5]) ? 4'b0011 : 4'b0111;
											assign node2336 = (inp[5]) ? 4'b0001 : 4'b0001;
									assign node2339 = (inp[9]) ? node2347 : node2340;
										assign node2340 = (inp[12]) ? node2344 : node2341;
											assign node2341 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node2344 = (inp[5]) ? 4'b0111 : 4'b0011;
										assign node2347 = (inp[12]) ? 4'b0101 : 4'b0111;
							assign node2350 = (inp[1]) ? node2372 : node2351;
								assign node2351 = (inp[13]) ? node2359 : node2352;
									assign node2352 = (inp[9]) ? node2354 : 4'b0011;
										assign node2354 = (inp[2]) ? 4'b0001 : node2355;
											assign node2355 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node2359 = (inp[5]) ? node2365 : node2360;
										assign node2360 = (inp[15]) ? node2362 : 4'b1001;
											assign node2362 = (inp[2]) ? 4'b1111 : 4'b1011;
										assign node2365 = (inp[15]) ? node2369 : node2366;
											assign node2366 = (inp[12]) ? 4'b1111 : 4'b1001;
											assign node2369 = (inp[10]) ? 4'b1001 : 4'b1101;
								assign node2372 = (inp[2]) ? node2384 : node2373;
									assign node2373 = (inp[15]) ? node2379 : node2374;
										assign node2374 = (inp[9]) ? node2376 : 4'b1001;
											assign node2376 = (inp[12]) ? 4'b1111 : 4'b1011;
										assign node2379 = (inp[12]) ? 4'b1101 : node2380;
											assign node2380 = (inp[13]) ? 4'b1101 : 4'b1011;
									assign node2384 = (inp[15]) ? node2390 : node2385;
										assign node2385 = (inp[5]) ? 4'b1011 : node2386;
											assign node2386 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node2390 = (inp[3]) ? node2392 : 4'b1011;
											assign node2392 = (inp[4]) ? 4'b1001 : 4'b1011;
						assign node2395 = (inp[6]) ? node2451 : node2396;
							assign node2396 = (inp[13]) ? node2424 : node2397;
								assign node2397 = (inp[1]) ? node2411 : node2398;
									assign node2398 = (inp[15]) ? node2404 : node2399;
										assign node2399 = (inp[3]) ? 4'b0111 : node2400;
											assign node2400 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node2404 = (inp[5]) ? node2408 : node2405;
											assign node2405 = (inp[3]) ? 4'b0011 : 4'b0111;
											assign node2408 = (inp[10]) ? 4'b0001 : 4'b0101;
									assign node2411 = (inp[12]) ? node2419 : node2412;
										assign node2412 = (inp[5]) ? node2416 : node2413;
											assign node2413 = (inp[15]) ? 4'b1111 : 4'b1001;
											assign node2416 = (inp[10]) ? 4'b1111 : 4'b1011;
										assign node2419 = (inp[2]) ? 4'b1111 : node2420;
											assign node2420 = (inp[15]) ? 4'b1101 : 4'b1111;
								assign node2424 = (inp[1]) ? node2438 : node2425;
									assign node2425 = (inp[2]) ? node2433 : node2426;
										assign node2426 = (inp[12]) ? node2430 : node2427;
											assign node2427 = (inp[9]) ? 4'b1101 : 4'b1111;
											assign node2430 = (inp[15]) ? 4'b1101 : 4'b1001;
										assign node2433 = (inp[9]) ? 4'b1011 : node2434;
											assign node2434 = (inp[10]) ? 4'b1111 : 4'b1101;
									assign node2438 = (inp[9]) ? node2444 : node2439;
										assign node2439 = (inp[10]) ? 4'b1011 : node2440;
											assign node2440 = (inp[2]) ? 4'b1011 : 4'b1001;
										assign node2444 = (inp[3]) ? node2448 : node2445;
											assign node2445 = (inp[12]) ? 4'b1011 : 4'b1001;
											assign node2448 = (inp[15]) ? 4'b1101 : 4'b1111;
							assign node2451 = (inp[13]) ? node2475 : node2452;
								assign node2452 = (inp[1]) ? node2464 : node2453;
									assign node2453 = (inp[9]) ? node2459 : node2454;
										assign node2454 = (inp[5]) ? node2456 : 4'b1101;
											assign node2456 = (inp[2]) ? 4'b1101 : 4'b1001;
										assign node2459 = (inp[3]) ? node2461 : 4'b1111;
											assign node2461 = (inp[15]) ? 4'b1001 : 4'b1011;
									assign node2464 = (inp[12]) ? node2470 : node2465;
										assign node2465 = (inp[4]) ? 4'b0111 : node2466;
											assign node2466 = (inp[2]) ? 4'b0001 : 4'b0101;
										assign node2470 = (inp[10]) ? 4'b0001 : node2471;
											assign node2471 = (inp[2]) ? 4'b0001 : 4'b0111;
								assign node2475 = (inp[10]) ? node2491 : node2476;
									assign node2476 = (inp[5]) ? node2484 : node2477;
										assign node2477 = (inp[2]) ? node2481 : node2478;
											assign node2478 = (inp[12]) ? 4'b0101 : 4'b0101;
											assign node2481 = (inp[4]) ? 4'b0001 : 4'b0001;
										assign node2484 = (inp[15]) ? node2488 : node2485;
											assign node2485 = (inp[1]) ? 4'b0111 : 4'b0101;
											assign node2488 = (inp[12]) ? 4'b0001 : 4'b0101;
									assign node2491 = (inp[5]) ? node2499 : node2492;
										assign node2492 = (inp[12]) ? node2496 : node2493;
											assign node2493 = (inp[3]) ? 4'b0111 : 4'b0011;
											assign node2496 = (inp[3]) ? 4'b0001 : 4'b0001;
										assign node2499 = (inp[15]) ? node2503 : node2500;
											assign node2500 = (inp[1]) ? 4'b0001 : 4'b0111;
											assign node2503 = (inp[12]) ? 4'b0101 : 4'b0001;
			assign node2506 = (inp[8]) ? node2900 : node2507;
				assign node2507 = (inp[14]) ? node2695 : node2508;
					assign node2508 = (inp[2]) ? node2604 : node2509;
						assign node2509 = (inp[6]) ? node2553 : node2510;
							assign node2510 = (inp[11]) ? node2532 : node2511;
								assign node2511 = (inp[1]) ? node2521 : node2512;
									assign node2512 = (inp[5]) ? node2516 : node2513;
										assign node2513 = (inp[13]) ? 4'b1000 : 4'b1100;
										assign node2516 = (inp[15]) ? 4'b1100 : node2517;
											assign node2517 = (inp[3]) ? 4'b1010 : 4'b1000;
									assign node2521 = (inp[13]) ? node2527 : node2522;
										assign node2522 = (inp[9]) ? node2524 : 4'b1010;
											assign node2524 = (inp[12]) ? 4'b1100 : 4'b1110;
										assign node2527 = (inp[4]) ? 4'b0100 : node2528;
											assign node2528 = (inp[3]) ? 4'b0000 : 4'b0110;
								assign node2532 = (inp[13]) ? node2544 : node2533;
									assign node2533 = (inp[15]) ? node2541 : node2534;
										assign node2534 = (inp[9]) ? node2538 : node2535;
											assign node2535 = (inp[12]) ? 4'b0100 : 4'b0000;
											assign node2538 = (inp[10]) ? 4'b0010 : 4'b0010;
										assign node2541 = (inp[5]) ? 4'b0100 : 4'b0010;
									assign node2544 = (inp[1]) ? node2548 : node2545;
										assign node2545 = (inp[10]) ? 4'b0000 : 4'b0010;
										assign node2548 = (inp[9]) ? 4'b1010 : node2549;
											assign node2549 = (inp[3]) ? 4'b1010 : 4'b1100;
							assign node2553 = (inp[11]) ? node2575 : node2554;
								assign node2554 = (inp[13]) ? node2566 : node2555;
									assign node2555 = (inp[4]) ? node2561 : node2556;
										assign node2556 = (inp[3]) ? 4'b0000 : node2557;
											assign node2557 = (inp[10]) ? 4'b0000 : 4'b0100;
										assign node2561 = (inp[12]) ? 4'b0010 : node2562;
											assign node2562 = (inp[9]) ? 4'b0100 : 4'b0010;
									assign node2566 = (inp[1]) ? node2570 : node2567;
										assign node2567 = (inp[12]) ? 4'b0100 : 4'b0010;
										assign node2570 = (inp[4]) ? 4'b1000 : node2571;
											assign node2571 = (inp[3]) ? 4'b1100 : 4'b1110;
								assign node2575 = (inp[15]) ? node2591 : node2576;
									assign node2576 = (inp[5]) ? node2584 : node2577;
										assign node2577 = (inp[13]) ? node2581 : node2578;
											assign node2578 = (inp[3]) ? 4'b1110 : 4'b1100;
											assign node2581 = (inp[4]) ? 4'b0000 : 4'b1000;
										assign node2584 = (inp[1]) ? node2588 : node2585;
											assign node2585 = (inp[4]) ? 4'b1110 : 4'b1010;
											assign node2588 = (inp[13]) ? 4'b0110 : 4'b1110;
									assign node2591 = (inp[3]) ? node2599 : node2592;
										assign node2592 = (inp[13]) ? node2596 : node2593;
											assign node2593 = (inp[1]) ? 4'b1000 : 4'b1010;
											assign node2596 = (inp[4]) ? 4'b1010 : 4'b1110;
										assign node2599 = (inp[4]) ? 4'b1100 : node2600;
											assign node2600 = (inp[12]) ? 4'b1000 : 4'b1010;
						assign node2604 = (inp[9]) ? node2650 : node2605;
							assign node2605 = (inp[15]) ? node2629 : node2606;
								assign node2606 = (inp[4]) ? node2620 : node2607;
									assign node2607 = (inp[11]) ? node2615 : node2608;
										assign node2608 = (inp[3]) ? node2612 : node2609;
											assign node2609 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node2612 = (inp[5]) ? 4'b1011 : 4'b1101;
										assign node2615 = (inp[5]) ? node2617 : 4'b1001;
											assign node2617 = (inp[13]) ? 4'b0001 : 4'b1011;
									assign node2620 = (inp[5]) ? node2626 : node2621;
										assign node2621 = (inp[10]) ? node2623 : 4'b0001;
											assign node2623 = (inp[13]) ? 4'b0001 : 4'b0101;
										assign node2626 = (inp[11]) ? 4'b0111 : 4'b1111;
								assign node2629 = (inp[4]) ? node2639 : node2630;
									assign node2630 = (inp[3]) ? node2636 : node2631;
										assign node2631 = (inp[13]) ? 4'b1011 : node2632;
											assign node2632 = (inp[11]) ? 4'b0011 : 4'b0111;
										assign node2636 = (inp[5]) ? 4'b0101 : 4'b0111;
									assign node2639 = (inp[13]) ? node2645 : node2640;
										assign node2640 = (inp[11]) ? node2642 : 4'b0101;
											assign node2642 = (inp[6]) ? 4'b1111 : 4'b0011;
										assign node2645 = (inp[12]) ? node2647 : 4'b0101;
											assign node2647 = (inp[10]) ? 4'b1101 : 4'b1101;
							assign node2650 = (inp[10]) ? node2674 : node2651;
								assign node2651 = (inp[15]) ? node2663 : node2652;
									assign node2652 = (inp[5]) ? node2658 : node2653;
										assign node2653 = (inp[1]) ? node2655 : 4'b1101;
											assign node2655 = (inp[4]) ? 4'b1011 : 4'b1001;
										assign node2658 = (inp[12]) ? 4'b1111 : node2659;
											assign node2659 = (inp[1]) ? 4'b0111 : 4'b1111;
									assign node2663 = (inp[1]) ? node2669 : node2664;
										assign node2664 = (inp[4]) ? 4'b1001 : node2665;
											assign node2665 = (inp[6]) ? 4'b1111 : 4'b1011;
										assign node2669 = (inp[12]) ? node2671 : 4'b1101;
											assign node2671 = (inp[3]) ? 4'b0001 : 4'b1101;
								assign node2674 = (inp[15]) ? node2682 : node2675;
									assign node2675 = (inp[1]) ? node2679 : node2676;
										assign node2676 = (inp[3]) ? 4'b0111 : 4'b1111;
										assign node2679 = (inp[3]) ? 4'b0011 : 4'b0111;
									assign node2682 = (inp[12]) ? node2690 : node2683;
										assign node2683 = (inp[6]) ? node2687 : node2684;
											assign node2684 = (inp[4]) ? 4'b0101 : 4'b1001;
											assign node2687 = (inp[11]) ? 4'b0001 : 4'b1001;
										assign node2690 = (inp[3]) ? 4'b0001 : node2691;
											assign node2691 = (inp[13]) ? 4'b0011 : 4'b0011;
					assign node2695 = (inp[10]) ? node2799 : node2696;
						assign node2696 = (inp[3]) ? node2752 : node2697;
							assign node2697 = (inp[15]) ? node2725 : node2698;
								assign node2698 = (inp[5]) ? node2712 : node2699;
									assign node2699 = (inp[11]) ? node2705 : node2700;
										assign node2700 = (inp[13]) ? node2702 : 4'b0001;
											assign node2702 = (inp[6]) ? 4'b1101 : 4'b0101;
										assign node2705 = (inp[6]) ? node2709 : node2706;
											assign node2706 = (inp[1]) ? 4'b1101 : 4'b0101;
											assign node2709 = (inp[13]) ? 4'b0001 : 4'b0101;
									assign node2712 = (inp[4]) ? node2720 : node2713;
										assign node2713 = (inp[2]) ? node2717 : node2714;
											assign node2714 = (inp[11]) ? 4'b1101 : 4'b0001;
											assign node2717 = (inp[6]) ? 4'b1111 : 4'b0101;
										assign node2720 = (inp[9]) ? 4'b0111 : node2721;
											assign node2721 = (inp[13]) ? 4'b1111 : 4'b0001;
								assign node2725 = (inp[1]) ? node2741 : node2726;
									assign node2726 = (inp[11]) ? node2734 : node2727;
										assign node2727 = (inp[2]) ? node2731 : node2728;
											assign node2728 = (inp[5]) ? 4'b0011 : 4'b1011;
											assign node2731 = (inp[12]) ? 4'b0111 : 4'b0011;
										assign node2734 = (inp[9]) ? node2738 : node2735;
											assign node2735 = (inp[5]) ? 4'b1011 : 4'b1111;
											assign node2738 = (inp[5]) ? 4'b0101 : 4'b0111;
									assign node2741 = (inp[12]) ? node2747 : node2742;
										assign node2742 = (inp[5]) ? 4'b0111 : node2743;
											assign node2743 = (inp[2]) ? 4'b1011 : 4'b0011;
										assign node2747 = (inp[4]) ? node2749 : 4'b0011;
											assign node2749 = (inp[5]) ? 4'b1001 : 4'b1011;
							assign node2752 = (inp[15]) ? node2774 : node2753;
								assign node2753 = (inp[5]) ? node2765 : node2754;
									assign node2754 = (inp[13]) ? node2760 : node2755;
										assign node2755 = (inp[11]) ? 4'b1111 : node2756;
											assign node2756 = (inp[9]) ? 4'b1111 : 4'b0101;
										assign node2760 = (inp[9]) ? 4'b1001 : node2761;
											assign node2761 = (inp[11]) ? 4'b0001 : 4'b0001;
									assign node2765 = (inp[4]) ? node2769 : node2766;
										assign node2766 = (inp[13]) ? 4'b1011 : 4'b1111;
										assign node2769 = (inp[2]) ? 4'b1111 : node2770;
											assign node2770 = (inp[11]) ? 4'b0011 : 4'b0111;
								assign node2774 = (inp[9]) ? node2786 : node2775;
									assign node2775 = (inp[5]) ? node2779 : node2776;
										assign node2776 = (inp[4]) ? 4'b1101 : 4'b1111;
										assign node2779 = (inp[4]) ? node2783 : node2780;
											assign node2780 = (inp[1]) ? 4'b1101 : 4'b0101;
											assign node2783 = (inp[6]) ? 4'b1001 : 4'b0001;
									assign node2786 = (inp[4]) ? node2792 : node2787;
										assign node2787 = (inp[6]) ? node2789 : 4'b0011;
											assign node2789 = (inp[11]) ? 4'b0101 : 4'b1101;
										assign node2792 = (inp[12]) ? node2796 : node2793;
											assign node2793 = (inp[2]) ? 4'b0101 : 4'b0101;
											assign node2796 = (inp[11]) ? 4'b0001 : 4'b0101;
						assign node2799 = (inp[11]) ? node2847 : node2800;
							assign node2800 = (inp[2]) ? node2824 : node2801;
								assign node2801 = (inp[12]) ? node2815 : node2802;
									assign node2802 = (inp[15]) ? node2808 : node2803;
										assign node2803 = (inp[6]) ? node2805 : 4'b1001;
											assign node2805 = (inp[1]) ? 4'b1001 : 4'b1101;
										assign node2808 = (inp[4]) ? node2812 : node2809;
											assign node2809 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node2812 = (inp[5]) ? 4'b0011 : 4'b1111;
									assign node2815 = (inp[3]) ? node2819 : node2816;
										assign node2816 = (inp[1]) ? 4'b1001 : 4'b1111;
										assign node2819 = (inp[15]) ? node2821 : 4'b0111;
											assign node2821 = (inp[5]) ? 4'b1101 : 4'b0101;
								assign node2824 = (inp[4]) ? node2838 : node2825;
									assign node2825 = (inp[6]) ? node2833 : node2826;
										assign node2826 = (inp[1]) ? node2830 : node2827;
											assign node2827 = (inp[13]) ? 4'b0111 : 4'b1001;
											assign node2830 = (inp[9]) ? 4'b0111 : 4'b0101;
										assign node2833 = (inp[1]) ? node2835 : 4'b1111;
											assign node2835 = (inp[15]) ? 4'b1011 : 4'b1001;
									assign node2838 = (inp[13]) ? node2844 : node2839;
										assign node2839 = (inp[6]) ? 4'b0001 : node2840;
											assign node2840 = (inp[12]) ? 4'b0001 : 4'b1001;
										assign node2844 = (inp[6]) ? 4'b1001 : 4'b0001;
							assign node2847 = (inp[6]) ? node2875 : node2848;
								assign node2848 = (inp[3]) ? node2862 : node2849;
									assign node2849 = (inp[15]) ? node2857 : node2850;
										assign node2850 = (inp[5]) ? node2854 : node2851;
											assign node2851 = (inp[2]) ? 4'b1001 : 4'b1001;
											assign node2854 = (inp[4]) ? 4'b1011 : 4'b1001;
										assign node2857 = (inp[4]) ? node2859 : 4'b1011;
											assign node2859 = (inp[12]) ? 4'b1111 : 4'b1101;
									assign node2862 = (inp[1]) ? node2870 : node2863;
										assign node2863 = (inp[13]) ? node2867 : node2864;
											assign node2864 = (inp[9]) ? 4'b0001 : 4'b0011;
											assign node2867 = (inp[2]) ? 4'b1111 : 4'b1101;
										assign node2870 = (inp[15]) ? 4'b1001 : node2871;
											assign node2871 = (inp[13]) ? 4'b1011 : 4'b1111;
								assign node2875 = (inp[1]) ? node2887 : node2876;
									assign node2876 = (inp[13]) ? node2884 : node2877;
										assign node2877 = (inp[12]) ? node2881 : node2878;
											assign node2878 = (inp[5]) ? 4'b1011 : 4'b1111;
											assign node2881 = (inp[5]) ? 4'b1001 : 4'b1011;
										assign node2884 = (inp[15]) ? 4'b0101 : 4'b0011;
									assign node2887 = (inp[15]) ? node2895 : node2888;
										assign node2888 = (inp[9]) ? node2892 : node2889;
											assign node2889 = (inp[4]) ? 4'b0111 : 4'b0001;
											assign node2892 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node2895 = (inp[5]) ? 4'b0001 : node2896;
											assign node2896 = (inp[4]) ? 4'b0001 : 4'b0101;
				assign node2900 = (inp[14]) ? node3102 : node2901;
					assign node2901 = (inp[2]) ? node3001 : node2902;
						assign node2902 = (inp[13]) ? node2952 : node2903;
							assign node2903 = (inp[3]) ? node2925 : node2904;
								assign node2904 = (inp[6]) ? node2916 : node2905;
									assign node2905 = (inp[5]) ? node2911 : node2906;
										assign node2906 = (inp[4]) ? node2908 : 4'b1001;
											assign node2908 = (inp[1]) ? 4'b0111 : 4'b1111;
										assign node2911 = (inp[15]) ? node2913 : 4'b0111;
											assign node2913 = (inp[4]) ? 4'b0101 : 4'b0111;
									assign node2916 = (inp[9]) ? node2920 : node2917;
										assign node2917 = (inp[10]) ? 4'b0111 : 4'b0101;
										assign node2920 = (inp[4]) ? node2922 : 4'b1111;
											assign node2922 = (inp[12]) ? 4'b1001 : 4'b1001;
								assign node2925 = (inp[6]) ? node2937 : node2926;
									assign node2926 = (inp[15]) ? node2934 : node2927;
										assign node2927 = (inp[11]) ? node2931 : node2928;
											assign node2928 = (inp[5]) ? 4'b0011 : 4'b1001;
											assign node2931 = (inp[4]) ? 4'b0111 : 4'b1111;
										assign node2934 = (inp[5]) ? 4'b1001 : 4'b1011;
									assign node2937 = (inp[4]) ? node2945 : node2938;
										assign node2938 = (inp[15]) ? node2942 : node2939;
											assign node2939 = (inp[12]) ? 4'b1111 : 4'b0111;
											assign node2942 = (inp[5]) ? 4'b0101 : 4'b0011;
										assign node2945 = (inp[5]) ? node2949 : node2946;
											assign node2946 = (inp[12]) ? 4'b0001 : 4'b0011;
											assign node2949 = (inp[11]) ? 4'b0011 : 4'b1011;
							assign node2952 = (inp[9]) ? node2976 : node2953;
								assign node2953 = (inp[11]) ? node2967 : node2954;
									assign node2954 = (inp[6]) ? node2962 : node2955;
										assign node2955 = (inp[15]) ? node2959 : node2956;
											assign node2956 = (inp[3]) ? 4'b0101 : 4'b0001;
											assign node2959 = (inp[1]) ? 4'b0111 : 4'b0011;
										assign node2962 = (inp[12]) ? 4'b1001 : node2963;
											assign node2963 = (inp[5]) ? 4'b1101 : 4'b1011;
									assign node2967 = (inp[6]) ? node2971 : node2968;
										assign node2968 = (inp[4]) ? 4'b1111 : 4'b1011;
										assign node2971 = (inp[4]) ? node2973 : 4'b0011;
											assign node2973 = (inp[15]) ? 4'b0101 : 4'b0111;
								assign node2976 = (inp[5]) ? node2988 : node2977;
									assign node2977 = (inp[12]) ? node2983 : node2978;
										assign node2978 = (inp[4]) ? 4'b0101 : node2979;
											assign node2979 = (inp[15]) ? 4'b0111 : 4'b0001;
										assign node2983 = (inp[4]) ? 4'b0001 : node2984;
											assign node2984 = (inp[6]) ? 4'b0101 : 4'b1101;
									assign node2988 = (inp[15]) ? node2994 : node2989;
										assign node2989 = (inp[6]) ? 4'b1111 : node2990;
											assign node2990 = (inp[11]) ? 4'b1111 : 4'b0111;
										assign node2994 = (inp[4]) ? node2998 : node2995;
											assign node2995 = (inp[10]) ? 4'b0101 : 4'b1101;
											assign node2998 = (inp[10]) ? 4'b1001 : 4'b1101;
						assign node3001 = (inp[15]) ? node3055 : node3002;
							assign node3002 = (inp[3]) ? node3026 : node3003;
								assign node3003 = (inp[10]) ? node3017 : node3004;
									assign node3004 = (inp[13]) ? node3010 : node3005;
										assign node3005 = (inp[11]) ? node3007 : 4'b1000;
											assign node3007 = (inp[6]) ? 4'b1000 : 4'b0000;
										assign node3010 = (inp[1]) ? node3014 : node3011;
											assign node3011 = (inp[9]) ? 4'b0000 : 4'b0100;
											assign node3014 = (inp[5]) ? 4'b0110 : 4'b1100;
									assign node3017 = (inp[5]) ? 4'b1110 : node3018;
										assign node3018 = (inp[6]) ? node3022 : node3019;
											assign node3019 = (inp[11]) ? 4'b1100 : 4'b0000;
											assign node3022 = (inp[1]) ? 4'b1100 : 4'b0100;
								assign node3026 = (inp[12]) ? node3042 : node3027;
									assign node3027 = (inp[5]) ? node3035 : node3028;
										assign node3028 = (inp[9]) ? node3032 : node3029;
											assign node3029 = (inp[4]) ? 4'b0110 : 4'b0100;
											assign node3032 = (inp[11]) ? 4'b1110 : 4'b1110;
										assign node3035 = (inp[13]) ? node3039 : node3036;
											assign node3036 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node3039 = (inp[9]) ? 4'b0110 : 4'b1110;
									assign node3042 = (inp[6]) ? node3048 : node3043;
										assign node3043 = (inp[10]) ? 4'b1010 : node3044;
											assign node3044 = (inp[1]) ? 4'b1110 : 4'b1010;
										assign node3048 = (inp[11]) ? node3052 : node3049;
											assign node3049 = (inp[13]) ? 4'b1010 : 4'b1110;
											assign node3052 = (inp[5]) ? 4'b1110 : 4'b0110;
							assign node3055 = (inp[3]) ? node3075 : node3056;
								assign node3056 = (inp[5]) ? node3068 : node3057;
									assign node3057 = (inp[6]) ? node3061 : node3058;
										assign node3058 = (inp[11]) ? 4'b1110 : 4'b0110;
										assign node3061 = (inp[13]) ? node3065 : node3062;
											assign node3062 = (inp[4]) ? 4'b1110 : 4'b1010;
											assign node3065 = (inp[12]) ? 4'b0110 : 4'b0010;
									assign node3068 = (inp[11]) ? 4'b1100 : node3069;
										assign node3069 = (inp[4]) ? node3071 : 4'b0110;
											assign node3071 = (inp[9]) ? 4'b0000 : 4'b0100;
								assign node3075 = (inp[1]) ? node3091 : node3076;
									assign node3076 = (inp[9]) ? node3084 : node3077;
										assign node3077 = (inp[4]) ? node3081 : node3078;
											assign node3078 = (inp[6]) ? 4'b0100 : 4'b0100;
											assign node3081 = (inp[11]) ? 4'b1100 : 4'b0000;
										assign node3084 = (inp[5]) ? node3088 : node3085;
											assign node3085 = (inp[4]) ? 4'b0000 : 4'b0010;
											assign node3088 = (inp[4]) ? 4'b1000 : 4'b0000;
									assign node3091 = (inp[9]) ? node3097 : node3092;
										assign node3092 = (inp[10]) ? 4'b0100 : node3093;
											assign node3093 = (inp[11]) ? 4'b1000 : 4'b0000;
										assign node3097 = (inp[4]) ? 4'b0100 : node3098;
											assign node3098 = (inp[13]) ? 4'b1100 : 4'b0100;
					assign node3102 = (inp[11]) ? node3194 : node3103;
						assign node3103 = (inp[6]) ? node3149 : node3104;
							assign node3104 = (inp[1]) ? node3126 : node3105;
								assign node3105 = (inp[13]) ? node3115 : node3106;
									assign node3106 = (inp[10]) ? node3110 : node3107;
										assign node3107 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node3110 = (inp[3]) ? node3112 : 4'b1110;
											assign node3112 = (inp[12]) ? 4'b1000 : 4'b1100;
									assign node3115 = (inp[3]) ? node3119 : node3116;
										assign node3116 = (inp[15]) ? 4'b0010 : 4'b0000;
										assign node3119 = (inp[2]) ? node3123 : node3120;
											assign node3120 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node3123 = (inp[10]) ? 4'b0100 : 4'b0100;
								assign node3126 = (inp[15]) ? node3138 : node3127;
									assign node3127 = (inp[5]) ? node3131 : node3128;
										assign node3128 = (inp[13]) ? 4'b0000 : 4'b0100;
										assign node3131 = (inp[3]) ? node3135 : node3132;
											assign node3132 = (inp[2]) ? 4'b0100 : 4'b0110;
											assign node3135 = (inp[2]) ? 4'b0110 : 4'b0010;
									assign node3138 = (inp[3]) ? node3144 : node3139;
										assign node3139 = (inp[9]) ? 4'b0010 : node3140;
											assign node3140 = (inp[4]) ? 4'b0010 : 4'b0110;
										assign node3144 = (inp[5]) ? 4'b0000 : node3145;
											assign node3145 = (inp[9]) ? 4'b0000 : 4'b0010;
							assign node3149 = (inp[13]) ? node3173 : node3150;
								assign node3150 = (inp[1]) ? node3164 : node3151;
									assign node3151 = (inp[3]) ? node3157 : node3152;
										assign node3152 = (inp[15]) ? 4'b0110 : node3153;
											assign node3153 = (inp[10]) ? 4'b0100 : 4'b0000;
										assign node3157 = (inp[12]) ? node3161 : node3158;
											assign node3158 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node3161 = (inp[2]) ? 4'b0010 : 4'b0000;
									assign node3164 = (inp[15]) ? node3170 : node3165;
										assign node3165 = (inp[5]) ? 4'b1110 : node3166;
											assign node3166 = (inp[10]) ? 4'b1000 : 4'b1110;
										assign node3170 = (inp[12]) ? 4'b1110 : 4'b1100;
								assign node3173 = (inp[3]) ? node3183 : node3174;
									assign node3174 = (inp[5]) ? 4'b1100 : node3175;
										assign node3175 = (inp[15]) ? node3179 : node3176;
											assign node3176 = (inp[10]) ? 4'b1000 : 4'b1000;
											assign node3179 = (inp[4]) ? 4'b1110 : 4'b1010;
									assign node3183 = (inp[15]) ? node3189 : node3184;
										assign node3184 = (inp[4]) ? 4'b1010 : node3185;
											assign node3185 = (inp[9]) ? 4'b1110 : 4'b1010;
										assign node3189 = (inp[10]) ? 4'b1010 : node3190;
											assign node3190 = (inp[2]) ? 4'b1100 : 4'b1000;
						assign node3194 = (inp[6]) ? node3246 : node3195;
							assign node3195 = (inp[1]) ? node3223 : node3196;
								assign node3196 = (inp[13]) ? node3210 : node3197;
									assign node3197 = (inp[5]) ? node3203 : node3198;
										assign node3198 = (inp[2]) ? node3200 : 4'b0000;
											assign node3200 = (inp[9]) ? 4'b0100 : 4'b0000;
										assign node3203 = (inp[12]) ? node3207 : node3204;
											assign node3204 = (inp[10]) ? 4'b0110 : 4'b0010;
											assign node3207 = (inp[9]) ? 4'b0010 : 4'b0000;
									assign node3210 = (inp[4]) ? node3218 : node3211;
										assign node3211 = (inp[10]) ? node3215 : node3212;
											assign node3212 = (inp[3]) ? 4'b1110 : 4'b1100;
											assign node3215 = (inp[9]) ? 4'b1100 : 4'b1000;
										assign node3218 = (inp[3]) ? 4'b1000 : node3219;
											assign node3219 = (inp[2]) ? 4'b1010 : 4'b1000;
								assign node3223 = (inp[5]) ? node3235 : node3224;
									assign node3224 = (inp[15]) ? node3230 : node3225;
										assign node3225 = (inp[2]) ? node3227 : 4'b1100;
											assign node3227 = (inp[10]) ? 4'b1100 : 4'b1000;
										assign node3230 = (inp[3]) ? node3232 : 4'b1010;
											assign node3232 = (inp[9]) ? 4'b1100 : 4'b1110;
									assign node3235 = (inp[15]) ? node3241 : node3236;
										assign node3236 = (inp[3]) ? 4'b1010 : node3237;
											assign node3237 = (inp[2]) ? 4'b1010 : 4'b1110;
										assign node3241 = (inp[2]) ? node3243 : 4'b1100;
											assign node3243 = (inp[10]) ? 4'b1000 : 4'b1100;
							assign node3246 = (inp[1]) ? node3274 : node3247;
								assign node3247 = (inp[13]) ? node3261 : node3248;
									assign node3248 = (inp[15]) ? node3254 : node3249;
										assign node3249 = (inp[5]) ? 4'b1010 : node3250;
											assign node3250 = (inp[10]) ? 4'b1100 : 4'b1110;
										assign node3254 = (inp[12]) ? node3258 : node3255;
											assign node3255 = (inp[4]) ? 4'b1100 : 4'b1110;
											assign node3258 = (inp[9]) ? 4'b1000 : 4'b1100;
									assign node3261 = (inp[4]) ? node3267 : node3262;
										assign node3262 = (inp[9]) ? 4'b0100 : node3263;
											assign node3263 = (inp[12]) ? 4'b0000 : 4'b0100;
										assign node3267 = (inp[5]) ? node3271 : node3268;
											assign node3268 = (inp[10]) ? 4'b0110 : 4'b0010;
											assign node3271 = (inp[15]) ? 4'b0100 : 4'b0110;
								assign node3274 = (inp[15]) ? node3288 : node3275;
									assign node3275 = (inp[3]) ? node3283 : node3276;
										assign node3276 = (inp[5]) ? node3280 : node3277;
											assign node3277 = (inp[12]) ? 4'b0000 : 4'b0000;
											assign node3280 = (inp[12]) ? 4'b0110 : 4'b0000;
										assign node3283 = (inp[9]) ? node3285 : 4'b0010;
											assign node3285 = (inp[2]) ? 4'b0010 : 4'b0110;
									assign node3288 = (inp[4]) ? node3292 : node3289;
										assign node3289 = (inp[9]) ? 4'b0100 : 4'b0000;
										assign node3292 = (inp[5]) ? node3296 : node3293;
											assign node3293 = (inp[3]) ? 4'b0100 : 4'b0010;
											assign node3296 = (inp[3]) ? 4'b0000 : 4'b0100;

endmodule