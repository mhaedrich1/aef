module dtc_split66_bm75 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node227;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node270;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node317;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node334;
	wire [3-1:0] node337;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node368;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node399;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node408;
	wire [3-1:0] node411;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node426;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node436;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node451;
	wire [3-1:0] node454;
	wire [3-1:0] node456;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node480;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node495;
	wire [3-1:0] node497;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node510;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node519;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node526;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node534;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node541;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node558;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node572;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node585;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node604;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node640;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node646;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node663;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node670;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node681;
	wire [3-1:0] node683;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node692;
	wire [3-1:0] node695;
	wire [3-1:0] node697;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node705;
	wire [3-1:0] node708;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node723;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node730;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node735;
	wire [3-1:0] node738;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node745;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node759;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node764;
	wire [3-1:0] node767;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node774;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node784;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node791;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node799;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node806;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node815;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node822;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node830;
	wire [3-1:0] node833;
	wire [3-1:0] node835;
	wire [3-1:0] node838;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node849;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node864;
	wire [3-1:0] node867;
	wire [3-1:0] node868;
	wire [3-1:0] node871;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node885;
	wire [3-1:0] node888;
	wire [3-1:0] node889;
	wire [3-1:0] node891;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node898;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node908;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node916;
	wire [3-1:0] node917;
	wire [3-1:0] node918;
	wire [3-1:0] node921;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node928;
	wire [3-1:0] node931;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node937;
	wire [3-1:0] node940;
	wire [3-1:0] node942;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node950;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node957;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node968;
	wire [3-1:0] node971;
	wire [3-1:0] node972;
	wire [3-1:0] node975;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node983;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node990;
	wire [3-1:0] node993;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node999;
	wire [3-1:0] node1002;
	wire [3-1:0] node1004;
	wire [3-1:0] node1007;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1012;
	wire [3-1:0] node1015;
	wire [3-1:0] node1016;
	wire [3-1:0] node1019;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1029;
	wire [3-1:0] node1032;
	wire [3-1:0] node1033;
	wire [3-1:0] node1036;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1044;
	wire [3-1:0] node1047;
	wire [3-1:0] node1048;
	wire [3-1:0] node1051;
	wire [3-1:0] node1054;
	wire [3-1:0] node1055;
	wire [3-1:0] node1056;
	wire [3-1:0] node1057;
	wire [3-1:0] node1060;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1067;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1076;
	wire [3-1:0] node1077;
	wire [3-1:0] node1080;
	wire [3-1:0] node1083;
	wire [3-1:0] node1084;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1087;
	wire [3-1:0] node1088;
	wire [3-1:0] node1090;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1097;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1110;
	wire [3-1:0] node1112;
	wire [3-1:0] node1115;
	wire [3-1:0] node1116;
	wire [3-1:0] node1118;
	wire [3-1:0] node1121;
	wire [3-1:0] node1122;
	wire [3-1:0] node1125;
	wire [3-1:0] node1128;
	wire [3-1:0] node1129;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1134;
	wire [3-1:0] node1137;
	wire [3-1:0] node1139;
	wire [3-1:0] node1142;
	wire [3-1:0] node1144;
	wire [3-1:0] node1146;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1152;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1157;
	wire [3-1:0] node1160;
	wire [3-1:0] node1161;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1168;
	wire [3-1:0] node1171;
	wire [3-1:0] node1172;
	wire [3-1:0] node1175;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1180;
	wire [3-1:0] node1181;
	wire [3-1:0] node1185;
	wire [3-1:0] node1186;
	wire [3-1:0] node1189;
	wire [3-1:0] node1192;
	wire [3-1:0] node1194;
	wire [3-1:0] node1196;
	wire [3-1:0] node1199;
	wire [3-1:0] node1200;
	wire [3-1:0] node1201;
	wire [3-1:0] node1202;
	wire [3-1:0] node1203;
	wire [3-1:0] node1206;
	wire [3-1:0] node1209;
	wire [3-1:0] node1210;
	wire [3-1:0] node1213;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1221;
	wire [3-1:0] node1224;
	wire [3-1:0] node1225;
	wire [3-1:0] node1228;
	wire [3-1:0] node1231;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1234;
	wire [3-1:0] node1237;
	wire [3-1:0] node1240;
	wire [3-1:0] node1241;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1250;
	wire [3-1:0] node1253;
	wire [3-1:0] node1254;
	wire [3-1:0] node1257;
	wire [3-1:0] node1260;
	wire [3-1:0] node1261;
	wire [3-1:0] node1262;
	wire [3-1:0] node1263;
	wire [3-1:0] node1265;
	wire [3-1:0] node1266;
	wire [3-1:0] node1267;
	wire [3-1:0] node1269;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1276;
	wire [3-1:0] node1279;
	wire [3-1:0] node1280;
	wire [3-1:0] node1282;
	wire [3-1:0] node1286;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1289;
	wire [3-1:0] node1291;
	wire [3-1:0] node1294;
	wire [3-1:0] node1295;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1302;
	wire [3-1:0] node1305;
	wire [3-1:0] node1306;
	wire [3-1:0] node1309;
	wire [3-1:0] node1312;
	wire [3-1:0] node1313;
	wire [3-1:0] node1314;
	wire [3-1:0] node1316;
	wire [3-1:0] node1319;
	wire [3-1:0] node1320;
	wire [3-1:0] node1323;
	wire [3-1:0] node1326;
	wire [3-1:0] node1328;
	wire [3-1:0] node1330;
	wire [3-1:0] node1333;
	wire [3-1:0] node1334;
	wire [3-1:0] node1335;
	wire [3-1:0] node1336;
	wire [3-1:0] node1337;
	wire [3-1:0] node1338;
	wire [3-1:0] node1341;
	wire [3-1:0] node1344;
	wire [3-1:0] node1346;
	wire [3-1:0] node1349;
	wire [3-1:0] node1350;
	wire [3-1:0] node1351;
	wire [3-1:0] node1354;
	wire [3-1:0] node1357;
	wire [3-1:0] node1359;
	wire [3-1:0] node1362;
	wire [3-1:0] node1363;
	wire [3-1:0] node1364;
	wire [3-1:0] node1366;
	wire [3-1:0] node1369;
	wire [3-1:0] node1370;
	wire [3-1:0] node1373;
	wire [3-1:0] node1376;
	wire [3-1:0] node1378;
	wire [3-1:0] node1380;
	wire [3-1:0] node1383;
	wire [3-1:0] node1384;
	wire [3-1:0] node1385;
	wire [3-1:0] node1386;
	wire [3-1:0] node1387;
	wire [3-1:0] node1390;
	wire [3-1:0] node1393;
	wire [3-1:0] node1394;
	wire [3-1:0] node1397;
	wire [3-1:0] node1400;
	wire [3-1:0] node1401;
	wire [3-1:0] node1402;
	wire [3-1:0] node1405;
	wire [3-1:0] node1408;
	wire [3-1:0] node1409;
	wire [3-1:0] node1412;
	wire [3-1:0] node1415;
	wire [3-1:0] node1416;
	wire [3-1:0] node1417;
	wire [3-1:0] node1418;
	wire [3-1:0] node1421;
	wire [3-1:0] node1424;
	wire [3-1:0] node1425;
	wire [3-1:0] node1428;
	wire [3-1:0] node1431;
	wire [3-1:0] node1432;
	wire [3-1:0] node1435;
	wire [3-1:0] node1437;
	wire [3-1:0] node1440;
	wire [3-1:0] node1441;
	wire [3-1:0] node1443;
	wire [3-1:0] node1444;
	wire [3-1:0] node1446;
	wire [3-1:0] node1447;
	wire [3-1:0] node1449;
	wire [3-1:0] node1454;
	wire [3-1:0] node1455;
	wire [3-1:0] node1457;
	wire [3-1:0] node1459;
	wire [3-1:0] node1460;
	wire [3-1:0] node1461;
	wire [3-1:0] node1466;
	wire [3-1:0] node1467;
	wire [3-1:0] node1468;
	wire [3-1:0] node1469;
	wire [3-1:0] node1470;
	wire [3-1:0] node1474;
	wire [3-1:0] node1475;
	wire [3-1:0] node1479;
	wire [3-1:0] node1480;
	wire [3-1:0] node1481;
	wire [3-1:0] node1485;
	wire [3-1:0] node1486;
	wire [3-1:0] node1489;
	wire [3-1:0] node1492;
	wire [3-1:0] node1493;
	wire [3-1:0] node1495;
	wire [3-1:0] node1496;
	wire [3-1:0] node1500;
	wire [3-1:0] node1501;
	wire [3-1:0] node1502;
	wire [3-1:0] node1505;
	wire [3-1:0] node1508;
	wire [3-1:0] node1509;

	assign outp = (inp[3]) ? node838 : node1;
		assign node1 = (inp[9]) ? node371 : node2;
			assign node2 = (inp[4]) ? node144 : node3;
				assign node3 = (inp[6]) ? node101 : node4;
					assign node4 = (inp[0]) ? node66 : node5;
						assign node5 = (inp[10]) ? node35 : node6;
							assign node6 = (inp[5]) ? node20 : node7;
								assign node7 = (inp[7]) ? node15 : node8;
									assign node8 = (inp[1]) ? node12 : node9;
										assign node9 = (inp[8]) ? 3'b011 : 3'b101;
										assign node12 = (inp[2]) ? 3'b111 : 3'b011;
									assign node15 = (inp[1]) ? 3'b111 : node16;
										assign node16 = (inp[8]) ? 3'b111 : 3'b011;
								assign node20 = (inp[7]) ? node28 : node21;
									assign node21 = (inp[2]) ? node25 : node22;
										assign node22 = (inp[8]) ? 3'b001 : 3'b101;
										assign node25 = (inp[11]) ? 3'b001 : 3'b011;
									assign node28 = (inp[11]) ? node32 : node29;
										assign node29 = (inp[1]) ? 3'b111 : 3'b011;
										assign node32 = (inp[2]) ? 3'b011 : 3'b001;
							assign node35 = (inp[5]) ? node51 : node36;
								assign node36 = (inp[1]) ? node44 : node37;
									assign node37 = (inp[2]) ? node41 : node38;
										assign node38 = (inp[7]) ? 3'b101 : 3'b001;
										assign node41 = (inp[7]) ? 3'b011 : 3'b101;
									assign node44 = (inp[2]) ? node48 : node45;
										assign node45 = (inp[8]) ? 3'b011 : 3'b101;
										assign node48 = (inp[7]) ? 3'b111 : 3'b011;
								assign node51 = (inp[1]) ? node59 : node52;
									assign node52 = (inp[7]) ? node56 : node53;
										assign node53 = (inp[11]) ? 3'b000 : 3'b001;
										assign node56 = (inp[11]) ? 3'b001 : 3'b101;
									assign node59 = (inp[11]) ? node63 : node60;
										assign node60 = (inp[7]) ? 3'b001 : 3'b101;
										assign node63 = (inp[7]) ? 3'b101 : 3'b001;
						assign node66 = (inp[10]) ? node78 : node67;
							assign node67 = (inp[5]) ? node69 : 3'b111;
								assign node69 = (inp[11]) ? node71 : 3'b111;
									assign node71 = (inp[1]) ? node75 : node72;
										assign node72 = (inp[7]) ? 3'b111 : 3'b011;
										assign node75 = (inp[8]) ? 3'b111 : 3'b111;
							assign node78 = (inp[5]) ? node88 : node79;
								assign node79 = (inp[7]) ? 3'b111 : node80;
									assign node80 = (inp[1]) ? node84 : node81;
										assign node81 = (inp[11]) ? 3'b011 : 3'b011;
										assign node84 = (inp[2]) ? 3'b111 : 3'b011;
								assign node88 = (inp[8]) ? node94 : node89;
									assign node89 = (inp[1]) ? 3'b011 : node90;
										assign node90 = (inp[11]) ? 3'b001 : 3'b011;
									assign node94 = (inp[1]) ? node98 : node95;
										assign node95 = (inp[7]) ? 3'b011 : 3'b101;
										assign node98 = (inp[7]) ? 3'b111 : 3'b011;
					assign node101 = (inp[0]) ? node133 : node102;
						assign node102 = (inp[10]) ? node112 : node103;
							assign node103 = (inp[1]) ? 3'b111 : node104;
								assign node104 = (inp[5]) ? node106 : 3'b111;
									assign node106 = (inp[8]) ? 3'b111 : node107;
										assign node107 = (inp[7]) ? 3'b111 : 3'b011;
							assign node112 = (inp[7]) ? node126 : node113;
								assign node113 = (inp[5]) ? node121 : node114;
									assign node114 = (inp[11]) ? node118 : node115;
										assign node115 = (inp[2]) ? 3'b111 : 3'b111;
										assign node118 = (inp[2]) ? 3'b011 : 3'b011;
									assign node121 = (inp[2]) ? 3'b011 : node122;
										assign node122 = (inp[11]) ? 3'b101 : 3'b011;
								assign node126 = (inp[1]) ? 3'b111 : node127;
									assign node127 = (inp[5]) ? node129 : 3'b111;
										assign node129 = (inp[2]) ? 3'b011 : 3'b001;
						assign node133 = (inp[2]) ? 3'b111 : node134;
							assign node134 = (inp[1]) ? 3'b111 : node135;
								assign node135 = (inp[7]) ? 3'b111 : node136;
									assign node136 = (inp[5]) ? node138 : 3'b111;
										assign node138 = (inp[8]) ? 3'b111 : 3'b011;
				assign node144 = (inp[6]) ? node264 : node145;
					assign node145 = (inp[5]) ? node205 : node146;
						assign node146 = (inp[0]) ? node176 : node147;
							assign node147 = (inp[7]) ? node163 : node148;
								assign node148 = (inp[10]) ? node156 : node149;
									assign node149 = (inp[11]) ? node153 : node150;
										assign node150 = (inp[1]) ? 3'b001 : 3'b001;
										assign node153 = (inp[1]) ? 3'b001 : 3'b110;
									assign node156 = (inp[1]) ? node160 : node157;
										assign node157 = (inp[11]) ? 3'b010 : 3'b110;
										assign node160 = (inp[11]) ? 3'b110 : 3'b001;
								assign node163 = (inp[10]) ? node171 : node164;
									assign node164 = (inp[8]) ? node168 : node165;
										assign node165 = (inp[1]) ? 3'b101 : 3'b001;
										assign node168 = (inp[1]) ? 3'b011 : 3'b101;
									assign node171 = (inp[1]) ? 3'b001 : node172;
										assign node172 = (inp[2]) ? 3'b001 : 3'b110;
							assign node176 = (inp[10]) ? node190 : node177;
								assign node177 = (inp[1]) ? node185 : node178;
									assign node178 = (inp[7]) ? node182 : node179;
										assign node179 = (inp[8]) ? 3'b001 : 3'b101;
										assign node182 = (inp[2]) ? 3'b011 : 3'b001;
									assign node185 = (inp[7]) ? node187 : 3'b011;
										assign node187 = (inp[8]) ? 3'b111 : 3'b011;
								assign node190 = (inp[11]) ? node198 : node191;
									assign node191 = (inp[8]) ? node195 : node192;
										assign node192 = (inp[1]) ? 3'b101 : 3'b001;
										assign node195 = (inp[2]) ? 3'b011 : 3'b001;
									assign node198 = (inp[1]) ? node202 : node199;
										assign node199 = (inp[8]) ? 3'b001 : 3'b000;
										assign node202 = (inp[8]) ? 3'b101 : 3'b101;
						assign node205 = (inp[0]) ? node235 : node206;
							assign node206 = (inp[10]) ? node222 : node207;
								assign node207 = (inp[7]) ? node215 : node208;
									assign node208 = (inp[1]) ? node212 : node209;
										assign node209 = (inp[11]) ? 3'b010 : 3'b110;
										assign node212 = (inp[2]) ? 3'b001 : 3'b110;
									assign node215 = (inp[1]) ? node219 : node216;
										assign node216 = (inp[2]) ? 3'b001 : 3'b110;
										assign node219 = (inp[8]) ? 3'b001 : 3'b001;
								assign node222 = (inp[11]) ? node230 : node223;
									assign node223 = (inp[7]) ? node227 : node224;
										assign node224 = (inp[1]) ? 3'b110 : 3'b010;
										assign node227 = (inp[8]) ? 3'b110 : 3'b110;
									assign node230 = (inp[1]) ? node232 : 3'b010;
										assign node232 = (inp[7]) ? 3'b110 : 3'b010;
							assign node235 = (inp[7]) ? node251 : node236;
								assign node236 = (inp[10]) ? node244 : node237;
									assign node237 = (inp[1]) ? node241 : node238;
										assign node238 = (inp[8]) ? 3'b001 : 3'b000;
										assign node241 = (inp[11]) ? 3'b101 : 3'b101;
									assign node244 = (inp[1]) ? node248 : node245;
										assign node245 = (inp[11]) ? 3'b110 : 3'b110;
										assign node248 = (inp[11]) ? 3'b110 : 3'b001;
								assign node251 = (inp[11]) ? node257 : node252;
									assign node252 = (inp[10]) ? 3'b101 : node253;
										assign node253 = (inp[1]) ? 3'b011 : 3'b101;
									assign node257 = (inp[10]) ? node261 : node258;
										assign node258 = (inp[8]) ? 3'b101 : 3'b001;
										assign node261 = (inp[1]) ? 3'b001 : 3'b001;
					assign node264 = (inp[0]) ? node320 : node265;
						assign node265 = (inp[7]) ? node291 : node266;
							assign node266 = (inp[5]) ? node280 : node267;
								assign node267 = (inp[10]) ? node273 : node268;
									assign node268 = (inp[11]) ? node270 : 3'b011;
										assign node270 = (inp[1]) ? 3'b011 : 3'b101;
									assign node273 = (inp[11]) ? node277 : node274;
										assign node274 = (inp[2]) ? 3'b101 : 3'b101;
										assign node277 = (inp[1]) ? 3'b101 : 3'b001;
								assign node280 = (inp[10]) ? node286 : node281;
									assign node281 = (inp[8]) ? 3'b101 : node282;
										assign node282 = (inp[1]) ? 3'b101 : 3'b001;
									assign node286 = (inp[1]) ? 3'b001 : node287;
										assign node287 = (inp[8]) ? 3'b001 : 3'b110;
							assign node291 = (inp[5]) ? node307 : node292;
								assign node292 = (inp[1]) ? node300 : node293;
									assign node293 = (inp[10]) ? node297 : node294;
										assign node294 = (inp[11]) ? 3'b011 : 3'b011;
										assign node297 = (inp[8]) ? 3'b001 : 3'b101;
									assign node300 = (inp[10]) ? node304 : node301;
										assign node301 = (inp[11]) ? 3'b111 : 3'b111;
										assign node304 = (inp[2]) ? 3'b011 : 3'b011;
								assign node307 = (inp[10]) ? node315 : node308;
									assign node308 = (inp[1]) ? node312 : node309;
										assign node309 = (inp[11]) ? 3'b101 : 3'b101;
										assign node312 = (inp[8]) ? 3'b011 : 3'b011;
									assign node315 = (inp[11]) ? node317 : 3'b101;
										assign node317 = (inp[1]) ? 3'b101 : 3'b001;
						assign node320 = (inp[10]) ? node342 : node321;
							assign node321 = (inp[5]) ? node329 : node322;
								assign node322 = (inp[11]) ? node324 : 3'b111;
									assign node324 = (inp[1]) ? 3'b111 : node325;
										assign node325 = (inp[2]) ? 3'b111 : 3'b011;
								assign node329 = (inp[7]) ? node337 : node330;
									assign node330 = (inp[1]) ? node334 : node331;
										assign node331 = (inp[2]) ? 3'b011 : 3'b011;
										assign node334 = (inp[8]) ? 3'b111 : 3'b011;
									assign node337 = (inp[11]) ? node339 : 3'b111;
										assign node339 = (inp[1]) ? 3'b111 : 3'b011;
							assign node342 = (inp[5]) ? node356 : node343;
								assign node343 = (inp[7]) ? node351 : node344;
									assign node344 = (inp[2]) ? node348 : node345;
										assign node345 = (inp[11]) ? 3'b011 : 3'b011;
										assign node348 = (inp[1]) ? 3'b011 : 3'b011;
									assign node351 = (inp[1]) ? 3'b111 : node352;
										assign node352 = (inp[8]) ? 3'b111 : 3'b011;
								assign node356 = (inp[1]) ? node364 : node357;
									assign node357 = (inp[2]) ? node361 : node358;
										assign node358 = (inp[8]) ? 3'b101 : 3'b001;
										assign node361 = (inp[7]) ? 3'b011 : 3'b101;
									assign node364 = (inp[2]) ? node368 : node365;
										assign node365 = (inp[7]) ? 3'b011 : 3'b101;
										assign node368 = (inp[11]) ? 3'b011 : 3'b011;
			assign node371 = (inp[4]) ? node595 : node372;
				assign node372 = (inp[6]) ? node488 : node373;
					assign node373 = (inp[0]) ? node429 : node374;
						assign node374 = (inp[10]) ? node402 : node375;
							assign node375 = (inp[5]) ? node389 : node376;
								assign node376 = (inp[7]) ? node384 : node377;
									assign node377 = (inp[1]) ? node381 : node378;
										assign node378 = (inp[2]) ? 3'b001 : 3'b110;
										assign node381 = (inp[11]) ? 3'b001 : 3'b101;
									assign node384 = (inp[1]) ? 3'b101 : node385;
										assign node385 = (inp[2]) ? 3'b101 : 3'b001;
								assign node389 = (inp[11]) ? node397 : node390;
									assign node390 = (inp[1]) ? node394 : node391;
										assign node391 = (inp[7]) ? 3'b001 : 3'b110;
										assign node394 = (inp[8]) ? 3'b001 : 3'b001;
									assign node397 = (inp[8]) ? node399 : 3'b110;
										assign node399 = (inp[1]) ? 3'b110 : 3'b110;
							assign node402 = (inp[5]) ? node416 : node403;
								assign node403 = (inp[7]) ? node411 : node404;
									assign node404 = (inp[1]) ? node408 : node405;
										assign node405 = (inp[8]) ? 3'b110 : 3'b010;
										assign node408 = (inp[11]) ? 3'b110 : 3'b001;
									assign node411 = (inp[8]) ? node413 : 3'b110;
										assign node413 = (inp[11]) ? 3'b000 : 3'b001;
								assign node416 = (inp[11]) ? node424 : node417;
									assign node417 = (inp[7]) ? node421 : node418;
										assign node418 = (inp[1]) ? 3'b010 : 3'b000;
										assign node421 = (inp[2]) ? 3'b110 : 3'b110;
									assign node424 = (inp[8]) ? node426 : 3'b010;
										assign node426 = (inp[7]) ? 3'b110 : 3'b010;
						assign node429 = (inp[10]) ? node459 : node430;
							assign node430 = (inp[7]) ? node446 : node431;
								assign node431 = (inp[2]) ? node439 : node432;
									assign node432 = (inp[1]) ? node436 : node433;
										assign node433 = (inp[5]) ? 3'b001 : 3'b101;
										assign node436 = (inp[5]) ? 3'b001 : 3'b011;
									assign node439 = (inp[5]) ? node443 : node440;
										assign node440 = (inp[1]) ? 3'b011 : 3'b101;
										assign node443 = (inp[1]) ? 3'b101 : 3'b001;
								assign node446 = (inp[8]) ? node454 : node447;
									assign node447 = (inp[5]) ? node451 : node448;
										assign node448 = (inp[2]) ? 3'b011 : 3'b111;
										assign node451 = (inp[11]) ? 3'b101 : 3'b011;
									assign node454 = (inp[1]) ? node456 : 3'b011;
										assign node456 = (inp[11]) ? 3'b011 : 3'b111;
							assign node459 = (inp[5]) ? node475 : node460;
								assign node460 = (inp[1]) ? node468 : node461;
									assign node461 = (inp[7]) ? node465 : node462;
										assign node462 = (inp[2]) ? 3'b001 : 3'b000;
										assign node465 = (inp[8]) ? 3'b101 : 3'b101;
									assign node468 = (inp[7]) ? node472 : node469;
										assign node469 = (inp[11]) ? 3'b001 : 3'b101;
										assign node472 = (inp[11]) ? 3'b101 : 3'b011;
								assign node475 = (inp[11]) ? node483 : node476;
									assign node476 = (inp[7]) ? node480 : node477;
										assign node477 = (inp[2]) ? 3'b001 : 3'b000;
										assign node480 = (inp[1]) ? 3'b101 : 3'b001;
									assign node483 = (inp[1]) ? node485 : 3'b110;
										assign node485 = (inp[7]) ? 3'b001 : 3'b000;
					assign node488 = (inp[0]) ? node544 : node489;
						assign node489 = (inp[5]) ? node513 : node490;
							assign node490 = (inp[1]) ? node500 : node491;
								assign node491 = (inp[7]) ? node495 : node492;
									assign node492 = (inp[10]) ? 3'b001 : 3'b101;
									assign node495 = (inp[11]) ? node497 : 3'b011;
										assign node497 = (inp[8]) ? 3'b011 : 3'b001;
								assign node500 = (inp[2]) ? node506 : node501;
									assign node501 = (inp[10]) ? 3'b011 : node502;
										assign node502 = (inp[7]) ? 3'b111 : 3'b011;
									assign node506 = (inp[8]) ? node510 : node507;
										assign node507 = (inp[10]) ? 3'b101 : 3'b011;
										assign node510 = (inp[10]) ? 3'b011 : 3'b111;
							assign node513 = (inp[10]) ? node529 : node514;
								assign node514 = (inp[1]) ? node522 : node515;
									assign node515 = (inp[8]) ? node519 : node516;
										assign node516 = (inp[7]) ? 3'b001 : 3'b001;
										assign node519 = (inp[7]) ? 3'b101 : 3'b001;
									assign node522 = (inp[7]) ? node526 : node523;
										assign node523 = (inp[8]) ? 3'b001 : 3'b101;
										assign node526 = (inp[11]) ? 3'b011 : 3'b011;
								assign node529 = (inp[1]) ? node537 : node530;
									assign node530 = (inp[7]) ? node534 : node531;
										assign node531 = (inp[11]) ? 3'b110 : 3'b000;
										assign node534 = (inp[8]) ? 3'b001 : 3'b000;
									assign node537 = (inp[11]) ? node541 : node538;
										assign node538 = (inp[7]) ? 3'b101 : 3'b001;
										assign node541 = (inp[8]) ? 3'b001 : 3'b000;
						assign node544 = (inp[10]) ? node566 : node545;
							assign node545 = (inp[5]) ? node553 : node546;
								assign node546 = (inp[11]) ? node548 : 3'b111;
									assign node548 = (inp[1]) ? 3'b111 : node549;
										assign node549 = (inp[8]) ? 3'b111 : 3'b011;
								assign node553 = (inp[7]) ? node561 : node554;
									assign node554 = (inp[1]) ? node558 : node555;
										assign node555 = (inp[8]) ? 3'b011 : 3'b101;
										assign node558 = (inp[8]) ? 3'b111 : 3'b011;
									assign node561 = (inp[1]) ? 3'b111 : node562;
										assign node562 = (inp[2]) ? 3'b111 : 3'b011;
							assign node566 = (inp[5]) ? node582 : node567;
								assign node567 = (inp[2]) ? node575 : node568;
									assign node568 = (inp[11]) ? node572 : node569;
										assign node569 = (inp[7]) ? 3'b111 : 3'b011;
										assign node572 = (inp[1]) ? 3'b011 : 3'b101;
									assign node575 = (inp[1]) ? node579 : node576;
										assign node576 = (inp[8]) ? 3'b111 : 3'b011;
										assign node579 = (inp[8]) ? 3'b111 : 3'b111;
								assign node582 = (inp[1]) ? node588 : node583;
									assign node583 = (inp[2]) ? node585 : 3'b101;
										assign node585 = (inp[7]) ? 3'b011 : 3'b101;
									assign node588 = (inp[8]) ? node592 : node589;
										assign node589 = (inp[7]) ? 3'b011 : 3'b101;
										assign node592 = (inp[7]) ? 3'b011 : 3'b011;
				assign node595 = (inp[6]) ? node715 : node596;
					assign node596 = (inp[0]) ? node656 : node597;
						assign node597 = (inp[10]) ? node627 : node598;
							assign node598 = (inp[7]) ? node614 : node599;
								assign node599 = (inp[5]) ? node607 : node600;
									assign node600 = (inp[1]) ? node604 : node601;
										assign node601 = (inp[2]) ? 3'b010 : 3'b100;
										assign node604 = (inp[11]) ? 3'b010 : 3'b010;
									assign node607 = (inp[1]) ? node611 : node608;
										assign node608 = (inp[8]) ? 3'b100 : 3'b000;
										assign node611 = (inp[2]) ? 3'b000 : 3'b100;
								assign node614 = (inp[5]) ? node622 : node615;
									assign node615 = (inp[1]) ? node619 : node616;
										assign node616 = (inp[11]) ? 3'b010 : 3'b110;
										assign node619 = (inp[8]) ? 3'b000 : 3'b110;
									assign node622 = (inp[1]) ? 3'b010 : node623;
										assign node623 = (inp[11]) ? 3'b100 : 3'b010;
							assign node627 = (inp[5]) ? node643 : node628;
								assign node628 = (inp[7]) ? node636 : node629;
									assign node629 = (inp[8]) ? node633 : node630;
										assign node630 = (inp[11]) ? 3'b000 : 3'b100;
										assign node633 = (inp[11]) ? 3'b100 : 3'b000;
									assign node636 = (inp[11]) ? node640 : node637;
										assign node637 = (inp[8]) ? 3'b010 : 3'b000;
										assign node640 = (inp[1]) ? 3'b010 : 3'b100;
								assign node643 = (inp[1]) ? node649 : node644;
									assign node644 = (inp[8]) ? node646 : 3'b000;
										assign node646 = (inp[2]) ? 3'b000 : 3'b000;
									assign node649 = (inp[7]) ? node653 : node650;
										assign node650 = (inp[2]) ? 3'b000 : 3'b000;
										assign node653 = (inp[2]) ? 3'b100 : 3'b100;
						assign node656 = (inp[5]) ? node686 : node657;
							assign node657 = (inp[10]) ? node673 : node658;
								assign node658 = (inp[11]) ? node666 : node659;
									assign node659 = (inp[1]) ? node663 : node660;
										assign node660 = (inp[7]) ? 3'b001 : 3'b110;
										assign node663 = (inp[7]) ? 3'b101 : 3'b001;
									assign node666 = (inp[7]) ? node670 : node667;
										assign node667 = (inp[2]) ? 3'b110 : 3'b110;
										assign node670 = (inp[8]) ? 3'b001 : 3'b000;
								assign node673 = (inp[1]) ? node681 : node674;
									assign node674 = (inp[11]) ? node678 : node675;
										assign node675 = (inp[7]) ? 3'b110 : 3'b010;
										assign node678 = (inp[8]) ? 3'b010 : 3'b000;
									assign node681 = (inp[7]) ? node683 : 3'b110;
										assign node683 = (inp[8]) ? 3'b001 : 3'b110;
							assign node686 = (inp[10]) ? node700 : node687;
								assign node687 = (inp[1]) ? node695 : node688;
									assign node688 = (inp[7]) ? node692 : node689;
										assign node689 = (inp[11]) ? 3'b010 : 3'b010;
										assign node692 = (inp[8]) ? 3'b110 : 3'b010;
									assign node695 = (inp[7]) ? node697 : 3'b110;
										assign node697 = (inp[11]) ? 3'b110 : 3'b001;
								assign node700 = (inp[7]) ? node708 : node701;
									assign node701 = (inp[1]) ? node705 : node702;
										assign node702 = (inp[2]) ? 3'b100 : 3'b100;
										assign node705 = (inp[11]) ? 3'b100 : 3'b010;
									assign node708 = (inp[1]) ? node712 : node709;
										assign node709 = (inp[11]) ? 3'b100 : 3'b010;
										assign node712 = (inp[2]) ? 3'b110 : 3'b010;
					assign node715 = (inp[0]) ? node777 : node716;
						assign node716 = (inp[10]) ? node748 : node717;
							assign node717 = (inp[5]) ? node733 : node718;
								assign node718 = (inp[1]) ? node726 : node719;
									assign node719 = (inp[7]) ? node723 : node720;
										assign node720 = (inp[2]) ? 3'b110 : 3'b010;
										assign node723 = (inp[11]) ? 3'b110 : 3'b001;
									assign node726 = (inp[7]) ? node730 : node727;
										assign node727 = (inp[11]) ? 3'b001 : 3'b001;
										assign node730 = (inp[8]) ? 3'b101 : 3'b001;
								assign node733 = (inp[7]) ? node741 : node734;
									assign node734 = (inp[1]) ? node738 : node735;
										assign node735 = (inp[11]) ? 3'b000 : 3'b010;
										assign node738 = (inp[2]) ? 3'b110 : 3'b110;
									assign node741 = (inp[11]) ? node745 : node742;
										assign node742 = (inp[1]) ? 3'b001 : 3'b110;
										assign node745 = (inp[2]) ? 3'b110 : 3'b010;
							assign node748 = (inp[5]) ? node762 : node749;
								assign node749 = (inp[7]) ? node755 : node750;
									assign node750 = (inp[8]) ? 3'b110 : node751;
										assign node751 = (inp[1]) ? 3'b110 : 3'b010;
									assign node755 = (inp[1]) ? node759 : node756;
										assign node756 = (inp[11]) ? 3'b110 : 3'b110;
										assign node759 = (inp[2]) ? 3'b001 : 3'b000;
								assign node762 = (inp[7]) ? node770 : node763;
									assign node763 = (inp[11]) ? node767 : node764;
										assign node764 = (inp[1]) ? 3'b010 : 3'b000;
										assign node767 = (inp[8]) ? 3'b100 : 3'b100;
									assign node770 = (inp[2]) ? node774 : node771;
										assign node771 = (inp[1]) ? 3'b010 : 3'b010;
										assign node774 = (inp[8]) ? 3'b110 : 3'b010;
						assign node777 = (inp[5]) ? node809 : node778;
							assign node778 = (inp[10]) ? node794 : node779;
								assign node779 = (inp[7]) ? node787 : node780;
									assign node780 = (inp[1]) ? node784 : node781;
										assign node781 = (inp[11]) ? 3'b001 : 3'b101;
										assign node784 = (inp[2]) ? 3'b011 : 3'b101;
									assign node787 = (inp[8]) ? node791 : node788;
										assign node788 = (inp[1]) ? 3'b011 : 3'b101;
										assign node791 = (inp[11]) ? 3'b011 : 3'b011;
								assign node794 = (inp[11]) ? node802 : node795;
									assign node795 = (inp[2]) ? node799 : node796;
										assign node796 = (inp[7]) ? 3'b101 : 3'b001;
										assign node799 = (inp[8]) ? 3'b001 : 3'b101;
									assign node802 = (inp[7]) ? node806 : node803;
										assign node803 = (inp[1]) ? 3'b001 : 3'b110;
										assign node806 = (inp[8]) ? 3'b001 : 3'b001;
							assign node809 = (inp[7]) ? node825 : node810;
								assign node810 = (inp[8]) ? node818 : node811;
									assign node811 = (inp[10]) ? node815 : node812;
										assign node812 = (inp[1]) ? 3'b001 : 3'b110;
										assign node815 = (inp[1]) ? 3'b110 : 3'b010;
									assign node818 = (inp[11]) ? node822 : node819;
										assign node819 = (inp[1]) ? 3'b101 : 3'b001;
										assign node822 = (inp[2]) ? 3'b000 : 3'b110;
								assign node825 = (inp[10]) ? node833 : node826;
									assign node826 = (inp[2]) ? node830 : node827;
										assign node827 = (inp[1]) ? 3'b001 : 3'b001;
										assign node830 = (inp[1]) ? 3'b101 : 3'b101;
									assign node833 = (inp[11]) ? node835 : 3'b001;
										assign node835 = (inp[2]) ? 3'b001 : 3'b110;
		assign node838 = (inp[9]) ? node1260 : node839;
			assign node839 = (inp[4]) ? node1083 : node840;
				assign node840 = (inp[6]) ? node960 : node841;
					assign node841 = (inp[0]) ? node901 : node842;
						assign node842 = (inp[5]) ? node874 : node843;
							assign node843 = (inp[10]) ? node859 : node844;
								assign node844 = (inp[11]) ? node852 : node845;
									assign node845 = (inp[2]) ? node849 : node846;
										assign node846 = (inp[1]) ? 3'b110 : 3'b010;
										assign node849 = (inp[1]) ? 3'b000 : 3'b110;
									assign node852 = (inp[1]) ? node856 : node853;
										assign node853 = (inp[7]) ? 3'b010 : 3'b100;
										assign node856 = (inp[2]) ? 3'b010 : 3'b010;
								assign node859 = (inp[1]) ? node867 : node860;
									assign node860 = (inp[11]) ? node864 : node861;
										assign node861 = (inp[7]) ? 3'b000 : 3'b100;
										assign node864 = (inp[7]) ? 3'b100 : 3'b000;
									assign node867 = (inp[7]) ? node871 : node868;
										assign node868 = (inp[8]) ? 3'b010 : 3'b100;
										assign node871 = (inp[11]) ? 3'b010 : 3'b010;
							assign node874 = (inp[10]) ? node888 : node875;
								assign node875 = (inp[7]) ? node881 : node876;
									assign node876 = (inp[2]) ? 3'b100 : node877;
										assign node877 = (inp[1]) ? 3'b100 : 3'b000;
									assign node881 = (inp[2]) ? node885 : node882;
										assign node882 = (inp[1]) ? 3'b010 : 3'b100;
										assign node885 = (inp[1]) ? 3'b010 : 3'b010;
								assign node888 = (inp[7]) ? node894 : node889;
									assign node889 = (inp[8]) ? node891 : 3'b000;
										assign node891 = (inp[11]) ? 3'b000 : 3'b000;
									assign node894 = (inp[1]) ? node898 : node895;
										assign node895 = (inp[8]) ? 3'b000 : 3'b000;
										assign node898 = (inp[2]) ? 3'b100 : 3'b100;
						assign node901 = (inp[10]) ? node931 : node902;
							assign node902 = (inp[1]) ? node916 : node903;
								assign node903 = (inp[11]) ? node911 : node904;
									assign node904 = (inp[2]) ? node908 : node905;
										assign node905 = (inp[7]) ? 3'b110 : 3'b010;
										assign node908 = (inp[5]) ? 3'b001 : 3'b001;
									assign node911 = (inp[7]) ? 3'b110 : node912;
										assign node912 = (inp[5]) ? 3'b010 : 3'b110;
								assign node916 = (inp[5]) ? node924 : node917;
									assign node917 = (inp[7]) ? node921 : node918;
										assign node918 = (inp[11]) ? 3'b001 : 3'b001;
										assign node921 = (inp[2]) ? 3'b101 : 3'b001;
									assign node924 = (inp[7]) ? node928 : node925;
										assign node925 = (inp[8]) ? 3'b110 : 3'b010;
										assign node928 = (inp[11]) ? 3'b110 : 3'b001;
							assign node931 = (inp[5]) ? node945 : node932;
								assign node932 = (inp[7]) ? node940 : node933;
									assign node933 = (inp[1]) ? node937 : node934;
										assign node934 = (inp[11]) ? 3'b010 : 3'b010;
										assign node937 = (inp[11]) ? 3'b010 : 3'b110;
									assign node940 = (inp[1]) ? node942 : 3'b110;
										assign node942 = (inp[8]) ? 3'b001 : 3'b110;
								assign node945 = (inp[11]) ? node953 : node946;
									assign node946 = (inp[1]) ? node950 : node947;
										assign node947 = (inp[2]) ? 3'b010 : 3'b100;
										assign node950 = (inp[8]) ? 3'b010 : 3'b010;
									assign node953 = (inp[7]) ? node957 : node954;
										assign node954 = (inp[2]) ? 3'b100 : 3'b100;
										assign node957 = (inp[2]) ? 3'b010 : 3'b100;
					assign node960 = (inp[0]) ? node1022 : node961;
						assign node961 = (inp[10]) ? node993 : node962;
							assign node962 = (inp[5]) ? node978 : node963;
								assign node963 = (inp[1]) ? node971 : node964;
									assign node964 = (inp[11]) ? node968 : node965;
										assign node965 = (inp[8]) ? 3'b101 : 3'b001;
										assign node968 = (inp[8]) ? 3'b001 : 3'b110;
									assign node971 = (inp[7]) ? node975 : node972;
										assign node972 = (inp[11]) ? 3'b001 : 3'b001;
										assign node975 = (inp[2]) ? 3'b101 : 3'b101;
								assign node978 = (inp[11]) ? node986 : node979;
									assign node979 = (inp[7]) ? node983 : node980;
										assign node980 = (inp[8]) ? 3'b010 : 3'b110;
										assign node983 = (inp[1]) ? 3'b001 : 3'b110;
									assign node986 = (inp[7]) ? node990 : node987;
										assign node987 = (inp[1]) ? 3'b110 : 3'b010;
										assign node990 = (inp[1]) ? 3'b110 : 3'b110;
							assign node993 = (inp[8]) ? node1007 : node994;
								assign node994 = (inp[7]) ? node1002 : node995;
									assign node995 = (inp[5]) ? node999 : node996;
										assign node996 = (inp[1]) ? 3'b110 : 3'b010;
										assign node999 = (inp[11]) ? 3'b000 : 3'b010;
									assign node1002 = (inp[5]) ? node1004 : 3'b110;
										assign node1004 = (inp[11]) ? 3'b010 : 3'b110;
								assign node1007 = (inp[5]) ? node1015 : node1008;
									assign node1008 = (inp[11]) ? node1012 : node1009;
										assign node1009 = (inp[7]) ? 3'b001 : 3'b000;
										assign node1012 = (inp[7]) ? 3'b110 : 3'b010;
									assign node1015 = (inp[2]) ? node1019 : node1016;
										assign node1016 = (inp[1]) ? 3'b010 : 3'b000;
										assign node1019 = (inp[11]) ? 3'b100 : 3'b110;
						assign node1022 = (inp[7]) ? node1054 : node1023;
							assign node1023 = (inp[5]) ? node1039 : node1024;
								assign node1024 = (inp[8]) ? node1032 : node1025;
									assign node1025 = (inp[10]) ? node1029 : node1026;
										assign node1026 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1029 = (inp[2]) ? 3'b001 : 3'b001;
									assign node1032 = (inp[1]) ? node1036 : node1033;
										assign node1033 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1036 = (inp[10]) ? 3'b101 : 3'b011;
								assign node1039 = (inp[10]) ? node1047 : node1040;
									assign node1040 = (inp[1]) ? node1044 : node1041;
										assign node1041 = (inp[8]) ? 3'b001 : 3'b110;
										assign node1044 = (inp[8]) ? 3'b101 : 3'b001;
									assign node1047 = (inp[11]) ? node1051 : node1048;
										assign node1048 = (inp[1]) ? 3'b001 : 3'b110;
										assign node1051 = (inp[1]) ? 3'b110 : 3'b010;
							assign node1054 = (inp[10]) ? node1070 : node1055;
								assign node1055 = (inp[5]) ? node1063 : node1056;
									assign node1056 = (inp[1]) ? node1060 : node1057;
										assign node1057 = (inp[11]) ? 3'b101 : 3'b011;
										assign node1060 = (inp[11]) ? 3'b011 : 3'b111;
									assign node1063 = (inp[11]) ? node1067 : node1064;
										assign node1064 = (inp[2]) ? 3'b011 : 3'b101;
										assign node1067 = (inp[1]) ? 3'b101 : 3'b001;
								assign node1070 = (inp[8]) ? node1076 : node1071;
									assign node1071 = (inp[5]) ? 3'b001 : node1072;
										assign node1072 = (inp[1]) ? 3'b101 : 3'b001;
									assign node1076 = (inp[1]) ? node1080 : node1077;
										assign node1077 = (inp[5]) ? 3'b110 : 3'b101;
										assign node1080 = (inp[5]) ? 3'b001 : 3'b011;
				assign node1083 = (inp[6]) ? node1149 : node1084;
					assign node1084 = (inp[0]) ? node1102 : node1085;
						assign node1085 = (inp[10]) ? 3'b000 : node1086;
							assign node1086 = (inp[5]) ? 3'b000 : node1087;
								assign node1087 = (inp[1]) ? node1093 : node1088;
									assign node1088 = (inp[8]) ? node1090 : 3'b000;
										assign node1090 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1093 = (inp[7]) ? node1097 : node1094;
										assign node1094 = (inp[2]) ? 3'b000 : 3'b000;
										assign node1097 = (inp[2]) ? 3'b100 : 3'b100;
						assign node1102 = (inp[5]) ? node1128 : node1103;
							assign node1103 = (inp[10]) ? node1115 : node1104;
								assign node1104 = (inp[7]) ? node1110 : node1105;
									assign node1105 = (inp[11]) ? 3'b100 : node1106;
										assign node1106 = (inp[1]) ? 3'b010 : 3'b100;
									assign node1110 = (inp[11]) ? node1112 : 3'b010;
										assign node1112 = (inp[8]) ? 3'b010 : 3'b010;
								assign node1115 = (inp[7]) ? node1121 : node1116;
									assign node1116 = (inp[8]) ? node1118 : 3'b000;
										assign node1118 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1121 = (inp[2]) ? node1125 : node1122;
										assign node1122 = (inp[8]) ? 3'b100 : 3'b100;
										assign node1125 = (inp[1]) ? 3'b010 : 3'b000;
							assign node1128 = (inp[11]) ? node1142 : node1129;
								assign node1129 = (inp[10]) ? node1137 : node1130;
									assign node1130 = (inp[7]) ? node1134 : node1131;
										assign node1131 = (inp[1]) ? 3'b100 : 3'b000;
										assign node1134 = (inp[1]) ? 3'b010 : 3'b100;
									assign node1137 = (inp[7]) ? node1139 : 3'b000;
										assign node1139 = (inp[2]) ? 3'b100 : 3'b000;
								assign node1142 = (inp[8]) ? node1144 : 3'b000;
									assign node1144 = (inp[1]) ? node1146 : 3'b000;
										assign node1146 = (inp[7]) ? 3'b100 : 3'b000;
					assign node1149 = (inp[0]) ? node1199 : node1150;
						assign node1150 = (inp[10]) ? node1178 : node1151;
							assign node1151 = (inp[7]) ? node1165 : node1152;
								assign node1152 = (inp[8]) ? node1160 : node1153;
									assign node1153 = (inp[5]) ? node1157 : node1154;
										assign node1154 = (inp[1]) ? 3'b010 : 3'b100;
										assign node1157 = (inp[1]) ? 3'b000 : 3'b000;
									assign node1160 = (inp[5]) ? 3'b100 : node1161;
										assign node1161 = (inp[1]) ? 3'b010 : 3'b100;
								assign node1165 = (inp[5]) ? node1171 : node1166;
									assign node1166 = (inp[1]) ? node1168 : 3'b010;
										assign node1168 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1171 = (inp[11]) ? node1175 : node1172;
										assign node1172 = (inp[1]) ? 3'b010 : 3'b000;
										assign node1175 = (inp[8]) ? 3'b100 : 3'b100;
							assign node1178 = (inp[5]) ? node1192 : node1179;
								assign node1179 = (inp[7]) ? node1185 : node1180;
									assign node1180 = (inp[8]) ? 3'b100 : node1181;
										assign node1181 = (inp[1]) ? 3'b000 : 3'b000;
									assign node1185 = (inp[2]) ? node1189 : node1186;
										assign node1186 = (inp[11]) ? 3'b100 : 3'b100;
										assign node1189 = (inp[8]) ? 3'b010 : 3'b100;
								assign node1192 = (inp[7]) ? node1194 : 3'b000;
									assign node1194 = (inp[2]) ? node1196 : 3'b000;
										assign node1196 = (inp[1]) ? 3'b100 : 3'b000;
						assign node1199 = (inp[5]) ? node1231 : node1200;
							assign node1200 = (inp[10]) ? node1216 : node1201;
								assign node1201 = (inp[1]) ? node1209 : node1202;
									assign node1202 = (inp[7]) ? node1206 : node1203;
										assign node1203 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1206 = (inp[2]) ? 3'b001 : 3'b110;
									assign node1209 = (inp[8]) ? node1213 : node1210;
										assign node1210 = (inp[7]) ? 3'b001 : 3'b110;
										assign node1213 = (inp[2]) ? 3'b001 : 3'b001;
								assign node1216 = (inp[11]) ? node1224 : node1217;
									assign node1217 = (inp[7]) ? node1221 : node1218;
										assign node1218 = (inp[1]) ? 3'b110 : 3'b010;
										assign node1221 = (inp[8]) ? 3'b110 : 3'b110;
									assign node1224 = (inp[7]) ? node1228 : node1225;
										assign node1225 = (inp[1]) ? 3'b010 : 3'b100;
										assign node1228 = (inp[1]) ? 3'b110 : 3'b010;
							assign node1231 = (inp[10]) ? node1245 : node1232;
								assign node1232 = (inp[11]) ? node1240 : node1233;
									assign node1233 = (inp[7]) ? node1237 : node1234;
										assign node1234 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1237 = (inp[1]) ? 3'b110 : 3'b110;
									assign node1240 = (inp[1]) ? 3'b010 : node1241;
										assign node1241 = (inp[7]) ? 3'b010 : 3'b100;
								assign node1245 = (inp[11]) ? node1253 : node1246;
									assign node1246 = (inp[7]) ? node1250 : node1247;
										assign node1247 = (inp[1]) ? 3'b010 : 3'b100;
										assign node1250 = (inp[8]) ? 3'b010 : 3'b010;
									assign node1253 = (inp[1]) ? node1257 : node1254;
										assign node1254 = (inp[7]) ? 3'b100 : 3'b000;
										assign node1257 = (inp[8]) ? 3'b000 : 3'b100;
			assign node1260 = (inp[4]) ? node1440 : node1261;
				assign node1261 = (inp[6]) ? node1333 : node1262;
					assign node1262 = (inp[0]) ? node1286 : node1263;
						assign node1263 = (inp[1]) ? node1265 : 3'b000;
							assign node1265 = (inp[10]) ? node1279 : node1266;
								assign node1266 = (inp[8]) ? node1272 : node1267;
									assign node1267 = (inp[7]) ? node1269 : 3'b000;
										assign node1269 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1272 = (inp[5]) ? node1276 : node1273;
										assign node1273 = (inp[11]) ? 3'b100 : 3'b100;
										assign node1276 = (inp[2]) ? 3'b100 : 3'b000;
								assign node1279 = (inp[5]) ? 3'b000 : node1280;
									assign node1280 = (inp[7]) ? node1282 : 3'b000;
										assign node1282 = (inp[11]) ? 3'b000 : 3'b000;
						assign node1286 = (inp[5]) ? node1312 : node1287;
							assign node1287 = (inp[10]) ? node1299 : node1288;
								assign node1288 = (inp[2]) ? node1294 : node1289;
									assign node1289 = (inp[7]) ? node1291 : 3'b100;
										assign node1291 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1294 = (inp[8]) ? 3'b010 : node1295;
										assign node1295 = (inp[1]) ? 3'b010 : 3'b100;
								assign node1299 = (inp[7]) ? node1305 : node1300;
									assign node1300 = (inp[1]) ? node1302 : 3'b000;
										assign node1302 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1305 = (inp[11]) ? node1309 : node1306;
										assign node1306 = (inp[1]) ? 3'b010 : 3'b100;
										assign node1309 = (inp[1]) ? 3'b100 : 3'b000;
							assign node1312 = (inp[10]) ? node1326 : node1313;
								assign node1313 = (inp[7]) ? node1319 : node1314;
									assign node1314 = (inp[1]) ? node1316 : 3'b000;
										assign node1316 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1319 = (inp[2]) ? node1323 : node1320;
										assign node1320 = (inp[8]) ? 3'b000 : 3'b100;
										assign node1323 = (inp[11]) ? 3'b100 : 3'b010;
								assign node1326 = (inp[1]) ? node1328 : 3'b000;
									assign node1328 = (inp[2]) ? node1330 : 3'b000;
										assign node1330 = (inp[11]) ? 3'b000 : 3'b100;
					assign node1333 = (inp[0]) ? node1383 : node1334;
						assign node1334 = (inp[5]) ? node1362 : node1335;
							assign node1335 = (inp[10]) ? node1349 : node1336;
								assign node1336 = (inp[8]) ? node1344 : node1337;
									assign node1337 = (inp[7]) ? node1341 : node1338;
										assign node1338 = (inp[1]) ? 3'b000 : 3'b100;
										assign node1341 = (inp[2]) ? 3'b010 : 3'b110;
									assign node1344 = (inp[7]) ? node1346 : 3'b010;
										assign node1346 = (inp[1]) ? 3'b110 : 3'b010;
								assign node1349 = (inp[7]) ? node1357 : node1350;
									assign node1350 = (inp[11]) ? node1354 : node1351;
										assign node1351 = (inp[1]) ? 3'b100 : 3'b000;
										assign node1354 = (inp[8]) ? 3'b000 : 3'b000;
									assign node1357 = (inp[2]) ? node1359 : 3'b100;
										assign node1359 = (inp[1]) ? 3'b000 : 3'b100;
							assign node1362 = (inp[10]) ? node1376 : node1363;
								assign node1363 = (inp[7]) ? node1369 : node1364;
									assign node1364 = (inp[1]) ? node1366 : 3'b000;
										assign node1366 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1369 = (inp[1]) ? node1373 : node1370;
										assign node1370 = (inp[2]) ? 3'b100 : 3'b100;
										assign node1373 = (inp[2]) ? 3'b010 : 3'b100;
								assign node1376 = (inp[8]) ? node1378 : 3'b000;
									assign node1378 = (inp[1]) ? node1380 : 3'b000;
										assign node1380 = (inp[7]) ? 3'b100 : 3'b000;
						assign node1383 = (inp[5]) ? node1415 : node1384;
							assign node1384 = (inp[10]) ? node1400 : node1385;
								assign node1385 = (inp[11]) ? node1393 : node1386;
									assign node1386 = (inp[1]) ? node1390 : node1387;
										assign node1387 = (inp[7]) ? 3'b001 : 3'b110;
										assign node1390 = (inp[2]) ? 3'b001 : 3'b001;
									assign node1393 = (inp[8]) ? node1397 : node1394;
										assign node1394 = (inp[7]) ? 3'b110 : 3'b010;
										assign node1397 = (inp[7]) ? 3'b000 : 3'b110;
								assign node1400 = (inp[7]) ? node1408 : node1401;
									assign node1401 = (inp[1]) ? node1405 : node1402;
										assign node1402 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1405 = (inp[11]) ? 3'b010 : 3'b010;
									assign node1408 = (inp[11]) ? node1412 : node1409;
										assign node1409 = (inp[8]) ? 3'b110 : 3'b110;
										assign node1412 = (inp[1]) ? 3'b010 : 3'b010;
							assign node1415 = (inp[7]) ? node1431 : node1416;
								assign node1416 = (inp[10]) ? node1424 : node1417;
									assign node1417 = (inp[1]) ? node1421 : node1418;
										assign node1418 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1421 = (inp[11]) ? 3'b010 : 3'b010;
									assign node1424 = (inp[1]) ? node1428 : node1425;
										assign node1425 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1428 = (inp[11]) ? 3'b100 : 3'b000;
								assign node1431 = (inp[10]) ? node1435 : node1432;
									assign node1432 = (inp[1]) ? 3'b110 : 3'b010;
									assign node1435 = (inp[2]) ? node1437 : 3'b010;
										assign node1437 = (inp[1]) ? 3'b010 : 3'b000;
				assign node1440 = (inp[6]) ? node1454 : node1441;
					assign node1441 = (inp[1]) ? node1443 : 3'b000;
						assign node1443 = (inp[10]) ? 3'b000 : node1444;
							assign node1444 = (inp[0]) ? node1446 : 3'b000;
								assign node1446 = (inp[11]) ? 3'b000 : node1447;
									assign node1447 = (inp[7]) ? node1449 : 3'b000;
										assign node1449 = (inp[5]) ? 3'b000 : 3'b100;
					assign node1454 = (inp[0]) ? node1466 : node1455;
						assign node1455 = (inp[7]) ? node1457 : 3'b000;
							assign node1457 = (inp[1]) ? node1459 : 3'b000;
								assign node1459 = (inp[11]) ? 3'b000 : node1460;
									assign node1460 = (inp[5]) ? 3'b000 : node1461;
										assign node1461 = (inp[8]) ? 3'b100 : 3'b000;
						assign node1466 = (inp[10]) ? node1492 : node1467;
							assign node1467 = (inp[5]) ? node1479 : node1468;
								assign node1468 = (inp[7]) ? node1474 : node1469;
									assign node1469 = (inp[1]) ? 3'b100 : node1470;
										assign node1470 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1474 = (inp[11]) ? 3'b100 : node1475;
										assign node1475 = (inp[2]) ? 3'b010 : 3'b010;
								assign node1479 = (inp[7]) ? node1485 : node1480;
									assign node1480 = (inp[11]) ? 3'b000 : node1481;
										assign node1481 = (inp[2]) ? 3'b000 : 3'b000;
									assign node1485 = (inp[1]) ? node1489 : node1486;
										assign node1486 = (inp[11]) ? 3'b000 : 3'b000;
										assign node1489 = (inp[8]) ? 3'b100 : 3'b100;
							assign node1492 = (inp[7]) ? node1500 : node1493;
								assign node1493 = (inp[1]) ? node1495 : 3'b000;
									assign node1495 = (inp[11]) ? 3'b000 : node1496;
										assign node1496 = (inp[8]) ? 3'b000 : 3'b000;
								assign node1500 = (inp[5]) ? node1508 : node1501;
									assign node1501 = (inp[1]) ? node1505 : node1502;
										assign node1502 = (inp[11]) ? 3'b000 : 3'b000;
										assign node1505 = (inp[11]) ? 3'b100 : 3'b100;
									assign node1508 = (inp[11]) ? 3'b000 : node1509;
										assign node1509 = (inp[8]) ? 3'b000 : 3'b000;

endmodule