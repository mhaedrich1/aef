module dtc_split875_bm64 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node15;
	wire [4-1:0] node17;
	wire [4-1:0] node18;
	wire [4-1:0] node22;
	wire [4-1:0] node24;
	wire [4-1:0] node28;
	wire [4-1:0] node30;
	wire [4-1:0] node31;
	wire [4-1:0] node33;
	wire [4-1:0] node34;
	wire [4-1:0] node38;
	wire [4-1:0] node40;
	wire [4-1:0] node42;
	wire [4-1:0] node46;
	wire [4-1:0] node48;
	wire [4-1:0] node49;
	wire [4-1:0] node50;
	wire [4-1:0] node51;
	wire [4-1:0] node52;
	wire [4-1:0] node54;
	wire [4-1:0] node58;
	wire [4-1:0] node60;
	wire [4-1:0] node62;
	wire [4-1:0] node66;
	wire [4-1:0] node68;
	wire [4-1:0] node69;
	wire [4-1:0] node71;
	wire [4-1:0] node72;
	wire [4-1:0] node76;
	wire [4-1:0] node78;
	wire [4-1:0] node79;
	wire [4-1:0] node84;
	wire [4-1:0] node86;
	wire [4-1:0] node87;
	wire [4-1:0] node88;
	wire [4-1:0] node89;
	wire [4-1:0] node90;
	wire [4-1:0] node91;
	wire [4-1:0] node92;
	wire [4-1:0] node94;
	wire [4-1:0] node98;
	wire [4-1:0] node100;
	wire [4-1:0] node101;
	wire [4-1:0] node106;
	wire [4-1:0] node108;
	wire [4-1:0] node109;
	wire [4-1:0] node110;
	wire [4-1:0] node112;
	wire [4-1:0] node116;
	wire [4-1:0] node118;
	wire [4-1:0] node119;
	wire [4-1:0] node124;
	wire [4-1:0] node126;
	wire [4-1:0] node127;
	wire [4-1:0] node128;
	wire [4-1:0] node130;
	wire [4-1:0] node132;
	wire [4-1:0] node134;
	wire [4-1:0] node138;
	wire [4-1:0] node140;
	wire [4-1:0] node141;
	wire [4-1:0] node142;
	wire [4-1:0] node144;
	wire [4-1:0] node148;
	wire [4-1:0] node150;
	wire [4-1:0] node152;
	wire [4-1:0] node156;
	wire [4-1:0] node157;
	wire [4-1:0] node158;
	wire [4-1:0] node159;
	wire [4-1:0] node160;
	wire [4-1:0] node161;
	wire [4-1:0] node162;
	wire [4-1:0] node163;
	wire [4-1:0] node164;
	wire [4-1:0] node165;
	wire [4-1:0] node170;
	wire [4-1:0] node172;
	wire [4-1:0] node174;
	wire [4-1:0] node178;
	wire [4-1:0] node180;
	wire [4-1:0] node181;
	wire [4-1:0] node182;
	wire [4-1:0] node183;
	wire [4-1:0] node188;
	wire [4-1:0] node190;
	wire [4-1:0] node192;
	wire [4-1:0] node196;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node200;
	wire [4-1:0] node201;
	wire [4-1:0] node203;
	wire [4-1:0] node204;
	wire [4-1:0] node208;
	wire [4-1:0] node210;
	wire [4-1:0] node212;
	wire [4-1:0] node216;
	wire [4-1:0] node218;
	wire [4-1:0] node219;
	wire [4-1:0] node220;
	wire [4-1:0] node222;
	wire [4-1:0] node226;
	wire [4-1:0] node228;
	wire [4-1:0] node229;
	wire [4-1:0] node233;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node237;
	wire [4-1:0] node238;
	wire [4-1:0] node239;
	wire [4-1:0] node241;
	wire [4-1:0] node242;
	wire [4-1:0] node246;
	wire [4-1:0] node248;
	wire [4-1:0] node249;
	wire [4-1:0] node250;
	wire [4-1:0] node257;
	wire [4-1:0] node258;
	wire [4-1:0] node260;
	wire [4-1:0] node261;
	wire [4-1:0] node262;
	wire [4-1:0] node263;
	wire [4-1:0] node265;
	wire [4-1:0] node266;
	wire [4-1:0] node270;
	wire [4-1:0] node271;
	wire [4-1:0] node277;
	wire [4-1:0] node278;
	wire [4-1:0] node279;
	wire [4-1:0] node281;
	wire [4-1:0] node282;
	wire [4-1:0] node283;
	wire [4-1:0] node284;
	wire [4-1:0] node291;
	wire [4-1:0] node292;
	wire [4-1:0] node294;
	wire [4-1:0] node296;
	wire [4-1:0] node297;
	wire [4-1:0] node299;
	wire [4-1:0] node303;
	wire [4-1:0] node304;
	wire [4-1:0] node305;
	wire [4-1:0] node307;
	wire [4-1:0] node311;
	wire [4-1:0] node312;
	wire [4-1:0] node314;
	wire [4-1:0] node315;
	wire [4-1:0] node320;
	wire [4-1:0] node322;
	wire [4-1:0] node323;
	wire [4-1:0] node324;
	wire [4-1:0] node325;
	wire [4-1:0] node326;
	wire [4-1:0] node327;
	wire [4-1:0] node329;
	wire [4-1:0] node330;
	wire [4-1:0] node334;
	wire [4-1:0] node336;
	wire [4-1:0] node337;
	wire [4-1:0] node342;
	wire [4-1:0] node344;
	wire [4-1:0] node345;
	wire [4-1:0] node346;
	wire [4-1:0] node348;
	wire [4-1:0] node352;
	wire [4-1:0] node354;
	wire [4-1:0] node356;
	wire [4-1:0] node360;
	wire [4-1:0] node362;
	wire [4-1:0] node363;
	wire [4-1:0] node364;
	wire [4-1:0] node365;
	wire [4-1:0] node366;
	wire [4-1:0] node367;
	wire [4-1:0] node372;
	wire [4-1:0] node374;
	wire [4-1:0] node376;
	wire [4-1:0] node380;
	wire [4-1:0] node382;
	wire [4-1:0] node383;
	wire [4-1:0] node385;
	wire [4-1:0] node386;
	wire [4-1:0] node390;
	wire [4-1:0] node392;
	wire [4-1:0] node394;
	wire [4-1:0] node397;
	wire [4-1:0] node398;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node403;
	wire [4-1:0] node404;
	wire [4-1:0] node405;
	wire [4-1:0] node406;
	wire [4-1:0] node407;
	wire [4-1:0] node408;
	wire [4-1:0] node409;
	wire [4-1:0] node414;
	wire [4-1:0] node416;
	wire [4-1:0] node417;
	wire [4-1:0] node422;
	wire [4-1:0] node424;
	wire [4-1:0] node425;
	wire [4-1:0] node426;
	wire [4-1:0] node428;
	wire [4-1:0] node432;
	wire [4-1:0] node434;
	wire [4-1:0] node435;
	wire [4-1:0] node440;
	wire [4-1:0] node442;
	wire [4-1:0] node443;
	wire [4-1:0] node444;
	wire [4-1:0] node445;
	wire [4-1:0] node447;
	wire [4-1:0] node448;
	wire [4-1:0] node452;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node460;
	wire [4-1:0] node462;
	wire [4-1:0] node463;
	wire [4-1:0] node464;
	wire [4-1:0] node466;
	wire [4-1:0] node470;
	wire [4-1:0] node472;
	wire [4-1:0] node473;
	wire [4-1:0] node478;
	wire [4-1:0] node480;
	wire [4-1:0] node481;
	wire [4-1:0] node482;
	wire [4-1:0] node483;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node486;
	wire [4-1:0] node488;
	wire [4-1:0] node492;
	wire [4-1:0] node494;
	wire [4-1:0] node496;
	wire [4-1:0] node500;
	wire [4-1:0] node502;
	wire [4-1:0] node503;
	wire [4-1:0] node504;
	wire [4-1:0] node506;
	wire [4-1:0] node510;
	wire [4-1:0] node511;
	wire [4-1:0] node513;
	wire [4-1:0] node518;
	wire [4-1:0] node520;
	wire [4-1:0] node521;
	wire [4-1:0] node522;
	wire [4-1:0] node523;
	wire [4-1:0] node524;
	wire [4-1:0] node526;
	wire [4-1:0] node530;
	wire [4-1:0] node532;
	wire [4-1:0] node534;
	wire [4-1:0] node538;
	wire [4-1:0] node540;
	wire [4-1:0] node541;
	wire [4-1:0] node543;
	wire [4-1:0] node544;
	wire [4-1:0] node548;
	wire [4-1:0] node550;
	wire [4-1:0] node553;
	wire [4-1:0] node554;
	wire [4-1:0] node555;
	wire [4-1:0] node556;
	wire [4-1:0] node557;
	wire [4-1:0] node558;
	wire [4-1:0] node559;
	wire [4-1:0] node560;
	wire [4-1:0] node562;
	wire [4-1:0] node566;
	wire [4-1:0] node568;
	wire [4-1:0] node569;
	wire [4-1:0] node573;
	wire [4-1:0] node575;
	wire [4-1:0] node576;
	wire [4-1:0] node577;
	wire [4-1:0] node578;
	wire [4-1:0] node580;
	wire [4-1:0] node586;
	wire [4-1:0] node588;
	wire [4-1:0] node589;
	wire [4-1:0] node590;
	wire [4-1:0] node592;
	wire [4-1:0] node596;
	wire [4-1:0] node598;
	wire [4-1:0] node600;
	wire [4-1:0] node603;
	wire [4-1:0] node604;
	wire [4-1:0] node605;
	wire [4-1:0] node606;
	wire [4-1:0] node607;
	wire [4-1:0] node608;
	wire [4-1:0] node609;
	wire [4-1:0] node611;
	wire [4-1:0] node615;
	wire [4-1:0] node617;
	wire [4-1:0] node621;
	wire [4-1:0] node622;
	wire [4-1:0] node624;
	wire [4-1:0] node625;
	wire [4-1:0] node626;
	wire [4-1:0] node632;
	wire [4-1:0] node633;
	wire [4-1:0] node634;
	wire [4-1:0] node636;
	wire [4-1:0] node638;
	wire [4-1:0] node640;
	wire [4-1:0] node645;
	wire [4-1:0] node647;
	wire [4-1:0] node648;
	wire [4-1:0] node649;
	wire [4-1:0] node651;
	wire [4-1:0] node652;
	wire [4-1:0] node656;
	wire [4-1:0] node657;
	wire [4-1:0] node659;
	wire [4-1:0] node660;
	wire [4-1:0] node666;
	wire [4-1:0] node667;
	wire [4-1:0] node668;
	wire [4-1:0] node669;
	wire [4-1:0] node670;
	wire [4-1:0] node671;
	wire [4-1:0] node674;
	wire [4-1:0] node675;
	wire [4-1:0] node676;
	wire [4-1:0] node681;
	wire [4-1:0] node682;
	wire [4-1:0] node684;
	wire [4-1:0] node685;
	wire [4-1:0] node689;
	wire [4-1:0] node691;
	wire [4-1:0] node693;
	wire [4-1:0] node696;
	wire [4-1:0] node697;
	wire [4-1:0] node698;
	wire [4-1:0] node699;
	wire [4-1:0] node702;
	wire [4-1:0] node703;
	wire [4-1:0] node705;
	wire [4-1:0] node709;
	wire [4-1:0] node710;
	wire [4-1:0] node711;
	wire [4-1:0] node712;
	wire [4-1:0] node715;
	wire [4-1:0] node718;
	wire [4-1:0] node719;
	wire [4-1:0] node722;
	wire [4-1:0] node725;
	wire [4-1:0] node726;
	wire [4-1:0] node727;
	wire [4-1:0] node730;
	wire [4-1:0] node733;
	wire [4-1:0] node734;
	wire [4-1:0] node735;
	wire [4-1:0] node738;
	wire [4-1:0] node741;
	wire [4-1:0] node742;
	wire [4-1:0] node745;
	wire [4-1:0] node748;
	wire [4-1:0] node749;
	wire [4-1:0] node751;
	wire [4-1:0] node754;
	wire [4-1:0] node757;
	wire [4-1:0] node758;
	wire [4-1:0] node759;
	wire [4-1:0] node760;
	wire [4-1:0] node762;
	wire [4-1:0] node764;
	wire [4-1:0] node767;
	wire [4-1:0] node769;
	wire [4-1:0] node770;
	wire [4-1:0] node771;
	wire [4-1:0] node776;
	wire [4-1:0] node777;
	wire [4-1:0] node779;
	wire [4-1:0] node782;
	wire [4-1:0] node783;
	wire [4-1:0] node784;
	wire [4-1:0] node789;
	wire [4-1:0] node790;
	wire [4-1:0] node791;
	wire [4-1:0] node792;
	wire [4-1:0] node795;
	wire [4-1:0] node796;
	wire [4-1:0] node800;
	wire [4-1:0] node801;
	wire [4-1:0] node805;
	wire [4-1:0] node806;
	wire [4-1:0] node807;
	wire [4-1:0] node808;
	wire [4-1:0] node809;
	wire [4-1:0] node815;
	wire [4-1:0] node816;
	wire [4-1:0] node818;
	wire [4-1:0] node820;
	wire [4-1:0] node823;
	wire [4-1:0] node826;
	wire [4-1:0] node827;
	wire [4-1:0] node828;
	wire [4-1:0] node829;
	wire [4-1:0] node830;
	wire [4-1:0] node831;
	wire [4-1:0] node832;
	wire [4-1:0] node836;
	wire [4-1:0] node838;
	wire [4-1:0] node840;
	wire [4-1:0] node843;
	wire [4-1:0] node844;
	wire [4-1:0] node846;
	wire [4-1:0] node849;
	wire [4-1:0] node852;
	wire [4-1:0] node853;
	wire [4-1:0] node855;
	wire [4-1:0] node856;
	wire [4-1:0] node858;
	wire [4-1:0] node862;
	wire [4-1:0] node864;
	wire [4-1:0] node865;
	wire [4-1:0] node869;
	wire [4-1:0] node870;
	wire [4-1:0] node871;
	wire [4-1:0] node873;
	wire [4-1:0] node874;
	wire [4-1:0] node879;
	wire [4-1:0] node880;
	wire [4-1:0] node881;
	wire [4-1:0] node883;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node890;
	wire [4-1:0] node891;
	wire [4-1:0] node893;
	wire [4-1:0] node894;
	wire [4-1:0] node896;
	wire [4-1:0] node900;
	wire [4-1:0] node902;
	wire [4-1:0] node903;
	wire [4-1:0] node907;
	wire [4-1:0] node908;
	wire [4-1:0] node910;
	wire [4-1:0] node912;
	wire [4-1:0] node915;
	wire [4-1:0] node916;
	wire [4-1:0] node918;
	wire [4-1:0] node920;
	wire [4-1:0] node924;
	wire [4-1:0] node925;
	wire [4-1:0] node926;
	wire [4-1:0] node928;
	wire [4-1:0] node931;
	wire [4-1:0] node933;
	wire [4-1:0] node934;
	wire [4-1:0] node938;
	wire [4-1:0] node941;
	wire [4-1:0] node942;
	wire [4-1:0] node943;
	wire [4-1:0] node944;
	wire [4-1:0] node945;
	wire [4-1:0] node946;
	wire [4-1:0] node948;
	wire [4-1:0] node949;
	wire [4-1:0] node950;
	wire [4-1:0] node955;
	wire [4-1:0] node957;
	wire [4-1:0] node958;
	wire [4-1:0] node959;
	wire [4-1:0] node960;
	wire [4-1:0] node966;
	wire [4-1:0] node967;
	wire [4-1:0] node968;
	wire [4-1:0] node970;
	wire [4-1:0] node972;
	wire [4-1:0] node975;
	wire [4-1:0] node976;
	wire [4-1:0] node977;
	wire [4-1:0] node982;
	wire [4-1:0] node983;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node987;
	wire [4-1:0] node993;
	wire [4-1:0] node994;
	wire [4-1:0] node995;
	wire [4-1:0] node996;
	wire [4-1:0] node997;
	wire [4-1:0] node999;
	wire [4-1:0] node1004;
	wire [4-1:0] node1005;
	wire [4-1:0] node1007;
	wire [4-1:0] node1009;
	wire [4-1:0] node1010;
	wire [4-1:0] node1014;
	wire [4-1:0] node1015;
	wire [4-1:0] node1019;
	wire [4-1:0] node1020;
	wire [4-1:0] node1021;
	wire [4-1:0] node1023;
	wire [4-1:0] node1027;
	wire [4-1:0] node1029;
	wire [4-1:0] node1030;
	wire [4-1:0] node1031;
	wire [4-1:0] node1036;
	wire [4-1:0] node1037;
	wire [4-1:0] node1038;
	wire [4-1:0] node1039;
	wire [4-1:0] node1040;
	wire [4-1:0] node1042;
	wire [4-1:0] node1046;
	wire [4-1:0] node1047;
	wire [4-1:0] node1049;
	wire [4-1:0] node1053;
	wire [4-1:0] node1055;
	wire [4-1:0] node1056;
	wire [4-1:0] node1057;
	wire [4-1:0] node1059;
	wire [4-1:0] node1061;
	wire [4-1:0] node1064;
	wire [4-1:0] node1065;
	wire [4-1:0] node1070;
	wire [4-1:0] node1071;
	wire [4-1:0] node1072;
	wire [4-1:0] node1073;
	wire [4-1:0] node1074;
	wire [4-1:0] node1075;
	wire [4-1:0] node1076;
	wire [4-1:0] node1081;
	wire [4-1:0] node1083;
	wire [4-1:0] node1087;
	wire [4-1:0] node1089;
	wire [4-1:0] node1090;
	wire [4-1:0] node1091;
	wire [4-1:0] node1093;
	wire [4-1:0] node1098;
	wire [4-1:0] node1099;
	wire [4-1:0] node1101;
	wire [4-1:0] node1102;
	wire [4-1:0] node1106;
	wire [4-1:0] node1108;
	wire [4-1:0] node1109;
	wire [4-1:0] node1113;
	wire [4-1:0] node1114;
	wire [4-1:0] node1115;
	wire [4-1:0] node1116;
	wire [4-1:0] node1117;
	wire [4-1:0] node1118;
	wire [4-1:0] node1119;
	wire [4-1:0] node1120;
	wire [4-1:0] node1124;
	wire [4-1:0] node1125;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1133;
	wire [4-1:0] node1134;
	wire [4-1:0] node1136;
	wire [4-1:0] node1138;
	wire [4-1:0] node1141;
	wire [4-1:0] node1143;
	wire [4-1:0] node1146;
	wire [4-1:0] node1147;
	wire [4-1:0] node1148;
	wire [4-1:0] node1149;
	wire [4-1:0] node1153;
	wire [4-1:0] node1155;
	wire [4-1:0] node1158;
	wire [4-1:0] node1159;
	wire [4-1:0] node1162;
	wire [4-1:0] node1163;
	wire [4-1:0] node1167;
	wire [4-1:0] node1168;
	wire [4-1:0] node1169;
	wire [4-1:0] node1170;
	wire [4-1:0] node1171;
	wire [4-1:0] node1173;
	wire [4-1:0] node1177;
	wire [4-1:0] node1178;
	wire [4-1:0] node1182;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1187;
	wire [4-1:0] node1190;
	wire [4-1:0] node1191;
	wire [4-1:0] node1192;
	wire [4-1:0] node1197;
	wire [4-1:0] node1198;
	wire [4-1:0] node1199;
	wire [4-1:0] node1201;
	wire [4-1:0] node1206;
	wire [4-1:0] node1207;
	wire [4-1:0] node1208;
	wire [4-1:0] node1209;
	wire [4-1:0] node1211;
	wire [4-1:0] node1212;
	wire [4-1:0] node1213;
	wire [4-1:0] node1218;
	wire [4-1:0] node1220;
	wire [4-1:0] node1223;
	wire [4-1:0] node1224;
	wire [4-1:0] node1225;
	wire [4-1:0] node1226;
	wire [4-1:0] node1228;
	wire [4-1:0] node1232;
	wire [4-1:0] node1233;
	wire [4-1:0] node1237;
	wire [4-1:0] node1238;
	wire [4-1:0] node1239;
	wire [4-1:0] node1243;
	wire [4-1:0] node1245;
	wire [4-1:0] node1248;
	wire [4-1:0] node1249;
	wire [4-1:0] node1250;
	wire [4-1:0] node1251;
	wire [4-1:0] node1252;
	wire [4-1:0] node1254;
	wire [4-1:0] node1258;
	wire [4-1:0] node1259;
	wire [4-1:0] node1263;
	wire [4-1:0] node1266;
	wire [4-1:0] node1267;
	wire [4-1:0] node1268;
	wire [4-1:0] node1270;
	wire [4-1:0] node1273;
	wire [4-1:0] node1274;
	wire [4-1:0] node1276;
	wire [4-1:0] node1279;
	wire [4-1:0] node1280;
	wire [4-1:0] node1284;
	wire [4-1:0] node1287;
	wire [4-1:0] node1288;
	wire [4-1:0] node1289;
	wire [4-1:0] node1290;
	wire [4-1:0] node1291;
	wire [4-1:0] node1292;
	wire [4-1:0] node1293;
	wire [4-1:0] node1294;
	wire [4-1:0] node1297;
	wire [4-1:0] node1300;
	wire [4-1:0] node1302;
	wire [4-1:0] node1305;
	wire [4-1:0] node1306;
	wire [4-1:0] node1308;
	wire [4-1:0] node1311;
	wire [4-1:0] node1312;
	wire [4-1:0] node1315;
	wire [4-1:0] node1318;
	wire [4-1:0] node1319;
	wire [4-1:0] node1320;
	wire [4-1:0] node1322;
	wire [4-1:0] node1325;
	wire [4-1:0] node1327;
	wire [4-1:0] node1330;
	wire [4-1:0] node1331;
	wire [4-1:0] node1332;
	wire [4-1:0] node1333;
	wire [4-1:0] node1336;
	wire [4-1:0] node1339;
	wire [4-1:0] node1340;
	wire [4-1:0] node1343;
	wire [4-1:0] node1346;
	wire [4-1:0] node1347;
	wire [4-1:0] node1351;
	wire [4-1:0] node1352;
	wire [4-1:0] node1353;
	wire [4-1:0] node1354;
	wire [4-1:0] node1357;
	wire [4-1:0] node1359;
	wire [4-1:0] node1362;
	wire [4-1:0] node1363;
	wire [4-1:0] node1366;
	wire [4-1:0] node1367;
	wire [4-1:0] node1371;
	wire [4-1:0] node1372;
	wire [4-1:0] node1373;
	wire [4-1:0] node1374;
	wire [4-1:0] node1378;
	wire [4-1:0] node1380;
	wire [4-1:0] node1383;
	wire [4-1:0] node1384;
	wire [4-1:0] node1386;
	wire [4-1:0] node1389;
	wire [4-1:0] node1392;
	wire [4-1:0] node1393;
	wire [4-1:0] node1394;
	wire [4-1:0] node1397;
	wire [4-1:0] node1400;
	wire [4-1:0] node1401;
	wire [4-1:0] node1404;
	wire [4-1:0] node1407;
	wire [4-1:0] node1408;
	wire [4-1:0] node1409;
	wire [4-1:0] node1410;
	wire [4-1:0] node1413;
	wire [4-1:0] node1416;
	wire [4-1:0] node1417;
	wire [4-1:0] node1420;
	wire [4-1:0] node1424;
	wire [4-1:0] node1426;
	wire [4-1:0] node1427;
	wire [4-1:0] node1428;
	wire [4-1:0] node1429;
	wire [4-1:0] node1430;
	wire [4-1:0] node1431;
	wire [4-1:0] node1432;
	wire [4-1:0] node1433;
	wire [4-1:0] node1434;
	wire [4-1:0] node1435;
	wire [4-1:0] node1436;
	wire [4-1:0] node1437;
	wire [4-1:0] node1442;
	wire [4-1:0] node1444;
	wire [4-1:0] node1448;
	wire [4-1:0] node1450;
	wire [4-1:0] node1451;
	wire [4-1:0] node1453;
	wire [4-1:0] node1454;
	wire [4-1:0] node1458;
	wire [4-1:0] node1460;
	wire [4-1:0] node1462;
	wire [4-1:0] node1466;
	wire [4-1:0] node1468;
	wire [4-1:0] node1469;
	wire [4-1:0] node1470;
	wire [4-1:0] node1471;
	wire [4-1:0] node1472;
	wire [4-1:0] node1474;
	wire [4-1:0] node1478;
	wire [4-1:0] node1480;
	wire [4-1:0] node1481;
	wire [4-1:0] node1486;
	wire [4-1:0] node1488;
	wire [4-1:0] node1489;
	wire [4-1:0] node1491;
	wire [4-1:0] node1492;
	wire [4-1:0] node1496;
	wire [4-1:0] node1498;
	wire [4-1:0] node1499;
	wire [4-1:0] node1504;
	wire [4-1:0] node1505;
	wire [4-1:0] node1506;
	wire [4-1:0] node1507;
	wire [4-1:0] node1508;
	wire [4-1:0] node1509;
	wire [4-1:0] node1510;
	wire [4-1:0] node1512;
	wire [4-1:0] node1516;
	wire [4-1:0] node1517;
	wire [4-1:0] node1519;
	wire [4-1:0] node1524;
	wire [4-1:0] node1525;
	wire [4-1:0] node1526;
	wire [4-1:0] node1528;
	wire [4-1:0] node1529;
	wire [4-1:0] node1530;
	wire [4-1:0] node1537;
	wire [4-1:0] node1538;
	wire [4-1:0] node1540;
	wire [4-1:0] node1541;
	wire [4-1:0] node1542;
	wire [4-1:0] node1543;
	wire [4-1:0] node1548;
	wire [4-1:0] node1550;
	wire [4-1:0] node1552;
	wire [4-1:0] node1555;
	wire [4-1:0] node1556;
	wire [4-1:0] node1558;
	wire [4-1:0] node1560;
	wire [4-1:0] node1561;
	wire [4-1:0] node1562;
	wire [4-1:0] node1567;
	wire [4-1:0] node1568;
	wire [4-1:0] node1570;
	wire [4-1:0] node1571;
	wire [4-1:0] node1575;
	wire [4-1:0] node1577;
	wire [4-1:0] node1578;
	wire [4-1:0] node1579;
	wire [4-1:0] node1584;
	wire [4-1:0] node1586;
	wire [4-1:0] node1587;
	wire [4-1:0] node1588;
	wire [4-1:0] node1589;
	wire [4-1:0] node1590;
	wire [4-1:0] node1592;
	wire [4-1:0] node1596;
	wire [4-1:0] node1598;
	wire [4-1:0] node1600;
	wire [4-1:0] node1604;
	wire [4-1:0] node1606;
	wire [4-1:0] node1607;
	wire [4-1:0] node1608;
	wire [4-1:0] node1610;
	wire [4-1:0] node1614;
	wire [4-1:0] node1616;
	wire [4-1:0] node1617;
	wire [4-1:0] node1621;
	wire [4-1:0] node1622;
	wire [4-1:0] node1624;
	wire [4-1:0] node1625;
	wire [4-1:0] node1626;
	wire [4-1:0] node1627;
	wire [4-1:0] node1628;
	wire [4-1:0] node1629;
	wire [4-1:0] node1630;
	wire [4-1:0] node1632;
	wire [4-1:0] node1636;
	wire [4-1:0] node1638;
	wire [4-1:0] node1640;
	wire [4-1:0] node1644;
	wire [4-1:0] node1646;
	wire [4-1:0] node1647;
	wire [4-1:0] node1648;
	wire [4-1:0] node1649;
	wire [4-1:0] node1654;
	wire [4-1:0] node1656;
	wire [4-1:0] node1657;
	wire [4-1:0] node1662;
	wire [4-1:0] node1664;
	wire [4-1:0] node1665;
	wire [4-1:0] node1666;
	wire [4-1:0] node1667;
	wire [4-1:0] node1668;
	wire [4-1:0] node1669;
	wire [4-1:0] node1674;
	wire [4-1:0] node1676;
	wire [4-1:0] node1677;
	wire [4-1:0] node1682;
	wire [4-1:0] node1684;
	wire [4-1:0] node1685;
	wire [4-1:0] node1686;
	wire [4-1:0] node1687;
	wire [4-1:0] node1692;
	wire [4-1:0] node1694;
	wire [4-1:0] node1695;
	wire [4-1:0] node1699;
	wire [4-1:0] node1700;
	wire [4-1:0] node1701;
	wire [4-1:0] node1702;
	wire [4-1:0] node1703;
	wire [4-1:0] node1704;
	wire [4-1:0] node1705;
	wire [4-1:0] node1709;
	wire [4-1:0] node1710;
	wire [4-1:0] node1711;
	wire [4-1:0] node1712;
	wire [4-1:0] node1717;
	wire [4-1:0] node1720;
	wire [4-1:0] node1722;
	wire [4-1:0] node1723;
	wire [4-1:0] node1725;
	wire [4-1:0] node1727;
	wire [4-1:0] node1730;
	wire [4-1:0] node1731;
	wire [4-1:0] node1735;
	wire [4-1:0] node1736;
	wire [4-1:0] node1737;
	wire [4-1:0] node1739;
	wire [4-1:0] node1741;
	wire [4-1:0] node1742;
	wire [4-1:0] node1746;
	wire [4-1:0] node1747;
	wire [4-1:0] node1750;
	wire [4-1:0] node1752;
	wire [4-1:0] node1755;
	wire [4-1:0] node1756;
	wire [4-1:0] node1758;
	wire [4-1:0] node1762;
	wire [4-1:0] node1763;
	wire [4-1:0] node1764;
	wire [4-1:0] node1765;
	wire [4-1:0] node1766;
	wire [4-1:0] node1767;
	wire [4-1:0] node1769;
	wire [4-1:0] node1773;
	wire [4-1:0] node1775;
	wire [4-1:0] node1779;
	wire [4-1:0] node1781;
	wire [4-1:0] node1782;
	wire [4-1:0] node1783;
	wire [4-1:0] node1784;
	wire [4-1:0] node1790;
	wire [4-1:0] node1791;
	wire [4-1:0] node1792;
	wire [4-1:0] node1793;
	wire [4-1:0] node1795;
	wire [4-1:0] node1798;
	wire [4-1:0] node1800;
	wire [4-1:0] node1801;
	wire [4-1:0] node1805;
	wire [4-1:0] node1806;
	wire [4-1:0] node1809;
	wire [4-1:0] node1811;
	wire [4-1:0] node1814;
	wire [4-1:0] node1815;
	wire [4-1:0] node1816;
	wire [4-1:0] node1820;
	wire [4-1:0] node1821;
	wire [4-1:0] node1823;
	wire [4-1:0] node1824;
	wire [4-1:0] node1829;
	wire [4-1:0] node1830;
	wire [4-1:0] node1831;
	wire [4-1:0] node1832;
	wire [4-1:0] node1833;
	wire [4-1:0] node1834;
	wire [4-1:0] node1838;
	wire [4-1:0] node1839;
	wire [4-1:0] node1840;
	wire [4-1:0] node1841;
	wire [4-1:0] node1847;
	wire [4-1:0] node1848;
	wire [4-1:0] node1849;
	wire [4-1:0] node1850;
	wire [4-1:0] node1851;
	wire [4-1:0] node1856;
	wire [4-1:0] node1857;
	wire [4-1:0] node1861;
	wire [4-1:0] node1862;
	wire [4-1:0] node1865;
	wire [4-1:0] node1866;
	wire [4-1:0] node1870;
	wire [4-1:0] node1871;
	wire [4-1:0] node1872;
	wire [4-1:0] node1874;
	wire [4-1:0] node1877;
	wire [4-1:0] node1878;
	wire [4-1:0] node1880;
	wire [4-1:0] node1882;
	wire [4-1:0] node1886;
	wire [4-1:0] node1887;
	wire [4-1:0] node1888;
	wire [4-1:0] node1889;
	wire [4-1:0] node1891;
	wire [4-1:0] node1896;
	wire [4-1:0] node1897;
	wire [4-1:0] node1901;
	wire [4-1:0] node1902;
	wire [4-1:0] node1903;
	wire [4-1:0] node1904;
	wire [4-1:0] node1905;
	wire [4-1:0] node1906;
	wire [4-1:0] node1907;
	wire [4-1:0] node1911;
	wire [4-1:0] node1913;
	wire [4-1:0] node1916;
	wire [4-1:0] node1917;
	wire [4-1:0] node1920;
	wire [4-1:0] node1921;
	wire [4-1:0] node1925;
	wire [4-1:0] node1928;
	wire [4-1:0] node1929;
	wire [4-1:0] node1930;
	wire [4-1:0] node1931;
	wire [4-1:0] node1932;
	wire [4-1:0] node1933;
	wire [4-1:0] node1937;
	wire [4-1:0] node1939;
	wire [4-1:0] node1942;
	wire [4-1:0] node1943;
	wire [4-1:0] node1947;
	wire [4-1:0] node1948;
	wire [4-1:0] node1949;
	wire [4-1:0] node1953;
	wire [4-1:0] node1955;
	wire [4-1:0] node1958;
	wire [4-1:0] node1961;
	wire [4-1:0] node1962;
	wire [4-1:0] node1963;
	wire [4-1:0] node1964;
	wire [4-1:0] node1967;
	wire [4-1:0] node1970;
	wire [4-1:0] node1971;
	wire [4-1:0] node1974;
	wire [4-1:0] node1978;
	wire [4-1:0] node1980;
	wire [4-1:0] node1981;
	wire [4-1:0] node1982;
	wire [4-1:0] node1983;
	wire [4-1:0] node1984;
	wire [4-1:0] node1985;
	wire [4-1:0] node1986;
	wire [4-1:0] node1987;
	wire [4-1:0] node1988;
	wire [4-1:0] node1989;
	wire [4-1:0] node1994;
	wire [4-1:0] node1995;
	wire [4-1:0] node1997;
	wire [4-1:0] node2002;
	wire [4-1:0] node2004;
	wire [4-1:0] node2005;
	wire [4-1:0] node2006;
	wire [4-1:0] node2007;
	wire [4-1:0] node2012;
	wire [4-1:0] node2013;
	wire [4-1:0] node2015;
	wire [4-1:0] node2020;
	wire [4-1:0] node2021;
	wire [4-1:0] node2022;
	wire [4-1:0] node2023;
	wire [4-1:0] node2024;
	wire [4-1:0] node2025;
	wire [4-1:0] node2030;
	wire [4-1:0] node2031;
	wire [4-1:0] node2032;
	wire [4-1:0] node2037;
	wire [4-1:0] node2038;
	wire [4-1:0] node2040;
	wire [4-1:0] node2041;
	wire [4-1:0] node2045;
	wire [4-1:0] node2047;
	wire [4-1:0] node2048;
	wire [4-1:0] node2049;
	wire [4-1:0] node2054;
	wire [4-1:0] node2056;
	wire [4-1:0] node2057;
	wire [4-1:0] node2058;
	wire [4-1:0] node2060;
	wire [4-1:0] node2064;
	wire [4-1:0] node2066;
	wire [4-1:0] node2068;
	wire [4-1:0] node2071;
	wire [4-1:0] node2072;
	wire [4-1:0] node2074;
	wire [4-1:0] node2075;
	wire [4-1:0] node2076;
	wire [4-1:0] node2077;
	wire [4-1:0] node2078;
	wire [4-1:0] node2079;
	wire [4-1:0] node2084;
	wire [4-1:0] node2086;
	wire [4-1:0] node2088;
	wire [4-1:0] node2092;
	wire [4-1:0] node2094;
	wire [4-1:0] node2095;
	wire [4-1:0] node2097;
	wire [4-1:0] node2098;
	wire [4-1:0] node2102;
	wire [4-1:0] node2104;
	wire [4-1:0] node2105;
	wire [4-1:0] node2109;
	wire [4-1:0] node2110;
	wire [4-1:0] node2111;
	wire [4-1:0] node2112;
	wire [4-1:0] node2113;
	wire [4-1:0] node2114;
	wire [4-1:0] node2118;
	wire [4-1:0] node2121;
	wire [4-1:0] node2122;
	wire [4-1:0] node2123;
	wire [4-1:0] node2127;
	wire [4-1:0] node2128;
	wire [4-1:0] node2130;
	wire [4-1:0] node2134;
	wire [4-1:0] node2135;
	wire [4-1:0] node2136;
	wire [4-1:0] node2138;
	wire [4-1:0] node2139;
	wire [4-1:0] node2143;
	wire [4-1:0] node2144;
	wire [4-1:0] node2148;
	wire [4-1:0] node2149;
	wire [4-1:0] node2152;
	wire [4-1:0] node2155;
	wire [4-1:0] node2156;
	wire [4-1:0] node2157;
	wire [4-1:0] node2158;
	wire [4-1:0] node2159;
	wire [4-1:0] node2162;
	wire [4-1:0] node2163;
	wire [4-1:0] node2167;
	wire [4-1:0] node2168;
	wire [4-1:0] node2169;
	wire [4-1:0] node2173;
	wire [4-1:0] node2174;
	wire [4-1:0] node2176;
	wire [4-1:0] node2180;
	wire [4-1:0] node2181;
	wire [4-1:0] node2184;
	wire [4-1:0] node2187;
	wire [4-1:0] node2188;
	wire [4-1:0] node2189;
	wire [4-1:0] node2192;
	wire [4-1:0] node2196;
	wire [4-1:0] node2198;
	wire [4-1:0] node2199;
	wire [4-1:0] node2200;
	wire [4-1:0] node2201;
	wire [4-1:0] node2202;
	wire [4-1:0] node2203;
	wire [4-1:0] node2204;
	wire [4-1:0] node2205;
	wire [4-1:0] node2210;
	wire [4-1:0] node2211;
	wire [4-1:0] node2215;
	wire [4-1:0] node2216;
	wire [4-1:0] node2217;
	wire [4-1:0] node2219;
	wire [4-1:0] node2222;
	wire [4-1:0] node2223;
	wire [4-1:0] node2228;
	wire [4-1:0] node2230;
	wire [4-1:0] node2232;
	wire [4-1:0] node2234;
	wire [4-1:0] node2237;
	wire [4-1:0] node2238;
	wire [4-1:0] node2240;
	wire [4-1:0] node2241;
	wire [4-1:0] node2242;
	wire [4-1:0] node2243;
	wire [4-1:0] node2248;
	wire [4-1:0] node2250;
	wire [4-1:0] node2252;
	wire [4-1:0] node2255;
	wire [4-1:0] node2256;
	wire [4-1:0] node2257;
	wire [4-1:0] node2258;
	wire [4-1:0] node2259;
	wire [4-1:0] node2264;
	wire [4-1:0] node2265;
	wire [4-1:0] node2267;
	wire [4-1:0] node2271;
	wire [4-1:0] node2272;
	wire [4-1:0] node2273;
	wire [4-1:0] node2276;
	wire [4-1:0] node2280;
	wire [4-1:0] node2282;
	wire [4-1:0] node2283;
	wire [4-1:0] node2284;
	wire [4-1:0] node2285;
	wire [4-1:0] node2286;
	wire [4-1:0] node2288;
	wire [4-1:0] node2292;
	wire [4-1:0] node2294;
	wire [4-1:0] node2296;
	wire [4-1:0] node2299;
	wire [4-1:0] node2300;
	wire [4-1:0] node2301;
	wire [4-1:0] node2304;
	wire [4-1:0] node2307;
	wire [4-1:0] node2308;
	wire [4-1:0] node2312;
	wire [4-1:0] node2314;
	wire [4-1:0] node2315;
	wire [4-1:0] node2316;
	wire [4-1:0] node2318;
	wire [4-1:0] node2321;
	wire [4-1:0] node2323;
	wire [4-1:0] node2326;
	wire [4-1:0] node2328;
	wire [4-1:0] node2329;

	assign outp = (inp[14]) ? node2 : 4'b0000;
		assign node2 = (inp[12]) ? node1424 : node3;
			assign node3 = (inp[3]) ? node397 : node4;
				assign node4 = (inp[0]) ? node156 : node5;
					assign node5 = (inp[4]) ? 4'b0000 : node6;
						assign node6 = (inp[11]) ? node84 : node7;
							assign node7 = (inp[7]) ? 4'b0010 : node8;
								assign node8 = (inp[5]) ? node46 : node9;
									assign node9 = (inp[9]) ? 4'b0010 : node10;
										assign node10 = (inp[13]) ? node28 : node11;
											assign node11 = (inp[15]) ? 4'b0000 : node12;
												assign node12 = (inp[8]) ? node22 : node13;
													assign node13 = (inp[2]) ? node15 : 4'b0010;
														assign node15 = (inp[10]) ? node17 : 4'b0010;
															assign node17 = (inp[6]) ? 4'b0010 : node18;
																assign node18 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node22 = (inp[1]) ? node24 : 4'b0000;
														assign node24 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node28 = (inp[15]) ? node30 : 4'b0010;
												assign node30 = (inp[8]) ? node38 : node31;
													assign node31 = (inp[10]) ? node33 : 4'b0010;
														assign node33 = (inp[1]) ? 4'b0010 : node34;
															assign node34 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node38 = (inp[1]) ? node40 : 4'b0000;
														assign node40 = (inp[10]) ? node42 : 4'b0010;
															assign node42 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node46 = (inp[9]) ? node48 : 4'b0000;
										assign node48 = (inp[13]) ? node66 : node49;
											assign node49 = (inp[15]) ? 4'b0000 : node50;
												assign node50 = (inp[1]) ? node58 : node51;
													assign node51 = (inp[8]) ? 4'b0000 : node52;
														assign node52 = (inp[10]) ? node54 : 4'b0010;
															assign node54 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node58 = (inp[8]) ? node60 : 4'b0010;
														assign node60 = (inp[10]) ? node62 : 4'b0010;
															assign node62 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node66 = (inp[15]) ? node68 : 4'b0010;
												assign node68 = (inp[8]) ? node76 : node69;
													assign node69 = (inp[10]) ? node71 : 4'b0010;
														assign node71 = (inp[1]) ? 4'b0010 : node72;
															assign node72 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node76 = (inp[1]) ? node78 : 4'b0000;
														assign node78 = (inp[6]) ? 4'b0010 : node79;
															assign node79 = (inp[10]) ? 4'b0000 : 4'b0010;
							assign node84 = (inp[7]) ? node86 : 4'b0000;
								assign node86 = (inp[9]) ? node124 : node87;
									assign node87 = (inp[5]) ? 4'b0000 : node88;
										assign node88 = (inp[13]) ? node106 : node89;
											assign node89 = (inp[15]) ? 4'b0000 : node90;
												assign node90 = (inp[8]) ? node98 : node91;
													assign node91 = (inp[6]) ? 4'b0010 : node92;
														assign node92 = (inp[10]) ? node94 : 4'b0010;
															assign node94 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node98 = (inp[1]) ? node100 : 4'b0000;
														assign node100 = (inp[6]) ? 4'b0010 : node101;
															assign node101 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node106 = (inp[15]) ? node108 : 4'b0010;
												assign node108 = (inp[8]) ? node116 : node109;
													assign node109 = (inp[1]) ? 4'b0010 : node110;
														assign node110 = (inp[10]) ? node112 : 4'b0010;
															assign node112 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node116 = (inp[1]) ? node118 : 4'b0000;
														assign node118 = (inp[6]) ? 4'b0010 : node119;
															assign node119 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node124 = (inp[5]) ? node126 : 4'b0010;
										assign node126 = (inp[15]) ? node138 : node127;
											assign node127 = (inp[13]) ? 4'b0010 : node128;
												assign node128 = (inp[8]) ? node130 : 4'b0010;
													assign node130 = (inp[1]) ? node132 : 4'b0000;
														assign node132 = (inp[10]) ? node134 : 4'b0010;
															assign node134 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node138 = (inp[13]) ? node140 : 4'b0000;
												assign node140 = (inp[1]) ? node148 : node141;
													assign node141 = (inp[8]) ? 4'b0000 : node142;
														assign node142 = (inp[10]) ? node144 : 4'b0010;
															assign node144 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node148 = (inp[8]) ? node150 : 4'b0010;
														assign node150 = (inp[10]) ? node152 : 4'b0010;
															assign node152 = (inp[2]) ? 4'b0000 : 4'b0010;
					assign node156 = (inp[4]) ? node320 : node157;
						assign node157 = (inp[7]) ? node233 : node158;
							assign node158 = (inp[9]) ? node196 : node159;
								assign node159 = (inp[11]) ? 4'b0010 : node160;
									assign node160 = (inp[13]) ? node178 : node161;
										assign node161 = (inp[5]) ? 4'b0010 : node162;
											assign node162 = (inp[1]) ? node170 : node163;
												assign node163 = (inp[15]) ? 4'b0010 : node164;
													assign node164 = (inp[6]) ? 4'b0000 : node165;
														assign node165 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node170 = (inp[15]) ? node172 : 4'b0000;
													assign node172 = (inp[8]) ? node174 : 4'b0000;
														assign node174 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node178 = (inp[5]) ? node180 : 4'b0000;
											assign node180 = (inp[1]) ? node188 : node181;
												assign node181 = (inp[15]) ? 4'b0010 : node182;
													assign node182 = (inp[6]) ? 4'b0000 : node183;
														assign node183 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node188 = (inp[8]) ? node190 : 4'b0000;
													assign node190 = (inp[15]) ? node192 : 4'b0000;
														assign node192 = (inp[6]) ? 4'b0000 : 4'b0010;
								assign node196 = (inp[11]) ? node198 : 4'b0000;
									assign node198 = (inp[5]) ? node216 : node199;
										assign node199 = (inp[13]) ? 4'b0000 : node200;
											assign node200 = (inp[15]) ? node208 : node201;
												assign node201 = (inp[8]) ? node203 : 4'b0000;
													assign node203 = (inp[1]) ? 4'b0000 : node204;
														assign node204 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node208 = (inp[1]) ? node210 : 4'b0010;
													assign node210 = (inp[8]) ? node212 : 4'b0000;
														assign node212 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node216 = (inp[13]) ? node218 : 4'b0010;
											assign node218 = (inp[1]) ? node226 : node219;
												assign node219 = (inp[15]) ? 4'b0010 : node220;
													assign node220 = (inp[8]) ? node222 : 4'b0000;
														assign node222 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node226 = (inp[8]) ? node228 : 4'b0000;
													assign node228 = (inp[6]) ? 4'b0000 : node229;
														assign node229 = (inp[15]) ? 4'b0010 : 4'b0000;
							assign node233 = (inp[9]) ? node257 : node234;
								assign node234 = (inp[5]) ? 4'b0000 : node235;
									assign node235 = (inp[13]) ? node237 : 4'b0000;
										assign node237 = (inp[11]) ? 4'b0000 : node238;
											assign node238 = (inp[1]) ? node246 : node239;
												assign node239 = (inp[6]) ? node241 : 4'b0000;
													assign node241 = (inp[15]) ? 4'b0000 : node242;
														assign node242 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node246 = (inp[15]) ? node248 : 4'b0010;
													assign node248 = (inp[6]) ? 4'b0010 : node249;
														assign node249 = (inp[10]) ? 4'b0000 : node250;
															assign node250 = (inp[8]) ? 4'b0000 : 4'b0010;
								assign node257 = (inp[11]) ? node277 : node258;
									assign node258 = (inp[5]) ? node260 : 4'b0010;
										assign node260 = (inp[13]) ? 4'b0010 : node261;
											assign node261 = (inp[1]) ? 4'b0010 : node262;
												assign node262 = (inp[15]) ? node270 : node263;
													assign node263 = (inp[10]) ? node265 : 4'b0010;
														assign node265 = (inp[6]) ? 4'b0010 : node266;
															assign node266 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node270 = (inp[8]) ? 4'b0000 : node271;
														assign node271 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node277 = (inp[13]) ? node291 : node278;
										assign node278 = (inp[5]) ? 4'b0000 : node279;
											assign node279 = (inp[1]) ? node281 : 4'b0000;
												assign node281 = (inp[15]) ? 4'b0000 : node282;
													assign node282 = (inp[6]) ? 4'b0010 : node283;
														assign node283 = (inp[10]) ? 4'b0000 : node284;
															assign node284 = (inp[8]) ? 4'b0000 : 4'b0010;
										assign node291 = (inp[5]) ? node303 : node292;
											assign node292 = (inp[15]) ? node294 : 4'b0010;
												assign node294 = (inp[8]) ? node296 : 4'b0010;
													assign node296 = (inp[6]) ? 4'b0010 : node297;
														assign node297 = (inp[10]) ? node299 : 4'b0010;
															assign node299 = (inp[1]) ? 4'b0010 : 4'b0000;
											assign node303 = (inp[1]) ? node311 : node304;
												assign node304 = (inp[15]) ? 4'b0000 : node305;
													assign node305 = (inp[6]) ? node307 : 4'b0000;
														assign node307 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node311 = (inp[6]) ? 4'b0010 : node312;
													assign node312 = (inp[15]) ? node314 : 4'b0010;
														assign node314 = (inp[8]) ? 4'b0000 : node315;
															assign node315 = (inp[10]) ? 4'b0000 : 4'b0010;
						assign node320 = (inp[7]) ? node322 : 4'b0010;
							assign node322 = (inp[11]) ? node360 : node323;
								assign node323 = (inp[9]) ? 4'b0000 : node324;
									assign node324 = (inp[5]) ? node342 : node325;
										assign node325 = (inp[13]) ? 4'b0000 : node326;
											assign node326 = (inp[15]) ? node334 : node327;
												assign node327 = (inp[8]) ? node329 : 4'b0000;
													assign node329 = (inp[1]) ? 4'b0000 : node330;
														assign node330 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node334 = (inp[1]) ? node336 : 4'b0010;
													assign node336 = (inp[6]) ? 4'b0000 : node337;
														assign node337 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node342 = (inp[13]) ? node344 : 4'b0010;
											assign node344 = (inp[15]) ? node352 : node345;
												assign node345 = (inp[6]) ? 4'b0000 : node346;
													assign node346 = (inp[8]) ? node348 : 4'b0000;
														assign node348 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node352 = (inp[1]) ? node354 : 4'b0010;
													assign node354 = (inp[8]) ? node356 : 4'b0000;
														assign node356 = (inp[6]) ? 4'b0000 : 4'b0010;
								assign node360 = (inp[9]) ? node362 : 4'b0010;
									assign node362 = (inp[13]) ? node380 : node363;
										assign node363 = (inp[5]) ? 4'b0010 : node364;
											assign node364 = (inp[15]) ? node372 : node365;
												assign node365 = (inp[6]) ? 4'b0000 : node366;
													assign node366 = (inp[1]) ? 4'b0000 : node367;
														assign node367 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node372 = (inp[1]) ? node374 : 4'b0010;
													assign node374 = (inp[8]) ? node376 : 4'b0000;
														assign node376 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node380 = (inp[5]) ? node382 : 4'b0000;
											assign node382 = (inp[15]) ? node390 : node383;
												assign node383 = (inp[8]) ? node385 : 4'b0000;
													assign node385 = (inp[6]) ? 4'b0000 : node386;
														assign node386 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node390 = (inp[1]) ? node392 : 4'b0010;
													assign node392 = (inp[8]) ? node394 : 4'b0000;
														assign node394 = (inp[6]) ? 4'b0000 : 4'b0010;
				assign node397 = (inp[0]) ? node553 : node398;
					assign node398 = (inp[4]) ? node400 : 4'b0010;
						assign node400 = (inp[7]) ? node478 : node401;
							assign node401 = (inp[11]) ? 4'b0000 : node402;
								assign node402 = (inp[9]) ? node440 : node403;
									assign node403 = (inp[5]) ? 4'b0000 : node404;
										assign node404 = (inp[15]) ? node422 : node405;
											assign node405 = (inp[13]) ? 4'b0010 : node406;
												assign node406 = (inp[8]) ? node414 : node407;
													assign node407 = (inp[6]) ? 4'b0010 : node408;
														assign node408 = (inp[1]) ? 4'b0010 : node409;
															assign node409 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node414 = (inp[1]) ? node416 : 4'b0000;
														assign node416 = (inp[6]) ? 4'b0010 : node417;
															assign node417 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node422 = (inp[13]) ? node424 : 4'b0000;
												assign node424 = (inp[1]) ? node432 : node425;
													assign node425 = (inp[8]) ? 4'b0000 : node426;
														assign node426 = (inp[10]) ? node428 : 4'b0010;
															assign node428 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node432 = (inp[10]) ? node434 : 4'b0010;
														assign node434 = (inp[6]) ? 4'b0010 : node435;
															assign node435 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node440 = (inp[5]) ? node442 : 4'b0010;
										assign node442 = (inp[15]) ? node460 : node443;
											assign node443 = (inp[13]) ? 4'b0010 : node444;
												assign node444 = (inp[8]) ? node452 : node445;
													assign node445 = (inp[10]) ? node447 : 4'b0010;
														assign node447 = (inp[1]) ? 4'b0010 : node448;
															assign node448 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node452 = (inp[1]) ? node454 : 4'b0000;
														assign node454 = (inp[6]) ? 4'b0010 : node455;
															assign node455 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node460 = (inp[13]) ? node462 : 4'b0000;
												assign node462 = (inp[8]) ? node470 : node463;
													assign node463 = (inp[1]) ? 4'b0010 : node464;
														assign node464 = (inp[10]) ? node466 : 4'b0010;
															assign node466 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node470 = (inp[1]) ? node472 : 4'b0000;
														assign node472 = (inp[6]) ? 4'b0010 : node473;
															assign node473 = (inp[10]) ? 4'b0000 : 4'b0010;
							assign node478 = (inp[11]) ? node480 : 4'b0010;
								assign node480 = (inp[9]) ? node518 : node481;
									assign node481 = (inp[5]) ? 4'b0000 : node482;
										assign node482 = (inp[15]) ? node500 : node483;
											assign node483 = (inp[13]) ? 4'b0010 : node484;
												assign node484 = (inp[1]) ? node492 : node485;
													assign node485 = (inp[8]) ? 4'b0000 : node486;
														assign node486 = (inp[10]) ? node488 : 4'b0010;
															assign node488 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node492 = (inp[10]) ? node494 : 4'b0010;
														assign node494 = (inp[8]) ? node496 : 4'b0010;
															assign node496 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node500 = (inp[13]) ? node502 : 4'b0000;
												assign node502 = (inp[1]) ? node510 : node503;
													assign node503 = (inp[8]) ? 4'b0000 : node504;
														assign node504 = (inp[10]) ? node506 : 4'b0010;
															assign node506 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node510 = (inp[6]) ? 4'b0010 : node511;
														assign node511 = (inp[8]) ? node513 : 4'b0010;
															assign node513 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node518 = (inp[5]) ? node520 : 4'b0010;
										assign node520 = (inp[15]) ? node538 : node521;
											assign node521 = (inp[13]) ? 4'b0010 : node522;
												assign node522 = (inp[8]) ? node530 : node523;
													assign node523 = (inp[6]) ? 4'b0010 : node524;
														assign node524 = (inp[10]) ? node526 : 4'b0010;
															assign node526 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node530 = (inp[1]) ? node532 : 4'b0000;
														assign node532 = (inp[10]) ? node534 : 4'b0010;
															assign node534 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node538 = (inp[13]) ? node540 : 4'b0000;
												assign node540 = (inp[8]) ? node548 : node541;
													assign node541 = (inp[10]) ? node543 : 4'b0010;
														assign node543 = (inp[6]) ? 4'b0010 : node544;
															assign node544 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node548 = (inp[1]) ? node550 : 4'b0000;
														assign node550 = (inp[6]) ? 4'b0010 : 4'b0000;
					assign node553 = (inp[9]) ? node941 : node554;
						assign node554 = (inp[7]) ? node666 : node555;
							assign node555 = (inp[4]) ? node603 : node556;
								assign node556 = (inp[11]) ? node586 : node557;
									assign node557 = (inp[13]) ? node573 : node558;
										assign node558 = (inp[1]) ? node566 : node559;
											assign node559 = (inp[5]) ? 4'b0010 : node560;
												assign node560 = (inp[15]) ? node562 : 4'b1000;
													assign node562 = (inp[6]) ? 4'b1000 : 4'b0010;
											assign node566 = (inp[15]) ? node568 : 4'b1000;
												assign node568 = (inp[6]) ? 4'b1000 : node569;
													assign node569 = (inp[5]) ? 4'b0010 : 4'b1000;
										assign node573 = (inp[1]) ? node575 : 4'b1000;
											assign node575 = (inp[5]) ? 4'b1000 : node576;
												assign node576 = (inp[6]) ? 4'b1010 : node577;
													assign node577 = (inp[15]) ? 4'b1000 : node578;
														assign node578 = (inp[10]) ? node580 : 4'b1010;
															assign node580 = (inp[8]) ? 4'b1000 : 4'b1010;
									assign node586 = (inp[13]) ? node588 : 4'b0010;
										assign node588 = (inp[5]) ? node596 : node589;
											assign node589 = (inp[1]) ? 4'b1000 : node590;
												assign node590 = (inp[15]) ? node592 : 4'b1000;
													assign node592 = (inp[6]) ? 4'b1000 : 4'b0010;
											assign node596 = (inp[1]) ? node598 : 4'b0010;
												assign node598 = (inp[15]) ? node600 : 4'b1000;
													assign node600 = (inp[6]) ? 4'b1000 : 4'b0010;
								assign node603 = (inp[11]) ? node645 : node604;
									assign node604 = (inp[13]) ? node632 : node605;
										assign node605 = (inp[5]) ? node621 : node606;
											assign node606 = (inp[1]) ? 4'b0010 : node607;
												assign node607 = (inp[15]) ? node615 : node608;
													assign node608 = (inp[6]) ? 4'b0010 : node609;
														assign node609 = (inp[10]) ? node611 : 4'b0010;
															assign node611 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node615 = (inp[6]) ? node617 : 4'b0000;
														assign node617 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node621 = (inp[15]) ? 4'b0000 : node622;
												assign node622 = (inp[1]) ? node624 : 4'b0000;
													assign node624 = (inp[6]) ? 4'b0010 : node625;
														assign node625 = (inp[8]) ? 4'b0000 : node626;
															assign node626 = (inp[10]) ? 4'b0000 : 4'b0010;
										assign node632 = (inp[6]) ? 4'b0010 : node633;
											assign node633 = (inp[1]) ? 4'b0010 : node634;
												assign node634 = (inp[15]) ? node636 : 4'b0010;
													assign node636 = (inp[10]) ? node638 : 4'b0010;
														assign node638 = (inp[5]) ? node640 : 4'b0010;
															assign node640 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node645 = (inp[13]) ? node647 : 4'b0000;
										assign node647 = (inp[5]) ? 4'b0000 : node648;
											assign node648 = (inp[1]) ? node656 : node649;
												assign node649 = (inp[6]) ? node651 : 4'b0000;
													assign node651 = (inp[8]) ? 4'b0000 : node652;
														assign node652 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node656 = (inp[6]) ? 4'b0010 : node657;
													assign node657 = (inp[15]) ? node659 : 4'b0010;
														assign node659 = (inp[10]) ? 4'b0000 : node660;
															assign node660 = (inp[8]) ? 4'b0000 : 4'b0010;
							assign node666 = (inp[13]) ? node826 : node667;
								assign node667 = (inp[4]) ? node757 : node668;
									assign node668 = (inp[1]) ? node696 : node669;
										assign node669 = (inp[11]) ? node681 : node670;
											assign node670 = (inp[6]) ? node674 : node671;
												assign node671 = (inp[5]) ? 4'b1010 : 4'b0000;
												assign node674 = (inp[8]) ? 4'b0000 : node675;
													assign node675 = (inp[15]) ? 4'b0000 : node676;
														assign node676 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node681 = (inp[5]) ? node689 : node682;
												assign node682 = (inp[15]) ? node684 : 4'b1010;
													assign node684 = (inp[6]) ? 4'b1010 : node685;
														assign node685 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node689 = (inp[6]) ? node691 : 4'b1000;
													assign node691 = (inp[15]) ? node693 : 4'b1010;
														assign node693 = (inp[8]) ? 4'b1000 : 4'b1010;
										assign node696 = (inp[11]) ? node748 : node697;
											assign node697 = (inp[15]) ? node709 : node698;
												assign node698 = (inp[5]) ? node702 : node699;
													assign node699 = (inp[6]) ? 4'b0000 : 4'b0010;
													assign node702 = (inp[6]) ? 4'b0010 : node703;
														assign node703 = (inp[8]) ? node705 : 4'b0010;
															assign node705 = (inp[10]) ? 4'b0000 : 4'b0010;
												assign node709 = (inp[10]) ? node725 : node710;
													assign node710 = (inp[8]) ? node718 : node711;
														assign node711 = (inp[5]) ? node715 : node712;
															assign node712 = (inp[6]) ? 4'b0000 : 4'b0010;
															assign node715 = (inp[6]) ? 4'b0010 : 4'b0000;
														assign node718 = (inp[5]) ? node722 : node719;
															assign node719 = (inp[6]) ? 4'b0000 : 4'b0010;
															assign node722 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node725 = (inp[2]) ? node733 : node726;
														assign node726 = (inp[5]) ? node730 : node727;
															assign node727 = (inp[6]) ? 4'b0000 : 4'b0010;
															assign node730 = (inp[6]) ? 4'b0010 : 4'b0000;
														assign node733 = (inp[8]) ? node741 : node734;
															assign node734 = (inp[5]) ? node738 : node735;
																assign node735 = (inp[6]) ? 4'b0000 : 4'b0010;
																assign node738 = (inp[6]) ? 4'b0010 : 4'b0000;
															assign node741 = (inp[5]) ? node745 : node742;
																assign node742 = (inp[6]) ? 4'b0000 : 4'b0010;
																assign node745 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node748 = (inp[5]) ? node754 : node749;
												assign node749 = (inp[6]) ? node751 : 4'b0000;
													assign node751 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node754 = (inp[6]) ? 4'b0000 : 4'b1010;
									assign node757 = (inp[1]) ? node789 : node758;
										assign node758 = (inp[5]) ? node776 : node759;
											assign node759 = (inp[11]) ? node767 : node760;
												assign node760 = (inp[15]) ? node762 : 4'b1000;
													assign node762 = (inp[8]) ? node764 : 4'b1000;
														assign node764 = (inp[6]) ? 4'b1000 : 4'b1010;
												assign node767 = (inp[15]) ? node769 : 4'b1010;
													assign node769 = (inp[6]) ? 4'b1010 : node770;
														assign node770 = (inp[8]) ? 4'b1000 : node771;
															assign node771 = (inp[2]) ? 4'b1000 : 4'b1010;
											assign node776 = (inp[11]) ? node782 : node777;
												assign node777 = (inp[6]) ? node779 : 4'b1010;
													assign node779 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node782 = (inp[15]) ? 4'b1000 : node783;
													assign node783 = (inp[8]) ? 4'b1000 : node784;
														assign node784 = (inp[6]) ? 4'b1010 : 4'b1000;
										assign node789 = (inp[15]) ? node805 : node790;
											assign node790 = (inp[6]) ? node800 : node791;
												assign node791 = (inp[11]) ? node795 : node792;
													assign node792 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node795 = (inp[5]) ? 4'b1010 : node796;
														assign node796 = (inp[8]) ? 4'b1010 : 4'b1000;
												assign node800 = (inp[5]) ? 4'b1010 : node801;
													assign node801 = (inp[11]) ? 4'b1000 : 4'b1010;
											assign node805 = (inp[11]) ? node815 : node806;
												assign node806 = (inp[5]) ? 4'b1000 : node807;
													assign node807 = (inp[6]) ? 4'b1010 : node808;
														assign node808 = (inp[10]) ? 4'b1000 : node809;
															assign node809 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node815 = (inp[6]) ? node823 : node816;
													assign node816 = (inp[5]) ? node818 : 4'b1010;
														assign node818 = (inp[10]) ? node820 : 4'b1010;
															assign node820 = (inp[8]) ? 4'b1000 : 4'b1010;
													assign node823 = (inp[5]) ? 4'b1010 : 4'b1000;
								assign node826 = (inp[5]) ? node888 : node827;
									assign node827 = (inp[6]) ? node869 : node828;
										assign node828 = (inp[4]) ? node852 : node829;
											assign node829 = (inp[1]) ? node843 : node830;
												assign node830 = (inp[8]) ? node836 : node831;
													assign node831 = (inp[15]) ? 4'b0010 : node832;
														assign node832 = (inp[11]) ? 4'b0000 : 4'b0010;
													assign node836 = (inp[15]) ? node838 : 4'b0010;
														assign node838 = (inp[10]) ? node840 : 4'b0010;
															assign node840 = (inp[11]) ? 4'b0010 : 4'b0000;
												assign node843 = (inp[15]) ? node849 : node844;
													assign node844 = (inp[8]) ? node846 : 4'b1000;
														assign node846 = (inp[11]) ? 4'b1000 : 4'b1010;
													assign node849 = (inp[11]) ? 4'b0010 : 4'b1010;
											assign node852 = (inp[1]) ? node862 : node853;
												assign node853 = (inp[11]) ? node855 : 4'b0000;
													assign node855 = (inp[15]) ? 4'b1000 : node856;
														assign node856 = (inp[8]) ? node858 : 4'b1010;
															assign node858 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node862 = (inp[8]) ? node864 : 4'b0000;
													assign node864 = (inp[11]) ? 4'b0000 : node865;
														assign node865 = (inp[15]) ? 4'b0010 : 4'b0000;
										assign node869 = (inp[4]) ? node879 : node870;
											assign node870 = (inp[1]) ? 4'b1010 : node871;
												assign node871 = (inp[11]) ? node873 : 4'b1000;
													assign node873 = (inp[8]) ? 4'b0000 : node874;
														assign node874 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node879 = (inp[1]) ? 4'b0010 : node880;
												assign node880 = (inp[11]) ? 4'b1010 : node881;
													assign node881 = (inp[8]) ? node883 : 4'b0010;
														assign node883 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node888 = (inp[6]) ? node924 : node889;
										assign node889 = (inp[4]) ? node907 : node890;
											assign node890 = (inp[11]) ? node900 : node891;
												assign node891 = (inp[1]) ? node893 : 4'b0000;
													assign node893 = (inp[15]) ? 4'b1000 : node894;
														assign node894 = (inp[8]) ? node896 : 4'b1010;
															assign node896 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node900 = (inp[15]) ? node902 : 4'b0010;
													assign node902 = (inp[8]) ? 4'b0000 : node903;
														assign node903 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node907 = (inp[1]) ? node915 : node908;
												assign node908 = (inp[11]) ? node910 : 4'b1010;
													assign node910 = (inp[15]) ? node912 : 4'b1000;
														assign node912 = (inp[8]) ? 4'b1010 : 4'b1000;
												assign node915 = (inp[11]) ? 4'b1010 : node916;
													assign node916 = (inp[10]) ? node918 : 4'b0010;
														assign node918 = (inp[8]) ? node920 : 4'b0010;
															assign node920 = (inp[15]) ? 4'b0000 : 4'b0010;
										assign node924 = (inp[1]) ? node938 : node925;
											assign node925 = (inp[4]) ? node931 : node926;
												assign node926 = (inp[11]) ? node928 : 4'b0010;
													assign node928 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node931 = (inp[11]) ? node933 : 4'b0000;
													assign node933 = (inp[8]) ? 4'b1000 : node934;
														assign node934 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node938 = (inp[4]) ? 4'b0000 : 4'b1000;
						assign node941 = (inp[7]) ? node1113 : node942;
							assign node942 = (inp[4]) ? node1036 : node943;
								assign node943 = (inp[11]) ? node993 : node944;
									assign node944 = (inp[13]) ? node966 : node945;
										assign node945 = (inp[5]) ? node955 : node946;
											assign node946 = (inp[1]) ? node948 : 4'b1010;
												assign node948 = (inp[6]) ? 4'b1000 : node949;
													assign node949 = (inp[8]) ? 4'b1010 : node950;
														assign node950 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node955 = (inp[15]) ? node957 : 4'b1010;
												assign node957 = (inp[1]) ? 4'b1010 : node958;
													assign node958 = (inp[6]) ? 4'b1010 : node959;
														assign node959 = (inp[10]) ? 4'b1000 : node960;
															assign node960 = (inp[8]) ? 4'b1000 : 4'b1010;
										assign node966 = (inp[1]) ? node982 : node967;
											assign node967 = (inp[6]) ? node975 : node968;
												assign node968 = (inp[15]) ? node970 : 4'b1000;
													assign node970 = (inp[5]) ? node972 : 4'b1000;
														assign node972 = (inp[8]) ? 4'b1010 : 4'b1000;
												assign node975 = (inp[8]) ? 4'b1000 : node976;
													assign node976 = (inp[15]) ? 4'b1000 : node977;
														assign node977 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node982 = (inp[6]) ? 4'b1010 : node983;
												assign node983 = (inp[5]) ? node985 : 4'b1010;
													assign node985 = (inp[8]) ? 4'b1000 : node986;
														assign node986 = (inp[15]) ? 4'b1000 : node987;
															assign node987 = (inp[10]) ? 4'b1000 : 4'b1010;
									assign node993 = (inp[13]) ? node1019 : node994;
										assign node994 = (inp[1]) ? node1004 : node995;
											assign node995 = (inp[8]) ? 4'b1000 : node996;
												assign node996 = (inp[15]) ? 4'b1000 : node997;
													assign node997 = (inp[6]) ? node999 : 4'b1000;
														assign node999 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node1004 = (inp[5]) ? node1014 : node1005;
												assign node1005 = (inp[15]) ? node1007 : 4'b1010;
													assign node1007 = (inp[10]) ? node1009 : 4'b1010;
														assign node1009 = (inp[6]) ? 4'b1010 : node1010;
															assign node1010 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node1014 = (inp[15]) ? 4'b1000 : node1015;
													assign node1015 = (inp[6]) ? 4'b1010 : 4'b1000;
										assign node1019 = (inp[1]) ? node1027 : node1020;
											assign node1020 = (inp[5]) ? 4'b1010 : node1021;
												assign node1021 = (inp[6]) ? node1023 : 4'b1010;
													assign node1023 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node1027 = (inp[5]) ? node1029 : 4'b1000;
												assign node1029 = (inp[6]) ? 4'b1000 : node1030;
													assign node1030 = (inp[15]) ? 4'b1010 : node1031;
														assign node1031 = (inp[8]) ? 4'b1010 : 4'b1000;
								assign node1036 = (inp[13]) ? node1070 : node1037;
									assign node1037 = (inp[11]) ? node1053 : node1038;
										assign node1038 = (inp[1]) ? node1046 : node1039;
											assign node1039 = (inp[5]) ? 4'b0010 : node1040;
												assign node1040 = (inp[15]) ? node1042 : 4'b1000;
													assign node1042 = (inp[6]) ? 4'b1000 : 4'b0010;
											assign node1046 = (inp[6]) ? 4'b1000 : node1047;
												assign node1047 = (inp[15]) ? node1049 : 4'b1000;
													assign node1049 = (inp[5]) ? 4'b0010 : 4'b1000;
										assign node1053 = (inp[5]) ? node1055 : 4'b0010;
											assign node1055 = (inp[1]) ? 4'b0010 : node1056;
												assign node1056 = (inp[15]) ? node1064 : node1057;
													assign node1057 = (inp[10]) ? node1059 : 4'b0010;
														assign node1059 = (inp[8]) ? node1061 : 4'b0010;
															assign node1061 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1064 = (inp[8]) ? 4'b0000 : node1065;
														assign node1065 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node1070 = (inp[11]) ? node1098 : node1071;
										assign node1071 = (inp[1]) ? node1087 : node1072;
											assign node1072 = (inp[5]) ? 4'b1000 : node1073;
												assign node1073 = (inp[6]) ? node1081 : node1074;
													assign node1074 = (inp[10]) ? 4'b1000 : node1075;
														assign node1075 = (inp[8]) ? 4'b1000 : node1076;
															assign node1076 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node1081 = (inp[8]) ? node1083 : 4'b1010;
														assign node1083 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node1087 = (inp[5]) ? node1089 : 4'b1010;
												assign node1089 = (inp[6]) ? 4'b1010 : node1090;
													assign node1090 = (inp[15]) ? 4'b1000 : node1091;
														assign node1091 = (inp[10]) ? node1093 : 4'b1010;
															assign node1093 = (inp[8]) ? 4'b1000 : 4'b1010;
										assign node1098 = (inp[5]) ? node1106 : node1099;
											assign node1099 = (inp[15]) ? node1101 : 4'b1000;
												assign node1101 = (inp[6]) ? 4'b1000 : node1102;
													assign node1102 = (inp[1]) ? 4'b1000 : 4'b0010;
											assign node1106 = (inp[1]) ? node1108 : 4'b0010;
												assign node1108 = (inp[6]) ? 4'b1000 : node1109;
													assign node1109 = (inp[15]) ? 4'b0010 : 4'b1000;
							assign node1113 = (inp[13]) ? node1287 : node1114;
								assign node1114 = (inp[4]) ? node1206 : node1115;
									assign node1115 = (inp[1]) ? node1167 : node1116;
										assign node1116 = (inp[6]) ? node1146 : node1117;
											assign node1117 = (inp[11]) ? node1133 : node1118;
												assign node1118 = (inp[5]) ? node1124 : node1119;
													assign node1119 = (inp[8]) ? 4'b0011 : node1120;
														assign node1120 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node1124 = (inp[10]) ? 4'b0001 : node1125;
														assign node1125 = (inp[2]) ? 4'b0001 : node1126;
															assign node1126 = (inp[8]) ? 4'b0001 : node1127;
																assign node1127 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node1133 = (inp[5]) ? node1141 : node1134;
													assign node1134 = (inp[8]) ? node1136 : 4'b1010;
														assign node1136 = (inp[15]) ? node1138 : 4'b1010;
															assign node1138 = (inp[10]) ? 4'b1000 : 4'b1010;
													assign node1141 = (inp[8]) ? node1143 : 4'b1000;
														assign node1143 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node1146 = (inp[11]) ? node1158 : node1147;
												assign node1147 = (inp[5]) ? node1153 : node1148;
													assign node1148 = (inp[8]) ? 4'b1001 : node1149;
														assign node1149 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node1153 = (inp[8]) ? node1155 : 4'b0011;
														assign node1155 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node1158 = (inp[5]) ? node1162 : node1159;
													assign node1159 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node1162 = (inp[15]) ? 4'b0001 : node1163;
														assign node1163 = (inp[8]) ? 4'b0001 : 4'b0011;
										assign node1167 = (inp[15]) ? node1185 : node1168;
											assign node1168 = (inp[6]) ? node1182 : node1169;
												assign node1169 = (inp[11]) ? node1177 : node1170;
													assign node1170 = (inp[5]) ? 4'b1011 : node1171;
														assign node1171 = (inp[10]) ? node1173 : 4'b0011;
															assign node1173 = (inp[8]) ? 4'b0001 : 4'b0011;
													assign node1177 = (inp[5]) ? 4'b1001 : node1178;
														assign node1178 = (inp[8]) ? 4'b1011 : 4'b1001;
												assign node1182 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node1185 = (inp[11]) ? node1197 : node1186;
												assign node1186 = (inp[5]) ? node1190 : node1187;
													assign node1187 = (inp[6]) ? 4'b1001 : 4'b0001;
													assign node1190 = (inp[6]) ? 4'b1001 : node1191;
														assign node1191 = (inp[8]) ? 4'b1001 : node1192;
															assign node1192 = (inp[10]) ? 4'b1001 : 4'b1011;
												assign node1197 = (inp[6]) ? 4'b0001 : node1198;
													assign node1198 = (inp[5]) ? 4'b0011 : node1199;
														assign node1199 = (inp[8]) ? node1201 : 4'b1011;
															assign node1201 = (inp[10]) ? 4'b1001 : 4'b1011;
									assign node1206 = (inp[1]) ? node1248 : node1207;
										assign node1207 = (inp[11]) ? node1223 : node1208;
											assign node1208 = (inp[5]) ? node1218 : node1209;
												assign node1209 = (inp[15]) ? node1211 : 4'b1010;
													assign node1211 = (inp[8]) ? 4'b1000 : node1212;
														assign node1212 = (inp[6]) ? 4'b1010 : node1213;
															assign node1213 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node1218 = (inp[15]) ? node1220 : 4'b1000;
													assign node1220 = (inp[6]) ? 4'b1010 : 4'b0010;
											assign node1223 = (inp[5]) ? node1237 : node1224;
												assign node1224 = (inp[6]) ? node1232 : node1225;
													assign node1225 = (inp[15]) ? 4'b0000 : node1226;
														assign node1226 = (inp[8]) ? node1228 : 4'b0010;
															assign node1228 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1232 = (inp[8]) ? 4'b1000 : node1233;
														assign node1233 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node1237 = (inp[15]) ? node1243 : node1238;
													assign node1238 = (inp[6]) ? 4'b0010 : node1239;
														assign node1239 = (inp[8]) ? 4'b0010 : 4'b0000;
													assign node1243 = (inp[8]) ? node1245 : 4'b0010;
														assign node1245 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node1248 = (inp[15]) ? node1266 : node1249;
											assign node1249 = (inp[6]) ? node1263 : node1250;
												assign node1250 = (inp[11]) ? node1258 : node1251;
													assign node1251 = (inp[8]) ? 4'b0001 : node1252;
														assign node1252 = (inp[10]) ? node1254 : 4'b0011;
															assign node1254 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node1258 = (inp[8]) ? 4'b1010 : node1259;
														assign node1259 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node1263 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node1266 = (inp[6]) ? node1284 : node1267;
												assign node1267 = (inp[11]) ? node1273 : node1268;
													assign node1268 = (inp[8]) ? node1270 : 4'b0001;
														assign node1270 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node1273 = (inp[10]) ? node1279 : node1274;
														assign node1274 = (inp[8]) ? node1276 : 4'b1010;
															assign node1276 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node1279 = (inp[8]) ? 4'b1000 : node1280;
															assign node1280 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node1284 = (inp[11]) ? 4'b0001 : 4'b1001;
								assign node1287 = (inp[6]) ? node1407 : node1288;
									assign node1288 = (inp[1]) ? node1392 : node1289;
										assign node1289 = (inp[4]) ? node1351 : node1290;
											assign node1290 = (inp[10]) ? node1318 : node1291;
												assign node1291 = (inp[5]) ? node1305 : node1292;
													assign node1292 = (inp[15]) ? node1300 : node1293;
														assign node1293 = (inp[11]) ? node1297 : node1294;
															assign node1294 = (inp[8]) ? 4'b0010 : 4'b0000;
															assign node1297 = (inp[8]) ? 4'b1000 : 4'b1010;
														assign node1300 = (inp[8]) ? node1302 : 4'b0010;
															assign node1302 = (inp[11]) ? 4'b0010 : 4'b0000;
													assign node1305 = (inp[11]) ? node1311 : node1306;
														assign node1306 = (inp[15]) ? node1308 : 4'b1010;
															assign node1308 = (inp[8]) ? 4'b1010 : 4'b1000;
														assign node1311 = (inp[15]) ? node1315 : node1312;
															assign node1312 = (inp[8]) ? 4'b0010 : 4'b0000;
															assign node1315 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node1318 = (inp[5]) ? node1330 : node1319;
													assign node1319 = (inp[11]) ? node1325 : node1320;
														assign node1320 = (inp[8]) ? node1322 : 4'b0000;
															assign node1322 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node1325 = (inp[15]) ? node1327 : 4'b1000;
															assign node1327 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1330 = (inp[11]) ? node1346 : node1331;
														assign node1331 = (inp[2]) ? node1339 : node1332;
															assign node1332 = (inp[15]) ? node1336 : node1333;
																assign node1333 = (inp[8]) ? 4'b1000 : 4'b1010;
																assign node1336 = (inp[8]) ? 4'b1010 : 4'b1000;
															assign node1339 = (inp[8]) ? node1343 : node1340;
																assign node1340 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node1343 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node1346 = (inp[15]) ? 4'b0000 : node1347;
															assign node1347 = (inp[8]) ? 4'b0010 : 4'b0000;
											assign node1351 = (inp[5]) ? node1371 : node1352;
												assign node1352 = (inp[11]) ? node1362 : node1353;
													assign node1353 = (inp[8]) ? node1357 : node1354;
														assign node1354 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node1357 = (inp[10]) ? node1359 : 4'b1011;
															assign node1359 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node1362 = (inp[15]) ? node1366 : node1363;
														assign node1363 = (inp[8]) ? 4'b0011 : 4'b0001;
														assign node1366 = (inp[8]) ? 4'b0001 : node1367;
															assign node1367 = (inp[10]) ? 4'b0001 : 4'b0011;
												assign node1371 = (inp[11]) ? node1383 : node1372;
													assign node1372 = (inp[15]) ? node1378 : node1373;
														assign node1373 = (inp[8]) ? 4'b1001 : node1374;
															assign node1374 = (inp[10]) ? 4'b1001 : 4'b1011;
														assign node1378 = (inp[10]) ? node1380 : 4'b0011;
															assign node1380 = (inp[8]) ? 4'b0001 : 4'b0011;
													assign node1383 = (inp[15]) ? node1389 : node1384;
														assign node1384 = (inp[8]) ? node1386 : 4'b1011;
															assign node1386 = (inp[10]) ? 4'b1001 : 4'b1011;
														assign node1389 = (inp[8]) ? 4'b1011 : 4'b1001;
										assign node1392 = (inp[11]) ? node1400 : node1393;
											assign node1393 = (inp[10]) ? node1397 : node1394;
												assign node1394 = (inp[15]) ? 4'b0111 : 4'b1111;
												assign node1397 = (inp[15]) ? 4'b0101 : 4'b1101;
											assign node1400 = (inp[10]) ? node1404 : node1401;
												assign node1401 = (inp[15]) ? 4'b0110 : 4'b1110;
												assign node1404 = (inp[15]) ? 4'b0100 : 4'b1100;
									assign node1407 = (inp[1]) ? 4'b0000 : node1408;
										assign node1408 = (inp[4]) ? node1416 : node1409;
											assign node1409 = (inp[5]) ? node1413 : node1410;
												assign node1410 = (inp[8]) ? 4'b1001 : 4'b1011;
												assign node1413 = (inp[8]) ? 4'b0001 : 4'b0011;
											assign node1416 = (inp[8]) ? node1420 : node1417;
												assign node1417 = (inp[5]) ? 4'b0010 : 4'b1010;
												assign node1420 = (inp[5]) ? 4'b0000 : 4'b1000;
			assign node1424 = (inp[0]) ? node1426 : 4'b0000;
				assign node1426 = (inp[4]) ? node1978 : node1427;
					assign node1427 = (inp[7]) ? node1621 : node1428;
						assign node1428 = (inp[3]) ? node1504 : node1429;
							assign node1429 = (inp[11]) ? 4'b0000 : node1430;
								assign node1430 = (inp[9]) ? node1466 : node1431;
									assign node1431 = (inp[5]) ? 4'b0000 : node1432;
										assign node1432 = (inp[13]) ? node1448 : node1433;
											assign node1433 = (inp[15]) ? 4'b0000 : node1434;
												assign node1434 = (inp[8]) ? node1442 : node1435;
													assign node1435 = (inp[1]) ? 4'b0010 : node1436;
														assign node1436 = (inp[6]) ? 4'b0010 : node1437;
															assign node1437 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1442 = (inp[1]) ? node1444 : 4'b0000;
														assign node1444 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node1448 = (inp[15]) ? node1450 : 4'b0010;
												assign node1450 = (inp[8]) ? node1458 : node1451;
													assign node1451 = (inp[10]) ? node1453 : 4'b0010;
														assign node1453 = (inp[6]) ? 4'b0010 : node1454;
															assign node1454 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node1458 = (inp[1]) ? node1460 : 4'b0000;
														assign node1460 = (inp[10]) ? node1462 : 4'b0010;
															assign node1462 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node1466 = (inp[5]) ? node1468 : 4'b0010;
										assign node1468 = (inp[13]) ? node1486 : node1469;
											assign node1469 = (inp[15]) ? 4'b0000 : node1470;
												assign node1470 = (inp[1]) ? node1478 : node1471;
													assign node1471 = (inp[8]) ? 4'b0000 : node1472;
														assign node1472 = (inp[10]) ? node1474 : 4'b0010;
															assign node1474 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1478 = (inp[10]) ? node1480 : 4'b0010;
														assign node1480 = (inp[6]) ? 4'b0010 : node1481;
															assign node1481 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node1486 = (inp[15]) ? node1488 : 4'b0010;
												assign node1488 = (inp[8]) ? node1496 : node1489;
													assign node1489 = (inp[10]) ? node1491 : 4'b0010;
														assign node1491 = (inp[6]) ? 4'b0010 : node1492;
															assign node1492 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node1496 = (inp[1]) ? node1498 : 4'b0000;
														assign node1498 = (inp[6]) ? 4'b0010 : node1499;
															assign node1499 = (inp[10]) ? 4'b0000 : 4'b0010;
							assign node1504 = (inp[11]) ? node1584 : node1505;
								assign node1505 = (inp[13]) ? node1537 : node1506;
									assign node1506 = (inp[9]) ? node1524 : node1507;
										assign node1507 = (inp[5]) ? 4'b0010 : node1508;
											assign node1508 = (inp[1]) ? node1516 : node1509;
												assign node1509 = (inp[15]) ? 4'b0010 : node1510;
													assign node1510 = (inp[8]) ? node1512 : 4'b0000;
														assign node1512 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node1516 = (inp[6]) ? 4'b0000 : node1517;
													assign node1517 = (inp[15]) ? node1519 : 4'b0000;
														assign node1519 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node1524 = (inp[5]) ? 4'b0000 : node1525;
											assign node1525 = (inp[15]) ? 4'b0000 : node1526;
												assign node1526 = (inp[1]) ? node1528 : 4'b0000;
													assign node1528 = (inp[6]) ? 4'b0010 : node1529;
														assign node1529 = (inp[10]) ? 4'b0000 : node1530;
															assign node1530 = (inp[2]) ? 4'b0010 : 4'b0000;
									assign node1537 = (inp[9]) ? node1555 : node1538;
										assign node1538 = (inp[5]) ? node1540 : 4'b0000;
											assign node1540 = (inp[1]) ? node1548 : node1541;
												assign node1541 = (inp[15]) ? 4'b0010 : node1542;
													assign node1542 = (inp[6]) ? 4'b0000 : node1543;
														assign node1543 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node1548 = (inp[15]) ? node1550 : 4'b0000;
													assign node1550 = (inp[8]) ? node1552 : 4'b0000;
														assign node1552 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node1555 = (inp[5]) ? node1567 : node1556;
											assign node1556 = (inp[15]) ? node1558 : 4'b0010;
												assign node1558 = (inp[8]) ? node1560 : 4'b0010;
													assign node1560 = (inp[1]) ? 4'b0010 : node1561;
														assign node1561 = (inp[6]) ? 4'b0010 : node1562;
															assign node1562 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node1567 = (inp[1]) ? node1575 : node1568;
												assign node1568 = (inp[6]) ? node1570 : 4'b0000;
													assign node1570 = (inp[15]) ? 4'b0000 : node1571;
														assign node1571 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node1575 = (inp[15]) ? node1577 : 4'b0010;
													assign node1577 = (inp[6]) ? 4'b0010 : node1578;
														assign node1578 = (inp[10]) ? 4'b0000 : node1579;
															assign node1579 = (inp[8]) ? 4'b0000 : 4'b0010;
								assign node1584 = (inp[9]) ? node1586 : 4'b0010;
									assign node1586 = (inp[13]) ? node1604 : node1587;
										assign node1587 = (inp[5]) ? 4'b0010 : node1588;
											assign node1588 = (inp[15]) ? node1596 : node1589;
												assign node1589 = (inp[6]) ? 4'b0000 : node1590;
													assign node1590 = (inp[8]) ? node1592 : 4'b0000;
														assign node1592 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node1596 = (inp[1]) ? node1598 : 4'b0010;
													assign node1598 = (inp[8]) ? node1600 : 4'b0000;
														assign node1600 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node1604 = (inp[5]) ? node1606 : 4'b0000;
											assign node1606 = (inp[15]) ? node1614 : node1607;
												assign node1607 = (inp[1]) ? 4'b0000 : node1608;
													assign node1608 = (inp[8]) ? node1610 : 4'b0000;
														assign node1610 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node1614 = (inp[1]) ? node1616 : 4'b0010;
													assign node1616 = (inp[6]) ? 4'b0000 : node1617;
														assign node1617 = (inp[8]) ? 4'b0010 : 4'b0000;
						assign node1621 = (inp[3]) ? node1699 : node1622;
							assign node1622 = (inp[11]) ? node1624 : 4'b0010;
								assign node1624 = (inp[5]) ? node1662 : node1625;
									assign node1625 = (inp[9]) ? 4'b0010 : node1626;
										assign node1626 = (inp[13]) ? node1644 : node1627;
											assign node1627 = (inp[15]) ? 4'b0000 : node1628;
												assign node1628 = (inp[1]) ? node1636 : node1629;
													assign node1629 = (inp[8]) ? 4'b0000 : node1630;
														assign node1630 = (inp[10]) ? node1632 : 4'b0010;
															assign node1632 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1636 = (inp[10]) ? node1638 : 4'b0010;
														assign node1638 = (inp[8]) ? node1640 : 4'b0010;
															assign node1640 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node1644 = (inp[15]) ? node1646 : 4'b0010;
												assign node1646 = (inp[1]) ? node1654 : node1647;
													assign node1647 = (inp[8]) ? 4'b0000 : node1648;
														assign node1648 = (inp[6]) ? 4'b0010 : node1649;
															assign node1649 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1654 = (inp[8]) ? node1656 : 4'b0010;
														assign node1656 = (inp[6]) ? 4'b0010 : node1657;
															assign node1657 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node1662 = (inp[9]) ? node1664 : 4'b0000;
										assign node1664 = (inp[13]) ? node1682 : node1665;
											assign node1665 = (inp[15]) ? 4'b0000 : node1666;
												assign node1666 = (inp[8]) ? node1674 : node1667;
													assign node1667 = (inp[6]) ? 4'b0010 : node1668;
														assign node1668 = (inp[1]) ? 4'b0010 : node1669;
															assign node1669 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1674 = (inp[1]) ? node1676 : 4'b0000;
														assign node1676 = (inp[6]) ? 4'b0010 : node1677;
															assign node1677 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node1682 = (inp[15]) ? node1684 : 4'b0010;
												assign node1684 = (inp[8]) ? node1692 : node1685;
													assign node1685 = (inp[1]) ? 4'b0010 : node1686;
														assign node1686 = (inp[6]) ? 4'b0010 : node1687;
															assign node1687 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1692 = (inp[1]) ? node1694 : 4'b0000;
														assign node1694 = (inp[6]) ? 4'b0010 : node1695;
															assign node1695 = (inp[10]) ? 4'b0000 : 4'b0010;
							assign node1699 = (inp[13]) ? node1829 : node1700;
								assign node1700 = (inp[11]) ? node1762 : node1701;
									assign node1701 = (inp[1]) ? node1735 : node1702;
										assign node1702 = (inp[5]) ? node1720 : node1703;
											assign node1703 = (inp[9]) ? node1709 : node1704;
												assign node1704 = (inp[6]) ? 4'b1000 : node1705;
													assign node1705 = (inp[15]) ? 4'b0010 : 4'b1000;
												assign node1709 = (inp[6]) ? node1717 : node1710;
													assign node1710 = (inp[10]) ? 4'b0000 : node1711;
														assign node1711 = (inp[8]) ? 4'b0000 : node1712;
															assign node1712 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node1717 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node1720 = (inp[9]) ? node1722 : 4'b0010;
												assign node1722 = (inp[6]) ? node1730 : node1723;
													assign node1723 = (inp[10]) ? node1725 : 4'b1010;
														assign node1725 = (inp[8]) ? node1727 : 4'b1010;
															assign node1727 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node1730 = (inp[8]) ? 4'b0000 : node1731;
														assign node1731 = (inp[15]) ? 4'b0000 : 4'b0010;
										assign node1735 = (inp[6]) ? node1755 : node1736;
											assign node1736 = (inp[15]) ? node1746 : node1737;
												assign node1737 = (inp[9]) ? node1739 : 4'b1000;
													assign node1739 = (inp[5]) ? node1741 : 4'b1000;
														assign node1741 = (inp[8]) ? 4'b0000 : node1742;
															assign node1742 = (inp[10]) ? 4'b0000 : 4'b0010;
												assign node1746 = (inp[9]) ? node1750 : node1747;
													assign node1747 = (inp[5]) ? 4'b0010 : 4'b1000;
													assign node1750 = (inp[5]) ? node1752 : 4'b0010;
														assign node1752 = (inp[8]) ? 4'b0010 : 4'b0000;
											assign node1755 = (inp[15]) ? 4'b1000 : node1756;
												assign node1756 = (inp[5]) ? node1758 : 4'b1010;
													assign node1758 = (inp[9]) ? 4'b1010 : 4'b1000;
									assign node1762 = (inp[9]) ? node1790 : node1763;
										assign node1763 = (inp[5]) ? node1779 : node1764;
											assign node1764 = (inp[1]) ? 4'b0010 : node1765;
												assign node1765 = (inp[15]) ? node1773 : node1766;
													assign node1766 = (inp[6]) ? 4'b0010 : node1767;
														assign node1767 = (inp[10]) ? node1769 : 4'b0010;
															assign node1769 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1773 = (inp[6]) ? node1775 : 4'b0000;
														assign node1775 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node1779 = (inp[1]) ? node1781 : 4'b0000;
												assign node1781 = (inp[15]) ? 4'b0000 : node1782;
													assign node1782 = (inp[6]) ? 4'b0010 : node1783;
														assign node1783 = (inp[8]) ? 4'b0000 : node1784;
															assign node1784 = (inp[10]) ? 4'b0000 : 4'b0010;
										assign node1790 = (inp[1]) ? node1814 : node1791;
											assign node1791 = (inp[6]) ? node1805 : node1792;
												assign node1792 = (inp[5]) ? node1798 : node1793;
													assign node1793 = (inp[8]) ? node1795 : 4'b1000;
														assign node1795 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node1798 = (inp[15]) ? node1800 : 4'b1010;
														assign node1800 = (inp[8]) ? 4'b1000 : node1801;
															assign node1801 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node1805 = (inp[15]) ? node1809 : node1806;
													assign node1806 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node1809 = (inp[8]) ? node1811 : 4'b1010;
														assign node1811 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node1814 = (inp[15]) ? node1820 : node1815;
												assign node1815 = (inp[6]) ? 4'b0010 : node1816;
													assign node1816 = (inp[5]) ? 4'b1010 : 4'b0010;
												assign node1820 = (inp[6]) ? 4'b0000 : node1821;
													assign node1821 = (inp[5]) ? node1823 : 4'b0000;
														assign node1823 = (inp[8]) ? 4'b1000 : node1824;
															assign node1824 = (inp[10]) ? 4'b1000 : 4'b1010;
								assign node1829 = (inp[9]) ? node1901 : node1830;
									assign node1830 = (inp[11]) ? node1870 : node1831;
										assign node1831 = (inp[5]) ? node1847 : node1832;
											assign node1832 = (inp[1]) ? node1838 : node1833;
												assign node1833 = (inp[15]) ? 4'b1010 : node1834;
													assign node1834 = (inp[6]) ? 4'b1000 : 4'b1010;
												assign node1838 = (inp[6]) ? 4'b1010 : node1839;
													assign node1839 = (inp[15]) ? 4'b1000 : node1840;
														assign node1840 = (inp[10]) ? 4'b1000 : node1841;
															assign node1841 = (inp[8]) ? 4'b1000 : 4'b1010;
											assign node1847 = (inp[8]) ? node1861 : node1848;
												assign node1848 = (inp[1]) ? node1856 : node1849;
													assign node1849 = (inp[6]) ? 4'b1010 : node1850;
														assign node1850 = (inp[15]) ? 4'b1000 : node1851;
															assign node1851 = (inp[10]) ? 4'b1000 : 4'b1010;
													assign node1856 = (inp[6]) ? 4'b1000 : node1857;
														assign node1857 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node1861 = (inp[6]) ? node1865 : node1862;
													assign node1862 = (inp[1]) ? 4'b1010 : 4'b1000;
													assign node1865 = (inp[15]) ? 4'b1000 : node1866;
														assign node1866 = (inp[1]) ? 4'b1000 : 4'b1010;
										assign node1870 = (inp[1]) ? node1886 : node1871;
											assign node1871 = (inp[5]) ? node1877 : node1872;
												assign node1872 = (inp[15]) ? node1874 : 4'b1000;
													assign node1874 = (inp[6]) ? 4'b1000 : 4'b0010;
												assign node1877 = (inp[6]) ? 4'b0010 : node1878;
													assign node1878 = (inp[15]) ? node1880 : 4'b0010;
														assign node1880 = (inp[10]) ? node1882 : 4'b0010;
															assign node1882 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node1886 = (inp[5]) ? node1896 : node1887;
												assign node1887 = (inp[6]) ? 4'b1010 : node1888;
													assign node1888 = (inp[15]) ? 4'b1000 : node1889;
														assign node1889 = (inp[8]) ? node1891 : 4'b1010;
															assign node1891 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node1896 = (inp[6]) ? 4'b1000 : node1897;
													assign node1897 = (inp[15]) ? 4'b0010 : 4'b1000;
									assign node1901 = (inp[1]) ? node1961 : node1902;
										assign node1902 = (inp[5]) ? node1928 : node1903;
											assign node1903 = (inp[6]) ? node1925 : node1904;
												assign node1904 = (inp[11]) ? node1916 : node1905;
													assign node1905 = (inp[15]) ? node1911 : node1906;
														assign node1906 = (inp[8]) ? 4'b1001 : node1907;
															assign node1907 = (inp[10]) ? 4'b1001 : 4'b1011;
														assign node1911 = (inp[8]) ? node1913 : 4'b0011;
															assign node1913 = (inp[2]) ? 4'b0001 : 4'b0011;
													assign node1916 = (inp[8]) ? node1920 : node1917;
														assign node1917 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node1920 = (inp[15]) ? 4'b1010 : node1921;
															assign node1921 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node1925 = (inp[8]) ? 4'b1001 : 4'b1011;
											assign node1928 = (inp[6]) ? node1958 : node1929;
												assign node1929 = (inp[11]) ? node1947 : node1930;
													assign node1930 = (inp[10]) ? node1942 : node1931;
														assign node1931 = (inp[2]) ? node1937 : node1932;
															assign node1932 = (inp[15]) ? 4'b0011 : node1933;
																assign node1933 = (inp[8]) ? 4'b0011 : 4'b0001;
															assign node1937 = (inp[15]) ? node1939 : 4'b0011;
																assign node1939 = (inp[8]) ? 4'b0001 : 4'b0011;
														assign node1942 = (inp[15]) ? 4'b0001 : node1943;
															assign node1943 = (inp[8]) ? 4'b0011 : 4'b0001;
													assign node1947 = (inp[15]) ? node1953 : node1948;
														assign node1948 = (inp[10]) ? 4'b1000 : node1949;
															assign node1949 = (inp[8]) ? 4'b1000 : 4'b1010;
														assign node1953 = (inp[8]) ? node1955 : 4'b0010;
															assign node1955 = (inp[10]) ? 4'b0000 : 4'b0010;
												assign node1958 = (inp[8]) ? 4'b0001 : 4'b0011;
										assign node1961 = (inp[6]) ? 4'b0000 : node1962;
											assign node1962 = (inp[11]) ? node1970 : node1963;
												assign node1963 = (inp[15]) ? node1967 : node1964;
													assign node1964 = (inp[10]) ? 4'b1001 : 4'b1011;
													assign node1967 = (inp[10]) ? 4'b0001 : 4'b0011;
												assign node1970 = (inp[15]) ? node1974 : node1971;
													assign node1971 = (inp[10]) ? 4'b1000 : 4'b1010;
													assign node1974 = (inp[10]) ? 4'b0000 : 4'b0010;
					assign node1978 = (inp[3]) ? node1980 : 4'b0000;
						assign node1980 = (inp[11]) ? node2196 : node1981;
							assign node1981 = (inp[9]) ? node2071 : node1982;
								assign node1982 = (inp[7]) ? node2020 : node1983;
									assign node1983 = (inp[5]) ? 4'b0000 : node1984;
										assign node1984 = (inp[13]) ? node2002 : node1985;
											assign node1985 = (inp[15]) ? 4'b0000 : node1986;
												assign node1986 = (inp[1]) ? node1994 : node1987;
													assign node1987 = (inp[8]) ? 4'b0000 : node1988;
														assign node1988 = (inp[6]) ? 4'b0010 : node1989;
															assign node1989 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1994 = (inp[6]) ? 4'b0010 : node1995;
														assign node1995 = (inp[10]) ? node1997 : 4'b0010;
															assign node1997 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node2002 = (inp[15]) ? node2004 : 4'b0010;
												assign node2004 = (inp[1]) ? node2012 : node2005;
													assign node2005 = (inp[8]) ? 4'b0000 : node2006;
														assign node2006 = (inp[6]) ? 4'b0010 : node2007;
															assign node2007 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node2012 = (inp[6]) ? 4'b0010 : node2013;
														assign node2013 = (inp[10]) ? node2015 : 4'b0010;
															assign node2015 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node2020 = (inp[5]) ? node2054 : node2021;
										assign node2021 = (inp[15]) ? node2037 : node2022;
											assign node2022 = (inp[13]) ? node2030 : node2023;
												assign node2023 = (inp[6]) ? 4'b0000 : node2024;
													assign node2024 = (inp[1]) ? 4'b0000 : node2025;
														assign node2025 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node2030 = (inp[1]) ? 4'b0010 : node2031;
													assign node2031 = (inp[8]) ? 4'b0000 : node2032;
														assign node2032 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node2037 = (inp[13]) ? node2045 : node2038;
												assign node2038 = (inp[1]) ? node2040 : 4'b0010;
													assign node2040 = (inp[6]) ? 4'b0000 : node2041;
														assign node2041 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node2045 = (inp[1]) ? node2047 : 4'b0000;
													assign node2047 = (inp[6]) ? 4'b0010 : node2048;
														assign node2048 = (inp[8]) ? 4'b0000 : node2049;
															assign node2049 = (inp[10]) ? 4'b0000 : 4'b0010;
										assign node2054 = (inp[13]) ? node2056 : 4'b0010;
											assign node2056 = (inp[1]) ? node2064 : node2057;
												assign node2057 = (inp[15]) ? 4'b0010 : node2058;
													assign node2058 = (inp[8]) ? node2060 : 4'b0000;
														assign node2060 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node2064 = (inp[8]) ? node2066 : 4'b0000;
													assign node2066 = (inp[15]) ? node2068 : 4'b0000;
														assign node2068 = (inp[6]) ? 4'b0000 : 4'b0010;
								assign node2071 = (inp[7]) ? node2109 : node2072;
									assign node2072 = (inp[5]) ? node2074 : 4'b0010;
										assign node2074 = (inp[13]) ? node2092 : node2075;
											assign node2075 = (inp[15]) ? 4'b0000 : node2076;
												assign node2076 = (inp[1]) ? node2084 : node2077;
													assign node2077 = (inp[8]) ? 4'b0000 : node2078;
														assign node2078 = (inp[6]) ? 4'b0010 : node2079;
															assign node2079 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node2084 = (inp[8]) ? node2086 : 4'b0010;
														assign node2086 = (inp[10]) ? node2088 : 4'b0010;
															assign node2088 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node2092 = (inp[15]) ? node2094 : 4'b0010;
												assign node2094 = (inp[8]) ? node2102 : node2095;
													assign node2095 = (inp[10]) ? node2097 : 4'b0010;
														assign node2097 = (inp[1]) ? 4'b0010 : node2098;
															assign node2098 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node2102 = (inp[1]) ? node2104 : 4'b0000;
														assign node2104 = (inp[6]) ? 4'b0010 : node2105;
															assign node2105 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node2109 = (inp[13]) ? node2155 : node2110;
										assign node2110 = (inp[5]) ? node2134 : node2111;
											assign node2111 = (inp[1]) ? node2121 : node2112;
												assign node2112 = (inp[15]) ? node2118 : node2113;
													assign node2113 = (inp[8]) ? 4'b1000 : node2114;
														assign node2114 = (inp[6]) ? 4'b1010 : 4'b1000;
													assign node2118 = (inp[6]) ? 4'b1000 : 4'b0010;
												assign node2121 = (inp[15]) ? node2127 : node2122;
													assign node2122 = (inp[8]) ? 4'b1010 : node2123;
														assign node2123 = (inp[6]) ? 4'b1010 : 4'b1000;
													assign node2127 = (inp[6]) ? 4'b1000 : node2128;
														assign node2128 = (inp[10]) ? node2130 : 4'b1010;
															assign node2130 = (inp[8]) ? 4'b1000 : 4'b1010;
											assign node2134 = (inp[1]) ? node2148 : node2135;
												assign node2135 = (inp[15]) ? node2143 : node2136;
													assign node2136 = (inp[8]) ? node2138 : 4'b0010;
														assign node2138 = (inp[6]) ? 4'b0010 : node2139;
															assign node2139 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node2143 = (inp[8]) ? 4'b0000 : node2144;
														assign node2144 = (inp[6]) ? 4'b0010 : 4'b0000;
												assign node2148 = (inp[15]) ? node2152 : node2149;
													assign node2149 = (inp[6]) ? 4'b1010 : 4'b1000;
													assign node2152 = (inp[6]) ? 4'b1000 : 4'b0010;
										assign node2155 = (inp[6]) ? node2187 : node2156;
											assign node2156 = (inp[1]) ? node2180 : node2157;
												assign node2157 = (inp[5]) ? node2167 : node2158;
													assign node2158 = (inp[15]) ? node2162 : node2159;
														assign node2159 = (inp[8]) ? 4'b0010 : 4'b0000;
														assign node2162 = (inp[10]) ? 4'b0000 : node2163;
															assign node2163 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node2167 = (inp[10]) ? node2173 : node2168;
														assign node2168 = (inp[8]) ? 4'b1010 : node2169;
															assign node2169 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node2173 = (inp[2]) ? 4'b1000 : node2174;
															assign node2174 = (inp[15]) ? node2176 : 4'b1010;
																assign node2176 = (inp[8]) ? 4'b1010 : 4'b1000;
												assign node2180 = (inp[15]) ? node2184 : node2181;
													assign node2181 = (inp[10]) ? 4'b1001 : 4'b1011;
													assign node2184 = (inp[10]) ? 4'b0001 : 4'b0011;
											assign node2187 = (inp[1]) ? 4'b0000 : node2188;
												assign node2188 = (inp[5]) ? node2192 : node2189;
													assign node2189 = (inp[8]) ? 4'b1000 : 4'b1010;
													assign node2192 = (inp[8]) ? 4'b0000 : 4'b0010;
							assign node2196 = (inp[7]) ? node2198 : 4'b0000;
								assign node2198 = (inp[5]) ? node2280 : node2199;
									assign node2199 = (inp[13]) ? node2237 : node2200;
										assign node2200 = (inp[15]) ? node2228 : node2201;
											assign node2201 = (inp[1]) ? node2215 : node2202;
												assign node2202 = (inp[9]) ? node2210 : node2203;
													assign node2203 = (inp[8]) ? 4'b0000 : node2204;
														assign node2204 = (inp[6]) ? 4'b0010 : node2205;
															assign node2205 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node2210 = (inp[6]) ? 4'b0000 : node2211;
														assign node2211 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node2215 = (inp[6]) ? 4'b0010 : node2216;
													assign node2216 = (inp[9]) ? node2222 : node2217;
														assign node2217 = (inp[8]) ? node2219 : 4'b0010;
															assign node2219 = (inp[10]) ? 4'b0000 : 4'b0010;
														assign node2222 = (inp[8]) ? 4'b0000 : node2223;
															assign node2223 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node2228 = (inp[9]) ? node2230 : 4'b0000;
												assign node2230 = (inp[1]) ? node2232 : 4'b0010;
													assign node2232 = (inp[8]) ? node2234 : 4'b0000;
														assign node2234 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node2237 = (inp[9]) ? node2255 : node2238;
											assign node2238 = (inp[15]) ? node2240 : 4'b0010;
												assign node2240 = (inp[8]) ? node2248 : node2241;
													assign node2241 = (inp[6]) ? 4'b0010 : node2242;
														assign node2242 = (inp[1]) ? 4'b0010 : node2243;
															assign node2243 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node2248 = (inp[1]) ? node2250 : 4'b0000;
														assign node2250 = (inp[10]) ? node2252 : 4'b0010;
															assign node2252 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node2255 = (inp[1]) ? node2271 : node2256;
												assign node2256 = (inp[8]) ? node2264 : node2257;
													assign node2257 = (inp[6]) ? 4'b1010 : node2258;
														assign node2258 = (inp[15]) ? 4'b0010 : node2259;
															assign node2259 = (inp[10]) ? 4'b1000 : 4'b1010;
													assign node2264 = (inp[6]) ? 4'b1000 : node2265;
														assign node2265 = (inp[15]) ? node2267 : 4'b1000;
															assign node2267 = (inp[10]) ? 4'b0000 : 4'b0010;
												assign node2271 = (inp[6]) ? 4'b0000 : node2272;
													assign node2272 = (inp[10]) ? node2276 : node2273;
														assign node2273 = (inp[15]) ? 4'b0010 : 4'b1010;
														assign node2276 = (inp[15]) ? 4'b0000 : 4'b1000;
									assign node2280 = (inp[9]) ? node2282 : 4'b0000;
										assign node2282 = (inp[15]) ? node2312 : node2283;
											assign node2283 = (inp[13]) ? node2299 : node2284;
												assign node2284 = (inp[1]) ? node2292 : node2285;
													assign node2285 = (inp[8]) ? 4'b0000 : node2286;
														assign node2286 = (inp[10]) ? node2288 : 4'b0010;
															assign node2288 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node2292 = (inp[10]) ? node2294 : 4'b0010;
														assign node2294 = (inp[8]) ? node2296 : 4'b0010;
															assign node2296 = (inp[6]) ? 4'b0010 : 4'b0000;
												assign node2299 = (inp[6]) ? node2307 : node2300;
													assign node2300 = (inp[1]) ? node2304 : node2301;
														assign node2301 = (inp[8]) ? 4'b0010 : 4'b0000;
														assign node2304 = (inp[10]) ? 4'b1000 : 4'b1010;
													assign node2307 = (inp[8]) ? 4'b0000 : node2308;
														assign node2308 = (inp[1]) ? 4'b0000 : 4'b0010;
											assign node2312 = (inp[13]) ? node2314 : 4'b0000;
												assign node2314 = (inp[10]) ? node2326 : node2315;
													assign node2315 = (inp[8]) ? node2321 : node2316;
														assign node2316 = (inp[6]) ? node2318 : 4'b0010;
															assign node2318 = (inp[1]) ? 4'b0000 : 4'b0010;
														assign node2321 = (inp[1]) ? node2323 : 4'b0000;
															assign node2323 = (inp[6]) ? 4'b0000 : 4'b0010;
													assign node2326 = (inp[6]) ? node2328 : 4'b0000;
														assign node2328 = (inp[1]) ? 4'b0000 : node2329;
															assign node2329 = (inp[8]) ? 4'b0000 : 4'b0010;

endmodule