module dtc_split75_bm84 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node47;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node197;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node256;
	wire [3-1:0] node260;
	wire [3-1:0] node263;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node273;
	wire [3-1:0] node275;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node284;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node295;
	wire [3-1:0] node297;
	wire [3-1:0] node299;
	wire [3-1:0] node302;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node309;

	assign outp = (inp[9]) ? node234 : node1;
		assign node1 = (inp[6]) ? node147 : node2;
			assign node2 = (inp[10]) ? node54 : node3;
				assign node3 = (inp[7]) ? node11 : node4;
					assign node4 = (inp[3]) ? node6 : 3'b111;
						assign node6 = (inp[8]) ? node8 : 3'b111;
							assign node8 = (inp[11]) ? 3'b011 : 3'b111;
					assign node11 = (inp[11]) ? node27 : node12;
						assign node12 = (inp[3]) ? node20 : node13;
							assign node13 = (inp[8]) ? node15 : 3'b111;
								assign node15 = (inp[1]) ? node17 : 3'b111;
									assign node17 = (inp[2]) ? 3'b111 : 3'b011;
							assign node20 = (inp[8]) ? 3'b011 : node21;
								assign node21 = (inp[4]) ? node23 : 3'b111;
									assign node23 = (inp[5]) ? 3'b011 : 3'b111;
						assign node27 = (inp[3]) ? node37 : node28;
							assign node28 = (inp[2]) ? 3'b011 : node29;
								assign node29 = (inp[8]) ? node33 : node30;
									assign node30 = (inp[4]) ? 3'b011 : 3'b111;
									assign node33 = (inp[1]) ? 3'b001 : 3'b011;
							assign node37 = (inp[8]) ? node43 : node38;
								assign node38 = (inp[4]) ? node40 : 3'b011;
									assign node40 = (inp[5]) ? 3'b101 : 3'b111;
								assign node43 = (inp[2]) ? node45 : 3'b101;
									assign node45 = (inp[5]) ? node47 : 3'b101;
										assign node47 = (inp[4]) ? node49 : 3'b001;
											assign node49 = (inp[1]) ? node51 : 3'b101;
												assign node51 = (inp[0]) ? 3'b001 : 3'b101;
				assign node54 = (inp[11]) ? node116 : node55;
					assign node55 = (inp[8]) ? node79 : node56;
						assign node56 = (inp[3]) ? node66 : node57;
							assign node57 = (inp[4]) ? node63 : node58;
								assign node58 = (inp[2]) ? 3'b111 : node59;
									assign node59 = (inp[7]) ? 3'b011 : 3'b111;
								assign node63 = (inp[7]) ? 3'b101 : 3'b111;
							assign node66 = (inp[4]) ? node76 : node67;
								assign node67 = (inp[7]) ? 3'b111 : node68;
									assign node68 = (inp[1]) ? 3'b011 : node69;
										assign node69 = (inp[5]) ? 3'b011 : node70;
											assign node70 = (inp[2]) ? 3'b011 : 3'b111;
								assign node76 = (inp[7]) ? 3'b001 : 3'b011;
						assign node79 = (inp[3]) ? node97 : node80;
							assign node80 = (inp[7]) ? node82 : 3'b011;
								assign node82 = (inp[2]) ? node90 : node83;
									assign node83 = (inp[4]) ? 3'b001 : node84;
										assign node84 = (inp[0]) ? node86 : 3'b101;
											assign node86 = (inp[5]) ? 3'b110 : 3'b101;
									assign node90 = (inp[5]) ? node92 : 3'b001;
										assign node92 = (inp[1]) ? node94 : 3'b001;
											assign node94 = (inp[0]) ? 3'b010 : 3'b001;
							assign node97 = (inp[4]) ? node107 : node98;
								assign node98 = (inp[7]) ? node100 : 3'b001;
									assign node100 = (inp[1]) ? node102 : 3'b001;
										assign node102 = (inp[5]) ? node104 : 3'b001;
											assign node104 = (inp[0]) ? 3'b110 : 3'b001;
								assign node107 = (inp[7]) ? node109 : 3'b101;
									assign node109 = (inp[1]) ? node111 : 3'b001;
										assign node111 = (inp[5]) ? node113 : 3'b001;
											assign node113 = (inp[0]) ? 3'b110 : 3'b001;
					assign node116 = (inp[7]) ? node126 : node117;
						assign node117 = (inp[3]) ? node121 : node118;
							assign node118 = (inp[8]) ? 3'b101 : 3'b011;
							assign node121 = (inp[8]) ? node123 : 3'b101;
								assign node123 = (inp[4]) ? 3'b001 : 3'b101;
						assign node126 = (inp[8]) ? node134 : node127;
							assign node127 = (inp[5]) ? node129 : 3'b101;
								assign node129 = (inp[4]) ? node131 : 3'b101;
									assign node131 = (inp[3]) ? 3'b110 : 3'b101;
							assign node134 = (inp[3]) ? node140 : node135;
								assign node135 = (inp[1]) ? node137 : 3'b101;
									assign node137 = (inp[2]) ? 3'b101 : 3'b110;
								assign node140 = (inp[5]) ? node142 : 3'b110;
									assign node142 = (inp[4]) ? node144 : 3'b110;
										assign node144 = (inp[0]) ? 3'b010 : 3'b110;
			assign node147 = (inp[10]) ? node213 : node148;
				assign node148 = (inp[11]) ? node194 : node149;
					assign node149 = (inp[7]) ? node173 : node150;
						assign node150 = (inp[4]) ? node162 : node151;
							assign node151 = (inp[8]) ? node153 : 3'b011;
								assign node153 = (inp[5]) ? node155 : 3'b011;
									assign node155 = (inp[2]) ? 3'b001 : node156;
										assign node156 = (inp[1]) ? 3'b001 : node157;
											assign node157 = (inp[3]) ? 3'b001 : 3'b101;
							assign node162 = (inp[3]) ? node170 : node163;
								assign node163 = (inp[8]) ? node165 : 3'b011;
									assign node165 = (inp[1]) ? 3'b001 : node166;
										assign node166 = (inp[2]) ? 3'b001 : 3'b101;
								assign node170 = (inp[8]) ? 3'b001 : 3'b101;
						assign node173 = (inp[8]) ? node183 : node174;
							assign node174 = (inp[3]) ? node180 : node175;
								assign node175 = (inp[4]) ? 3'b001 : node176;
									assign node176 = (inp[2]) ? 3'b001 : 3'b101;
								assign node180 = (inp[4]) ? 3'b110 : 3'b001;
							assign node183 = (inp[3]) ? node187 : node184;
								assign node184 = (inp[4]) ? 3'b110 : 3'b001;
								assign node187 = (inp[5]) ? node189 : 3'b110;
									assign node189 = (inp[4]) ? node191 : 3'b110;
										assign node191 = (inp[0]) ? 3'b010 : 3'b110;
					assign node194 = (inp[8]) ? node202 : node195;
						assign node195 = (inp[7]) ? node197 : 3'b001;
							assign node197 = (inp[3]) ? node199 : 3'b110;
								assign node199 = (inp[4]) ? 3'b010 : 3'b110;
						assign node202 = (inp[7]) ? node204 : 3'b110;
							assign node204 = (inp[5]) ? node206 : 3'b010;
								assign node206 = (inp[4]) ? node208 : 3'b010;
									assign node208 = (inp[3]) ? node210 : 3'b010;
										assign node210 = (inp[0]) ? 3'b100 : 3'b010;
				assign node213 = (inp[7]) ? node221 : node214;
					assign node214 = (inp[8]) ? node218 : node215;
						assign node215 = (inp[11]) ? 3'b010 : 3'b110;
						assign node218 = (inp[11]) ? 3'b100 : 3'b010;
					assign node221 = (inp[11]) ? 3'b000 : node222;
						assign node222 = (inp[5]) ? node224 : 3'b100;
							assign node224 = (inp[0]) ? node226 : 3'b100;
								assign node226 = (inp[8]) ? node228 : 3'b100;
									assign node228 = (inp[3]) ? node230 : 3'b100;
										assign node230 = (inp[4]) ? 3'b000 : 3'b100;
		assign node234 = (inp[6]) ? node306 : node235;
			assign node235 = (inp[10]) ? node291 : node236;
				assign node236 = (inp[8]) ? node266 : node237;
					assign node237 = (inp[7]) ? node263 : node238;
						assign node238 = (inp[4]) ? node250 : node239;
							assign node239 = (inp[11]) ? 3'b001 : node240;
								assign node240 = (inp[3]) ? node242 : 3'b101;
									assign node242 = (inp[2]) ? 3'b001 : node243;
										assign node243 = (inp[5]) ? node245 : 3'b101;
											assign node245 = (inp[0]) ? 3'b001 : 3'b101;
							assign node250 = (inp[11]) ? node260 : node251;
								assign node251 = (inp[3]) ? node253 : 3'b101;
									assign node253 = (inp[2]) ? 3'b001 : node254;
										assign node254 = (inp[5]) ? node256 : 3'b101;
											assign node256 = (inp[0]) ? 3'b001 : 3'b101;
								assign node260 = (inp[3]) ? 3'b110 : 3'b101;
						assign node263 = (inp[11]) ? 3'b100 : 3'b010;
					assign node266 = (inp[7]) ? node278 : node267;
						assign node267 = (inp[11]) ? node269 : 3'b000;
							assign node269 = (inp[5]) ? node271 : 3'b010;
								assign node271 = (inp[4]) ? node273 : 3'b010;
									assign node273 = (inp[0]) ? node275 : 3'b010;
										assign node275 = (inp[3]) ? 3'b101 : 3'b110;
						assign node278 = (inp[11]) ? node288 : node279;
							assign node279 = (inp[3]) ? node281 : 3'b010;
								assign node281 = (inp[2]) ? 3'b100 : node282;
									assign node282 = (inp[5]) ? node284 : 3'b010;
										assign node284 = (inp[0]) ? 3'b100 : 3'b010;
							assign node288 = (inp[4]) ? 3'b000 : 3'b100;
				assign node291 = (inp[7]) ? 3'b000 : node292;
					assign node292 = (inp[8]) ? node302 : node293;
						assign node293 = (inp[11]) ? node295 : 3'b010;
							assign node295 = (inp[0]) ? node297 : 3'b100;
								assign node297 = (inp[5]) ? node299 : 3'b100;
									assign node299 = (inp[4]) ? 3'b000 : 3'b100;
						assign node302 = (inp[11]) ? 3'b000 : 3'b100;
			assign node306 = (inp[8]) ? 3'b000 : node307;
				assign node307 = (inp[10]) ? 3'b000 : node308;
					assign node308 = (inp[11]) ? 3'b000 : node309;
						assign node309 = (inp[7]) ? 3'b000 : 3'b100;

endmodule