module dtc_split125_bm30 (
	input  wire [14-1:0] inp,
	output wire [8-1:0] outp
);

	wire [8-1:0] node1;
	wire [8-1:0] node2;
	wire [8-1:0] node3;
	wire [8-1:0] node4;
	wire [8-1:0] node5;
	wire [8-1:0] node6;
	wire [8-1:0] node7;
	wire [8-1:0] node9;
	wire [8-1:0] node11;
	wire [8-1:0] node14;
	wire [8-1:0] node15;
	wire [8-1:0] node18;
	wire [8-1:0] node19;
	wire [8-1:0] node21;
	wire [8-1:0] node25;
	wire [8-1:0] node26;
	wire [8-1:0] node28;
	wire [8-1:0] node30;
	wire [8-1:0] node31;
	wire [8-1:0] node34;
	wire [8-1:0] node37;
	wire [8-1:0] node39;
	wire [8-1:0] node41;
	wire [8-1:0] node43;
	wire [8-1:0] node44;
	wire [8-1:0] node48;
	wire [8-1:0] node49;
	wire [8-1:0] node50;
	wire [8-1:0] node51;
	wire [8-1:0] node53;
	wire [8-1:0] node56;
	wire [8-1:0] node58;
	wire [8-1:0] node60;
	wire [8-1:0] node63;
	wire [8-1:0] node64;
	wire [8-1:0] node66;
	wire [8-1:0] node68;
	wire [8-1:0] node71;
	wire [8-1:0] node72;
	wire [8-1:0] node75;
	wire [8-1:0] node79;
	wire [8-1:0] node80;
	wire [8-1:0] node81;
	wire [8-1:0] node82;
	wire [8-1:0] node85;
	wire [8-1:0] node86;
	wire [8-1:0] node87;
	wire [8-1:0] node88;
	wire [8-1:0] node93;
	wire [8-1:0] node94;
	wire [8-1:0] node96;
	wire [8-1:0] node99;
	wire [8-1:0] node100;
	wire [8-1:0] node104;
	wire [8-1:0] node105;
	wire [8-1:0] node107;
	wire [8-1:0] node110;
	wire [8-1:0] node111;
	wire [8-1:0] node112;
	wire [8-1:0] node115;
	wire [8-1:0] node116;
	wire [8-1:0] node120;
	wire [8-1:0] node121;
	wire [8-1:0] node122;
	wire [8-1:0] node126;
	wire [8-1:0] node129;
	wire [8-1:0] node130;
	wire [8-1:0] node131;
	wire [8-1:0] node132;
	wire [8-1:0] node133;
	wire [8-1:0] node136;
	wire [8-1:0] node138;
	wire [8-1:0] node139;
	wire [8-1:0] node143;
	wire [8-1:0] node144;
	wire [8-1:0] node146;
	wire [8-1:0] node149;
	wire [8-1:0] node152;
	wire [8-1:0] node153;
	wire [8-1:0] node154;
	wire [8-1:0] node156;
	wire [8-1:0] node160;
	wire [8-1:0] node161;
	wire [8-1:0] node162;
	wire [8-1:0] node166;
	wire [8-1:0] node167;
	wire [8-1:0] node170;
	wire [8-1:0] node171;
	wire [8-1:0] node175;
	wire [8-1:0] node176;
	wire [8-1:0] node177;
	wire [8-1:0] node178;
	wire [8-1:0] node179;
	wire [8-1:0] node183;
	wire [8-1:0] node186;
	wire [8-1:0] node189;
	wire [8-1:0] node190;
	wire [8-1:0] node191;
	wire [8-1:0] node193;
	wire [8-1:0] node194;
	wire [8-1:0] node197;
	wire [8-1:0] node200;
	wire [8-1:0] node201;
	wire [8-1:0] node202;
	wire [8-1:0] node203;
	wire [8-1:0] node209;
	wire [8-1:0] node210;
	wire [8-1:0] node211;
	wire [8-1:0] node212;
	wire [8-1:0] node215;
	wire [8-1:0] node217;
	wire [8-1:0] node221;
	wire [8-1:0] node224;
	wire [8-1:0] node225;
	wire [8-1:0] node226;
	wire [8-1:0] node227;
	wire [8-1:0] node228;
	wire [8-1:0] node229;
	wire [8-1:0] node230;
	wire [8-1:0] node231;
	wire [8-1:0] node234;
	wire [8-1:0] node237;
	wire [8-1:0] node240;
	wire [8-1:0] node242;
	wire [8-1:0] node244;
	wire [8-1:0] node247;
	wire [8-1:0] node248;
	wire [8-1:0] node250;
	wire [8-1:0] node252;
	wire [8-1:0] node255;
	wire [8-1:0] node256;
	wire [8-1:0] node259;
	wire [8-1:0] node262;
	wire [8-1:0] node263;
	wire [8-1:0] node264;
	wire [8-1:0] node265;
	wire [8-1:0] node266;
	wire [8-1:0] node268;
	wire [8-1:0] node271;
	wire [8-1:0] node273;
	wire [8-1:0] node277;
	wire [8-1:0] node278;
	wire [8-1:0] node282;
	wire [8-1:0] node283;
	wire [8-1:0] node284;
	wire [8-1:0] node285;
	wire [8-1:0] node290;
	wire [8-1:0] node291;
	wire [8-1:0] node292;
	wire [8-1:0] node294;
	wire [8-1:0] node295;
	wire [8-1:0] node300;
	wire [8-1:0] node303;
	wire [8-1:0] node304;
	wire [8-1:0] node305;
	wire [8-1:0] node306;
	wire [8-1:0] node309;
	wire [8-1:0] node310;
	wire [8-1:0] node313;
	wire [8-1:0] node315;
	wire [8-1:0] node317;
	wire [8-1:0] node320;
	wire [8-1:0] node321;
	wire [8-1:0] node322;
	wire [8-1:0] node323;
	wire [8-1:0] node326;
	wire [8-1:0] node329;
	wire [8-1:0] node332;
	wire [8-1:0] node333;
	wire [8-1:0] node334;
	wire [8-1:0] node337;
	wire [8-1:0] node340;
	wire [8-1:0] node341;
	wire [8-1:0] node343;
	wire [8-1:0] node347;
	wire [8-1:0] node348;
	wire [8-1:0] node349;
	wire [8-1:0] node350;
	wire [8-1:0] node351;
	wire [8-1:0] node354;
	wire [8-1:0] node357;
	wire [8-1:0] node358;
	wire [8-1:0] node361;
	wire [8-1:0] node364;
	wire [8-1:0] node365;
	wire [8-1:0] node366;
	wire [8-1:0] node368;
	wire [8-1:0] node373;
	wire [8-1:0] node374;
	wire [8-1:0] node375;
	wire [8-1:0] node376;
	wire [8-1:0] node380;
	wire [8-1:0] node382;
	wire [8-1:0] node385;
	wire [8-1:0] node387;
	wire [8-1:0] node388;
	wire [8-1:0] node389;
	wire [8-1:0] node391;
	wire [8-1:0] node395;
	wire [8-1:0] node398;
	wire [8-1:0] node399;
	wire [8-1:0] node400;
	wire [8-1:0] node401;
	wire [8-1:0] node402;
	wire [8-1:0] node404;
	wire [8-1:0] node407;
	wire [8-1:0] node408;
	wire [8-1:0] node409;
	wire [8-1:0] node411;
	wire [8-1:0] node415;
	wire [8-1:0] node418;
	wire [8-1:0] node419;
	wire [8-1:0] node420;
	wire [8-1:0] node421;
	wire [8-1:0] node424;
	wire [8-1:0] node427;
	wire [8-1:0] node430;
	wire [8-1:0] node431;
	wire [8-1:0] node434;
	wire [8-1:0] node436;
	wire [8-1:0] node438;
	wire [8-1:0] node441;
	wire [8-1:0] node442;
	wire [8-1:0] node443;
	wire [8-1:0] node444;
	wire [8-1:0] node445;
	wire [8-1:0] node448;
	wire [8-1:0] node451;
	wire [8-1:0] node454;
	wire [8-1:0] node455;
	wire [8-1:0] node457;
	wire [8-1:0] node461;
	wire [8-1:0] node462;
	wire [8-1:0] node463;
	wire [8-1:0] node466;
	wire [8-1:0] node469;
	wire [8-1:0] node470;
	wire [8-1:0] node472;
	wire [8-1:0] node473;
	wire [8-1:0] node476;
	wire [8-1:0] node479;
	wire [8-1:0] node480;
	wire [8-1:0] node481;
	wire [8-1:0] node484;
	wire [8-1:0] node488;
	wire [8-1:0] node489;
	wire [8-1:0] node490;
	wire [8-1:0] node491;
	wire [8-1:0] node492;
	wire [8-1:0] node494;
	wire [8-1:0] node497;
	wire [8-1:0] node500;
	wire [8-1:0] node501;
	wire [8-1:0] node504;
	wire [8-1:0] node507;
	wire [8-1:0] node508;
	wire [8-1:0] node510;
	wire [8-1:0] node511;
	wire [8-1:0] node512;
	wire [8-1:0] node517;
	wire [8-1:0] node518;
	wire [8-1:0] node520;
	wire [8-1:0] node523;
	wire [8-1:0] node524;
	wire [8-1:0] node528;
	wire [8-1:0] node529;
	wire [8-1:0] node530;
	wire [8-1:0] node532;
	wire [8-1:0] node533;
	wire [8-1:0] node534;
	wire [8-1:0] node538;
	wire [8-1:0] node541;
	wire [8-1:0] node542;
	wire [8-1:0] node545;
	wire [8-1:0] node547;
	wire [8-1:0] node550;
	wire [8-1:0] node551;
	wire [8-1:0] node552;
	wire [8-1:0] node553;
	wire [8-1:0] node557;
	wire [8-1:0] node560;
	wire [8-1:0] node561;
	wire [8-1:0] node563;
	wire [8-1:0] node566;
	wire [8-1:0] node567;
	wire [8-1:0] node570;
	wire [8-1:0] node573;
	wire [8-1:0] node574;
	wire [8-1:0] node575;
	wire [8-1:0] node576;
	wire [8-1:0] node577;
	wire [8-1:0] node578;
	wire [8-1:0] node579;
	wire [8-1:0] node580;
	wire [8-1:0] node584;
	wire [8-1:0] node586;
	wire [8-1:0] node589;
	wire [8-1:0] node590;
	wire [8-1:0] node591;
	wire [8-1:0] node596;
	wire [8-1:0] node597;
	wire [8-1:0] node598;
	wire [8-1:0] node599;
	wire [8-1:0] node600;
	wire [8-1:0] node603;
	wire [8-1:0] node605;
	wire [8-1:0] node609;
	wire [8-1:0] node612;
	wire [8-1:0] node613;
	wire [8-1:0] node615;
	wire [8-1:0] node616;
	wire [8-1:0] node620;
	wire [8-1:0] node623;
	wire [8-1:0] node624;
	wire [8-1:0] node625;
	wire [8-1:0] node626;
	wire [8-1:0] node627;
	wire [8-1:0] node628;
	wire [8-1:0] node633;
	wire [8-1:0] node634;
	wire [8-1:0] node637;
	wire [8-1:0] node640;
	wire [8-1:0] node641;
	wire [8-1:0] node642;
	wire [8-1:0] node643;
	wire [8-1:0] node648;
	wire [8-1:0] node649;
	wire [8-1:0] node651;
	wire [8-1:0] node655;
	wire [8-1:0] node656;
	wire [8-1:0] node657;
	wire [8-1:0] node658;
	wire [8-1:0] node662;
	wire [8-1:0] node663;
	wire [8-1:0] node666;
	wire [8-1:0] node669;
	wire [8-1:0] node670;
	wire [8-1:0] node674;
	wire [8-1:0] node675;
	wire [8-1:0] node676;
	wire [8-1:0] node677;
	wire [8-1:0] node678;
	wire [8-1:0] node680;
	wire [8-1:0] node682;
	wire [8-1:0] node683;
	wire [8-1:0] node687;
	wire [8-1:0] node688;
	wire [8-1:0] node690;
	wire [8-1:0] node693;
	wire [8-1:0] node696;
	wire [8-1:0] node697;
	wire [8-1:0] node698;
	wire [8-1:0] node700;
	wire [8-1:0] node703;
	wire [8-1:0] node704;
	wire [8-1:0] node708;
	wire [8-1:0] node710;
	wire [8-1:0] node713;
	wire [8-1:0] node714;
	wire [8-1:0] node715;
	wire [8-1:0] node716;
	wire [8-1:0] node719;
	wire [8-1:0] node722;
	wire [8-1:0] node723;
	wire [8-1:0] node724;
	wire [8-1:0] node725;
	wire [8-1:0] node729;
	wire [8-1:0] node732;
	wire [8-1:0] node733;
	wire [8-1:0] node734;
	wire [8-1:0] node739;
	wire [8-1:0] node740;
	wire [8-1:0] node741;
	wire [8-1:0] node742;
	wire [8-1:0] node745;
	wire [8-1:0] node748;
	wire [8-1:0] node750;
	wire [8-1:0] node753;
	wire [8-1:0] node754;
	wire [8-1:0] node757;
	wire [8-1:0] node760;
	wire [8-1:0] node761;
	wire [8-1:0] node762;
	wire [8-1:0] node763;
	wire [8-1:0] node764;
	wire [8-1:0] node765;
	wire [8-1:0] node769;
	wire [8-1:0] node771;
	wire [8-1:0] node774;
	wire [8-1:0] node775;
	wire [8-1:0] node776;
	wire [8-1:0] node779;
	wire [8-1:0] node782;
	wire [8-1:0] node783;
	wire [8-1:0] node787;
	wire [8-1:0] node788;
	wire [8-1:0] node789;
	wire [8-1:0] node790;
	wire [8-1:0] node792;
	wire [8-1:0] node797;
	wire [8-1:0] node798;
	wire [8-1:0] node800;
	wire [8-1:0] node801;
	wire [8-1:0] node805;
	wire [8-1:0] node807;
	wire [8-1:0] node810;
	wire [8-1:0] node811;
	wire [8-1:0] node812;
	wire [8-1:0] node813;
	wire [8-1:0] node814;
	wire [8-1:0] node817;
	wire [8-1:0] node820;
	wire [8-1:0] node822;
	wire [8-1:0] node823;
	wire [8-1:0] node827;
	wire [8-1:0] node828;
	wire [8-1:0] node829;
	wire [8-1:0] node830;
	wire [8-1:0] node834;
	wire [8-1:0] node837;
	wire [8-1:0] node838;
	wire [8-1:0] node842;
	wire [8-1:0] node843;
	wire [8-1:0] node844;
	wire [8-1:0] node847;
	wire [8-1:0] node850;
	wire [8-1:0] node851;
	wire [8-1:0] node852;
	wire [8-1:0] node856;
	wire [8-1:0] node857;
	wire [8-1:0] node859;
	wire [8-1:0] node862;
	wire [8-1:0] node865;
	wire [8-1:0] node866;
	wire [8-1:0] node867;
	wire [8-1:0] node868;
	wire [8-1:0] node869;
	wire [8-1:0] node870;
	wire [8-1:0] node871;
	wire [8-1:0] node872;
	wire [8-1:0] node875;
	wire [8-1:0] node878;
	wire [8-1:0] node880;
	wire [8-1:0] node881;
	wire [8-1:0] node885;
	wire [8-1:0] node886;
	wire [8-1:0] node887;
	wire [8-1:0] node890;
	wire [8-1:0] node893;
	wire [8-1:0] node896;
	wire [8-1:0] node897;
	wire [8-1:0] node898;
	wire [8-1:0] node901;
	wire [8-1:0] node902;
	wire [8-1:0] node905;
	wire [8-1:0] node908;
	wire [8-1:0] node910;
	wire [8-1:0] node912;
	wire [8-1:0] node915;
	wire [8-1:0] node916;
	wire [8-1:0] node917;
	wire [8-1:0] node918;
	wire [8-1:0] node919;
	wire [8-1:0] node923;
	wire [8-1:0] node926;
	wire [8-1:0] node928;
	wire [8-1:0] node930;
	wire [8-1:0] node933;
	wire [8-1:0] node934;
	wire [8-1:0] node935;
	wire [8-1:0] node936;
	wire [8-1:0] node940;
	wire [8-1:0] node942;
	wire [8-1:0] node943;
	wire [8-1:0] node944;
	wire [8-1:0] node949;
	wire [8-1:0] node950;
	wire [8-1:0] node951;
	wire [8-1:0] node954;
	wire [8-1:0] node957;
	wire [8-1:0] node958;
	wire [8-1:0] node959;
	wire [8-1:0] node963;
	wire [8-1:0] node966;
	wire [8-1:0] node967;
	wire [8-1:0] node969;
	wire [8-1:0] node970;
	wire [8-1:0] node971;
	wire [8-1:0] node976;
	wire [8-1:0] node977;
	wire [8-1:0] node978;
	wire [8-1:0] node980;
	wire [8-1:0] node983;
	wire [8-1:0] node985;
	wire [8-1:0] node988;
	wire [8-1:0] node989;
	wire [8-1:0] node990;
	wire [8-1:0] node991;
	wire [8-1:0] node994;
	wire [8-1:0] node997;
	wire [8-1:0] node999;
	wire [8-1:0] node1001;
	wire [8-1:0] node1004;
	wire [8-1:0] node1005;
	wire [8-1:0] node1007;
	wire [8-1:0] node1010;
	wire [8-1:0] node1011;
	wire [8-1:0] node1015;
	wire [8-1:0] node1016;
	wire [8-1:0] node1017;
	wire [8-1:0] node1018;
	wire [8-1:0] node1019;
	wire [8-1:0] node1020;
	wire [8-1:0] node1021;
	wire [8-1:0] node1024;
	wire [8-1:0] node1027;
	wire [8-1:0] node1030;
	wire [8-1:0] node1031;
	wire [8-1:0] node1032;
	wire [8-1:0] node1036;
	wire [8-1:0] node1038;
	wire [8-1:0] node1041;
	wire [8-1:0] node1042;
	wire [8-1:0] node1043;
	wire [8-1:0] node1045;
	wire [8-1:0] node1048;
	wire [8-1:0] node1051;
	wire [8-1:0] node1053;
	wire [8-1:0] node1056;
	wire [8-1:0] node1057;
	wire [8-1:0] node1058;
	wire [8-1:0] node1059;
	wire [8-1:0] node1060;
	wire [8-1:0] node1064;
	wire [8-1:0] node1067;
	wire [8-1:0] node1068;
	wire [8-1:0] node1071;
	wire [8-1:0] node1072;
	wire [8-1:0] node1073;
	wire [8-1:0] node1076;
	wire [8-1:0] node1080;
	wire [8-1:0] node1081;
	wire [8-1:0] node1082;
	wire [8-1:0] node1084;
	wire [8-1:0] node1086;
	wire [8-1:0] node1089;
	wire [8-1:0] node1090;
	wire [8-1:0] node1091;
	wire [8-1:0] node1096;
	wire [8-1:0] node1097;
	wire [8-1:0] node1098;
	wire [8-1:0] node1101;
	wire [8-1:0] node1103;
	wire [8-1:0] node1106;
	wire [8-1:0] node1107;
	wire [8-1:0] node1111;
	wire [8-1:0] node1112;
	wire [8-1:0] node1113;
	wire [8-1:0] node1114;
	wire [8-1:0] node1116;
	wire [8-1:0] node1117;
	wire [8-1:0] node1118;
	wire [8-1:0] node1123;
	wire [8-1:0] node1124;
	wire [8-1:0] node1127;
	wire [8-1:0] node1130;
	wire [8-1:0] node1131;
	wire [8-1:0] node1132;
	wire [8-1:0] node1133;
	wire [8-1:0] node1136;
	wire [8-1:0] node1138;
	wire [8-1:0] node1141;
	wire [8-1:0] node1144;
	wire [8-1:0] node1145;
	wire [8-1:0] node1146;
	wire [8-1:0] node1149;
	wire [8-1:0] node1152;
	wire [8-1:0] node1153;
	wire [8-1:0] node1157;
	wire [8-1:0] node1158;
	wire [8-1:0] node1159;
	wire [8-1:0] node1160;
	wire [8-1:0] node1164;
	wire [8-1:0] node1165;
	wire [8-1:0] node1167;
	wire [8-1:0] node1168;
	wire [8-1:0] node1172;
	wire [8-1:0] node1173;
	wire [8-1:0] node1176;
	wire [8-1:0] node1179;
	wire [8-1:0] node1180;
	wire [8-1:0] node1181;
	wire [8-1:0] node1184;
	wire [8-1:0] node1185;
	wire [8-1:0] node1188;
	wire [8-1:0] node1189;
	wire [8-1:0] node1192;
	wire [8-1:0] node1195;
	wire [8-1:0] node1198;
	wire [8-1:0] node1199;
	wire [8-1:0] node1200;
	wire [8-1:0] node1201;
	wire [8-1:0] node1202;
	wire [8-1:0] node1203;
	wire [8-1:0] node1204;
	wire [8-1:0] node1205;
	wire [8-1:0] node1206;
	wire [8-1:0] node1209;
	wire [8-1:0] node1210;
	wire [8-1:0] node1213;
	wire [8-1:0] node1216;
	wire [8-1:0] node1217;
	wire [8-1:0] node1219;
	wire [8-1:0] node1220;
	wire [8-1:0] node1224;
	wire [8-1:0] node1225;
	wire [8-1:0] node1228;
	wire [8-1:0] node1231;
	wire [8-1:0] node1232;
	wire [8-1:0] node1234;
	wire [8-1:0] node1236;
	wire [8-1:0] node1239;
	wire [8-1:0] node1240;
	wire [8-1:0] node1242;
	wire [8-1:0] node1245;
	wire [8-1:0] node1248;
	wire [8-1:0] node1249;
	wire [8-1:0] node1250;
	wire [8-1:0] node1251;
	wire [8-1:0] node1255;
	wire [8-1:0] node1258;
	wire [8-1:0] node1259;
	wire [8-1:0] node1261;
	wire [8-1:0] node1263;
	wire [8-1:0] node1266;
	wire [8-1:0] node1267;
	wire [8-1:0] node1268;
	wire [8-1:0] node1269;
	wire [8-1:0] node1272;
	wire [8-1:0] node1273;
	wire [8-1:0] node1278;
	wire [8-1:0] node1279;
	wire [8-1:0] node1281;
	wire [8-1:0] node1284;
	wire [8-1:0] node1287;
	wire [8-1:0] node1288;
	wire [8-1:0] node1289;
	wire [8-1:0] node1290;
	wire [8-1:0] node1291;
	wire [8-1:0] node1293;
	wire [8-1:0] node1296;
	wire [8-1:0] node1299;
	wire [8-1:0] node1301;
	wire [8-1:0] node1302;
	wire [8-1:0] node1306;
	wire [8-1:0] node1307;
	wire [8-1:0] node1308;
	wire [8-1:0] node1310;
	wire [8-1:0] node1314;
	wire [8-1:0] node1317;
	wire [8-1:0] node1318;
	wire [8-1:0] node1319;
	wire [8-1:0] node1321;
	wire [8-1:0] node1323;
	wire [8-1:0] node1326;
	wire [8-1:0] node1327;
	wire [8-1:0] node1328;
	wire [8-1:0] node1332;
	wire [8-1:0] node1333;
	wire [8-1:0] node1334;
	wire [8-1:0] node1335;
	wire [8-1:0] node1340;
	wire [8-1:0] node1343;
	wire [8-1:0] node1344;
	wire [8-1:0] node1345;
	wire [8-1:0] node1346;
	wire [8-1:0] node1349;
	wire [8-1:0] node1352;
	wire [8-1:0] node1354;
	wire [8-1:0] node1356;
	wire [8-1:0] node1359;
	wire [8-1:0] node1360;
	wire [8-1:0] node1361;
	wire [8-1:0] node1363;
	wire [8-1:0] node1365;
	wire [8-1:0] node1368;
	wire [8-1:0] node1372;
	wire [8-1:0] node1373;
	wire [8-1:0] node1374;
	wire [8-1:0] node1375;
	wire [8-1:0] node1376;
	wire [8-1:0] node1378;
	wire [8-1:0] node1380;
	wire [8-1:0] node1383;
	wire [8-1:0] node1384;
	wire [8-1:0] node1387;
	wire [8-1:0] node1390;
	wire [8-1:0] node1391;
	wire [8-1:0] node1392;
	wire [8-1:0] node1395;
	wire [8-1:0] node1397;
	wire [8-1:0] node1398;
	wire [8-1:0] node1402;
	wire [8-1:0] node1404;
	wire [8-1:0] node1407;
	wire [8-1:0] node1408;
	wire [8-1:0] node1409;
	wire [8-1:0] node1411;
	wire [8-1:0] node1412;
	wire [8-1:0] node1413;
	wire [8-1:0] node1416;
	wire [8-1:0] node1419;
	wire [8-1:0] node1421;
	wire [8-1:0] node1424;
	wire [8-1:0] node1425;
	wire [8-1:0] node1426;
	wire [8-1:0] node1430;
	wire [8-1:0] node1432;
	wire [8-1:0] node1434;
	wire [8-1:0] node1437;
	wire [8-1:0] node1438;
	wire [8-1:0] node1441;
	wire [8-1:0] node1442;
	wire [8-1:0] node1444;
	wire [8-1:0] node1448;
	wire [8-1:0] node1449;
	wire [8-1:0] node1450;
	wire [8-1:0] node1451;
	wire [8-1:0] node1452;
	wire [8-1:0] node1454;
	wire [8-1:0] node1457;
	wire [8-1:0] node1459;
	wire [8-1:0] node1460;
	wire [8-1:0] node1463;
	wire [8-1:0] node1466;
	wire [8-1:0] node1467;
	wire [8-1:0] node1470;
	wire [8-1:0] node1473;
	wire [8-1:0] node1474;
	wire [8-1:0] node1475;
	wire [8-1:0] node1478;
	wire [8-1:0] node1479;
	wire [8-1:0] node1481;
	wire [8-1:0] node1485;
	wire [8-1:0] node1486;
	wire [8-1:0] node1489;
	wire [8-1:0] node1492;
	wire [8-1:0] node1493;
	wire [8-1:0] node1494;
	wire [8-1:0] node1495;
	wire [8-1:0] node1496;
	wire [8-1:0] node1499;
	wire [8-1:0] node1502;
	wire [8-1:0] node1503;
	wire [8-1:0] node1506;
	wire [8-1:0] node1508;
	wire [8-1:0] node1511;
	wire [8-1:0] node1513;
	wire [8-1:0] node1514;
	wire [8-1:0] node1515;
	wire [8-1:0] node1520;
	wire [8-1:0] node1521;
	wire [8-1:0] node1522;
	wire [8-1:0] node1525;
	wire [8-1:0] node1527;
	wire [8-1:0] node1530;
	wire [8-1:0] node1531;
	wire [8-1:0] node1532;
	wire [8-1:0] node1535;
	wire [8-1:0] node1538;
	wire [8-1:0] node1539;
	wire [8-1:0] node1541;
	wire [8-1:0] node1544;
	wire [8-1:0] node1546;
	wire [8-1:0] node1549;
	wire [8-1:0] node1550;
	wire [8-1:0] node1551;
	wire [8-1:0] node1552;
	wire [8-1:0] node1553;
	wire [8-1:0] node1554;
	wire [8-1:0] node1555;
	wire [8-1:0] node1558;
	wire [8-1:0] node1561;
	wire [8-1:0] node1562;
	wire [8-1:0] node1565;
	wire [8-1:0] node1568;
	wire [8-1:0] node1569;
	wire [8-1:0] node1570;
	wire [8-1:0] node1571;
	wire [8-1:0] node1572;
	wire [8-1:0] node1573;
	wire [8-1:0] node1579;
	wire [8-1:0] node1581;
	wire [8-1:0] node1582;
	wire [8-1:0] node1586;
	wire [8-1:0] node1587;
	wire [8-1:0] node1591;
	wire [8-1:0] node1592;
	wire [8-1:0] node1593;
	wire [8-1:0] node1594;
	wire [8-1:0] node1598;
	wire [8-1:0] node1600;
	wire [8-1:0] node1603;
	wire [8-1:0] node1604;
	wire [8-1:0] node1607;
	wire [8-1:0] node1609;
	wire [8-1:0] node1612;
	wire [8-1:0] node1613;
	wire [8-1:0] node1614;
	wire [8-1:0] node1615;
	wire [8-1:0] node1616;
	wire [8-1:0] node1617;
	wire [8-1:0] node1621;
	wire [8-1:0] node1623;
	wire [8-1:0] node1626;
	wire [8-1:0] node1628;
	wire [8-1:0] node1629;
	wire [8-1:0] node1631;
	wire [8-1:0] node1635;
	wire [8-1:0] node1636;
	wire [8-1:0] node1637;
	wire [8-1:0] node1638;
	wire [8-1:0] node1640;
	wire [8-1:0] node1644;
	wire [8-1:0] node1645;
	wire [8-1:0] node1646;
	wire [8-1:0] node1650;
	wire [8-1:0] node1653;
	wire [8-1:0] node1654;
	wire [8-1:0] node1655;
	wire [8-1:0] node1659;
	wire [8-1:0] node1660;
	wire [8-1:0] node1663;
	wire [8-1:0] node1665;
	wire [8-1:0] node1668;
	wire [8-1:0] node1669;
	wire [8-1:0] node1670;
	wire [8-1:0] node1671;
	wire [8-1:0] node1672;
	wire [8-1:0] node1676;
	wire [8-1:0] node1678;
	wire [8-1:0] node1679;
	wire [8-1:0] node1681;
	wire [8-1:0] node1685;
	wire [8-1:0] node1686;
	wire [8-1:0] node1687;
	wire [8-1:0] node1688;
	wire [8-1:0] node1693;
	wire [8-1:0] node1694;
	wire [8-1:0] node1696;
	wire [8-1:0] node1700;
	wire [8-1:0] node1701;
	wire [8-1:0] node1702;
	wire [8-1:0] node1703;
	wire [8-1:0] node1707;
	wire [8-1:0] node1708;
	wire [8-1:0] node1709;
	wire [8-1:0] node1713;
	wire [8-1:0] node1716;
	wire [8-1:0] node1717;
	wire [8-1:0] node1720;
	wire [8-1:0] node1721;
	wire [8-1:0] node1725;
	wire [8-1:0] node1726;
	wire [8-1:0] node1727;
	wire [8-1:0] node1728;
	wire [8-1:0] node1729;
	wire [8-1:0] node1730;
	wire [8-1:0] node1733;
	wire [8-1:0] node1735;
	wire [8-1:0] node1738;
	wire [8-1:0] node1739;
	wire [8-1:0] node1740;
	wire [8-1:0] node1744;
	wire [8-1:0] node1745;
	wire [8-1:0] node1749;
	wire [8-1:0] node1750;
	wire [8-1:0] node1751;
	wire [8-1:0] node1754;
	wire [8-1:0] node1755;
	wire [8-1:0] node1757;
	wire [8-1:0] node1760;
	wire [8-1:0] node1763;
	wire [8-1:0] node1764;
	wire [8-1:0] node1767;
	wire [8-1:0] node1769;
	wire [8-1:0] node1772;
	wire [8-1:0] node1773;
	wire [8-1:0] node1774;
	wire [8-1:0] node1775;
	wire [8-1:0] node1776;
	wire [8-1:0] node1777;
	wire [8-1:0] node1781;
	wire [8-1:0] node1784;
	wire [8-1:0] node1787;
	wire [8-1:0] node1789;
	wire [8-1:0] node1791;
	wire [8-1:0] node1794;
	wire [8-1:0] node1795;
	wire [8-1:0] node1796;
	wire [8-1:0] node1797;
	wire [8-1:0] node1801;
	wire [8-1:0] node1802;
	wire [8-1:0] node1803;
	wire [8-1:0] node1806;
	wire [8-1:0] node1810;
	wire [8-1:0] node1811;
	wire [8-1:0] node1812;
	wire [8-1:0] node1816;
	wire [8-1:0] node1819;
	wire [8-1:0] node1820;
	wire [8-1:0] node1821;
	wire [8-1:0] node1822;
	wire [8-1:0] node1823;
	wire [8-1:0] node1824;
	wire [8-1:0] node1827;
	wire [8-1:0] node1830;
	wire [8-1:0] node1831;
	wire [8-1:0] node1835;
	wire [8-1:0] node1836;
	wire [8-1:0] node1838;
	wire [8-1:0] node1841;
	wire [8-1:0] node1842;
	wire [8-1:0] node1845;
	wire [8-1:0] node1848;
	wire [8-1:0] node1849;
	wire [8-1:0] node1850;
	wire [8-1:0] node1852;
	wire [8-1:0] node1854;
	wire [8-1:0] node1858;
	wire [8-1:0] node1859;
	wire [8-1:0] node1860;
	wire [8-1:0] node1861;
	wire [8-1:0] node1866;
	wire [8-1:0] node1869;
	wire [8-1:0] node1870;
	wire [8-1:0] node1871;
	wire [8-1:0] node1872;
	wire [8-1:0] node1875;
	wire [8-1:0] node1878;
	wire [8-1:0] node1880;
	wire [8-1:0] node1881;
	wire [8-1:0] node1885;
	wire [8-1:0] node1886;
	wire [8-1:0] node1887;
	wire [8-1:0] node1889;
	wire [8-1:0] node1893;
	wire [8-1:0] node1894;
	wire [8-1:0] node1897;
	wire [8-1:0] node1898;
	wire [8-1:0] node1900;
	wire [8-1:0] node1901;
	wire [8-1:0] node1906;
	wire [8-1:0] node1907;
	wire [8-1:0] node1908;
	wire [8-1:0] node1909;
	wire [8-1:0] node1910;
	wire [8-1:0] node1911;
	wire [8-1:0] node1913;
	wire [8-1:0] node1915;
	wire [8-1:0] node1916;
	wire [8-1:0] node1919;
	wire [8-1:0] node1922;
	wire [8-1:0] node1923;
	wire [8-1:0] node1924;
	wire [8-1:0] node1925;
	wire [8-1:0] node1930;
	wire [8-1:0] node1933;
	wire [8-1:0] node1934;
	wire [8-1:0] node1936;
	wire [8-1:0] node1938;
	wire [8-1:0] node1939;
	wire [8-1:0] node1942;
	wire [8-1:0] node1943;
	wire [8-1:0] node1947;
	wire [8-1:0] node1948;
	wire [8-1:0] node1949;
	wire [8-1:0] node1952;
	wire [8-1:0] node1955;
	wire [8-1:0] node1956;
	wire [8-1:0] node1957;
	wire [8-1:0] node1961;
	wire [8-1:0] node1962;
	wire [8-1:0] node1966;
	wire [8-1:0] node1967;
	wire [8-1:0] node1969;
	wire [8-1:0] node1970;
	wire [8-1:0] node1971;
	wire [8-1:0] node1972;
	wire [8-1:0] node1976;
	wire [8-1:0] node1978;
	wire [8-1:0] node1981;
	wire [8-1:0] node1984;
	wire [8-1:0] node1985;
	wire [8-1:0] node1986;
	wire [8-1:0] node1987;
	wire [8-1:0] node1988;
	wire [8-1:0] node1992;
	wire [8-1:0] node1995;
	wire [8-1:0] node1997;
	wire [8-1:0] node1998;
	wire [8-1:0] node2002;
	wire [8-1:0] node2003;
	wire [8-1:0] node2005;
	wire [8-1:0] node2008;
	wire [8-1:0] node2010;
	wire [8-1:0] node2013;
	wire [8-1:0] node2014;
	wire [8-1:0] node2016;
	wire [8-1:0] node2017;
	wire [8-1:0] node2018;
	wire [8-1:0] node2019;
	wire [8-1:0] node2021;
	wire [8-1:0] node2024;
	wire [8-1:0] node2026;
	wire [8-1:0] node2029;
	wire [8-1:0] node2030;
	wire [8-1:0] node2032;
	wire [8-1:0] node2034;
	wire [8-1:0] node2037;
	wire [8-1:0] node2038;
	wire [8-1:0] node2042;
	wire [8-1:0] node2043;
	wire [8-1:0] node2045;
	wire [8-1:0] node2047;
	wire [8-1:0] node2050;
	wire [8-1:0] node2051;
	wire [8-1:0] node2052;
	wire [8-1:0] node2055;
	wire [8-1:0] node2058;
	wire [8-1:0] node2061;
	wire [8-1:0] node2062;
	wire [8-1:0] node2063;
	wire [8-1:0] node2064;
	wire [8-1:0] node2066;
	wire [8-1:0] node2069;
	wire [8-1:0] node2070;
	wire [8-1:0] node2073;
	wire [8-1:0] node2075;
	wire [8-1:0] node2078;
	wire [8-1:0] node2079;
	wire [8-1:0] node2081;
	wire [8-1:0] node2082;
	wire [8-1:0] node2086;
	wire [8-1:0] node2087;
	wire [8-1:0] node2091;
	wire [8-1:0] node2092;
	wire [8-1:0] node2093;
	wire [8-1:0] node2094;
	wire [8-1:0] node2095;
	wire [8-1:0] node2098;
	wire [8-1:0] node2102;
	wire [8-1:0] node2103;
	wire [8-1:0] node2105;
	wire [8-1:0] node2106;
	wire [8-1:0] node2109;
	wire [8-1:0] node2112;
	wire [8-1:0] node2113;
	wire [8-1:0] node2114;
	wire [8-1:0] node2118;
	wire [8-1:0] node2121;
	wire [8-1:0] node2122;
	wire [8-1:0] node2123;
	wire [8-1:0] node2124;
	wire [8-1:0] node2125;
	wire [8-1:0] node2129;
	wire [8-1:0] node2132;
	wire [8-1:0] node2133;
	wire [8-1:0] node2135;
	wire [8-1:0] node2138;
	wire [8-1:0] node2141;
	wire [8-1:0] node2142;
	wire [8-1:0] node2145;
	wire [8-1:0] node2148;
	wire [8-1:0] node2149;
	wire [8-1:0] node2151;
	wire [8-1:0] node2152;
	wire [8-1:0] node2153;
	wire [8-1:0] node2154;
	wire [8-1:0] node2155;
	wire [8-1:0] node2159;
	wire [8-1:0] node2162;
	wire [8-1:0] node2163;
	wire [8-1:0] node2164;
	wire [8-1:0] node2166;
	wire [8-1:0] node2169;
	wire [8-1:0] node2171;
	wire [8-1:0] node2173;
	wire [8-1:0] node2176;
	wire [8-1:0] node2177;
	wire [8-1:0] node2181;
	wire [8-1:0] node2182;
	wire [8-1:0] node2183;
	wire [8-1:0] node2186;
	wire [8-1:0] node2189;
	wire [8-1:0] node2190;
	wire [8-1:0] node2191;
	wire [8-1:0] node2192;
	wire [8-1:0] node2195;
	wire [8-1:0] node2199;
	wire [8-1:0] node2200;
	wire [8-1:0] node2202;
	wire [8-1:0] node2205;
	wire [8-1:0] node2208;
	wire [8-1:0] node2209;
	wire [8-1:0] node2210;
	wire [8-1:0] node2211;
	wire [8-1:0] node2212;
	wire [8-1:0] node2214;
	wire [8-1:0] node2217;
	wire [8-1:0] node2218;
	wire [8-1:0] node2222;
	wire [8-1:0] node2223;
	wire [8-1:0] node2225;
	wire [8-1:0] node2228;
	wire [8-1:0] node2229;
	wire [8-1:0] node2233;
	wire [8-1:0] node2234;
	wire [8-1:0] node2235;
	wire [8-1:0] node2238;
	wire [8-1:0] node2239;
	wire [8-1:0] node2241;
	wire [8-1:0] node2245;
	wire [8-1:0] node2246;
	wire [8-1:0] node2247;
	wire [8-1:0] node2249;
	wire [8-1:0] node2252;
	wire [8-1:0] node2253;
	wire [8-1:0] node2257;
	wire [8-1:0] node2258;
	wire [8-1:0] node2259;
	wire [8-1:0] node2263;
	wire [8-1:0] node2264;
	wire [8-1:0] node2267;
	wire [8-1:0] node2270;
	wire [8-1:0] node2271;
	wire [8-1:0] node2272;
	wire [8-1:0] node2273;
	wire [8-1:0] node2274;
	wire [8-1:0] node2275;
	wire [8-1:0] node2279;
	wire [8-1:0] node2280;
	wire [8-1:0] node2284;
	wire [8-1:0] node2285;
	wire [8-1:0] node2289;
	wire [8-1:0] node2290;
	wire [8-1:0] node2291;
	wire [8-1:0] node2295;
	wire [8-1:0] node2296;
	wire [8-1:0] node2298;
	wire [8-1:0] node2301;
	wire [8-1:0] node2302;
	wire [8-1:0] node2306;
	wire [8-1:0] node2307;
	wire [8-1:0] node2308;
	wire [8-1:0] node2309;
	wire [8-1:0] node2311;
	wire [8-1:0] node2312;
	wire [8-1:0] node2316;
	wire [8-1:0] node2317;
	wire [8-1:0] node2320;
	wire [8-1:0] node2321;
	wire [8-1:0] node2325;
	wire [8-1:0] node2327;
	wire [8-1:0] node2328;
	wire [8-1:0] node2329;
	wire [8-1:0] node2334;
	wire [8-1:0] node2335;
	wire [8-1:0] node2336;
	wire [8-1:0] node2337;
	wire [8-1:0] node2341;
	wire [8-1:0] node2344;
	wire [8-1:0] node2345;
	wire [8-1:0] node2347;

	assign outp = (inp[4]) ? node1198 : node1;
		assign node1 = (inp[13]) ? node573 : node2;
			assign node2 = (inp[7]) ? node224 : node3;
				assign node3 = (inp[11]) ? node79 : node4;
					assign node4 = (inp[0]) ? node48 : node5;
						assign node5 = (inp[8]) ? node25 : node6;
							assign node6 = (inp[1]) ? node14 : node7;
								assign node7 = (inp[2]) ? node9 : 8'b01111111;
									assign node9 = (inp[5]) ? node11 : 8'b00101111;
										assign node11 = (inp[6]) ? 8'b01111111 : 8'b00101111;
								assign node14 = (inp[5]) ? node18 : node15;
									assign node15 = (inp[2]) ? 8'b00101110 : 8'b00111110;
									assign node18 = (inp[3]) ? 8'b01111111 : node19;
										assign node19 = (inp[2]) ? node21 : 8'b00111110;
											assign node21 = (inp[6]) ? 8'b00111110 : 8'b00101110;
							assign node25 = (inp[2]) ? node37 : node26;
								assign node26 = (inp[1]) ? node28 : 8'b00111011;
									assign node28 = (inp[5]) ? node30 : 8'b00111010;
										assign node30 = (inp[10]) ? node34 : node31;
											assign node31 = (inp[9]) ? 8'b00111011 : 8'b00111010;
											assign node34 = (inp[3]) ? 8'b01111111 : 8'b00111110;
								assign node37 = (inp[1]) ? node39 : 8'b00101011;
									assign node39 = (inp[5]) ? node41 : 8'b00101010;
										assign node41 = (inp[12]) ? node43 : 8'b00111110;
											assign node43 = (inp[6]) ? 8'b00111011 : node44;
												assign node44 = (inp[9]) ? 8'b00101011 : 8'b00101010;
						assign node48 = (inp[5]) ? 8'b01111111 : node49;
							assign node49 = (inp[6]) ? node63 : node50;
								assign node50 = (inp[8]) ? node56 : node51;
									assign node51 = (inp[3]) ? node53 : 8'b01111111;
										assign node53 = (inp[1]) ? 8'b00111110 : 8'b01111111;
									assign node56 = (inp[10]) ? node58 : 8'b01111111;
										assign node58 = (inp[3]) ? node60 : 8'b00111011;
											assign node60 = (inp[12]) ? 8'b00111010 : 8'b00111011;
								assign node63 = (inp[2]) ? node71 : node64;
									assign node64 = (inp[3]) ? node66 : 8'b01111111;
										assign node66 = (inp[1]) ? node68 : 8'b01111111;
											assign node68 = (inp[10]) ? 8'b00111010 : 8'b00111110;
									assign node71 = (inp[12]) ? node75 : node72;
										assign node72 = (inp[1]) ? 8'b00101110 : 8'b00101111;
										assign node75 = (inp[8]) ? 8'b00101011 : 8'b00101111;
					assign node79 = (inp[8]) ? node129 : node80;
						assign node80 = (inp[1]) ? node104 : node81;
							assign node81 = (inp[2]) ? node85 : node82;
								assign node82 = (inp[12]) ? 8'b01111111 : 8'b00101111;
								assign node85 = (inp[12]) ? node93 : node86;
									assign node86 = (inp[9]) ? 8'b00111110 : node87;
										assign node87 = (inp[5]) ? 8'b00101110 : node88;
											assign node88 = (inp[0]) ? 8'b00101110 : 8'b00111110;
									assign node93 = (inp[10]) ? node99 : node94;
										assign node94 = (inp[0]) ? node96 : 8'b00101111;
											assign node96 = (inp[6]) ? 8'b00101111 : 8'b00111110;
										assign node99 = (inp[5]) ? 8'b00111110 : node100;
											assign node100 = (inp[6]) ? 8'b00101111 : 8'b00111110;
							assign node104 = (inp[2]) ? node110 : node105;
								assign node105 = (inp[12]) ? node107 : 8'b00101110;
									assign node107 = (inp[0]) ? 8'b00111011 : 8'b00111110;
								assign node110 = (inp[12]) ? node120 : node111;
									assign node111 = (inp[5]) ? node115 : node112;
										assign node112 = (inp[3]) ? 8'b00111011 : 8'b00111010;
										assign node115 = (inp[6]) ? 8'b00101010 : node116;
											assign node116 = (inp[3]) ? 8'b00111010 : 8'b00111011;
									assign node120 = (inp[0]) ? node126 : node121;
										assign node121 = (inp[9]) ? 8'b00101110 : node122;
											assign node122 = (inp[10]) ? 8'b00101110 : 8'b00111011;
										assign node126 = (inp[5]) ? 8'b00111010 : 8'b00111011;
						assign node129 = (inp[2]) ? node175 : node130;
							assign node130 = (inp[12]) ? node152 : node131;
								assign node131 = (inp[0]) ? node143 : node132;
									assign node132 = (inp[5]) ? node136 : node133;
										assign node133 = (inp[1]) ? 8'b00101010 : 8'b00101011;
										assign node136 = (inp[10]) ? node138 : 8'b00101010;
											assign node138 = (inp[3]) ? 8'b00001011 : node139;
												assign node139 = (inp[9]) ? 8'b00001111 : 8'b00001110;
									assign node143 = (inp[3]) ? node149 : node144;
										assign node144 = (inp[1]) ? node146 : 8'b00001111;
											assign node146 = (inp[10]) ? 8'b00001111 : 8'b00001011;
										assign node149 = (inp[1]) ? 8'b00001011 : 8'b00101011;
								assign node152 = (inp[5]) ? node160 : node153;
									assign node153 = (inp[1]) ? 8'b00111010 : node154;
										assign node154 = (inp[0]) ? node156 : 8'b00111011;
											assign node156 = (inp[10]) ? 8'b00111011 : 8'b00011111;
									assign node160 = (inp[1]) ? node166 : node161;
										assign node161 = (inp[0]) ? 8'b00011111 : node162;
											assign node162 = (inp[10]) ? 8'b00011111 : 8'b00111011;
										assign node166 = (inp[3]) ? node170 : node167;
											assign node167 = (inp[10]) ? 8'b00011011 : 8'b00111010;
											assign node170 = (inp[0]) ? 8'b00011011 : node171;
												assign node171 = (inp[10]) ? 8'b00011011 : 8'b00011111;
							assign node175 = (inp[1]) ? node189 : node176;
								assign node176 = (inp[5]) ? node186 : node177;
									assign node177 = (inp[9]) ? node183 : node178;
										assign node178 = (inp[3]) ? 8'b00001111 : node179;
											assign node179 = (inp[12]) ? 8'b00011110 : 8'b00001110;
										assign node183 = (inp[0]) ? 8'b00111010 : 8'b00101011;
									assign node186 = (inp[12]) ? 8'b00011110 : 8'b00001110;
								assign node189 = (inp[0]) ? node209 : node190;
									assign node190 = (inp[3]) ? node200 : node191;
										assign node191 = (inp[10]) ? node193 : 8'b00101010;
											assign node193 = (inp[12]) ? node197 : node194;
												assign node194 = (inp[6]) ? 8'b00001011 : 8'b00011011;
												assign node197 = (inp[6]) ? 8'b00011011 : 8'b00001110;
										assign node200 = (inp[10]) ? 8'b00011010 : node201;
											assign node201 = (inp[6]) ? 8'b00011110 : node202;
												assign node202 = (inp[12]) ? 8'b00001111 : node203;
													assign node203 = (inp[5]) ? 8'b00011110 : 8'b00011111;
									assign node209 = (inp[5]) ? node221 : node210;
										assign node210 = (inp[12]) ? 8'b00101010 : node211;
											assign node211 = (inp[10]) ? node215 : node212;
												assign node212 = (inp[9]) ? 8'b00001010 : 8'b00001011;
												assign node215 = (inp[9]) ? node217 : 8'b00001110;
													assign node217 = (inp[3]) ? 8'b00011111 : 8'b00011110;
										assign node221 = (inp[12]) ? 8'b00011010 : 8'b00001010;
				assign node224 = (inp[9]) ? node398 : node225;
					assign node225 = (inp[11]) ? node303 : node226;
						assign node226 = (inp[6]) ? node262 : node227;
							assign node227 = (inp[10]) ? node247 : node228;
								assign node228 = (inp[0]) ? node240 : node229;
									assign node229 = (inp[8]) ? node237 : node230;
										assign node230 = (inp[5]) ? node234 : node231;
											assign node231 = (inp[1]) ? 8'b00111110 : 8'b01111111;
											assign node234 = (inp[1]) ? 8'b00101111 : 8'b00101110;
										assign node237 = (inp[2]) ? 8'b00101010 : 8'b00111010;
									assign node240 = (inp[3]) ? node242 : 8'b01111111;
										assign node242 = (inp[5]) ? node244 : 8'b00111110;
											assign node244 = (inp[12]) ? 8'b00111110 : 8'b01111111;
								assign node247 = (inp[5]) ? node255 : node248;
									assign node248 = (inp[3]) ? node250 : 8'b00111011;
										assign node250 = (inp[2]) ? node252 : 8'b00111010;
											assign node252 = (inp[0]) ? 8'b00111010 : 8'b00101010;
									assign node255 = (inp[8]) ? node259 : node256;
										assign node256 = (inp[0]) ? 8'b00111011 : 8'b00101011;
										assign node259 = (inp[1]) ? 8'b01111111 : 8'b00101111;
							assign node262 = (inp[3]) ? node282 : node263;
								assign node263 = (inp[0]) ? node277 : node264;
									assign node264 = (inp[1]) ? 8'b00101010 : node265;
										assign node265 = (inp[12]) ? node271 : node266;
											assign node266 = (inp[5]) ? node268 : 8'b00101011;
												assign node268 = (inp[8]) ? 8'b01111111 : 8'b00101011;
											assign node271 = (inp[8]) ? node273 : 8'b00101111;
												assign node273 = (inp[5]) ? 8'b00101111 : 8'b00101011;
									assign node277 = (inp[1]) ? 8'b00101111 : node278;
										assign node278 = (inp[10]) ? 8'b00101011 : 8'b00101111;
								assign node282 = (inp[5]) ? node290 : node283;
									assign node283 = (inp[10]) ? 8'b00101010 : node284;
										assign node284 = (inp[1]) ? 8'b00101110 : node285;
											assign node285 = (inp[0]) ? 8'b00101110 : 8'b00101010;
									assign node290 = (inp[1]) ? node300 : node291;
										assign node291 = (inp[2]) ? 8'b00111110 : node292;
											assign node292 = (inp[12]) ? node294 : 8'b00101010;
												assign node294 = (inp[0]) ? 8'b00101110 : node295;
													assign node295 = (inp[8]) ? 8'b00101110 : 8'b00101010;
										assign node300 = (inp[8]) ? 8'b01111111 : 8'b00111011;
						assign node303 = (inp[8]) ? node347 : node304;
							assign node304 = (inp[10]) ? node320 : node305;
								assign node305 = (inp[1]) ? node309 : node306;
									assign node306 = (inp[5]) ? 8'b00111110 : 8'b00101111;
									assign node309 = (inp[5]) ? node313 : node310;
										assign node310 = (inp[0]) ? 8'b00111010 : 8'b00101110;
										assign node313 = (inp[0]) ? node315 : 8'b00111011;
											assign node315 = (inp[2]) ? node317 : 8'b00101011;
												assign node317 = (inp[3]) ? 8'b00111010 : 8'b00101010;
								assign node320 = (inp[12]) ? node332 : node321;
									assign node321 = (inp[3]) ? node329 : node322;
										assign node322 = (inp[1]) ? node326 : node323;
											assign node323 = (inp[0]) ? 8'b00101011 : 8'b00111010;
											assign node326 = (inp[0]) ? 8'b00001110 : 8'b00011111;
										assign node329 = (inp[6]) ? 8'b00011111 : 8'b00001111;
									assign node332 = (inp[6]) ? node340 : node333;
										assign node333 = (inp[3]) ? node337 : node334;
											assign node334 = (inp[2]) ? 8'b00011110 : 8'b00011111;
											assign node337 = (inp[2]) ? 8'b00011111 : 8'b00111010;
										assign node340 = (inp[3]) ? 8'b00101010 : node341;
											assign node341 = (inp[0]) ? node343 : 8'b00101010;
												assign node343 = (inp[2]) ? 8'b00001111 : 8'b00101011;
							assign node347 = (inp[5]) ? node373 : node348;
								assign node348 = (inp[3]) ? node364 : node349;
									assign node349 = (inp[1]) ? node357 : node350;
										assign node350 = (inp[10]) ? node354 : node351;
											assign node351 = (inp[12]) ? 8'b00011111 : 8'b00111010;
											assign node354 = (inp[12]) ? 8'b00111011 : 8'b00101011;
										assign node357 = (inp[10]) ? node361 : node358;
											assign node358 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node361 = (inp[0]) ? 8'b00011110 : 8'b00011111;
									assign node364 = (inp[10]) ? 8'b00101010 : node365;
										assign node365 = (inp[12]) ? 8'b00111010 : node366;
											assign node366 = (inp[0]) ? node368 : 8'b00011111;
												assign node368 = (inp[6]) ? 8'b00011011 : 8'b00001011;
								assign node373 = (inp[10]) ? node385 : node374;
									assign node374 = (inp[0]) ? node380 : node375;
										assign node375 = (inp[2]) ? 8'b00011111 : node376;
											assign node376 = (inp[6]) ? 8'b00011110 : 8'b00101010;
										assign node380 = (inp[12]) ? node382 : 8'b00001010;
											assign node382 = (inp[3]) ? 8'b00011110 : 8'b00011010;
									assign node385 = (inp[3]) ? node387 : 8'b00011010;
										assign node387 = (inp[12]) ? node395 : node388;
											assign node388 = (inp[0]) ? 8'b00001011 : node389;
												assign node389 = (inp[2]) ? node391 : 8'b00001011;
													assign node391 = (inp[6]) ? 8'b00001010 : 8'b00011010;
											assign node395 = (inp[1]) ? 8'b00001011 : 8'b00001110;
					assign node398 = (inp[8]) ? node488 : node399;
						assign node399 = (inp[10]) ? node441 : node400;
							assign node400 = (inp[11]) ? node418 : node401;
								assign node401 = (inp[3]) ? node407 : node402;
									assign node402 = (inp[0]) ? node404 : 8'b00001110;
										assign node404 = (inp[6]) ? 8'b00001111 : 8'b00011111;
									assign node407 = (inp[5]) ? node415 : node408;
										assign node408 = (inp[6]) ? 8'b00001110 : node409;
											assign node409 = (inp[2]) ? node411 : 8'b00011110;
												assign node411 = (inp[12]) ? 8'b00001110 : 8'b00011110;
										assign node415 = (inp[6]) ? 8'b00011110 : 8'b00011111;
								assign node418 = (inp[12]) ? node430 : node419;
									assign node419 = (inp[6]) ? node427 : node420;
										assign node420 = (inp[2]) ? node424 : node421;
											assign node421 = (inp[3]) ? 8'b00001110 : 8'b00001011;
											assign node424 = (inp[0]) ? 8'b00001011 : 8'b00011011;
										assign node427 = (inp[2]) ? 8'b00001010 : 8'b00011010;
									assign node430 = (inp[2]) ? node434 : node431;
										assign node431 = (inp[5]) ? 8'b00001011 : 8'b00001111;
										assign node434 = (inp[0]) ? node436 : 8'b00001011;
											assign node436 = (inp[5]) ? node438 : 8'b00001110;
												assign node438 = (inp[1]) ? 8'b00011010 : 8'b00011110;
							assign node441 = (inp[3]) ? node461 : node442;
								assign node442 = (inp[1]) ? node454 : node443;
									assign node443 = (inp[5]) ? node451 : node444;
										assign node444 = (inp[11]) ? node448 : node445;
											assign node445 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node448 = (inp[2]) ? 8'b00011010 : 8'b00001011;
										assign node451 = (inp[6]) ? 8'b00011010 : 8'b00011011;
									assign node454 = (inp[5]) ? 8'b11110111 : node455;
										assign node455 = (inp[2]) ? node457 : 8'b10000001;
											assign node457 = (inp[12]) ? 8'b00000010 : 8'b10000010;
								assign node461 = (inp[11]) ? node469 : node462;
									assign node462 = (inp[6]) ? node466 : node463;
										assign node463 = (inp[1]) ? 8'b10011001 : 8'b00011010;
										assign node466 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node469 = (inp[12]) ? node479 : node470;
										assign node470 = (inp[2]) ? node472 : 8'b11110111;
											assign node472 = (inp[1]) ? node476 : node473;
												assign node473 = (inp[6]) ? 8'b10100101 : 8'b11110111;
												assign node476 = (inp[5]) ? 8'b10110100 : 8'b10100101;
										assign node479 = (inp[6]) ? 8'b00000010 : node480;
											assign node480 = (inp[1]) ? node484 : node481;
												assign node481 = (inp[0]) ? 8'b11110101 : 8'b00000010;
												assign node484 = (inp[2]) ? 8'b11110101 : 8'b11111101;
						assign node488 = (inp[0]) ? node528 : node489;
							assign node489 = (inp[5]) ? node507 : node490;
								assign node490 = (inp[3]) ? node500 : node491;
									assign node491 = (inp[12]) ? node497 : node492;
										assign node492 = (inp[11]) ? node494 : 8'b00011010;
											assign node494 = (inp[2]) ? 8'b00011010 : 8'b00001011;
										assign node497 = (inp[10]) ? 8'b00001011 : 8'b00011011;
									assign node500 = (inp[12]) ? node504 : node501;
										assign node501 = (inp[11]) ? 8'b11110111 : 8'b10000010;
										assign node504 = (inp[6]) ? 8'b00000010 : 8'b00011010;
								assign node507 = (inp[3]) ? node517 : node508;
									assign node508 = (inp[10]) ? node510 : 8'b11110111;
										assign node510 = (inp[1]) ? 8'b10000100 : node511;
											assign node511 = (inp[6]) ? 8'b10101100 : node512;
												assign node512 = (inp[12]) ? 8'b10101101 : 8'b10001101;
									assign node517 = (inp[1]) ? node523 : node518;
										assign node518 = (inp[11]) ? node520 : 8'b00000010;
											assign node520 = (inp[12]) ? 8'b00011010 : 8'b00001010;
										assign node523 = (inp[11]) ? 8'b10110100 : node524;
											assign node524 = (inp[2]) ? 8'b10000001 : 8'b10011001;
							assign node528 = (inp[11]) ? node550 : node529;
								assign node529 = (inp[3]) ? node541 : node530;
									assign node530 = (inp[6]) ? node532 : 8'b10011101;
										assign node532 = (inp[10]) ? node538 : node533;
											assign node533 = (inp[5]) ? 8'b10011101 : node534;
												assign node534 = (inp[1]) ? 8'b10000101 : 8'b10001101;
											assign node538 = (inp[5]) ? 8'b10001101 : 8'b00001011;
									assign node541 = (inp[2]) ? node545 : node542;
										assign node542 = (inp[6]) ? 8'b10000100 : 8'b10011100;
										assign node545 = (inp[5]) ? node547 : 8'b10010000;
											assign node547 = (inp[1]) ? 8'b10010101 : 8'b10010100;
								assign node550 = (inp[2]) ? node560 : node551;
									assign node551 = (inp[1]) ? node557 : node552;
										assign node552 = (inp[10]) ? 8'b10101101 : node553;
											assign node553 = (inp[12]) ? 8'b10111100 : 8'b10101100;
										assign node557 = (inp[10]) ? 8'b10111001 : 8'b10100001;
									assign node560 = (inp[3]) ? node566 : node561;
										assign node561 = (inp[1]) ? node563 : 8'b10111100;
											assign node563 = (inp[10]) ? 8'b10110100 : 8'b10110000;
										assign node566 = (inp[10]) ? node570 : node567;
											assign node567 = (inp[6]) ? 8'b10100100 : 8'b10110001;
											assign node570 = (inp[6]) ? 8'b00000010 : 8'b10100000;
			assign node573 = (inp[5]) ? node865 : node574;
				assign node574 = (inp[0]) ? node674 : node575;
					assign node575 = (inp[8]) ? node623 : node576;
						assign node576 = (inp[7]) ? node596 : node577;
							assign node577 = (inp[1]) ? node589 : node578;
								assign node578 = (inp[2]) ? node584 : node579;
									assign node579 = (inp[12]) ? 8'b00011111 : node580;
										assign node580 = (inp[11]) ? 8'b00001111 : 8'b00011111;
									assign node584 = (inp[11]) ? node586 : 8'b00001111;
										assign node586 = (inp[12]) ? 8'b00001111 : 8'b00011110;
								assign node589 = (inp[2]) ? 8'b00001110 : node590;
									assign node590 = (inp[12]) ? 8'b00011110 : node591;
										assign node591 = (inp[10]) ? 8'b00001110 : 8'b00011110;
							assign node596 = (inp[10]) ? node612 : node597;
								assign node597 = (inp[12]) ? node609 : node598;
									assign node598 = (inp[9]) ? 8'b00011011 : node599;
										assign node599 = (inp[2]) ? node603 : node600;
											assign node600 = (inp[3]) ? 8'b00001110 : 8'b00001111;
											assign node603 = (inp[11]) ? node605 : 8'b00001110;
												assign node605 = (inp[1]) ? 8'b00011011 : 8'b00011110;
									assign node609 = (inp[1]) ? 8'b00001110 : 8'b00001111;
								assign node612 = (inp[2]) ? node620 : node613;
									assign node613 = (inp[3]) ? node615 : 8'b00001011;
										assign node615 = (inp[6]) ? 8'b00000010 : node616;
											assign node616 = (inp[9]) ? 8'b00001010 : 8'b00011010;
									assign node620 = (inp[12]) ? 8'b00000010 : 8'b11110111;
						assign node623 = (inp[1]) ? node655 : node624;
							assign node624 = (inp[7]) ? node640 : node625;
								assign node625 = (inp[3]) ? node633 : node626;
									assign node626 = (inp[6]) ? 8'b00001011 : node627;
										assign node627 = (inp[9]) ? 8'b00001011 : node628;
											assign node628 = (inp[12]) ? 8'b00011011 : 8'b00001011;
									assign node633 = (inp[11]) ? node637 : node634;
										assign node634 = (inp[2]) ? 8'b00001011 : 8'b00011011;
										assign node637 = (inp[2]) ? 8'b00011010 : 8'b00001011;
								assign node640 = (inp[3]) ? node648 : node641;
									assign node641 = (inp[12]) ? 8'b00001011 : node642;
										assign node642 = (inp[6]) ? 8'b00011010 : node643;
											assign node643 = (inp[9]) ? 8'b00001011 : 8'b00011011;
									assign node648 = (inp[12]) ? 8'b00000010 : node649;
										assign node649 = (inp[9]) ? node651 : 8'b11110111;
											assign node651 = (inp[2]) ? 8'b10000010 : 8'b00001010;
							assign node655 = (inp[2]) ? node669 : node656;
								assign node656 = (inp[6]) ? node662 : node657;
									assign node657 = (inp[7]) ? 8'b00011010 : node658;
										assign node658 = (inp[11]) ? 8'b00001010 : 8'b00011010;
									assign node662 = (inp[11]) ? node666 : node663;
										assign node663 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node666 = (inp[12]) ? 8'b00011010 : 8'b11110111;
								assign node669 = (inp[12]) ? 8'b00000010 : node670;
									assign node670 = (inp[11]) ? 8'b11110111 : 8'b10000010;
					assign node674 = (inp[9]) ? node760 : node675;
						assign node675 = (inp[11]) ? node713 : node676;
							assign node676 = (inp[10]) ? node696 : node677;
								assign node677 = (inp[6]) ? node687 : node678;
									assign node678 = (inp[3]) ? node680 : 8'b11111101;
										assign node680 = (inp[8]) ? node682 : 8'b10111100;
											assign node682 = (inp[7]) ? 8'b10110100 : node683;
												assign node683 = (inp[12]) ? 8'b11111101 : 8'b10111100;
									assign node687 = (inp[8]) ? node693 : node688;
										assign node688 = (inp[1]) ? node690 : 8'b11111101;
											assign node690 = (inp[3]) ? 8'b10111100 : 8'b10101101;
										assign node693 = (inp[7]) ? 8'b10100101 : 8'b10101101;
								assign node696 = (inp[1]) ? node708 : node697;
									assign node697 = (inp[7]) ? node703 : node698;
										assign node698 = (inp[6]) ? node700 : 8'b11111101;
											assign node700 = (inp[2]) ? 8'b10101101 : 8'b10111001;
										assign node703 = (inp[3]) ? 8'b10100000 : node704;
											assign node704 = (inp[6]) ? 8'b10101001 : 8'b10111001;
									assign node708 = (inp[6]) ? node710 : 8'b10110000;
										assign node710 = (inp[3]) ? 8'b10100000 : 8'b10100001;
							assign node713 = (inp[8]) ? node739 : node714;
								assign node714 = (inp[7]) ? node722 : node715;
									assign node715 = (inp[1]) ? node719 : node716;
										assign node716 = (inp[6]) ? 8'b10101101 : 8'b10101100;
										assign node719 = (inp[2]) ? 8'b10111001 : 8'b10101001;
									assign node722 = (inp[2]) ? node732 : node723;
										assign node723 = (inp[10]) ? node729 : node724;
											assign node724 = (inp[3]) ? 8'b10111001 : node725;
												assign node725 = (inp[12]) ? 8'b10111001 : 8'b10111000;
											assign node729 = (inp[12]) ? 8'b10101001 : 8'b10101000;
										assign node732 = (inp[3]) ? 8'b10100000 : node733;
											assign node733 = (inp[6]) ? 8'b10111000 : node734;
												assign node734 = (inp[1]) ? 8'b10101000 : 8'b10101100;
								assign node739 = (inp[2]) ? node753 : node740;
									assign node740 = (inp[3]) ? node748 : node741;
										assign node741 = (inp[6]) ? node745 : node742;
											assign node742 = (inp[7]) ? 8'b10001001 : 8'b10011001;
											assign node745 = (inp[7]) ? 8'b10011100 : 8'b10011101;
										assign node748 = (inp[6]) ? node750 : 8'b10001100;
											assign node750 = (inp[1]) ? 8'b10010001 : 8'b10000100;
									assign node753 = (inp[10]) ? node757 : node754;
										assign node754 = (inp[3]) ? 8'b10010001 : 8'b10010000;
										assign node757 = (inp[1]) ? 8'b10010100 : 8'b10101000;
						assign node760 = (inp[8]) ? node810 : node761;
							assign node761 = (inp[3]) ? node787 : node762;
								assign node762 = (inp[10]) ? node774 : node763;
									assign node763 = (inp[2]) ? node769 : node764;
										assign node764 = (inp[6]) ? 8'b00011111 : node765;
											assign node765 = (inp[12]) ? 8'b00011111 : 8'b00001111;
										assign node769 = (inp[6]) ? node771 : 8'b00011111;
											assign node771 = (inp[11]) ? 8'b00001011 : 8'b00001111;
									assign node774 = (inp[7]) ? node782 : node775;
										assign node775 = (inp[11]) ? node779 : node776;
											assign node776 = (inp[12]) ? 8'b00011111 : 8'b00001111;
											assign node779 = (inp[6]) ? 8'b00011011 : 8'b00011010;
										assign node782 = (inp[6]) ? 8'b00001011 : node783;
											assign node783 = (inp[2]) ? 8'b00001010 : 8'b00011011;
								assign node787 = (inp[7]) ? node797 : node788;
									assign node788 = (inp[1]) ? 8'b00011110 : node789;
										assign node789 = (inp[10]) ? 8'b00011111 : node790;
											assign node790 = (inp[2]) ? node792 : 8'b00001111;
												assign node792 = (inp[12]) ? 8'b00001111 : 8'b00011110;
									assign node797 = (inp[2]) ? node805 : node798;
										assign node798 = (inp[10]) ? node800 : 8'b00001110;
											assign node800 = (inp[6]) ? 8'b00000010 : node801;
												assign node801 = (inp[12]) ? 8'b00011010 : 8'b00001010;
										assign node805 = (inp[6]) ? node807 : 8'b10100101;
											assign node807 = (inp[10]) ? 8'b00000010 : 8'b00011011;
							assign node810 = (inp[10]) ? node842 : node811;
								assign node811 = (inp[11]) ? node827 : node812;
									assign node812 = (inp[3]) ? node820 : node813;
										assign node813 = (inp[1]) ? node817 : node814;
											assign node814 = (inp[2]) ? 8'b10011101 : 8'b10001101;
											assign node817 = (inp[6]) ? 8'b10000101 : 8'b10010101;
										assign node820 = (inp[7]) ? node822 : 8'b10011100;
											assign node822 = (inp[6]) ? 8'b10000100 : node823;
												assign node823 = (inp[1]) ? 8'b10011100 : 8'b10010100;
									assign node827 = (inp[1]) ? node837 : node828;
										assign node828 = (inp[6]) ? node834 : node829;
											assign node829 = (inp[2]) ? 8'b10100001 : node830;
												assign node830 = (inp[3]) ? 8'b11111101 : 8'b10101101;
											assign node834 = (inp[7]) ? 8'b10111100 : 8'b10101101;
										assign node837 = (inp[6]) ? 8'b10110000 : node838;
											assign node838 = (inp[7]) ? 8'b10100001 : 8'b10110001;
								assign node842 = (inp[6]) ? node850 : node843;
									assign node843 = (inp[11]) ? node847 : node844;
										assign node844 = (inp[2]) ? 8'b00011011 : 8'b00011010;
										assign node847 = (inp[12]) ? 8'b00011010 : 8'b00001010;
									assign node850 = (inp[1]) ? node856 : node851;
										assign node851 = (inp[3]) ? 8'b00000010 : node852;
											assign node852 = (inp[11]) ? 8'b00011010 : 8'b00001011;
										assign node856 = (inp[11]) ? node862 : node857;
											assign node857 = (inp[3]) ? node859 : 8'b10000001;
												assign node859 = (inp[12]) ? 8'b00011010 : 8'b10000010;
											assign node862 = (inp[12]) ? 8'b10100101 : 8'b11110111;
				assign node865 = (inp[11]) ? node1015 : node866;
					assign node866 = (inp[0]) ? node966 : node867;
						assign node867 = (inp[9]) ? node915 : node868;
							assign node868 = (inp[1]) ? node896 : node869;
								assign node869 = (inp[8]) ? node885 : node870;
									assign node870 = (inp[12]) ? node878 : node871;
										assign node871 = (inp[2]) ? node875 : node872;
											assign node872 = (inp[10]) ? 8'b00001011 : 8'b00011110;
											assign node875 = (inp[6]) ? 8'b00011111 : 8'b00001111;
										assign node878 = (inp[7]) ? node880 : 8'b00011111;
											assign node880 = (inp[3]) ? 8'b00011110 : node881;
												assign node881 = (inp[6]) ? 8'b00011111 : 8'b00011011;
									assign node885 = (inp[10]) ? node893 : node886;
										assign node886 = (inp[7]) ? node890 : node887;
											assign node887 = (inp[6]) ? 8'b00011011 : 8'b00001011;
											assign node890 = (inp[2]) ? 8'b10000010 : 8'b00001011;
										assign node893 = (inp[7]) ? 8'b10001101 : 8'b10011101;
								assign node896 = (inp[7]) ? node908 : node897;
									assign node897 = (inp[10]) ? node901 : node898;
										assign node898 = (inp[2]) ? 8'b00011110 : 8'b00011010;
										assign node901 = (inp[8]) ? node905 : node902;
											assign node902 = (inp[2]) ? 8'b00001110 : 8'b00011110;
											assign node905 = (inp[2]) ? 8'b10000100 : 8'b10011100;
									assign node908 = (inp[2]) ? node910 : 8'b10000100;
										assign node910 = (inp[3]) ? node912 : 8'b10010000;
											assign node912 = (inp[6]) ? 8'b10010001 : 8'b10000001;
							assign node915 = (inp[7]) ? node933 : node916;
								assign node916 = (inp[8]) ? node926 : node917;
									assign node917 = (inp[2]) ? node923 : node918;
										assign node918 = (inp[3]) ? 8'b11111101 : node919;
											assign node919 = (inp[10]) ? 8'b11111101 : 8'b10111100;
										assign node923 = (inp[6]) ? 8'b11111101 : 8'b10101101;
									assign node926 = (inp[10]) ? node928 : 8'b10111001;
										assign node928 = (inp[3]) ? node930 : 8'b10111100;
											assign node930 = (inp[6]) ? 8'b11111101 : 8'b10101101;
								assign node933 = (inp[10]) ? node949 : node934;
									assign node934 = (inp[6]) ? node940 : node935;
										assign node935 = (inp[1]) ? 8'b10111000 : node936;
											assign node936 = (inp[12]) ? 8'b10111000 : 8'b10111001;
										assign node940 = (inp[8]) ? node942 : 8'b10111100;
											assign node942 = (inp[2]) ? 8'b10110000 : node943;
												assign node943 = (inp[1]) ? 8'b10100000 : node944;
													assign node944 = (inp[3]) ? 8'b10100000 : 8'b10101001;
									assign node949 = (inp[8]) ? node957 : node950;
										assign node950 = (inp[3]) ? node954 : node951;
											assign node951 = (inp[6]) ? 8'b10111001 : 8'b10111000;
											assign node954 = (inp[6]) ? 8'b10110001 : 8'b10100001;
										assign node957 = (inp[1]) ? node963 : node958;
											assign node958 = (inp[3]) ? 8'b10100100 : node959;
												assign node959 = (inp[12]) ? 8'b10101101 : 8'b11111101;
											assign node963 = (inp[12]) ? 8'b11111101 : 8'b11110101;
						assign node966 = (inp[7]) ? node976 : node967;
							assign node967 = (inp[8]) ? node969 : 8'b11111101;
								assign node969 = (inp[12]) ? 8'b11111101 : node970;
									assign node970 = (inp[10]) ? 8'b11111101 : node971;
										assign node971 = (inp[9]) ? 8'b11111101 : 8'b11110101;
							assign node976 = (inp[6]) ? node988 : node977;
								assign node977 = (inp[8]) ? node983 : node978;
									assign node978 = (inp[10]) ? node980 : 8'b11111101;
										assign node980 = (inp[2]) ? 8'b10110001 : 8'b10111001;
									assign node983 = (inp[2]) ? node985 : 8'b11111101;
										assign node985 = (inp[1]) ? 8'b11110101 : 8'b11111101;
								assign node988 = (inp[2]) ? node1004 : node989;
									assign node989 = (inp[12]) ? node997 : node990;
										assign node990 = (inp[8]) ? node994 : node991;
											assign node991 = (inp[9]) ? 8'b10100001 : 8'b10100000;
											assign node994 = (inp[1]) ? 8'b10100101 : 8'b10100100;
										assign node997 = (inp[3]) ? node999 : 8'b10101101;
											assign node999 = (inp[8]) ? node1001 : 8'b10101101;
												assign node1001 = (inp[1]) ? 8'b10100101 : 8'b10100100;
									assign node1004 = (inp[12]) ? node1010 : node1005;
										assign node1005 = (inp[10]) ? node1007 : 8'b11111101;
											assign node1007 = (inp[1]) ? 8'b10110001 : 8'b10111001;
										assign node1010 = (inp[1]) ? 8'b11110101 : node1011;
											assign node1011 = (inp[8]) ? 8'b10110100 : 8'b10110000;
					assign node1015 = (inp[2]) ? node1111 : node1016;
						assign node1016 = (inp[12]) ? node1056 : node1017;
							assign node1017 = (inp[7]) ? node1041 : node1018;
								assign node1018 = (inp[9]) ? node1030 : node1019;
									assign node1019 = (inp[0]) ? node1027 : node1020;
										assign node1020 = (inp[1]) ? node1024 : node1021;
											assign node1021 = (inp[8]) ? 8'b00001011 : 8'b00001111;
											assign node1024 = (inp[8]) ? 8'b10101100 : 8'b00001110;
										assign node1027 = (inp[8]) ? 8'b10001101 : 8'b10101101;
									assign node1030 = (inp[8]) ? node1036 : node1031;
										assign node1031 = (inp[0]) ? 8'b10101001 : node1032;
											assign node1032 = (inp[10]) ? 8'b10101100 : 8'b10101101;
										assign node1036 = (inp[0]) ? node1038 : 8'b10101001;
											assign node1038 = (inp[1]) ? 8'b10001001 : 8'b10001101;
								assign node1041 = (inp[6]) ? node1051 : node1042;
									assign node1042 = (inp[3]) ? node1048 : node1043;
										assign node1043 = (inp[8]) ? node1045 : 8'b10001101;
											assign node1045 = (inp[1]) ? 8'b10001100 : 8'b10001101;
										assign node1048 = (inp[0]) ? 8'b10001001 : 8'b10101101;
									assign node1051 = (inp[3]) ? node1053 : 8'b10010101;
										assign node1053 = (inp[10]) ? 8'b10010100 : 8'b10111000;
							assign node1056 = (inp[1]) ? node1080 : node1057;
								assign node1057 = (inp[7]) ? node1067 : node1058;
									assign node1058 = (inp[8]) ? node1064 : node1059;
										assign node1059 = (inp[9]) ? 8'b11111101 : node1060;
											assign node1060 = (inp[0]) ? 8'b11111101 : 8'b00011111;
										assign node1064 = (inp[9]) ? 8'b10011101 : 8'b11111101;
									assign node1067 = (inp[6]) ? node1071 : node1068;
										assign node1068 = (inp[0]) ? 8'b11111101 : 8'b10011101;
										assign node1071 = (inp[3]) ? 8'b10100000 : node1072;
											assign node1072 = (inp[8]) ? node1076 : node1073;
												assign node1073 = (inp[10]) ? 8'b10101001 : 8'b10101101;
												assign node1076 = (inp[9]) ? 8'b10001101 : 8'b10101101;
								assign node1080 = (inp[3]) ? node1096 : node1081;
									assign node1081 = (inp[0]) ? node1089 : node1082;
										assign node1082 = (inp[9]) ? node1084 : 8'b00011010;
											assign node1084 = (inp[8]) ? node1086 : 8'b10111000;
												assign node1086 = (inp[6]) ? 8'b10000100 : 8'b10011100;
										assign node1089 = (inp[6]) ? 8'b10000101 : node1090;
											assign node1090 = (inp[8]) ? 8'b10011001 : node1091;
												assign node1091 = (inp[10]) ? 8'b10011101 : 8'b10111001;
									assign node1096 = (inp[10]) ? node1106 : node1097;
										assign node1097 = (inp[0]) ? node1101 : node1098;
											assign node1098 = (inp[9]) ? 8'b10111001 : 8'b11111101;
											assign node1101 = (inp[6]) ? node1103 : 8'b10011001;
												assign node1103 = (inp[7]) ? 8'b10101001 : 8'b10111001;
										assign node1106 = (inp[0]) ? 8'b10111001 : node1107;
											assign node1107 = (inp[9]) ? 8'b10011001 : 8'b00011011;
						assign node1111 = (inp[1]) ? node1157 : node1112;
							assign node1112 = (inp[7]) ? node1130 : node1113;
								assign node1113 = (inp[0]) ? node1123 : node1114;
									assign node1114 = (inp[3]) ? node1116 : 8'b10111100;
										assign node1116 = (inp[8]) ? 8'b10111100 : node1117;
											assign node1117 = (inp[12]) ? 8'b00001111 : node1118;
												assign node1118 = (inp[6]) ? 8'b00001110 : 8'b00011110;
									assign node1123 = (inp[12]) ? node1127 : node1124;
										assign node1124 = (inp[8]) ? 8'b10001100 : 8'b10101100;
										assign node1127 = (inp[8]) ? 8'b10011100 : 8'b10111100;
								assign node1130 = (inp[3]) ? node1144 : node1131;
									assign node1131 = (inp[8]) ? node1141 : node1132;
										assign node1132 = (inp[10]) ? node1136 : node1133;
											assign node1133 = (inp[9]) ? 8'b10101100 : 8'b10111100;
											assign node1136 = (inp[0]) ? node1138 : 8'b00011010;
												assign node1138 = (inp[12]) ? 8'b10111000 : 8'b10101000;
										assign node1141 = (inp[6]) ? 8'b10001100 : 8'b10101101;
									assign node1144 = (inp[10]) ? node1152 : node1145;
										assign node1145 = (inp[8]) ? node1149 : node1146;
											assign node1146 = (inp[9]) ? 8'b10111001 : 8'b10101001;
											assign node1149 = (inp[0]) ? 8'b10000001 : 8'b10100101;
										assign node1152 = (inp[6]) ? 8'b10010101 : node1153;
											assign node1153 = (inp[8]) ? 8'b10000001 : 8'b10000101;
							assign node1157 = (inp[8]) ? node1179 : node1158;
								assign node1158 = (inp[10]) ? node1164 : node1159;
									assign node1159 = (inp[0]) ? 8'b10111000 : node1160;
										assign node1160 = (inp[6]) ? 8'b10111000 : 8'b10101001;
									assign node1164 = (inp[7]) ? node1172 : node1165;
										assign node1165 = (inp[9]) ? node1167 : 8'b00011010;
											assign node1167 = (inp[12]) ? 8'b10101100 : node1168;
												assign node1168 = (inp[3]) ? 8'b10101000 : 8'b10101001;
										assign node1172 = (inp[0]) ? node1176 : node1173;
											assign node1173 = (inp[3]) ? 8'b10100101 : 8'b11110101;
											assign node1176 = (inp[12]) ? 8'b10010100 : 8'b10000100;
								assign node1179 = (inp[0]) ? node1195 : node1180;
									assign node1180 = (inp[12]) ? node1184 : node1181;
										assign node1181 = (inp[7]) ? 8'b10010101 : 8'b11110111;
										assign node1184 = (inp[6]) ? node1188 : node1185;
											assign node1185 = (inp[3]) ? 8'b10100001 : 8'b00000010;
											assign node1188 = (inp[7]) ? node1192 : node1189;
												assign node1189 = (inp[10]) ? 8'b10110000 : 8'b10110100;
												assign node1192 = (inp[3]) ? 8'b10010000 : 8'b10010001;
									assign node1195 = (inp[12]) ? 8'b10010000 : 8'b10000000;
		assign node1198 = (inp[7]) ? node1906 : node1199;
			assign node1199 = (inp[13]) ? node1549 : node1200;
				assign node1200 = (inp[9]) ? node1372 : node1201;
					assign node1201 = (inp[8]) ? node1287 : node1202;
						assign node1202 = (inp[10]) ? node1248 : node1203;
							assign node1203 = (inp[6]) ? node1231 : node1204;
								assign node1204 = (inp[11]) ? node1216 : node1205;
									assign node1205 = (inp[3]) ? node1209 : node1206;
										assign node1206 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node1209 = (inp[5]) ? node1213 : node1210;
											assign node1210 = (inp[2]) ? 8'b10010000 : 8'b00000010;
											assign node1213 = (inp[2]) ? 8'b10010001 : 8'b10000001;
									assign node1216 = (inp[3]) ? node1224 : node1217;
										assign node1217 = (inp[12]) ? node1219 : 8'b11110111;
											assign node1219 = (inp[2]) ? 8'b11110101 : node1220;
												assign node1220 = (inp[5]) ? 8'b10100101 : 8'b00000010;
										assign node1224 = (inp[2]) ? node1228 : node1225;
											assign node1225 = (inp[12]) ? 8'b00000010 : 8'b11110111;
											assign node1228 = (inp[5]) ? 8'b00011010 : 8'b00001010;
								assign node1231 = (inp[2]) ? node1239 : node1232;
									assign node1232 = (inp[11]) ? node1234 : 8'b00011010;
										assign node1234 = (inp[5]) ? node1236 : 8'b00001010;
											assign node1236 = (inp[0]) ? 8'b00001011 : 8'b00001010;
									assign node1239 = (inp[3]) ? node1245 : node1240;
										assign node1240 = (inp[5]) ? node1242 : 8'b00000010;
											assign node1242 = (inp[12]) ? 8'b10010000 : 8'b10010001;
										assign node1245 = (inp[11]) ? 8'b11110111 : 8'b00011011;
							assign node1248 = (inp[11]) ? node1258 : node1249;
								assign node1249 = (inp[6]) ? node1255 : node1250;
									assign node1250 = (inp[5]) ? 8'b00001111 : node1251;
										assign node1251 = (inp[2]) ? 8'b00011110 : 8'b00001110;
									assign node1255 = (inp[3]) ? 8'b00011111 : 8'b00011110;
								assign node1258 = (inp[5]) ? node1266 : node1259;
									assign node1259 = (inp[3]) ? node1261 : 8'b00001110;
										assign node1261 = (inp[1]) ? node1263 : 8'b00001111;
											assign node1263 = (inp[2]) ? 8'b00011011 : 8'b00011110;
									assign node1266 = (inp[3]) ? node1278 : node1267;
										assign node1267 = (inp[2]) ? 8'b00011011 : node1268;
											assign node1268 = (inp[1]) ? node1272 : node1269;
												assign node1269 = (inp[12]) ? 8'b00001110 : 8'b00011011;
												assign node1272 = (inp[0]) ? 8'b00011011 : node1273;
													assign node1273 = (inp[6]) ? 8'b00001110 : 8'b00011011;
										assign node1278 = (inp[1]) ? node1284 : node1279;
											assign node1279 = (inp[6]) ? node1281 : 8'b00011110;
												assign node1281 = (inp[2]) ? 8'b00011110 : 8'b00011111;
											assign node1284 = (inp[0]) ? 8'b00011010 : 8'b00001010;
						assign node1287 = (inp[0]) ? node1317 : node1288;
							assign node1288 = (inp[12]) ? node1306 : node1289;
								assign node1289 = (inp[1]) ? node1299 : node1290;
									assign node1290 = (inp[3]) ? node1296 : node1291;
										assign node1291 = (inp[10]) ? node1293 : 8'b11110111;
											assign node1293 = (inp[11]) ? 8'b10101100 : 8'b10000010;
										assign node1296 = (inp[2]) ? 8'b00011010 : 8'b00001011;
									assign node1299 = (inp[5]) ? node1301 : 8'b11110111;
										assign node1301 = (inp[6]) ? 8'b10101101 : node1302;
											assign node1302 = (inp[10]) ? 8'b10000101 : 8'b10000001;
								assign node1306 = (inp[3]) ? node1314 : node1307;
									assign node1307 = (inp[10]) ? 8'b10000100 : node1308;
										assign node1308 = (inp[6]) ? node1310 : 8'b00000010;
											assign node1310 = (inp[11]) ? 8'b00000010 : 8'b00011010;
									assign node1314 = (inp[6]) ? 8'b00011010 : 8'b00001011;
							assign node1317 = (inp[11]) ? node1343 : node1318;
								assign node1318 = (inp[6]) ? node1326 : node1319;
									assign node1319 = (inp[2]) ? node1321 : 8'b10000100;
										assign node1321 = (inp[12]) ? node1323 : 8'b10010100;
											assign node1323 = (inp[10]) ? 8'b10010000 : 8'b10010101;
									assign node1326 = (inp[2]) ? node1332 : node1327;
										assign node1327 = (inp[12]) ? 8'b10011100 : node1328;
											assign node1328 = (inp[5]) ? 8'b10011100 : 8'b10011101;
										assign node1332 = (inp[5]) ? node1340 : node1333;
											assign node1333 = (inp[12]) ? 8'b00000010 : node1334;
												assign node1334 = (inp[3]) ? 8'b10000100 : node1335;
													assign node1335 = (inp[1]) ? 8'b10000101 : 8'b10000100;
											assign node1340 = (inp[1]) ? 8'b10010101 : 8'b10011101;
								assign node1343 = (inp[6]) ? node1359 : node1344;
									assign node1344 = (inp[10]) ? node1352 : node1345;
										assign node1345 = (inp[5]) ? node1349 : node1346;
											assign node1346 = (inp[3]) ? 8'b10110001 : 8'b10100000;
											assign node1349 = (inp[1]) ? 8'b10110000 : 8'b10110001;
										assign node1352 = (inp[12]) ? node1354 : 8'b11110111;
											assign node1354 = (inp[2]) ? node1356 : 8'b00000010;
												assign node1356 = (inp[3]) ? 8'b10110000 : 8'b10110100;
									assign node1359 = (inp[10]) ? 8'b11111101 : node1360;
										assign node1360 = (inp[1]) ? node1368 : node1361;
											assign node1361 = (inp[2]) ? node1363 : 8'b10111100;
												assign node1363 = (inp[3]) ? node1365 : 8'b10100100;
													assign node1365 = (inp[5]) ? 8'b10101100 : 8'b10101101;
											assign node1368 = (inp[2]) ? 8'b10110000 : 8'b10101001;
					assign node1372 = (inp[11]) ? node1448 : node1373;
						assign node1373 = (inp[10]) ? node1407 : node1374;
							assign node1374 = (inp[3]) ? node1390 : node1375;
								assign node1375 = (inp[0]) ? node1383 : node1376;
									assign node1376 = (inp[6]) ? node1378 : 8'b00101010;
										assign node1378 = (inp[2]) ? node1380 : 8'b00111010;
											assign node1380 = (inp[5]) ? 8'b00111010 : 8'b00101010;
									assign node1383 = (inp[8]) ? node1387 : node1384;
										assign node1384 = (inp[5]) ? 8'b00111010 : 8'b00101010;
										assign node1387 = (inp[12]) ? 8'b01111111 : 8'b00101111;
								assign node1390 = (inp[6]) ? node1402 : node1391;
									assign node1391 = (inp[0]) ? node1395 : node1392;
										assign node1392 = (inp[12]) ? 8'b00101010 : 8'b00101011;
										assign node1395 = (inp[12]) ? node1397 : 8'b01111111;
											assign node1397 = (inp[8]) ? 8'b00101111 : node1398;
												assign node1398 = (inp[2]) ? 8'b00111011 : 8'b00101011;
									assign node1402 = (inp[8]) ? node1404 : 8'b00111011;
										assign node1404 = (inp[1]) ? 8'b00111110 : 8'b00111011;
							assign node1407 = (inp[5]) ? node1437 : node1408;
								assign node1408 = (inp[8]) ? node1424 : node1409;
									assign node1409 = (inp[1]) ? node1411 : 8'b00101111;
										assign node1411 = (inp[3]) ? node1419 : node1412;
											assign node1412 = (inp[0]) ? node1416 : node1413;
												assign node1413 = (inp[6]) ? 8'b00111110 : 8'b00101110;
												assign node1416 = (inp[2]) ? 8'b00101111 : 8'b01111111;
											assign node1419 = (inp[2]) ? node1421 : 8'b00111110;
												assign node1421 = (inp[6]) ? 8'b00101110 : 8'b00111110;
									assign node1424 = (inp[1]) ? node1430 : node1425;
										assign node1425 = (inp[0]) ? 8'b00111010 : node1426;
											assign node1426 = (inp[12]) ? 8'b00101010 : 8'b00111010;
										assign node1430 = (inp[2]) ? node1432 : 8'b00111010;
											assign node1432 = (inp[0]) ? node1434 : 8'b00101010;
												assign node1434 = (inp[3]) ? 8'b00101010 : 8'b00101011;
								assign node1437 = (inp[6]) ? node1441 : node1438;
									assign node1438 = (inp[3]) ? 8'b00101111 : 8'b00101110;
									assign node1441 = (inp[3]) ? 8'b01111111 : node1442;
										assign node1442 = (inp[1]) ? node1444 : 8'b00111110;
											assign node1444 = (inp[8]) ? 8'b01111111 : 8'b00111110;
						assign node1448 = (inp[0]) ? node1492 : node1449;
							assign node1449 = (inp[6]) ? node1473 : node1450;
								assign node1450 = (inp[12]) ? node1466 : node1451;
									assign node1451 = (inp[2]) ? node1457 : node1452;
										assign node1452 = (inp[5]) ? node1454 : 8'b00111010;
											assign node1454 = (inp[1]) ? 8'b00011010 : 8'b00011110;
										assign node1457 = (inp[5]) ? node1459 : 8'b00011111;
											assign node1459 = (inp[3]) ? node1463 : node1460;
												assign node1460 = (inp[10]) ? 8'b00111011 : 8'b00011111;
												assign node1463 = (inp[8]) ? 8'b00011110 : 8'b00111010;
									assign node1466 = (inp[1]) ? node1470 : node1467;
										assign node1467 = (inp[3]) ? 8'b00101011 : 8'b00101010;
										assign node1470 = (inp[3]) ? 8'b00001111 : 8'b00001110;
								assign node1473 = (inp[12]) ? node1485 : node1474;
									assign node1474 = (inp[5]) ? node1478 : node1475;
										assign node1475 = (inp[1]) ? 8'b00101010 : 8'b00101110;
										assign node1478 = (inp[2]) ? 8'b00101010 : node1479;
											assign node1479 = (inp[3]) ? node1481 : 8'b00101010;
												assign node1481 = (inp[1]) ? 8'b00001111 : 8'b00101011;
									assign node1485 = (inp[2]) ? node1489 : node1486;
										assign node1486 = (inp[8]) ? 8'b00111010 : 8'b00111011;
										assign node1489 = (inp[1]) ? 8'b00101110 : 8'b00101010;
							assign node1492 = (inp[10]) ? node1520 : node1493;
								assign node1493 = (inp[12]) ? node1511 : node1494;
									assign node1494 = (inp[8]) ? node1502 : node1495;
										assign node1495 = (inp[3]) ? node1499 : node1496;
											assign node1496 = (inp[6]) ? 8'b00001110 : 8'b00011110;
											assign node1499 = (inp[2]) ? 8'b00101010 : 8'b00111010;
										assign node1502 = (inp[2]) ? node1506 : node1503;
											assign node1503 = (inp[1]) ? 8'b00001011 : 8'b00001111;
											assign node1506 = (inp[6]) ? node1508 : 8'b00001010;
												assign node1508 = (inp[1]) ? 8'b00011010 : 8'b00011011;
									assign node1511 = (inp[8]) ? node1513 : 8'b00011111;
										assign node1513 = (inp[5]) ? 8'b00001111 : node1514;
											assign node1514 = (inp[6]) ? 8'b00001110 : node1515;
												assign node1515 = (inp[2]) ? 8'b00011010 : 8'b00001110;
								assign node1520 = (inp[1]) ? node1530 : node1521;
									assign node1521 = (inp[6]) ? node1525 : node1522;
										assign node1522 = (inp[3]) ? 8'b00111010 : 8'b00011011;
										assign node1525 = (inp[12]) ? node1527 : 8'b00001110;
											assign node1527 = (inp[3]) ? 8'b00011111 : 8'b00011110;
									assign node1530 = (inp[6]) ? node1538 : node1531;
										assign node1531 = (inp[2]) ? node1535 : node1532;
											assign node1532 = (inp[12]) ? 8'b00101010 : 8'b00111010;
											assign node1535 = (inp[12]) ? 8'b00011010 : 8'b00001010;
										assign node1538 = (inp[3]) ? node1544 : node1539;
											assign node1539 = (inp[2]) ? node1541 : 8'b00101011;
												assign node1541 = (inp[5]) ? 8'b00101010 : 8'b00101011;
											assign node1544 = (inp[2]) ? node1546 : 8'b00111110;
												assign node1546 = (inp[8]) ? 8'b00101010 : 8'b00101110;
				assign node1549 = (inp[5]) ? node1725 : node1550;
					assign node1550 = (inp[0]) ? node1612 : node1551;
						assign node1551 = (inp[2]) ? node1591 : node1552;
							assign node1552 = (inp[10]) ? node1568 : node1553;
								assign node1553 = (inp[6]) ? node1561 : node1554;
									assign node1554 = (inp[3]) ? node1558 : node1555;
										assign node1555 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node1558 = (inp[12]) ? 8'b00001011 : 8'b00011010;
									assign node1561 = (inp[3]) ? node1565 : node1562;
										assign node1562 = (inp[11]) ? 8'b00001010 : 8'b00011010;
										assign node1565 = (inp[1]) ? 8'b00011010 : 8'b00011011;
								assign node1568 = (inp[8]) ? node1586 : node1569;
									assign node1569 = (inp[1]) ? node1579 : node1570;
										assign node1570 = (inp[6]) ? 8'b00011111 : node1571;
											assign node1571 = (inp[3]) ? 8'b00011110 : node1572;
												assign node1572 = (inp[9]) ? 8'b00001110 : node1573;
													assign node1573 = (inp[12]) ? 8'b00001110 : 8'b00011011;
										assign node1579 = (inp[3]) ? node1581 : 8'b00001110;
											assign node1581 = (inp[11]) ? 8'b00001110 : node1582;
												assign node1582 = (inp[6]) ? 8'b00011110 : 8'b00001110;
									assign node1586 = (inp[6]) ? 8'b00011010 : node1587;
										assign node1587 = (inp[3]) ? 8'b00001011 : 8'b00000010;
							assign node1591 = (inp[11]) ? node1603 : node1592;
								assign node1592 = (inp[12]) ? node1598 : node1593;
									assign node1593 = (inp[8]) ? 8'b10000010 : node1594;
										assign node1594 = (inp[10]) ? 8'b00001110 : 8'b10000010;
									assign node1598 = (inp[6]) ? node1600 : 8'b00000010;
										assign node1600 = (inp[9]) ? 8'b00000010 : 8'b00001011;
								assign node1603 = (inp[12]) ? node1607 : node1604;
									assign node1604 = (inp[8]) ? 8'b11110111 : 8'b00011011;
									assign node1607 = (inp[1]) ? node1609 : 8'b00001011;
										assign node1609 = (inp[10]) ? 8'b00001110 : 8'b00000010;
						assign node1612 = (inp[9]) ? node1668 : node1613;
							assign node1613 = (inp[6]) ? node1635 : node1614;
								assign node1614 = (inp[8]) ? node1626 : node1615;
									assign node1615 = (inp[11]) ? node1621 : node1616;
										assign node1616 = (inp[10]) ? 8'b10101100 : node1617;
											assign node1617 = (inp[2]) ? 8'b10110000 : 8'b10100000;
										assign node1621 = (inp[10]) ? node1623 : 8'b10010101;
											assign node1623 = (inp[2]) ? 8'b10101001 : 8'b10111001;
									assign node1626 = (inp[11]) ? node1628 : 8'b11110101;
										assign node1628 = (inp[10]) ? 8'b10000101 : node1629;
											assign node1629 = (inp[1]) ? node1631 : 8'b10000100;
												assign node1631 = (inp[12]) ? 8'b10010001 : 8'b10010000;
								assign node1635 = (inp[8]) ? node1653 : node1636;
									assign node1636 = (inp[10]) ? node1644 : node1637;
										assign node1637 = (inp[2]) ? 8'b10101001 : node1638;
											assign node1638 = (inp[1]) ? node1640 : 8'b10111001;
												assign node1640 = (inp[3]) ? 8'b10111000 : 8'b10111001;
										assign node1644 = (inp[2]) ? node1650 : node1645;
											assign node1645 = (inp[11]) ? 8'b10111100 : node1646;
												assign node1646 = (inp[3]) ? 8'b10111100 : 8'b11111101;
											assign node1650 = (inp[11]) ? 8'b10111001 : 8'b10101101;
									assign node1653 = (inp[2]) ? node1659 : node1654;
										assign node1654 = (inp[10]) ? 8'b10111001 : node1655;
											assign node1655 = (inp[12]) ? 8'b10011001 : 8'b10001001;
										assign node1659 = (inp[12]) ? node1663 : node1660;
											assign node1660 = (inp[3]) ? 8'b10111000 : 8'b10010100;
											assign node1663 = (inp[1]) ? node1665 : 8'b10101001;
												assign node1665 = (inp[3]) ? 8'b10100000 : 8'b10100001;
							assign node1668 = (inp[10]) ? node1700 : node1669;
								assign node1669 = (inp[8]) ? node1685 : node1670;
									assign node1670 = (inp[1]) ? node1676 : node1671;
										assign node1671 = (inp[11]) ? 8'b00000010 : node1672;
											assign node1672 = (inp[3]) ? 8'b00011011 : 8'b00011010;
										assign node1676 = (inp[11]) ? node1678 : 8'b10000010;
											assign node1678 = (inp[3]) ? 8'b11110111 : node1679;
												assign node1679 = (inp[6]) ? node1681 : 8'b10110100;
													assign node1681 = (inp[12]) ? 8'b10100101 : 8'b10110100;
									assign node1685 = (inp[11]) ? node1693 : node1686;
										assign node1686 = (inp[2]) ? 8'b10011101 : node1687;
											assign node1687 = (inp[12]) ? 8'b10000100 : node1688;
												assign node1688 = (inp[3]) ? 8'b10001101 : 8'b10011100;
										assign node1693 = (inp[12]) ? 8'b10100100 : node1694;
											assign node1694 = (inp[6]) ? node1696 : 8'b10111100;
												assign node1696 = (inp[3]) ? 8'b10101101 : 8'b10101100;
								assign node1700 = (inp[3]) ? node1716 : node1701;
									assign node1701 = (inp[12]) ? node1707 : node1702;
										assign node1702 = (inp[11]) ? 8'b10100100 : node1703;
											assign node1703 = (inp[1]) ? 8'b10000001 : 8'b10010000;
										assign node1707 = (inp[1]) ? node1713 : node1708;
											assign node1708 = (inp[2]) ? 8'b00000010 : node1709;
												assign node1709 = (inp[6]) ? 8'b00011010 : 8'b00000010;
											assign node1713 = (inp[2]) ? 8'b10010001 : 8'b00001011;
									assign node1716 = (inp[11]) ? node1720 : node1717;
										assign node1717 = (inp[6]) ? 8'b00001110 : 8'b00011110;
										assign node1720 = (inp[2]) ? 8'b00001011 : node1721;
											assign node1721 = (inp[8]) ? 8'b00001010 : 8'b00001110;
					assign node1725 = (inp[3]) ? node1819 : node1726;
						assign node1726 = (inp[8]) ? node1772 : node1727;
							assign node1727 = (inp[10]) ? node1749 : node1728;
								assign node1728 = (inp[6]) ? node1738 : node1729;
									assign node1729 = (inp[9]) ? node1733 : node1730;
										assign node1730 = (inp[12]) ? 8'b00000010 : 8'b10010100;
										assign node1733 = (inp[11]) ? node1735 : 8'b10100001;
											assign node1735 = (inp[0]) ? 8'b10000101 : 8'b10010101;
									assign node1738 = (inp[2]) ? node1744 : node1739;
										assign node1739 = (inp[1]) ? 8'b10111001 : node1740;
											assign node1740 = (inp[12]) ? 8'b10111000 : 8'b10101000;
										assign node1744 = (inp[9]) ? 8'b10110000 : node1745;
											assign node1745 = (inp[0]) ? 8'b10110001 : 8'b10010000;
								assign node1749 = (inp[9]) ? node1763 : node1750;
									assign node1750 = (inp[0]) ? node1754 : node1751;
										assign node1751 = (inp[11]) ? 8'b00011110 : 8'b00001110;
										assign node1754 = (inp[1]) ? node1760 : node1755;
											assign node1755 = (inp[12]) ? node1757 : 8'b10101100;
												assign node1757 = (inp[6]) ? 8'b10111100 : 8'b10101100;
											assign node1760 = (inp[12]) ? 8'b11111101 : 8'b10101001;
									assign node1763 = (inp[11]) ? node1767 : node1764;
										assign node1764 = (inp[2]) ? 8'b10101100 : 8'b10101101;
										assign node1767 = (inp[6]) ? node1769 : 8'b10111001;
											assign node1769 = (inp[12]) ? 8'b10111001 : 8'b10101001;
							assign node1772 = (inp[2]) ? node1794 : node1773;
								assign node1773 = (inp[6]) ? node1787 : node1774;
									assign node1774 = (inp[12]) ? node1784 : node1775;
										assign node1775 = (inp[1]) ? node1781 : node1776;
											assign node1776 = (inp[0]) ? 8'b10010001 : node1777;
												assign node1777 = (inp[10]) ? 8'b10010001 : 8'b11110111;
											assign node1781 = (inp[0]) ? 8'b10010000 : 8'b10010001;
										assign node1784 = (inp[9]) ? 8'b10100101 : 8'b00000010;
									assign node1787 = (inp[12]) ? node1789 : 8'b00001010;
										assign node1789 = (inp[10]) ? node1791 : 8'b10011001;
											assign node1791 = (inp[9]) ? 8'b10011100 : 8'b10111100;
								assign node1794 = (inp[1]) ? node1810 : node1795;
									assign node1795 = (inp[11]) ? node1801 : node1796;
										assign node1796 = (inp[9]) ? 8'b10110000 : node1797;
											assign node1797 = (inp[0]) ? 8'b10110100 : 8'b10000100;
										assign node1801 = (inp[12]) ? 8'b10100000 : node1802;
											assign node1802 = (inp[10]) ? node1806 : node1803;
												assign node1803 = (inp[0]) ? 8'b10000001 : 8'b10010101;
												assign node1806 = (inp[6]) ? 8'b10100001 : 8'b10110001;
									assign node1810 = (inp[0]) ? node1816 : node1811;
										assign node1811 = (inp[6]) ? 8'b11110101 : node1812;
											assign node1812 = (inp[11]) ? 8'b10010101 : 8'b10000100;
										assign node1816 = (inp[11]) ? 8'b10010000 : 8'b11110101;
						assign node1819 = (inp[6]) ? node1869 : node1820;
							assign node1820 = (inp[1]) ? node1848 : node1821;
								assign node1821 = (inp[9]) ? node1835 : node1822;
									assign node1822 = (inp[0]) ? node1830 : node1823;
										assign node1823 = (inp[10]) ? node1827 : node1824;
											assign node1824 = (inp[8]) ? 8'b00011010 : 8'b00001011;
											assign node1827 = (inp[8]) ? 8'b10001101 : 8'b00001111;
										assign node1830 = (inp[2]) ? 8'b11111101 : node1831;
											assign node1831 = (inp[12]) ? 8'b10001101 : 8'b10101101;
									assign node1835 = (inp[10]) ? node1841 : node1836;
										assign node1836 = (inp[0]) ? node1838 : 8'b10101001;
											assign node1838 = (inp[2]) ? 8'b10011100 : 8'b10101001;
										assign node1841 = (inp[8]) ? node1845 : node1842;
											assign node1842 = (inp[2]) ? 8'b11111101 : 8'b10101101;
											assign node1845 = (inp[12]) ? 8'b10001101 : 8'b10101101;
								assign node1848 = (inp[10]) ? node1858 : node1849;
									assign node1849 = (inp[11]) ? 8'b10110100 : node1850;
										assign node1850 = (inp[9]) ? node1852 : 8'b10000001;
											assign node1852 = (inp[0]) ? node1854 : 8'b10100001;
												assign node1854 = (inp[2]) ? 8'b10110001 : 8'b10100101;
									assign node1858 = (inp[11]) ? node1866 : node1859;
										assign node1859 = (inp[2]) ? 8'b11111101 : node1860;
											assign node1860 = (inp[12]) ? 8'b10000101 : node1861;
												assign node1861 = (inp[8]) ? 8'b10100101 : 8'b10101101;
										assign node1866 = (inp[0]) ? 8'b10101000 : 8'b10101001;
							assign node1869 = (inp[11]) ? node1885 : node1870;
								assign node1870 = (inp[0]) ? node1878 : node1871;
									assign node1871 = (inp[10]) ? node1875 : node1872;
										assign node1872 = (inp[1]) ? 8'b10011001 : 8'b10111001;
										assign node1875 = (inp[9]) ? 8'b11111101 : 8'b10011101;
									assign node1878 = (inp[2]) ? node1880 : 8'b11111101;
										assign node1880 = (inp[10]) ? 8'b11111101 : node1881;
											assign node1881 = (inp[8]) ? 8'b11111101 : 8'b10111001;
								assign node1885 = (inp[12]) ? node1893 : node1886;
									assign node1886 = (inp[1]) ? 8'b10000000 : node1887;
										assign node1887 = (inp[10]) ? node1889 : 8'b10001101;
											assign node1889 = (inp[9]) ? 8'b10101100 : 8'b10001100;
									assign node1893 = (inp[2]) ? node1897 : node1894;
										assign node1894 = (inp[1]) ? 8'b10011101 : 8'b10111001;
										assign node1897 = (inp[1]) ? 8'b10110100 : node1898;
											assign node1898 = (inp[0]) ? node1900 : 8'b00011010;
												assign node1900 = (inp[8]) ? 8'b10011100 : node1901;
													assign node1901 = (inp[10]) ? 8'b10111100 : 8'b10111000;
			assign node1906 = (inp[12]) ? node2148 : node1907;
				assign node1907 = (inp[11]) ? node2013 : node1908;
					assign node1908 = (inp[1]) ? node1966 : node1909;
						assign node1909 = (inp[13]) ? node1933 : node1910;
							assign node1910 = (inp[8]) ? node1922 : node1911;
								assign node1911 = (inp[2]) ? node1913 : 8'b10000010;
									assign node1913 = (inp[9]) ? node1915 : 8'b10000010;
										assign node1915 = (inp[5]) ? node1919 : node1916;
											assign node1916 = (inp[6]) ? 8'b10000010 : 8'b10010000;
											assign node1919 = (inp[6]) ? 8'b10010000 : 8'b10000010;
								assign node1922 = (inp[2]) ? node1930 : node1923;
									assign node1923 = (inp[6]) ? 8'b10000010 : node1924;
										assign node1924 = (inp[9]) ? 8'b10000100 : node1925;
											assign node1925 = (inp[0]) ? 8'b10000100 : 8'b10000010;
									assign node1930 = (inp[0]) ? 8'b10010100 : 8'b10000100;
							assign node1933 = (inp[5]) ? node1947 : node1934;
								assign node1934 = (inp[0]) ? node1936 : 8'b10000010;
									assign node1936 = (inp[9]) ? node1938 : 8'b10100000;
										assign node1938 = (inp[10]) ? node1942 : node1939;
											assign node1939 = (inp[8]) ? 8'b10000100 : 8'b10000010;
											assign node1942 = (inp[8]) ? 8'b10000010 : node1943;
												assign node1943 = (inp[6]) ? 8'b10000010 : 8'b10010000;
								assign node1947 = (inp[2]) ? node1955 : node1948;
									assign node1948 = (inp[0]) ? node1952 : node1949;
										assign node1949 = (inp[10]) ? 8'b10000100 : 8'b10000010;
										assign node1952 = (inp[8]) ? 8'b10100100 : 8'b10100000;
									assign node1955 = (inp[8]) ? node1961 : node1956;
										assign node1956 = (inp[0]) ? 8'b10110000 : node1957;
											assign node1957 = (inp[6]) ? 8'b10110000 : 8'b10100000;
										assign node1961 = (inp[10]) ? 8'b10010100 : node1962;
											assign node1962 = (inp[0]) ? 8'b10110100 : 8'b10110000;
						assign node1966 = (inp[5]) ? node1984 : node1967;
							assign node1967 = (inp[0]) ? node1969 : 8'b10000010;
								assign node1969 = (inp[3]) ? node1981 : node1970;
									assign node1970 = (inp[10]) ? node1976 : node1971;
										assign node1971 = (inp[2]) ? 8'b10010101 : node1972;
											assign node1972 = (inp[8]) ? 8'b10000101 : 8'b10000001;
										assign node1976 = (inp[13]) ? node1978 : 8'b10000001;
											assign node1978 = (inp[2]) ? 8'b10000001 : 8'b10100001;
									assign node1981 = (inp[9]) ? 8'b10000010 : 8'b10100000;
							assign node1984 = (inp[13]) ? node2002 : node1985;
								assign node1985 = (inp[2]) ? node1995 : node1986;
									assign node1986 = (inp[8]) ? node1992 : node1987;
										assign node1987 = (inp[0]) ? 8'b10000001 : node1988;
											assign node1988 = (inp[3]) ? 8'b10000001 : 8'b10000010;
										assign node1992 = (inp[10]) ? 8'b10000101 : 8'b10000001;
									assign node1995 = (inp[6]) ? node1997 : 8'b10000010;
										assign node1997 = (inp[0]) ? 8'b10010101 : node1998;
											assign node1998 = (inp[3]) ? 8'b10010001 : 8'b10010000;
								assign node2002 = (inp[0]) ? node2008 : node2003;
									assign node2003 = (inp[9]) ? node2005 : 8'b10000001;
										assign node2005 = (inp[2]) ? 8'b10100000 : 8'b10100001;
									assign node2008 = (inp[8]) ? node2010 : 8'b10110001;
										assign node2010 = (inp[2]) ? 8'b11110101 : 8'b10100101;
					assign node2013 = (inp[0]) ? node2061 : node2014;
						assign node2014 = (inp[5]) ? node2016 : 8'b11110111;
							assign node2016 = (inp[2]) ? node2042 : node2017;
								assign node2017 = (inp[10]) ? node2029 : node2018;
									assign node2018 = (inp[9]) ? node2024 : node2019;
										assign node2019 = (inp[1]) ? node2021 : 8'b11110111;
											assign node2021 = (inp[3]) ? 8'b10110100 : 8'b11110111;
										assign node2024 = (inp[13]) ? node2026 : 8'b11110111;
											assign node2026 = (inp[3]) ? 8'b10010100 : 8'b10010101;
									assign node2029 = (inp[8]) ? node2037 : node2030;
										assign node2030 = (inp[3]) ? node2032 : 8'b11110111;
											assign node2032 = (inp[9]) ? node2034 : 8'b10110100;
												assign node2034 = (inp[1]) ? 8'b10010100 : 8'b10010101;
										assign node2037 = (inp[1]) ? 8'b10110000 : node2038;
											assign node2038 = (inp[13]) ? 8'b10010001 : 8'b10110001;
								assign node2042 = (inp[6]) ? node2050 : node2043;
									assign node2043 = (inp[1]) ? node2045 : 8'b11110111;
										assign node2045 = (inp[13]) ? node2047 : 8'b10110100;
											assign node2047 = (inp[9]) ? 8'b10010100 : 8'b10110100;
									assign node2050 = (inp[9]) ? node2058 : node2051;
										assign node2051 = (inp[10]) ? node2055 : node2052;
											assign node2052 = (inp[1]) ? 8'b10100100 : 8'b10100101;
											assign node2055 = (inp[1]) ? 8'b10100000 : 8'b10100001;
										assign node2058 = (inp[13]) ? 8'b10000101 : 8'b10100101;
						assign node2061 = (inp[1]) ? node2091 : node2062;
							assign node2062 = (inp[2]) ? node2078 : node2063;
								assign node2063 = (inp[8]) ? node2069 : node2064;
									assign node2064 = (inp[13]) ? node2066 : 8'b11110111;
										assign node2066 = (inp[5]) ? 8'b10010101 : 8'b11110111;
									assign node2069 = (inp[13]) ? node2073 : node2070;
										assign node2070 = (inp[10]) ? 8'b11110111 : 8'b10110001;
										assign node2073 = (inp[10]) ? node2075 : 8'b10010001;
											assign node2075 = (inp[5]) ? 8'b10010001 : 8'b10010101;
								assign node2078 = (inp[5]) ? node2086 : node2079;
									assign node2079 = (inp[6]) ? node2081 : 8'b10100101;
										assign node2081 = (inp[10]) ? 8'b11110111 : node2082;
											assign node2082 = (inp[3]) ? 8'b11110111 : 8'b10110001;
									assign node2086 = (inp[8]) ? 8'b10100001 : node2087;
										assign node2087 = (inp[13]) ? 8'b10000101 : 8'b10100101;
							assign node2091 = (inp[13]) ? node2121 : node2092;
								assign node2092 = (inp[2]) ? node2102 : node2093;
									assign node2093 = (inp[6]) ? 8'b10110001 : node2094;
										assign node2094 = (inp[5]) ? node2098 : node2095;
											assign node2095 = (inp[3]) ? 8'b11110111 : 8'b10110100;
											assign node2098 = (inp[8]) ? 8'b10110000 : 8'b10110100;
									assign node2102 = (inp[8]) ? node2112 : node2103;
										assign node2103 = (inp[10]) ? node2105 : 8'b10100100;
											assign node2105 = (inp[3]) ? node2109 : node2106;
												assign node2106 = (inp[6]) ? 8'b10110100 : 8'b10100100;
												assign node2109 = (inp[5]) ? 8'b10100100 : 8'b11110111;
										assign node2112 = (inp[10]) ? node2118 : node2113;
											assign node2113 = (inp[3]) ? 8'b10100001 : node2114;
												assign node2114 = (inp[6]) ? 8'b10110000 : 8'b10100000;
											assign node2118 = (inp[5]) ? 8'b10100000 : 8'b10100100;
								assign node2121 = (inp[5]) ? node2141 : node2122;
									assign node2122 = (inp[9]) ? node2132 : node2123;
										assign node2123 = (inp[10]) ? node2129 : node2124;
											assign node2124 = (inp[3]) ? 8'b10010001 : node2125;
												assign node2125 = (inp[2]) ? 8'b10000000 : 8'b10010000;
											assign node2129 = (inp[3]) ? 8'b10010101 : 8'b10010100;
										assign node2132 = (inp[3]) ? node2138 : node2133;
											assign node2133 = (inp[2]) ? node2135 : 8'b10110100;
												assign node2135 = (inp[10]) ? 8'b10110100 : 8'b10100000;
											assign node2138 = (inp[10]) ? 8'b11110111 : 8'b10100001;
									assign node2141 = (inp[8]) ? node2145 : node2142;
										assign node2142 = (inp[2]) ? 8'b10000100 : 8'b10010100;
										assign node2145 = (inp[3]) ? 8'b10000000 : 8'b10010000;
				assign node2148 = (inp[0]) ? node2208 : node2149;
					assign node2149 = (inp[5]) ? node2151 : 8'b00000010;
						assign node2151 = (inp[3]) ? node2181 : node2152;
							assign node2152 = (inp[6]) ? node2162 : node2153;
								assign node2153 = (inp[10]) ? node2159 : node2154;
									assign node2154 = (inp[1]) ? 8'b00000010 : node2155;
										assign node2155 = (inp[9]) ? 8'b10100000 : 8'b00000010;
									assign node2159 = (inp[8]) ? 8'b10000100 : 8'b00000010;
								assign node2162 = (inp[2]) ? node2176 : node2163;
									assign node2163 = (inp[9]) ? node2169 : node2164;
										assign node2164 = (inp[10]) ? node2166 : 8'b00000010;
											assign node2166 = (inp[13]) ? 8'b00000010 : 8'b10000100;
										assign node2169 = (inp[10]) ? node2171 : 8'b10100000;
											assign node2171 = (inp[8]) ? node2173 : 8'b10100000;
												assign node2173 = (inp[13]) ? 8'b10000100 : 8'b10100100;
									assign node2176 = (inp[11]) ? 8'b11110101 : node2177;
										assign node2177 = (inp[13]) ? 8'b10110000 : 8'b10010000;
							assign node2181 = (inp[1]) ? node2189 : node2182;
								assign node2182 = (inp[11]) ? node2186 : node2183;
									assign node2183 = (inp[6]) ? 8'b10010000 : 8'b10100000;
									assign node2186 = (inp[10]) ? 8'b10110001 : 8'b00000010;
								assign node2189 = (inp[11]) ? node2199 : node2190;
									assign node2190 = (inp[8]) ? 8'b10000101 : node2191;
										assign node2191 = (inp[2]) ? node2195 : node2192;
											assign node2192 = (inp[9]) ? 8'b10100001 : 8'b10000001;
											assign node2195 = (inp[13]) ? 8'b10000001 : 8'b10010001;
									assign node2199 = (inp[2]) ? node2205 : node2200;
										assign node2200 = (inp[13]) ? node2202 : 8'b10100101;
											assign node2202 = (inp[6]) ? 8'b10000001 : 8'b10100001;
										assign node2205 = (inp[6]) ? 8'b10110100 : 8'b10100101;
					assign node2208 = (inp[2]) ? node2270 : node2209;
						assign node2209 = (inp[5]) ? node2233 : node2210;
							assign node2210 = (inp[8]) ? node2222 : node2211;
								assign node2211 = (inp[3]) ? node2217 : node2212;
									assign node2212 = (inp[1]) ? node2214 : 8'b00000010;
										assign node2214 = (inp[13]) ? 8'b10100101 : 8'b10000001;
									assign node2217 = (inp[9]) ? 8'b00000010 : node2218;
										assign node2218 = (inp[13]) ? 8'b10100000 : 8'b00000010;
								assign node2222 = (inp[10]) ? node2228 : node2223;
									assign node2223 = (inp[9]) ? node2225 : 8'b10100100;
										assign node2225 = (inp[11]) ? 8'b10100100 : 8'b10000100;
									assign node2228 = (inp[3]) ? 8'b10100000 : node2229;
										assign node2229 = (inp[1]) ? 8'b10000001 : 8'b00000010;
							assign node2233 = (inp[1]) ? node2245 : node2234;
								assign node2234 = (inp[8]) ? node2238 : node2235;
									assign node2235 = (inp[13]) ? 8'b10100000 : 8'b00000010;
									assign node2238 = (inp[10]) ? 8'b10000100 : node2239;
										assign node2239 = (inp[11]) ? node2241 : 8'b10100100;
											assign node2241 = (inp[13]) ? 8'b10000100 : 8'b10100100;
								assign node2245 = (inp[6]) ? node2257 : node2246;
									assign node2246 = (inp[3]) ? node2252 : node2247;
										assign node2247 = (inp[11]) ? node2249 : 8'b10000101;
											assign node2249 = (inp[8]) ? 8'b10000001 : 8'b10000101;
										assign node2252 = (inp[8]) ? 8'b10100101 : node2253;
											assign node2253 = (inp[13]) ? 8'b10000101 : 8'b10100101;
									assign node2257 = (inp[13]) ? node2263 : node2258;
										assign node2258 = (inp[11]) ? 8'b10100001 : node2259;
											assign node2259 = (inp[8]) ? 8'b10000101 : 8'b10000001;
										assign node2263 = (inp[11]) ? node2267 : node2264;
											assign node2264 = (inp[10]) ? 8'b10100101 : 8'b10100001;
											assign node2267 = (inp[8]) ? 8'b10000001 : 8'b10000101;
						assign node2270 = (inp[6]) ? node2306 : node2271;
							assign node2271 = (inp[11]) ? node2289 : node2272;
								assign node2272 = (inp[13]) ? node2284 : node2273;
									assign node2273 = (inp[1]) ? node2279 : node2274;
										assign node2274 = (inp[10]) ? 8'b10010000 : node2275;
											assign node2275 = (inp[8]) ? 8'b10010100 : 8'b10010000;
										assign node2279 = (inp[8]) ? 8'b10010101 : node2280;
											assign node2280 = (inp[3]) ? 8'b10010000 : 8'b10010001;
									assign node2284 = (inp[1]) ? 8'b11110101 : node2285;
										assign node2285 = (inp[8]) ? 8'b10110100 : 8'b10110000;
								assign node2289 = (inp[9]) ? node2295 : node2290;
									assign node2290 = (inp[3]) ? 8'b10110100 : node2291;
										assign node2291 = (inp[5]) ? 8'b10010000 : 8'b10010101;
									assign node2295 = (inp[3]) ? node2301 : node2296;
										assign node2296 = (inp[1]) ? node2298 : 8'b11110101;
											assign node2298 = (inp[10]) ? 8'b10110000 : 8'b10110100;
										assign node2301 = (inp[10]) ? 8'b11110101 : node2302;
											assign node2302 = (inp[8]) ? 8'b10110001 : 8'b11110101;
							assign node2306 = (inp[5]) ? node2334 : node2307;
								assign node2307 = (inp[3]) ? node2325 : node2308;
									assign node2308 = (inp[1]) ? node2316 : node2309;
										assign node2309 = (inp[8]) ? node2311 : 8'b00000010;
											assign node2311 = (inp[10]) ? 8'b10100000 : node2312;
												assign node2312 = (inp[13]) ? 8'b10100100 : 8'b10000100;
										assign node2316 = (inp[8]) ? node2320 : node2317;
											assign node2317 = (inp[13]) ? 8'b10000101 : 8'b10000001;
											assign node2320 = (inp[13]) ? 8'b10100101 : node2321;
												assign node2321 = (inp[9]) ? 8'b10100101 : 8'b10000101;
									assign node2325 = (inp[13]) ? node2327 : 8'b00000010;
										assign node2327 = (inp[9]) ? 8'b00000010 : node2328;
											assign node2328 = (inp[11]) ? 8'b10100000 : node2329;
												assign node2329 = (inp[10]) ? 8'b10100000 : 8'b10100100;
								assign node2334 = (inp[11]) ? node2344 : node2335;
									assign node2335 = (inp[1]) ? node2341 : node2336;
										assign node2336 = (inp[8]) ? 8'b10010100 : node2337;
											assign node2337 = (inp[9]) ? 8'b10010000 : 8'b10110000;
										assign node2341 = (inp[10]) ? 8'b10010101 : 8'b10010001;
									assign node2344 = (inp[13]) ? 8'b10010101 : node2345;
										assign node2345 = (inp[9]) ? node2347 : 8'b10110100;
											assign node2347 = (inp[1]) ? 8'b10110000 : 8'b10110001;

endmodule