module dtc_split125_bm47 (
	input  wire [16-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node6;
	wire [1-1:0] node7;
	wire [1-1:0] node8;
	wire [1-1:0] node9;
	wire [1-1:0] node10;
	wire [1-1:0] node14;
	wire [1-1:0] node15;
	wire [1-1:0] node19;
	wire [1-1:0] node21;
	wire [1-1:0] node25;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node28;
	wire [1-1:0] node29;
	wire [1-1:0] node31;
	wire [1-1:0] node34;
	wire [1-1:0] node36;
	wire [1-1:0] node39;
	wire [1-1:0] node41;
	wire [1-1:0] node44;
	wire [1-1:0] node46;
	wire [1-1:0] node47;
	wire [1-1:0] node48;
	wire [1-1:0] node50;
	wire [1-1:0] node53;
	wire [1-1:0] node55;
	wire [1-1:0] node58;
	wire [1-1:0] node59;
	wire [1-1:0] node63;
	wire [1-1:0] node64;
	wire [1-1:0] node66;
	wire [1-1:0] node67;
	wire [1-1:0] node68;
	wire [1-1:0] node69;
	wire [1-1:0] node73;
	wire [1-1:0] node74;
	wire [1-1:0] node78;
	wire [1-1:0] node79;
	wire [1-1:0] node84;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node87;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node90;
	wire [1-1:0] node91;
	wire [1-1:0] node93;
	wire [1-1:0] node94;
	wire [1-1:0] node96;
	wire [1-1:0] node99;
	wire [1-1:0] node100;
	wire [1-1:0] node105;
	wire [1-1:0] node107;
	wire [1-1:0] node110;
	wire [1-1:0] node111;
	wire [1-1:0] node113;
	wire [1-1:0] node114;
	wire [1-1:0] node118;
	wire [1-1:0] node119;
	wire [1-1:0] node121;
	wire [1-1:0] node125;
	wire [1-1:0] node126;
	wire [1-1:0] node127;
	wire [1-1:0] node129;
	wire [1-1:0] node130;
	wire [1-1:0] node135;
	wire [1-1:0] node136;
	wire [1-1:0] node137;
	wire [1-1:0] node138;
	wire [1-1:0] node141;
	wire [1-1:0] node144;
	wire [1-1:0] node146;
	wire [1-1:0] node149;
	wire [1-1:0] node151;
	wire [1-1:0] node152;
	wire [1-1:0] node156;
	wire [1-1:0] node157;
	wire [1-1:0] node158;
	wire [1-1:0] node160;
	wire [1-1:0] node161;
	wire [1-1:0] node163;
	wire [1-1:0] node166;
	wire [1-1:0] node167;
	wire [1-1:0] node169;
	wire [1-1:0] node174;
	wire [1-1:0] node175;
	wire [1-1:0] node176;
	wire [1-1:0] node177;
	wire [1-1:0] node178;
	wire [1-1:0] node183;
	wire [1-1:0] node184;
	wire [1-1:0] node186;
	wire [1-1:0] node189;
	wire [1-1:0] node191;
	wire [1-1:0] node192;
	wire [1-1:0] node194;
	wire [1-1:0] node198;
	wire [1-1:0] node199;
	wire [1-1:0] node201;
	wire [1-1:0] node202;
	wire [1-1:0] node207;
	wire [1-1:0] node208;
	wire [1-1:0] node209;
	wire [1-1:0] node211;
	wire [1-1:0] node212;
	wire [1-1:0] node213;
	wire [1-1:0] node214;
	wire [1-1:0] node218;
	wire [1-1:0] node219;
	wire [1-1:0] node224;
	wire [1-1:0] node225;
	wire [1-1:0] node226;
	wire [1-1:0] node228;
	wire [1-1:0] node230;
	wire [1-1:0] node233;
	wire [1-1:0] node235;
	wire [1-1:0] node238;
	wire [1-1:0] node239;
	wire [1-1:0] node240;
	wire [1-1:0] node242;
	wire [1-1:0] node244;
	wire [1-1:0] node248;
	wire [1-1:0] node249;
	wire [1-1:0] node251;
	wire [1-1:0] node253;
	wire [1-1:0] node257;
	wire [1-1:0] node258;
	wire [1-1:0] node259;
	wire [1-1:0] node260;
	wire [1-1:0] node261;
	wire [1-1:0] node262;
	wire [1-1:0] node263;
	wire [1-1:0] node266;
	wire [1-1:0] node267;
	wire [1-1:0] node272;
	wire [1-1:0] node273;
	wire [1-1:0] node274;
	wire [1-1:0] node277;
	wire [1-1:0] node281;
	wire [1-1:0] node283;
	wire [1-1:0] node285;
	wire [1-1:0] node288;
	wire [1-1:0] node290;
	wire [1-1:0] node291;
	wire [1-1:0] node292;
	wire [1-1:0] node297;
	wire [1-1:0] node298;
	wire [1-1:0] node300;
	wire [1-1:0] node301;
	wire [1-1:0] node305;
	wire [1-1:0] node306;
	wire [1-1:0] node307;
	wire [1-1:0] node309;
	wire [1-1:0] node311;
	wire [1-1:0] node314;
	wire [1-1:0] node315;
	wire [1-1:0] node317;
	wire [1-1:0] node321;
	wire [1-1:0] node322;
	wire [1-1:0] node326;
	wire [1-1:0] node327;
	wire [1-1:0] node328;
	wire [1-1:0] node330;
	wire [1-1:0] node331;
	wire [1-1:0] node332;
	wire [1-1:0] node333;
	wire [1-1:0] node334;
	wire [1-1:0] node338;
	wire [1-1:0] node339;
	wire [1-1:0] node343;
	wire [1-1:0] node345;
	wire [1-1:0] node349;
	wire [1-1:0] node350;
	wire [1-1:0] node351;
	wire [1-1:0] node352;
	wire [1-1:0] node353;
	wire [1-1:0] node354;
	wire [1-1:0] node355;
	wire [1-1:0] node358;
	wire [1-1:0] node362;
	wire [1-1:0] node363;
	wire [1-1:0] node364;
	wire [1-1:0] node369;
	wire [1-1:0] node370;
	wire [1-1:0] node374;
	wire [1-1:0] node376;
	wire [1-1:0] node377;
	wire [1-1:0] node379;
	wire [1-1:0] node382;
	wire [1-1:0] node383;
	wire [1-1:0] node385;
	wire [1-1:0] node388;
	wire [1-1:0] node390;
	wire [1-1:0] node391;
	wire [1-1:0] node394;
	wire [1-1:0] node397;
	wire [1-1:0] node398;
	wire [1-1:0] node400;
	wire [1-1:0] node401;
	wire [1-1:0] node403;
	wire [1-1:0] node405;
	wire [1-1:0] node408;
	wire [1-1:0] node409;
	wire [1-1:0] node410;
	wire [1-1:0] node412;
	wire [1-1:0] node418;
	wire [1-1:0] node419;
	wire [1-1:0] node420;
	wire [1-1:0] node421;
	wire [1-1:0] node423;
	wire [1-1:0] node424;
	wire [1-1:0] node425;
	wire [1-1:0] node426;
	wire [1-1:0] node432;
	wire [1-1:0] node433;
	wire [1-1:0] node434;
	wire [1-1:0] node435;
	wire [1-1:0] node436;
	wire [1-1:0] node439;
	wire [1-1:0] node444;
	wire [1-1:0] node446;
	wire [1-1:0] node447;
	wire [1-1:0] node449;
	wire [1-1:0] node451;
	wire [1-1:0] node454;
	wire [1-1:0] node457;
	wire [1-1:0] node459;
	wire [1-1:0] node460;
	wire [1-1:0] node461;
	wire [1-1:0] node463;
	wire [1-1:0] node465;
	wire [1-1:0] node468;
	wire [1-1:0] node472;
	wire [1-1:0] node473;
	wire [1-1:0] node475;
	wire [1-1:0] node476;
	wire [1-1:0] node477;
	wire [1-1:0] node478;
	wire [1-1:0] node479;
	wire [1-1:0] node482;
	wire [1-1:0] node483;
	wire [1-1:0] node488;
	wire [1-1:0] node490;
	wire [1-1:0] node494;
	wire [1-1:0] node495;
	wire [1-1:0] node496;
	wire [1-1:0] node498;
	wire [1-1:0] node499;
	wire [1-1:0] node500;
	wire [1-1:0] node502;
	wire [1-1:0] node507;
	wire [1-1:0] node508;
	wire [1-1:0] node512;
	wire [1-1:0] node513;
	wire [1-1:0] node514;
	wire [1-1:0] node515;
	wire [1-1:0] node516;
	wire [1-1:0] node518;
	wire [1-1:0] node523;
	wire [1-1:0] node526;
	wire [1-1:0] node528;
	wire [1-1:0] node531;
	wire [1-1:0] node532;
	wire [1-1:0] node534;
	wire [1-1:0] node535;
	wire [1-1:0] node536;
	wire [1-1:0] node537;
	wire [1-1:0] node538;
	wire [1-1:0] node542;
	wire [1-1:0] node544;
	wire [1-1:0] node547;
	wire [1-1:0] node549;
	wire [1-1:0] node553;
	wire [1-1:0] node554;
	wire [1-1:0] node555;
	wire [1-1:0] node556;
	wire [1-1:0] node557;
	wire [1-1:0] node558;
	wire [1-1:0] node562;
	wire [1-1:0] node564;
	wire [1-1:0] node567;
	wire [1-1:0] node569;
	wire [1-1:0] node572;
	wire [1-1:0] node574;
	wire [1-1:0] node575;
	wire [1-1:0] node576;
	wire [1-1:0] node578;
	wire [1-1:0] node581;
	wire [1-1:0] node583;
	wire [1-1:0] node586;
	wire [1-1:0] node588;
	wire [1-1:0] node591;
	wire [1-1:0] node592;
	wire [1-1:0] node594;
	wire [1-1:0] node595;
	wire [1-1:0] node596;
	wire [1-1:0] node597;
	wire [1-1:0] node601;
	wire [1-1:0] node603;
	wire [1-1:0] node606;
	wire [1-1:0] node608;
	wire [1-1:0] node612;
	wire [1-1:0] node613;
	wire [1-1:0] node614;
	wire [1-1:0] node615;
	wire [1-1:0] node616;
	wire [1-1:0] node617;
	wire [1-1:0] node618;
	wire [1-1:0] node619;
	wire [1-1:0] node621;
	wire [1-1:0] node622;
	wire [1-1:0] node623;
	wire [1-1:0] node627;
	wire [1-1:0] node629;
	wire [1-1:0] node633;
	wire [1-1:0] node634;
	wire [1-1:0] node635;
	wire [1-1:0] node637;
	wire [1-1:0] node641;
	wire [1-1:0] node642;
	wire [1-1:0] node643;
	wire [1-1:0] node644;
	wire [1-1:0] node645;
	wire [1-1:0] node648;
	wire [1-1:0] node649;
	wire [1-1:0] node654;
	wire [1-1:0] node655;
	wire [1-1:0] node659;
	wire [1-1:0] node661;
	wire [1-1:0] node664;
	wire [1-1:0] node665;
	wire [1-1:0] node667;
	wire [1-1:0] node668;
	wire [1-1:0] node670;
	wire [1-1:0] node673;
	wire [1-1:0] node674;
	wire [1-1:0] node675;
	wire [1-1:0] node679;
	wire [1-1:0] node680;
	wire [1-1:0] node685;
	wire [1-1:0] node686;
	wire [1-1:0] node687;
	wire [1-1:0] node688;
	wire [1-1:0] node689;
	wire [1-1:0] node691;
	wire [1-1:0] node694;
	wire [1-1:0] node695;
	wire [1-1:0] node696;
	wire [1-1:0] node697;
	wire [1-1:0] node698;
	wire [1-1:0] node704;
	wire [1-1:0] node705;
	wire [1-1:0] node709;
	wire [1-1:0] node710;
	wire [1-1:0] node712;
	wire [1-1:0] node713;
	wire [1-1:0] node715;
	wire [1-1:0] node718;
	wire [1-1:0] node721;
	wire [1-1:0] node722;
	wire [1-1:0] node724;
	wire [1-1:0] node725;
	wire [1-1:0] node729;
	wire [1-1:0] node730;
	wire [1-1:0] node732;
	wire [1-1:0] node733;
	wire [1-1:0] node737;
	wire [1-1:0] node739;
	wire [1-1:0] node741;
	wire [1-1:0] node744;
	wire [1-1:0] node745;
	wire [1-1:0] node747;
	wire [1-1:0] node748;
	wire [1-1:0] node751;
	wire [1-1:0] node753;
	wire [1-1:0] node757;
	wire [1-1:0] node758;
	wire [1-1:0] node760;
	wire [1-1:0] node761;
	wire [1-1:0] node762;
	wire [1-1:0] node764;
	wire [1-1:0] node766;
	wire [1-1:0] node767;
	wire [1-1:0] node773;
	wire [1-1:0] node774;
	wire [1-1:0] node775;
	wire [1-1:0] node776;
	wire [1-1:0] node777;
	wire [1-1:0] node778;
	wire [1-1:0] node784;
	wire [1-1:0] node785;
	wire [1-1:0] node787;
	wire [1-1:0] node790;
	wire [1-1:0] node791;
	wire [1-1:0] node795;
	wire [1-1:0] node797;
	wire [1-1:0] node798;
	wire [1-1:0] node799;
	wire [1-1:0] node801;
	wire [1-1:0] node802;
	wire [1-1:0] node805;
	wire [1-1:0] node810;
	wire [1-1:0] node811;
	wire [1-1:0] node812;
	wire [1-1:0] node813;
	wire [1-1:0] node814;
	wire [1-1:0] node815;
	wire [1-1:0] node817;
	wire [1-1:0] node820;
	wire [1-1:0] node821;
	wire [1-1:0] node822;
	wire [1-1:0] node823;
	wire [1-1:0] node825;
	wire [1-1:0] node830;
	wire [1-1:0] node831;
	wire [1-1:0] node833;
	wire [1-1:0] node837;
	wire [1-1:0] node838;
	wire [1-1:0] node840;
	wire [1-1:0] node842;
	wire [1-1:0] node846;
	wire [1-1:0] node847;
	wire [1-1:0] node848;
	wire [1-1:0] node849;
	wire [1-1:0] node850;
	wire [1-1:0] node852;
	wire [1-1:0] node856;
	wire [1-1:0] node857;
	wire [1-1:0] node860;
	wire [1-1:0] node862;
	wire [1-1:0] node865;
	wire [1-1:0] node866;
	wire [1-1:0] node868;
	wire [1-1:0] node870;
	wire [1-1:0] node874;
	wire [1-1:0] node875;
	wire [1-1:0] node877;
	wire [1-1:0] node878;
	wire [1-1:0] node882;
	wire [1-1:0] node884;
	wire [1-1:0] node887;
	wire [1-1:0] node888;
	wire [1-1:0] node889;
	wire [1-1:0] node891;
	wire [1-1:0] node892;
	wire [1-1:0] node894;
	wire [1-1:0] node898;
	wire [1-1:0] node899;
	wire [1-1:0] node901;
	wire [1-1:0] node902;
	wire [1-1:0] node904;
	wire [1-1:0] node905;
	wire [1-1:0] node910;
	wire [1-1:0] node912;
	wire [1-1:0] node913;
	wire [1-1:0] node915;
	wire [1-1:0] node919;
	wire [1-1:0] node920;
	wire [1-1:0] node922;
	wire [1-1:0] node923;
	wire [1-1:0] node924;
	wire [1-1:0] node928;
	wire [1-1:0] node930;
	wire [1-1:0] node931;
	wire [1-1:0] node936;
	wire [1-1:0] node937;
	wire [1-1:0] node938;
	wire [1-1:0] node939;
	wire [1-1:0] node940;
	wire [1-1:0] node942;
	wire [1-1:0] node943;
	wire [1-1:0] node944;
	wire [1-1:0] node946;
	wire [1-1:0] node949;
	wire [1-1:0] node951;
	wire [1-1:0] node955;
	wire [1-1:0] node956;
	wire [1-1:0] node957;
	wire [1-1:0] node961;
	wire [1-1:0] node963;
	wire [1-1:0] node964;
	wire [1-1:0] node968;
	wire [1-1:0] node969;
	wire [1-1:0] node971;
	wire [1-1:0] node972;
	wire [1-1:0] node975;
	wire [1-1:0] node977;
	wire [1-1:0] node981;
	wire [1-1:0] node982;
	wire [1-1:0] node983;
	wire [1-1:0] node985;
	wire [1-1:0] node988;
	wire [1-1:0] node989;
	wire [1-1:0] node990;
	wire [1-1:0] node994;
	wire [1-1:0] node996;
	wire [1-1:0] node999;
	wire [1-1:0] node1000;
	wire [1-1:0] node1001;
	wire [1-1:0] node1003;
	wire [1-1:0] node1004;
	wire [1-1:0] node1010;
	wire [1-1:0] node1011;
	wire [1-1:0] node1012;
	wire [1-1:0] node1013;
	wire [1-1:0] node1015;
	wire [1-1:0] node1018;
	wire [1-1:0] node1020;
	wire [1-1:0] node1021;
	wire [1-1:0] node1024;
	wire [1-1:0] node1025;
	wire [1-1:0] node1029;
	wire [1-1:0] node1030;
	wire [1-1:0] node1032;
	wire [1-1:0] node1034;
	wire [1-1:0] node1038;
	wire [1-1:0] node1039;
	wire [1-1:0] node1040;
	wire [1-1:0] node1042;
	wire [1-1:0] node1044;
	wire [1-1:0] node1048;
	wire [1-1:0] node1049;
	wire [1-1:0] node1050;
	wire [1-1:0] node1051;
	wire [1-1:0] node1053;
	wire [1-1:0] node1054;
	wire [1-1:0] node1060;
	wire [1-1:0] node1062;
	wire [1-1:0] node1063;
	wire [1-1:0] node1067;
	wire [1-1:0] node1068;
	wire [1-1:0] node1069;
	wire [1-1:0] node1070;
	wire [1-1:0] node1072;
	wire [1-1:0] node1073;
	wire [1-1:0] node1074;
	wire [1-1:0] node1075;
	wire [1-1:0] node1079;
	wire [1-1:0] node1081;
	wire [1-1:0] node1085;
	wire [1-1:0] node1086;
	wire [1-1:0] node1087;
	wire [1-1:0] node1089;
	wire [1-1:0] node1092;
	wire [1-1:0] node1093;
	wire [1-1:0] node1094;
	wire [1-1:0] node1098;
	wire [1-1:0] node1100;
	wire [1-1:0] node1103;
	wire [1-1:0] node1105;
	wire [1-1:0] node1106;
	wire [1-1:0] node1107;
	wire [1-1:0] node1110;
	wire [1-1:0] node1111;
	wire [1-1:0] node1115;
	wire [1-1:0] node1117;
	wire [1-1:0] node1120;
	wire [1-1:0] node1122;
	wire [1-1:0] node1123;
	wire [1-1:0] node1124;
	wire [1-1:0] node1125;
	wire [1-1:0] node1129;
	wire [1-1:0] node1130;
	wire [1-1:0] node1131;
	wire [1-1:0] node1135;
	wire [1-1:0] node1136;
	wire [1-1:0] node1141;
	wire [1-1:0] node1142;
	wire [1-1:0] node1143;
	wire [1-1:0] node1144;
	wire [1-1:0] node1145;
	wire [1-1:0] node1146;
	wire [1-1:0] node1148;
	wire [1-1:0] node1149;
	wire [1-1:0] node1151;
	wire [1-1:0] node1155;
	wire [1-1:0] node1156;
	wire [1-1:0] node1157;
	wire [1-1:0] node1158;
	wire [1-1:0] node1163;
	wire [1-1:0] node1164;
	wire [1-1:0] node1166;
	wire [1-1:0] node1170;
	wire [1-1:0] node1171;
	wire [1-1:0] node1173;
	wire [1-1:0] node1175;
	wire [1-1:0] node1177;
	wire [1-1:0] node1180;
	wire [1-1:0] node1181;
	wire [1-1:0] node1183;
	wire [1-1:0] node1185;
	wire [1-1:0] node1186;
	wire [1-1:0] node1191;
	wire [1-1:0] node1192;
	wire [1-1:0] node1193;
	wire [1-1:0] node1194;
	wire [1-1:0] node1195;
	wire [1-1:0] node1201;
	wire [1-1:0] node1202;
	wire [1-1:0] node1203;
	wire [1-1:0] node1204;
	wire [1-1:0] node1206;
	wire [1-1:0] node1208;
	wire [1-1:0] node1212;
	wire [1-1:0] node1214;
	wire [1-1:0] node1215;
	wire [1-1:0] node1219;
	wire [1-1:0] node1220;
	wire [1-1:0] node1222;
	wire [1-1:0] node1224;
	wire [1-1:0] node1225;
	wire [1-1:0] node1230;
	wire [1-1:0] node1231;
	wire [1-1:0] node1232;
	wire [1-1:0] node1233;
	wire [1-1:0] node1235;
	wire [1-1:0] node1236;
	wire [1-1:0] node1238;
	wire [1-1:0] node1242;
	wire [1-1:0] node1243;
	wire [1-1:0] node1245;
	wire [1-1:0] node1246;
	wire [1-1:0] node1249;
	wire [1-1:0] node1253;
	wire [1-1:0] node1254;
	wire [1-1:0] node1256;
	wire [1-1:0] node1257;
	wire [1-1:0] node1258;
	wire [1-1:0] node1259;
	wire [1-1:0] node1264;
	wire [1-1:0] node1268;
	wire [1-1:0] node1269;
	wire [1-1:0] node1270;
	wire [1-1:0] node1271;
	wire [1-1:0] node1272;
	wire [1-1:0] node1276;
	wire [1-1:0] node1278;
	wire [1-1:0] node1281;
	wire [1-1:0] node1283;
	wire [1-1:0] node1284;
	wire [1-1:0] node1285;
	wire [1-1:0] node1290;
	wire [1-1:0] node1291;
	wire [1-1:0] node1292;
	wire [1-1:0] node1293;
	wire [1-1:0] node1297;
	wire [1-1:0] node1298;
	wire [1-1:0] node1299;
	wire [1-1:0] node1301;
	wire [1-1:0] node1305;
	wire [1-1:0] node1306;
	wire [1-1:0] node1310;
	wire [1-1:0] node1311;
	wire [1-1:0] node1313;
	wire [1-1:0] node1317;
	wire [1-1:0] node1318;
	wire [1-1:0] node1319;
	wire [1-1:0] node1320;
	wire [1-1:0] node1322;
	wire [1-1:0] node1323;
	wire [1-1:0] node1324;
	wire [1-1:0] node1326;
	wire [1-1:0] node1329;
	wire [1-1:0] node1330;
	wire [1-1:0] node1335;
	wire [1-1:0] node1336;
	wire [1-1:0] node1337;
	wire [1-1:0] node1338;
	wire [1-1:0] node1339;
	wire [1-1:0] node1345;
	wire [1-1:0] node1347;
	wire [1-1:0] node1348;
	wire [1-1:0] node1349;
	wire [1-1:0] node1354;
	wire [1-1:0] node1355;
	wire [1-1:0] node1356;
	wire [1-1:0] node1358;
	wire [1-1:0] node1359;
	wire [1-1:0] node1364;
	wire [1-1:0] node1365;
	wire [1-1:0] node1366;
	wire [1-1:0] node1368;
	wire [1-1:0] node1369;
	wire [1-1:0] node1372;
	wire [1-1:0] node1375;
	wire [1-1:0] node1378;
	wire [1-1:0] node1380;
	wire [1-1:0] node1383;
	wire [1-1:0] node1384;
	wire [1-1:0] node1386;
	wire [1-1:0] node1387;
	wire [1-1:0] node1389;
	wire [1-1:0] node1393;
	wire [1-1:0] node1394;
	wire [1-1:0] node1395;
	wire [1-1:0] node1396;
	wire [1-1:0] node1398;
	wire [1-1:0] node1400;
	wire [1-1:0] node1403;
	wire [1-1:0] node1406;
	wire [1-1:0] node1408;
	wire [1-1:0] node1409;
	wire [1-1:0] node1413;
	wire [1-1:0] node1415;
	wire [1-1:0] node1416;
	wire [1-1:0] node1420;
	wire [1-1:0] node1421;
	wire [1-1:0] node1422;
	wire [1-1:0] node1423;
	wire [1-1:0] node1425;
	wire [1-1:0] node1426;
	wire [1-1:0] node1427;
	wire [1-1:0] node1428;
	wire [1-1:0] node1432;
	wire [1-1:0] node1433;
	wire [1-1:0] node1434;
	wire [1-1:0] node1438;
	wire [1-1:0] node1440;
	wire [1-1:0] node1444;
	wire [1-1:0] node1445;
	wire [1-1:0] node1446;
	wire [1-1:0] node1447;
	wire [1-1:0] node1448;
	wire [1-1:0] node1452;
	wire [1-1:0] node1453;
	wire [1-1:0] node1457;
	wire [1-1:0] node1458;
	wire [1-1:0] node1462;
	wire [1-1:0] node1464;
	wire [1-1:0] node1465;
	wire [1-1:0] node1466;
	wire [1-1:0] node1467;
	wire [1-1:0] node1471;
	wire [1-1:0] node1472;
	wire [1-1:0] node1476;
	wire [1-1:0] node1477;
	wire [1-1:0] node1481;
	wire [1-1:0] node1483;
	wire [1-1:0] node1484;
	wire [1-1:0] node1485;
	wire [1-1:0] node1486;
	wire [1-1:0] node1490;
	wire [1-1:0] node1491;
	wire [1-1:0] node1493;
	wire [1-1:0] node1496;
	wire [1-1:0] node1498;
	wire [1-1:0] node1502;
	wire [1-1:0] node1503;
	wire [1-1:0] node1504;
	wire [1-1:0] node1505;
	wire [1-1:0] node1506;
	wire [1-1:0] node1507;
	wire [1-1:0] node1508;
	wire [1-1:0] node1512;
	wire [1-1:0] node1513;
	wire [1-1:0] node1515;
	wire [1-1:0] node1517;
	wire [1-1:0] node1521;
	wire [1-1:0] node1522;
	wire [1-1:0] node1523;
	wire [1-1:0] node1524;
	wire [1-1:0] node1526;
	wire [1-1:0] node1527;
	wire [1-1:0] node1528;
	wire [1-1:0] node1533;
	wire [1-1:0] node1534;
	wire [1-1:0] node1535;
	wire [1-1:0] node1539;
	wire [1-1:0] node1541;
	wire [1-1:0] node1542;
	wire [1-1:0] node1546;
	wire [1-1:0] node1547;
	wire [1-1:0] node1549;
	wire [1-1:0] node1552;
	wire [1-1:0] node1553;
	wire [1-1:0] node1556;
	wire [1-1:0] node1558;
	wire [1-1:0] node1561;
	wire [1-1:0] node1562;
	wire [1-1:0] node1563;
	wire [1-1:0] node1566;
	wire [1-1:0] node1567;
	wire [1-1:0] node1570;
	wire [1-1:0] node1572;
	wire [1-1:0] node1575;
	wire [1-1:0] node1576;
	wire [1-1:0] node1577;
	wire [1-1:0] node1582;
	wire [1-1:0] node1583;
	wire [1-1:0] node1584;
	wire [1-1:0] node1585;
	wire [1-1:0] node1586;
	wire [1-1:0] node1588;
	wire [1-1:0] node1592;
	wire [1-1:0] node1593;
	wire [1-1:0] node1595;
	wire [1-1:0] node1596;
	wire [1-1:0] node1600;
	wire [1-1:0] node1603;
	wire [1-1:0] node1605;
	wire [1-1:0] node1607;
	wire [1-1:0] node1608;
	wire [1-1:0] node1609;
	wire [1-1:0] node1614;
	wire [1-1:0] node1615;
	wire [1-1:0] node1616;
	wire [1-1:0] node1617;
	wire [1-1:0] node1618;
	wire [1-1:0] node1620;
	wire [1-1:0] node1625;
	wire [1-1:0] node1626;
	wire [1-1:0] node1627;
	wire [1-1:0] node1628;
	wire [1-1:0] node1631;
	wire [1-1:0] node1634;
	wire [1-1:0] node1636;
	wire [1-1:0] node1640;
	wire [1-1:0] node1641;
	wire [1-1:0] node1642;
	wire [1-1:0] node1643;
	wire [1-1:0] node1647;
	wire [1-1:0] node1649;
	wire [1-1:0] node1651;
	wire [1-1:0] node1655;
	wire [1-1:0] node1656;
	wire [1-1:0] node1657;
	wire [1-1:0] node1658;
	wire [1-1:0] node1659;
	wire [1-1:0] node1661;
	wire [1-1:0] node1662;
	wire [1-1:0] node1664;
	wire [1-1:0] node1665;
	wire [1-1:0] node1670;
	wire [1-1:0] node1671;
	wire [1-1:0] node1672;
	wire [1-1:0] node1676;
	wire [1-1:0] node1677;
	wire [1-1:0] node1678;
	wire [1-1:0] node1682;
	wire [1-1:0] node1685;
	wire [1-1:0] node1686;
	wire [1-1:0] node1687;
	wire [1-1:0] node1689;
	wire [1-1:0] node1690;
	wire [1-1:0] node1693;
	wire [1-1:0] node1694;
	wire [1-1:0] node1700;
	wire [1-1:0] node1701;
	wire [1-1:0] node1702;
	wire [1-1:0] node1703;
	wire [1-1:0] node1707;
	wire [1-1:0] node1709;
	wire [1-1:0] node1711;
	wire [1-1:0] node1714;
	wire [1-1:0] node1715;
	wire [1-1:0] node1716;
	wire [1-1:0] node1717;
	wire [1-1:0] node1720;
	wire [1-1:0] node1722;
	wire [1-1:0] node1725;
	wire [1-1:0] node1726;
	wire [1-1:0] node1727;
	wire [1-1:0] node1733;
	wire [1-1:0] node1734;
	wire [1-1:0] node1735;
	wire [1-1:0] node1736;
	wire [1-1:0] node1737;
	wire [1-1:0] node1738;
	wire [1-1:0] node1742;
	wire [1-1:0] node1745;
	wire [1-1:0] node1747;
	wire [1-1:0] node1750;
	wire [1-1:0] node1752;
	wire [1-1:0] node1754;
	wire [1-1:0] node1755;
	wire [1-1:0] node1757;
	wire [1-1:0] node1760;
	wire [1-1:0] node1763;
	wire [1-1:0] node1764;
	wire [1-1:0] node1765;
	wire [1-1:0] node1766;
	wire [1-1:0] node1771;
	wire [1-1:0] node1773;
	wire [1-1:0] node1775;
	wire [1-1:0] node1776;
	wire [1-1:0] node1780;
	wire [1-1:0] node1781;
	wire [1-1:0] node1782;
	wire [1-1:0] node1784;
	wire [1-1:0] node1785;
	wire [1-1:0] node1786;
	wire [1-1:0] node1788;
	wire [1-1:0] node1791;
	wire [1-1:0] node1792;
	wire [1-1:0] node1793;
	wire [1-1:0] node1797;
	wire [1-1:0] node1798;
	wire [1-1:0] node1803;
	wire [1-1:0] node1804;
	wire [1-1:0] node1805;
	wire [1-1:0] node1807;
	wire [1-1:0] node1810;
	wire [1-1:0] node1811;
	wire [1-1:0] node1812;
	wire [1-1:0] node1816;
	wire [1-1:0] node1817;
	wire [1-1:0] node1821;
	wire [1-1:0] node1823;
	wire [1-1:0] node1824;
	wire [1-1:0] node1826;
	wire [1-1:0] node1828;
	wire [1-1:0] node1830;
	wire [1-1:0] node1833;
	wire [1-1:0] node1834;
	wire [1-1:0] node1838;
	wire [1-1:0] node1840;
	wire [1-1:0] node1841;
	wire [1-1:0] node1842;
	wire [1-1:0] node1844;
	wire [1-1:0] node1847;
	wire [1-1:0] node1848;
	wire [1-1:0] node1850;
	wire [1-1:0] node1853;
	wire [1-1:0] node1854;
	wire [1-1:0] node1855;
	wire [1-1:0] node1857;
	wire [1-1:0] node1858;
	wire [1-1:0] node1861;
	wire [1-1:0] node1864;
	wire [1-1:0] node1866;
	wire [1-1:0] node1869;
	wire [1-1:0] node1870;

	assign outp = (inp[6]) ? node612 : node1;
		assign node1 = (inp[15]) ? node531 : node2;
			assign node2 = (inp[12]) ? node84 : node3;
				assign node3 = (inp[0]) ? node25 : node4;
					assign node4 = (inp[1]) ? node6 : 1'b1;
						assign node6 = (inp[8]) ? 1'b1 : node7;
							assign node7 = (inp[11]) ? node19 : node8;
								assign node8 = (inp[13]) ? node14 : node9;
									assign node9 = (inp[2]) ? 1'b0 : node10;
										assign node10 = (inp[14]) ? 1'b1 : 1'b0;
									assign node14 = (inp[2]) ? 1'b1 : node15;
										assign node15 = (inp[14]) ? 1'b0 : 1'b1;
								assign node19 = (inp[14]) ? node21 : 1'b0;
									assign node21 = (inp[2]) ? 1'b0 : 1'b1;
					assign node25 = (inp[4]) ? node63 : node26;
						assign node26 = (inp[1]) ? node44 : node27;
							assign node27 = (inp[11]) ? node39 : node28;
								assign node28 = (inp[13]) ? node34 : node29;
									assign node29 = (inp[14]) ? node31 : 1'b0;
										assign node31 = (inp[2]) ? 1'b0 : 1'b1;
									assign node34 = (inp[14]) ? node36 : 1'b1;
										assign node36 = (inp[2]) ? 1'b1 : 1'b0;
								assign node39 = (inp[14]) ? node41 : 1'b0;
									assign node41 = (inp[2]) ? 1'b0 : 1'b1;
							assign node44 = (inp[8]) ? node46 : 1'b1;
								assign node46 = (inp[2]) ? node58 : node47;
									assign node47 = (inp[14]) ? node53 : node48;
										assign node48 = (inp[13]) ? node50 : 1'b0;
											assign node50 = (inp[11]) ? 1'b0 : 1'b1;
										assign node53 = (inp[13]) ? node55 : 1'b1;
											assign node55 = (inp[11]) ? 1'b1 : 1'b0;
									assign node58 = (inp[11]) ? 1'b0 : node59;
										assign node59 = (inp[13]) ? 1'b1 : 1'b0;
						assign node63 = (inp[8]) ? 1'b1 : node64;
							assign node64 = (inp[1]) ? node66 : 1'b1;
								assign node66 = (inp[2]) ? node78 : node67;
									assign node67 = (inp[14]) ? node73 : node68;
										assign node68 = (inp[11]) ? 1'b0 : node69;
											assign node69 = (inp[13]) ? 1'b1 : 1'b0;
										assign node73 = (inp[11]) ? 1'b1 : node74;
											assign node74 = (inp[13]) ? 1'b0 : 1'b1;
									assign node78 = (inp[11]) ? 1'b0 : node79;
										assign node79 = (inp[13]) ? 1'b1 : 1'b0;
				assign node84 = (inp[10]) ? node326 : node85;
					assign node85 = (inp[9]) ? node207 : node86;
						assign node86 = (inp[7]) ? node156 : node87;
							assign node87 = (inp[3]) ? node125 : node88;
								assign node88 = (inp[13]) ? node110 : node89;
									assign node89 = (inp[4]) ? node105 : node90;
										assign node90 = (inp[8]) ? 1'b1 : node91;
											assign node91 = (inp[5]) ? node93 : 1'b0;
												assign node93 = (inp[2]) ? node99 : node94;
													assign node94 = (inp[1]) ? node96 : 1'b0;
														assign node96 = (inp[14]) ? 1'b0 : 1'b1;
													assign node99 = (inp[11]) ? 1'b0 : node100;
														assign node100 = (inp[1]) ? 1'b1 : 1'b0;
										assign node105 = (inp[1]) ? node107 : 1'b0;
											assign node107 = (inp[8]) ? 1'b0 : 1'b1;
									assign node110 = (inp[11]) ? node118 : node111;
										assign node111 = (inp[14]) ? node113 : 1'b0;
											assign node113 = (inp[2]) ? 1'b0 : node114;
												assign node114 = (inp[0]) ? 1'b1 : 1'b0;
										assign node118 = (inp[1]) ? 1'b1 : node119;
											assign node119 = (inp[0]) ? node121 : 1'b0;
												assign node121 = (inp[4]) ? 1'b0 : 1'b1;
								assign node125 = (inp[0]) ? node135 : node126;
									assign node126 = (inp[8]) ? 1'b1 : node127;
										assign node127 = (inp[1]) ? node129 : 1'b1;
											assign node129 = (inp[13]) ? 1'b0 : node130;
												assign node130 = (inp[4]) ? 1'b0 : 1'b1;
									assign node135 = (inp[4]) ? node149 : node136;
										assign node136 = (inp[1]) ? node144 : node137;
											assign node137 = (inp[14]) ? node141 : node138;
												assign node138 = (inp[2]) ? 1'b1 : 1'b0;
												assign node141 = (inp[2]) ? 1'b0 : 1'b1;
											assign node144 = (inp[5]) ? node146 : 1'b1;
												assign node146 = (inp[13]) ? 1'b1 : 1'b0;
										assign node149 = (inp[1]) ? node151 : 1'b1;
											assign node151 = (inp[8]) ? 1'b1 : node152;
												assign node152 = (inp[14]) ? 1'b1 : 1'b0;
							assign node156 = (inp[0]) ? node174 : node157;
								assign node157 = (inp[8]) ? 1'b0 : node158;
									assign node158 = (inp[1]) ? node160 : 1'b0;
										assign node160 = (inp[13]) ? node166 : node161;
											assign node161 = (inp[5]) ? node163 : 1'b1;
												assign node163 = (inp[14]) ? 1'b0 : 1'b1;
											assign node166 = (inp[3]) ? 1'b0 : node167;
												assign node167 = (inp[11]) ? node169 : 1'b0;
													assign node169 = (inp[2]) ? 1'b1 : 1'b0;
								assign node174 = (inp[4]) ? node198 : node175;
									assign node175 = (inp[13]) ? node183 : node176;
										assign node176 = (inp[5]) ? 1'b1 : node177;
											assign node177 = (inp[14]) ? 1'b0 : node178;
												assign node178 = (inp[8]) ? 1'b1 : 1'b0;
										assign node183 = (inp[1]) ? node189 : node184;
											assign node184 = (inp[2]) ? node186 : 1'b1;
												assign node186 = (inp[11]) ? 1'b1 : 1'b0;
											assign node189 = (inp[5]) ? node191 : 1'b1;
												assign node191 = (inp[14]) ? 1'b0 : node192;
													assign node192 = (inp[8]) ? node194 : 1'b0;
														assign node194 = (inp[11]) ? 1'b1 : 1'b0;
									assign node198 = (inp[8]) ? 1'b0 : node199;
										assign node199 = (inp[1]) ? node201 : 1'b0;
											assign node201 = (inp[2]) ? 1'b1 : node202;
												assign node202 = (inp[14]) ? 1'b0 : 1'b1;
						assign node207 = (inp[3]) ? node257 : node208;
							assign node208 = (inp[0]) ? node224 : node209;
								assign node209 = (inp[1]) ? node211 : 1'b1;
									assign node211 = (inp[8]) ? 1'b1 : node212;
										assign node212 = (inp[11]) ? node218 : node213;
											assign node213 = (inp[13]) ? 1'b1 : node214;
												assign node214 = (inp[4]) ? 1'b0 : 1'b1;
											assign node218 = (inp[2]) ? 1'b0 : node219;
												assign node219 = (inp[14]) ? 1'b1 : 1'b0;
								assign node224 = (inp[13]) ? node238 : node225;
									assign node225 = (inp[4]) ? node233 : node226;
										assign node226 = (inp[14]) ? node228 : 1'b0;
											assign node228 = (inp[2]) ? node230 : 1'b1;
												assign node230 = (inp[8]) ? 1'b0 : 1'b1;
										assign node233 = (inp[1]) ? node235 : 1'b1;
											assign node235 = (inp[8]) ? 1'b1 : 1'b0;
									assign node238 = (inp[5]) ? node248 : node239;
										assign node239 = (inp[4]) ? 1'b1 : node240;
											assign node240 = (inp[7]) ? node242 : 1'b0;
												assign node242 = (inp[14]) ? node244 : 1'b1;
													assign node244 = (inp[11]) ? 1'b1 : 1'b0;
										assign node248 = (inp[8]) ? 1'b1 : node249;
											assign node249 = (inp[4]) ? node251 : 1'b1;
												assign node251 = (inp[14]) ? node253 : 1'b1;
													assign node253 = (inp[2]) ? 1'b1 : 1'b0;
							assign node257 = (inp[7]) ? node297 : node258;
								assign node258 = (inp[8]) ? node288 : node259;
									assign node259 = (inp[14]) ? node281 : node260;
										assign node260 = (inp[11]) ? node272 : node261;
											assign node261 = (inp[13]) ? 1'b0 : node262;
												assign node262 = (inp[0]) ? node266 : node263;
													assign node263 = (inp[1]) ? 1'b1 : 1'b0;
													assign node266 = (inp[5]) ? 1'b0 : node267;
														assign node267 = (inp[4]) ? 1'b1 : 1'b0;
											assign node272 = (inp[5]) ? 1'b1 : node273;
												assign node273 = (inp[1]) ? node277 : node274;
													assign node274 = (inp[4]) ? 1'b0 : 1'b1;
													assign node277 = (inp[0]) ? 1'b0 : 1'b1;
										assign node281 = (inp[5]) ? node283 : 1'b0;
											assign node283 = (inp[0]) ? node285 : 1'b1;
												assign node285 = (inp[13]) ? 1'b0 : 1'b1;
									assign node288 = (inp[0]) ? node290 : 1'b0;
										assign node290 = (inp[1]) ? 1'b0 : node291;
											assign node291 = (inp[4]) ? 1'b0 : node292;
												assign node292 = (inp[2]) ? 1'b1 : 1'b0;
								assign node297 = (inp[0]) ? node305 : node298;
									assign node298 = (inp[1]) ? node300 : 1'b1;
										assign node300 = (inp[8]) ? 1'b1 : node301;
											assign node301 = (inp[11]) ? 1'b0 : 1'b1;
									assign node305 = (inp[4]) ? node321 : node306;
										assign node306 = (inp[1]) ? node314 : node307;
											assign node307 = (inp[8]) ? node309 : 1'b0;
												assign node309 = (inp[14]) ? node311 : 1'b0;
													assign node311 = (inp[2]) ? 1'b0 : 1'b1;
											assign node314 = (inp[11]) ? 1'b1 : node315;
												assign node315 = (inp[14]) ? node317 : 1'b1;
													assign node317 = (inp[5]) ? 1'b1 : 1'b0;
										assign node321 = (inp[8]) ? 1'b1 : node322;
											assign node322 = (inp[11]) ? 1'b0 : 1'b1;
					assign node326 = (inp[3]) ? node418 : node327;
						assign node327 = (inp[0]) ? node349 : node328;
							assign node328 = (inp[1]) ? node330 : 1'b0;
								assign node330 = (inp[8]) ? 1'b0 : node331;
									assign node331 = (inp[2]) ? node343 : node332;
										assign node332 = (inp[14]) ? node338 : node333;
											assign node333 = (inp[11]) ? 1'b1 : node334;
												assign node334 = (inp[9]) ? 1'b0 : 1'b1;
											assign node338 = (inp[11]) ? 1'b0 : node339;
												assign node339 = (inp[13]) ? 1'b1 : 1'b0;
										assign node343 = (inp[13]) ? node345 : 1'b1;
											assign node345 = (inp[11]) ? 1'b1 : 1'b0;
							assign node349 = (inp[4]) ? node397 : node350;
								assign node350 = (inp[1]) ? node374 : node351;
									assign node351 = (inp[2]) ? node369 : node352;
										assign node352 = (inp[7]) ? node362 : node353;
											assign node353 = (inp[9]) ? 1'b1 : node354;
												assign node354 = (inp[5]) ? node358 : node355;
													assign node355 = (inp[11]) ? 1'b1 : 1'b0;
													assign node358 = (inp[8]) ? 1'b1 : 1'b0;
											assign node362 = (inp[9]) ? 1'b0 : node363;
												assign node363 = (inp[11]) ? 1'b0 : node364;
													assign node364 = (inp[14]) ? 1'b1 : 1'b0;
										assign node369 = (inp[8]) ? 1'b1 : node370;
											assign node370 = (inp[13]) ? 1'b0 : 1'b1;
									assign node374 = (inp[8]) ? node376 : 1'b0;
										assign node376 = (inp[13]) ? node382 : node377;
											assign node377 = (inp[14]) ? node379 : 1'b1;
												assign node379 = (inp[5]) ? 1'b0 : 1'b1;
											assign node382 = (inp[7]) ? node388 : node383;
												assign node383 = (inp[14]) ? node385 : 1'b0;
													assign node385 = (inp[2]) ? 1'b1 : 1'b0;
												assign node388 = (inp[14]) ? node390 : 1'b1;
													assign node390 = (inp[2]) ? node394 : node391;
														assign node391 = (inp[11]) ? 1'b0 : 1'b1;
														assign node394 = (inp[11]) ? 1'b1 : 1'b0;
								assign node397 = (inp[8]) ? 1'b0 : node398;
									assign node398 = (inp[1]) ? node400 : 1'b0;
										assign node400 = (inp[7]) ? node408 : node401;
											assign node401 = (inp[2]) ? node403 : 1'b0;
												assign node403 = (inp[13]) ? node405 : 1'b1;
													assign node405 = (inp[11]) ? 1'b1 : 1'b0;
											assign node408 = (inp[9]) ? 1'b1 : node409;
												assign node409 = (inp[14]) ? 1'b0 : node410;
													assign node410 = (inp[13]) ? node412 : 1'b1;
														assign node412 = (inp[11]) ? 1'b1 : 1'b0;
						assign node418 = (inp[7]) ? node472 : node419;
							assign node419 = (inp[8]) ? node457 : node420;
								assign node420 = (inp[1]) ? node432 : node421;
									assign node421 = (inp[0]) ? node423 : 1'b1;
										assign node423 = (inp[13]) ? 1'b1 : node424;
											assign node424 = (inp[4]) ? 1'b1 : node425;
												assign node425 = (inp[2]) ? 1'b0 : node426;
													assign node426 = (inp[11]) ? 1'b1 : 1'b0;
									assign node432 = (inp[0]) ? node444 : node433;
										assign node433 = (inp[2]) ? 1'b0 : node434;
											assign node434 = (inp[11]) ? 1'b0 : node435;
												assign node435 = (inp[14]) ? node439 : node436;
													assign node436 = (inp[13]) ? 1'b1 : 1'b0;
													assign node439 = (inp[13]) ? 1'b0 : 1'b1;
										assign node444 = (inp[4]) ? node446 : 1'b1;
											assign node446 = (inp[11]) ? node454 : node447;
												assign node447 = (inp[9]) ? node449 : 1'b1;
													assign node449 = (inp[5]) ? node451 : 1'b1;
														assign node451 = (inp[14]) ? 1'b0 : 1'b1;
												assign node454 = (inp[5]) ? 1'b1 : 1'b0;
								assign node457 = (inp[0]) ? node459 : 1'b1;
									assign node459 = (inp[4]) ? 1'b1 : node460;
										assign node460 = (inp[2]) ? node468 : node461;
											assign node461 = (inp[1]) ? node463 : 1'b1;
												assign node463 = (inp[9]) ? node465 : 1'b1;
													assign node465 = (inp[11]) ? 1'b1 : 1'b0;
											assign node468 = (inp[5]) ? 1'b0 : 1'b1;
							assign node472 = (inp[1]) ? node494 : node473;
								assign node473 = (inp[0]) ? node475 : 1'b0;
									assign node475 = (inp[4]) ? 1'b0 : node476;
										assign node476 = (inp[8]) ? node488 : node477;
											assign node477 = (inp[5]) ? 1'b0 : node478;
												assign node478 = (inp[14]) ? node482 : node479;
													assign node479 = (inp[2]) ? 1'b0 : 1'b1;
													assign node482 = (inp[13]) ? 1'b1 : node483;
														assign node483 = (inp[2]) ? 1'b1 : 1'b0;
											assign node488 = (inp[9]) ? node490 : 1'b1;
												assign node490 = (inp[5]) ? 1'b1 : 1'b0;
								assign node494 = (inp[5]) ? node512 : node495;
									assign node495 = (inp[8]) ? node507 : node496;
										assign node496 = (inp[9]) ? node498 : 1'b1;
											assign node498 = (inp[14]) ? 1'b1 : node499;
												assign node499 = (inp[0]) ? 1'b0 : node500;
													assign node500 = (inp[4]) ? node502 : 1'b1;
														assign node502 = (inp[13]) ? 1'b0 : 1'b1;
										assign node507 = (inp[4]) ? 1'b0 : node508;
											assign node508 = (inp[0]) ? 1'b1 : 1'b0;
									assign node512 = (inp[9]) ? node526 : node513;
										assign node513 = (inp[4]) ? node523 : node514;
											assign node514 = (inp[11]) ? 1'b0 : node515;
												assign node515 = (inp[2]) ? 1'b0 : node516;
													assign node516 = (inp[0]) ? node518 : 1'b1;
														assign node518 = (inp[13]) ? 1'b0 : 1'b1;
											assign node523 = (inp[8]) ? 1'b0 : 1'b1;
										assign node526 = (inp[11]) ? node528 : 1'b0;
											assign node528 = (inp[8]) ? 1'b1 : 1'b0;
			assign node531 = (inp[1]) ? node553 : node532;
				assign node532 = (inp[0]) ? node534 : 1'b1;
					assign node534 = (inp[4]) ? 1'b1 : node535;
						assign node535 = (inp[2]) ? node547 : node536;
							assign node536 = (inp[14]) ? node542 : node537;
								assign node537 = (inp[11]) ? 1'b0 : node538;
									assign node538 = (inp[13]) ? 1'b1 : 1'b0;
								assign node542 = (inp[13]) ? node544 : 1'b1;
									assign node544 = (inp[11]) ? 1'b1 : 1'b0;
							assign node547 = (inp[13]) ? node549 : 1'b0;
								assign node549 = (inp[11]) ? 1'b0 : 1'b1;
				assign node553 = (inp[8]) ? node591 : node554;
					assign node554 = (inp[0]) ? node572 : node555;
						assign node555 = (inp[11]) ? node567 : node556;
							assign node556 = (inp[13]) ? node562 : node557;
								assign node557 = (inp[2]) ? 1'b0 : node558;
									assign node558 = (inp[14]) ? 1'b1 : 1'b0;
								assign node562 = (inp[14]) ? node564 : 1'b1;
									assign node564 = (inp[2]) ? 1'b1 : 1'b0;
							assign node567 = (inp[14]) ? node569 : 1'b0;
								assign node569 = (inp[2]) ? 1'b0 : 1'b1;
						assign node572 = (inp[4]) ? node574 : 1'b1;
							assign node574 = (inp[11]) ? node586 : node575;
								assign node575 = (inp[13]) ? node581 : node576;
									assign node576 = (inp[14]) ? node578 : 1'b0;
										assign node578 = (inp[2]) ? 1'b0 : 1'b1;
									assign node581 = (inp[14]) ? node583 : 1'b1;
										assign node583 = (inp[2]) ? 1'b1 : 1'b0;
								assign node586 = (inp[14]) ? node588 : 1'b0;
									assign node588 = (inp[2]) ? 1'b0 : 1'b1;
					assign node591 = (inp[4]) ? 1'b1 : node592;
						assign node592 = (inp[0]) ? node594 : 1'b1;
							assign node594 = (inp[11]) ? node606 : node595;
								assign node595 = (inp[13]) ? node601 : node596;
									assign node596 = (inp[2]) ? 1'b0 : node597;
										assign node597 = (inp[14]) ? 1'b1 : 1'b0;
									assign node601 = (inp[14]) ? node603 : 1'b1;
										assign node603 = (inp[2]) ? 1'b1 : 1'b0;
								assign node606 = (inp[14]) ? node608 : 1'b0;
									assign node608 = (inp[2]) ? 1'b0 : 1'b1;
		assign node612 = (inp[5]) ? node1420 : node613;
			assign node613 = (inp[12]) ? node1067 : node614;
				assign node614 = (inp[9]) ? node810 : node615;
					assign node615 = (inp[3]) ? node685 : node616;
						assign node616 = (inp[4]) ? node664 : node617;
							assign node617 = (inp[0]) ? node633 : node618;
								assign node618 = (inp[8]) ? 1'b0 : node619;
									assign node619 = (inp[1]) ? node621 : 1'b0;
										assign node621 = (inp[14]) ? node627 : node622;
											assign node622 = (inp[11]) ? 1'b1 : node623;
												assign node623 = (inp[13]) ? 1'b0 : 1'b1;
											assign node627 = (inp[2]) ? node629 : 1'b0;
												assign node629 = (inp[13]) ? 1'b0 : 1'b1;
								assign node633 = (inp[8]) ? node641 : node634;
									assign node634 = (inp[1]) ? 1'b0 : node635;
										assign node635 = (inp[13]) ? node637 : 1'b1;
											assign node637 = (inp[11]) ? 1'b1 : 1'b0;
									assign node641 = (inp[2]) ? node659 : node642;
										assign node642 = (inp[1]) ? node654 : node643;
											assign node643 = (inp[10]) ? 1'b0 : node644;
												assign node644 = (inp[14]) ? node648 : node645;
													assign node645 = (inp[13]) ? 1'b0 : 1'b1;
													assign node648 = (inp[11]) ? 1'b0 : node649;
														assign node649 = (inp[13]) ? 1'b1 : 1'b0;
											assign node654 = (inp[15]) ? 1'b1 : node655;
												assign node655 = (inp[11]) ? 1'b1 : 1'b0;
										assign node659 = (inp[13]) ? node661 : 1'b1;
											assign node661 = (inp[11]) ? 1'b1 : 1'b0;
							assign node664 = (inp[8]) ? 1'b0 : node665;
								assign node665 = (inp[1]) ? node667 : 1'b0;
									assign node667 = (inp[13]) ? node673 : node668;
										assign node668 = (inp[14]) ? node670 : 1'b1;
											assign node670 = (inp[2]) ? 1'b1 : 1'b0;
										assign node673 = (inp[11]) ? node679 : node674;
											assign node674 = (inp[0]) ? 1'b0 : node675;
												assign node675 = (inp[14]) ? 1'b1 : 1'b0;
											assign node679 = (inp[15]) ? 1'b1 : node680;
												assign node680 = (inp[14]) ? 1'b0 : 1'b1;
						assign node685 = (inp[7]) ? node757 : node686;
							assign node686 = (inp[8]) ? node744 : node687;
								assign node687 = (inp[13]) ? node709 : node688;
									assign node688 = (inp[15]) ? node694 : node689;
										assign node689 = (inp[14]) ? node691 : 1'b0;
											assign node691 = (inp[4]) ? 1'b0 : 1'b1;
										assign node694 = (inp[2]) ? node704 : node695;
											assign node695 = (inp[14]) ? 1'b1 : node696;
												assign node696 = (inp[10]) ? 1'b0 : node697;
													assign node697 = (inp[1]) ? 1'b1 : node698;
														assign node698 = (inp[4]) ? 1'b1 : 1'b0;
											assign node704 = (inp[1]) ? 1'b0 : node705;
												assign node705 = (inp[11]) ? 1'b1 : 1'b0;
									assign node709 = (inp[14]) ? node721 : node710;
										assign node710 = (inp[11]) ? node712 : 1'b1;
											assign node712 = (inp[2]) ? node718 : node713;
												assign node713 = (inp[1]) ? node715 : 1'b1;
													assign node715 = (inp[4]) ? 1'b0 : 1'b1;
												assign node718 = (inp[1]) ? 1'b1 : 1'b0;
										assign node721 = (inp[1]) ? node729 : node722;
											assign node722 = (inp[2]) ? node724 : 1'b1;
												assign node724 = (inp[4]) ? 1'b1 : node725;
													assign node725 = (inp[0]) ? 1'b0 : 1'b1;
											assign node729 = (inp[0]) ? node737 : node730;
												assign node730 = (inp[4]) ? node732 : 1'b0;
													assign node732 = (inp[10]) ? 1'b0 : node733;
														assign node733 = (inp[2]) ? 1'b1 : 1'b0;
												assign node737 = (inp[10]) ? node739 : 1'b1;
													assign node739 = (inp[4]) ? node741 : 1'b1;
														assign node741 = (inp[15]) ? 1'b0 : 1'b0;
								assign node744 = (inp[4]) ? 1'b1 : node745;
									assign node745 = (inp[0]) ? node747 : 1'b1;
										assign node747 = (inp[10]) ? node751 : node748;
											assign node748 = (inp[13]) ? 1'b1 : 1'b0;
											assign node751 = (inp[2]) ? node753 : 1'b1;
												assign node753 = (inp[1]) ? 1'b1 : 1'b0;
							assign node757 = (inp[0]) ? node773 : node758;
								assign node758 = (inp[1]) ? node760 : 1'b0;
									assign node760 = (inp[8]) ? 1'b0 : node761;
										assign node761 = (inp[11]) ? 1'b1 : node762;
											assign node762 = (inp[15]) ? node764 : 1'b0;
												assign node764 = (inp[13]) ? node766 : 1'b1;
													assign node766 = (inp[2]) ? 1'b0 : node767;
														assign node767 = (inp[14]) ? 1'b1 : 1'b0;
								assign node773 = (inp[4]) ? node795 : node774;
									assign node774 = (inp[8]) ? node784 : node775;
										assign node775 = (inp[1]) ? 1'b0 : node776;
											assign node776 = (inp[2]) ? 1'b1 : node777;
												assign node777 = (inp[14]) ? 1'b0 : node778;
													assign node778 = (inp[13]) ? 1'b0 : 1'b1;
										assign node784 = (inp[13]) ? node790 : node785;
											assign node785 = (inp[14]) ? node787 : 1'b1;
												assign node787 = (inp[2]) ? 1'b1 : 1'b0;
											assign node790 = (inp[11]) ? 1'b1 : node791;
												assign node791 = (inp[14]) ? 1'b1 : 1'b0;
									assign node795 = (inp[1]) ? node797 : 1'b0;
										assign node797 = (inp[8]) ? 1'b0 : node798;
											assign node798 = (inp[11]) ? 1'b0 : node799;
												assign node799 = (inp[14]) ? node801 : 1'b1;
													assign node801 = (inp[15]) ? node805 : node802;
														assign node802 = (inp[10]) ? 1'b0 : 1'b1;
														assign node805 = (inp[13]) ? 1'b0 : 1'b1;
					assign node810 = (inp[10]) ? node936 : node811;
						assign node811 = (inp[7]) ? node887 : node812;
							assign node812 = (inp[3]) ? node846 : node813;
								assign node813 = (inp[4]) ? node837 : node814;
									assign node814 = (inp[0]) ? node820 : node815;
										assign node815 = (inp[1]) ? node817 : 1'b1;
											assign node817 = (inp[8]) ? 1'b1 : 1'b0;
										assign node820 = (inp[8]) ? node830 : node821;
											assign node821 = (inp[1]) ? 1'b1 : node822;
												assign node822 = (inp[11]) ? 1'b0 : node823;
													assign node823 = (inp[14]) ? node825 : 1'b1;
														assign node825 = (inp[2]) ? 1'b1 : 1'b0;
											assign node830 = (inp[11]) ? 1'b0 : node831;
												assign node831 = (inp[15]) ? node833 : 1'b0;
													assign node833 = (inp[13]) ? 1'b1 : 1'b0;
									assign node837 = (inp[8]) ? 1'b1 : node838;
										assign node838 = (inp[11]) ? node840 : 1'b1;
											assign node840 = (inp[1]) ? node842 : 1'b1;
												assign node842 = (inp[2]) ? 1'b0 : 1'b1;
								assign node846 = (inp[14]) ? node874 : node847;
									assign node847 = (inp[4]) ? node865 : node848;
										assign node848 = (inp[11]) ? node856 : node849;
											assign node849 = (inp[13]) ? 1'b0 : node850;
												assign node850 = (inp[15]) ? node852 : 1'b1;
													assign node852 = (inp[0]) ? 1'b0 : 1'b1;
											assign node856 = (inp[0]) ? node860 : node857;
												assign node857 = (inp[1]) ? 1'b1 : 1'b0;
												assign node860 = (inp[2]) ? node862 : 1'b1;
													assign node862 = (inp[1]) ? 1'b0 : 1'b1;
										assign node865 = (inp[8]) ? 1'b0 : node866;
											assign node866 = (inp[1]) ? node868 : 1'b0;
												assign node868 = (inp[0]) ? node870 : 1'b1;
													assign node870 = (inp[15]) ? 1'b1 : 1'b0;
									assign node874 = (inp[2]) ? node882 : node875;
										assign node875 = (inp[4]) ? node877 : 1'b0;
											assign node877 = (inp[11]) ? 1'b0 : node878;
												assign node878 = (inp[13]) ? 1'b1 : 1'b0;
										assign node882 = (inp[15]) ? node884 : 1'b0;
											assign node884 = (inp[4]) ? 1'b0 : 1'b1;
							assign node887 = (inp[8]) ? node919 : node888;
								assign node888 = (inp[1]) ? node898 : node889;
									assign node889 = (inp[0]) ? node891 : 1'b1;
										assign node891 = (inp[4]) ? 1'b1 : node892;
											assign node892 = (inp[13]) ? node894 : 1'b0;
												assign node894 = (inp[11]) ? 1'b0 : 1'b1;
									assign node898 = (inp[0]) ? node910 : node899;
										assign node899 = (inp[15]) ? node901 : 1'b0;
											assign node901 = (inp[4]) ? 1'b0 : node902;
												assign node902 = (inp[13]) ? node904 : 1'b0;
													assign node904 = (inp[14]) ? 1'b0 : node905;
														assign node905 = (inp[3]) ? 1'b0 : 1'b1;
										assign node910 = (inp[4]) ? node912 : 1'b1;
											assign node912 = (inp[2]) ? 1'b0 : node913;
												assign node913 = (inp[13]) ? node915 : 1'b1;
													assign node915 = (inp[3]) ? 1'b0 : 1'b1;
								assign node919 = (inp[4]) ? 1'b1 : node920;
									assign node920 = (inp[0]) ? node922 : 1'b1;
										assign node922 = (inp[14]) ? node928 : node923;
											assign node923 = (inp[11]) ? 1'b0 : node924;
												assign node924 = (inp[13]) ? 1'b1 : 1'b0;
											assign node928 = (inp[2]) ? node930 : 1'b1;
												assign node930 = (inp[11]) ? 1'b0 : node931;
													assign node931 = (inp[13]) ? 1'b1 : 1'b0;
						assign node936 = (inp[7]) ? node1010 : node937;
							assign node937 = (inp[3]) ? node981 : node938;
								assign node938 = (inp[4]) ? node968 : node939;
									assign node939 = (inp[0]) ? node955 : node940;
										assign node940 = (inp[1]) ? node942 : 1'b0;
											assign node942 = (inp[8]) ? 1'b0 : node943;
												assign node943 = (inp[13]) ? node949 : node944;
													assign node944 = (inp[15]) ? node946 : 1'b1;
														assign node946 = (inp[14]) ? 1'b0 : 1'b1;
													assign node949 = (inp[11]) ? node951 : 1'b0;
														assign node951 = (inp[14]) ? 1'b0 : 1'b1;
										assign node955 = (inp[1]) ? node961 : node956;
											assign node956 = (inp[11]) ? 1'b1 : node957;
												assign node957 = (inp[8]) ? 1'b0 : 1'b1;
											assign node961 = (inp[8]) ? node963 : 1'b0;
												assign node963 = (inp[11]) ? 1'b1 : node964;
													assign node964 = (inp[2]) ? 1'b0 : 1'b1;
									assign node968 = (inp[8]) ? 1'b0 : node969;
										assign node969 = (inp[1]) ? node971 : 1'b0;
											assign node971 = (inp[13]) ? node975 : node972;
												assign node972 = (inp[11]) ? 1'b0 : 1'b1;
												assign node975 = (inp[11]) ? node977 : 1'b0;
													assign node977 = (inp[0]) ? 1'b1 : 1'b0;
								assign node981 = (inp[8]) ? node999 : node982;
									assign node982 = (inp[1]) ? node988 : node983;
										assign node983 = (inp[0]) ? node985 : 1'b1;
											assign node985 = (inp[4]) ? 1'b1 : 1'b0;
										assign node988 = (inp[11]) ? node994 : node989;
											assign node989 = (inp[0]) ? 1'b1 : node990;
												assign node990 = (inp[4]) ? 1'b0 : 1'b1;
											assign node994 = (inp[14]) ? node996 : 1'b0;
												assign node996 = (inp[4]) ? 1'b0 : 1'b1;
									assign node999 = (inp[2]) ? 1'b1 : node1000;
										assign node1000 = (inp[4]) ? 1'b1 : node1001;
											assign node1001 = (inp[14]) ? node1003 : 1'b0;
												assign node1003 = (inp[11]) ? 1'b1 : node1004;
													assign node1004 = (inp[13]) ? 1'b0 : 1'b1;
							assign node1010 = (inp[2]) ? node1038 : node1011;
								assign node1011 = (inp[4]) ? node1029 : node1012;
									assign node1012 = (inp[8]) ? node1018 : node1013;
										assign node1013 = (inp[13]) ? node1015 : 1'b0;
											assign node1015 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1018 = (inp[0]) ? node1020 : 1'b0;
											assign node1020 = (inp[3]) ? node1024 : node1021;
												assign node1021 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1024 = (inp[14]) ? 1'b1 : node1025;
													assign node1025 = (inp[15]) ? 1'b0 : 1'b1;
									assign node1029 = (inp[14]) ? 1'b0 : node1030;
										assign node1030 = (inp[11]) ? node1032 : 1'b0;
											assign node1032 = (inp[1]) ? node1034 : 1'b0;
												assign node1034 = (inp[8]) ? 1'b0 : 1'b1;
								assign node1038 = (inp[0]) ? node1048 : node1039;
									assign node1039 = (inp[8]) ? 1'b0 : node1040;
										assign node1040 = (inp[1]) ? node1042 : 1'b0;
											assign node1042 = (inp[13]) ? node1044 : 1'b1;
												assign node1044 = (inp[11]) ? 1'b1 : 1'b0;
									assign node1048 = (inp[11]) ? node1060 : node1049;
										assign node1049 = (inp[13]) ? 1'b0 : node1050;
											assign node1050 = (inp[15]) ? 1'b1 : node1051;
												assign node1051 = (inp[3]) ? node1053 : 1'b1;
													assign node1053 = (inp[4]) ? 1'b0 : node1054;
														assign node1054 = (inp[8]) ? 1'b1 : 1'b0;
										assign node1060 = (inp[4]) ? node1062 : 1'b1;
											assign node1062 = (inp[8]) ? 1'b0 : node1063;
												assign node1063 = (inp[1]) ? 1'b1 : 1'b0;
				assign node1067 = (inp[15]) ? node1141 : node1068;
					assign node1068 = (inp[4]) ? node1120 : node1069;
						assign node1069 = (inp[0]) ? node1085 : node1070;
							assign node1070 = (inp[1]) ? node1072 : 1'b1;
								assign node1072 = (inp[8]) ? 1'b1 : node1073;
									assign node1073 = (inp[11]) ? node1079 : node1074;
										assign node1074 = (inp[3]) ? 1'b1 : node1075;
											assign node1075 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1079 = (inp[14]) ? node1081 : 1'b0;
											assign node1081 = (inp[2]) ? 1'b0 : 1'b1;
							assign node1085 = (inp[1]) ? node1103 : node1086;
								assign node1086 = (inp[14]) ? node1092 : node1087;
									assign node1087 = (inp[13]) ? node1089 : 1'b0;
										assign node1089 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1092 = (inp[2]) ? node1098 : node1093;
										assign node1093 = (inp[11]) ? 1'b1 : node1094;
											assign node1094 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1098 = (inp[8]) ? node1100 : 1'b0;
											assign node1100 = (inp[13]) ? 1'b1 : 1'b0;
								assign node1103 = (inp[8]) ? node1105 : 1'b1;
									assign node1105 = (inp[11]) ? node1115 : node1106;
										assign node1106 = (inp[13]) ? node1110 : node1107;
											assign node1107 = (inp[2]) ? 1'b0 : 1'b1;
											assign node1110 = (inp[10]) ? 1'b1 : node1111;
												assign node1111 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1115 = (inp[14]) ? node1117 : 1'b0;
											assign node1117 = (inp[3]) ? 1'b1 : 1'b0;
						assign node1120 = (inp[1]) ? node1122 : 1'b1;
							assign node1122 = (inp[8]) ? 1'b1 : node1123;
								assign node1123 = (inp[14]) ? node1129 : node1124;
									assign node1124 = (inp[11]) ? 1'b0 : node1125;
										assign node1125 = (inp[13]) ? 1'b1 : 1'b0;
									assign node1129 = (inp[2]) ? node1135 : node1130;
										assign node1130 = (inp[11]) ? 1'b1 : node1131;
											assign node1131 = (inp[9]) ? 1'b1 : 1'b0;
										assign node1135 = (inp[11]) ? 1'b0 : node1136;
											assign node1136 = (inp[13]) ? 1'b1 : 1'b0;
					assign node1141 = (inp[7]) ? node1317 : node1142;
						assign node1142 = (inp[3]) ? node1230 : node1143;
							assign node1143 = (inp[10]) ? node1191 : node1144;
								assign node1144 = (inp[9]) ? node1170 : node1145;
									assign node1145 = (inp[2]) ? node1155 : node1146;
										assign node1146 = (inp[4]) ? node1148 : 1'b0;
											assign node1148 = (inp[8]) ? 1'b0 : node1149;
												assign node1149 = (inp[1]) ? node1151 : 1'b0;
													assign node1151 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1155 = (inp[13]) ? node1163 : node1156;
											assign node1156 = (inp[1]) ? 1'b1 : node1157;
												assign node1157 = (inp[11]) ? 1'b0 : node1158;
													assign node1158 = (inp[8]) ? 1'b1 : 1'b0;
											assign node1163 = (inp[4]) ? 1'b0 : node1164;
												assign node1164 = (inp[11]) ? node1166 : 1'b0;
													assign node1166 = (inp[0]) ? 1'b1 : 1'b0;
									assign node1170 = (inp[8]) ? node1180 : node1171;
										assign node1171 = (inp[1]) ? node1173 : 1'b1;
											assign node1173 = (inp[14]) ? node1175 : 1'b0;
												assign node1175 = (inp[11]) ? node1177 : 1'b1;
													assign node1177 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1180 = (inp[4]) ? 1'b1 : node1181;
											assign node1181 = (inp[0]) ? node1183 : 1'b1;
												assign node1183 = (inp[13]) ? node1185 : 1'b1;
													assign node1185 = (inp[14]) ? 1'b0 : node1186;
														assign node1186 = (inp[11]) ? 1'b0 : 1'b1;
								assign node1191 = (inp[1]) ? node1201 : node1192;
									assign node1192 = (inp[4]) ? 1'b0 : node1193;
										assign node1193 = (inp[13]) ? 1'b0 : node1194;
											assign node1194 = (inp[9]) ? 1'b0 : node1195;
												assign node1195 = (inp[0]) ? 1'b1 : 1'b0;
									assign node1201 = (inp[8]) ? node1219 : node1202;
										assign node1202 = (inp[4]) ? node1212 : node1203;
											assign node1203 = (inp[0]) ? 1'b0 : node1204;
												assign node1204 = (inp[9]) ? node1206 : 1'b0;
													assign node1206 = (inp[2]) ? node1208 : 1'b1;
														assign node1208 = (inp[13]) ? 1'b0 : 1'b1;
											assign node1212 = (inp[13]) ? node1214 : 1'b1;
												assign node1214 = (inp[11]) ? 1'b1 : node1215;
													assign node1215 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1219 = (inp[4]) ? 1'b0 : node1220;
											assign node1220 = (inp[0]) ? node1222 : 1'b0;
												assign node1222 = (inp[13]) ? node1224 : 1'b1;
													assign node1224 = (inp[14]) ? 1'b1 : node1225;
														assign node1225 = (inp[11]) ? 1'b1 : 1'b0;
							assign node1230 = (inp[9]) ? node1268 : node1231;
								assign node1231 = (inp[8]) ? node1253 : node1232;
									assign node1232 = (inp[1]) ? node1242 : node1233;
										assign node1233 = (inp[0]) ? node1235 : 1'b1;
											assign node1235 = (inp[4]) ? 1'b1 : node1236;
												assign node1236 = (inp[14]) ? node1238 : 1'b0;
													assign node1238 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1242 = (inp[0]) ? 1'b1 : node1243;
											assign node1243 = (inp[14]) ? node1245 : 1'b0;
												assign node1245 = (inp[2]) ? node1249 : node1246;
													assign node1246 = (inp[11]) ? 1'b1 : 1'b0;
													assign node1249 = (inp[13]) ? 1'b1 : 1'b0;
									assign node1253 = (inp[4]) ? 1'b1 : node1254;
										assign node1254 = (inp[0]) ? node1256 : 1'b1;
											assign node1256 = (inp[11]) ? node1264 : node1257;
												assign node1257 = (inp[2]) ? 1'b1 : node1258;
													assign node1258 = (inp[1]) ? 1'b1 : node1259;
														assign node1259 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1264 = (inp[2]) ? 1'b0 : 1'b1;
								assign node1268 = (inp[10]) ? node1290 : node1269;
									assign node1269 = (inp[8]) ? node1281 : node1270;
										assign node1270 = (inp[1]) ? node1276 : node1271;
											assign node1271 = (inp[13]) ? 1'b0 : node1272;
												assign node1272 = (inp[2]) ? 1'b0 : 1'b1;
											assign node1276 = (inp[0]) ? node1278 : 1'b1;
												assign node1278 = (inp[4]) ? 1'b1 : 1'b0;
										assign node1281 = (inp[0]) ? node1283 : 1'b0;
											assign node1283 = (inp[4]) ? 1'b0 : node1284;
												assign node1284 = (inp[11]) ? 1'b1 : node1285;
													assign node1285 = (inp[14]) ? 1'b1 : 1'b0;
									assign node1290 = (inp[8]) ? node1310 : node1291;
										assign node1291 = (inp[1]) ? node1297 : node1292;
											assign node1292 = (inp[13]) ? 1'b1 : node1293;
												assign node1293 = (inp[14]) ? 1'b1 : 1'b0;
											assign node1297 = (inp[4]) ? node1305 : node1298;
												assign node1298 = (inp[0]) ? 1'b1 : node1299;
													assign node1299 = (inp[11]) ? node1301 : 1'b0;
														assign node1301 = (inp[14]) ? 1'b1 : 1'b0;
												assign node1305 = (inp[11]) ? 1'b0 : node1306;
													assign node1306 = (inp[13]) ? 1'b1 : 1'b0;
										assign node1310 = (inp[4]) ? 1'b1 : node1311;
											assign node1311 = (inp[13]) ? node1313 : 1'b1;
												assign node1313 = (inp[11]) ? 1'b0 : 1'b1;
						assign node1317 = (inp[10]) ? node1383 : node1318;
							assign node1318 = (inp[9]) ? node1354 : node1319;
								assign node1319 = (inp[1]) ? node1335 : node1320;
									assign node1320 = (inp[0]) ? node1322 : 1'b0;
										assign node1322 = (inp[4]) ? 1'b0 : node1323;
											assign node1323 = (inp[13]) ? node1329 : node1324;
												assign node1324 = (inp[11]) ? node1326 : 1'b1;
													assign node1326 = (inp[2]) ? 1'b1 : 1'b0;
												assign node1329 = (inp[2]) ? 1'b0 : node1330;
													assign node1330 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1335 = (inp[8]) ? node1345 : node1336;
										assign node1336 = (inp[13]) ? 1'b1 : node1337;
											assign node1337 = (inp[2]) ? 1'b1 : node1338;
												assign node1338 = (inp[14]) ? 1'b0 : node1339;
													assign node1339 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1345 = (inp[0]) ? node1347 : 1'b0;
											assign node1347 = (inp[4]) ? 1'b0 : node1348;
												assign node1348 = (inp[11]) ? 1'b1 : node1349;
													assign node1349 = (inp[3]) ? 1'b1 : 1'b0;
								assign node1354 = (inp[1]) ? node1364 : node1355;
									assign node1355 = (inp[4]) ? 1'b1 : node1356;
										assign node1356 = (inp[0]) ? node1358 : 1'b1;
											assign node1358 = (inp[11]) ? 1'b0 : node1359;
												assign node1359 = (inp[13]) ? 1'b1 : 1'b0;
									assign node1364 = (inp[8]) ? node1378 : node1365;
										assign node1365 = (inp[2]) ? node1375 : node1366;
											assign node1366 = (inp[13]) ? node1368 : 1'b1;
												assign node1368 = (inp[0]) ? node1372 : node1369;
													assign node1369 = (inp[3]) ? 1'b1 : 1'b0;
													assign node1372 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1375 = (inp[0]) ? 1'b1 : 1'b0;
										assign node1378 = (inp[0]) ? node1380 : 1'b1;
											assign node1380 = (inp[4]) ? 1'b1 : 1'b0;
							assign node1383 = (inp[1]) ? node1393 : node1384;
								assign node1384 = (inp[0]) ? node1386 : 1'b0;
									assign node1386 = (inp[4]) ? 1'b0 : node1387;
										assign node1387 = (inp[13]) ? node1389 : 1'b1;
											assign node1389 = (inp[11]) ? 1'b1 : 1'b0;
								assign node1393 = (inp[8]) ? node1413 : node1394;
									assign node1394 = (inp[0]) ? node1406 : node1395;
										assign node1395 = (inp[9]) ? node1403 : node1396;
											assign node1396 = (inp[4]) ? node1398 : 1'b1;
												assign node1398 = (inp[3]) ? node1400 : 1'b1;
													assign node1400 = (inp[2]) ? 1'b1 : 1'b0;
											assign node1403 = (inp[3]) ? 1'b1 : 1'b0;
										assign node1406 = (inp[4]) ? node1408 : 1'b0;
											assign node1408 = (inp[11]) ? 1'b1 : node1409;
												assign node1409 = (inp[3]) ? 1'b1 : 1'b0;
									assign node1413 = (inp[0]) ? node1415 : 1'b0;
										assign node1415 = (inp[4]) ? 1'b0 : node1416;
											assign node1416 = (inp[13]) ? 1'b0 : 1'b1;
			assign node1420 = (inp[12]) ? node1502 : node1421;
				assign node1421 = (inp[4]) ? node1481 : node1422;
					assign node1422 = (inp[0]) ? node1444 : node1423;
						assign node1423 = (inp[1]) ? node1425 : 1'b1;
							assign node1425 = (inp[8]) ? 1'b1 : node1426;
								assign node1426 = (inp[14]) ? node1432 : node1427;
									assign node1427 = (inp[11]) ? 1'b0 : node1428;
										assign node1428 = (inp[13]) ? 1'b1 : 1'b0;
									assign node1432 = (inp[2]) ? node1438 : node1433;
										assign node1433 = (inp[11]) ? 1'b1 : node1434;
											assign node1434 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1438 = (inp[13]) ? node1440 : 1'b0;
											assign node1440 = (inp[11]) ? 1'b0 : 1'b1;
						assign node1444 = (inp[1]) ? node1462 : node1445;
							assign node1445 = (inp[11]) ? node1457 : node1446;
								assign node1446 = (inp[13]) ? node1452 : node1447;
									assign node1447 = (inp[2]) ? 1'b0 : node1448;
										assign node1448 = (inp[14]) ? 1'b1 : 1'b0;
									assign node1452 = (inp[2]) ? 1'b1 : node1453;
										assign node1453 = (inp[14]) ? 1'b0 : 1'b1;
								assign node1457 = (inp[2]) ? 1'b0 : node1458;
									assign node1458 = (inp[14]) ? 1'b1 : 1'b0;
							assign node1462 = (inp[8]) ? node1464 : 1'b1;
								assign node1464 = (inp[2]) ? node1476 : node1465;
									assign node1465 = (inp[14]) ? node1471 : node1466;
										assign node1466 = (inp[11]) ? 1'b0 : node1467;
											assign node1467 = (inp[13]) ? 1'b1 : 1'b0;
										assign node1471 = (inp[11]) ? 1'b1 : node1472;
											assign node1472 = (inp[13]) ? 1'b0 : 1'b1;
									assign node1476 = (inp[11]) ? 1'b0 : node1477;
										assign node1477 = (inp[13]) ? 1'b1 : 1'b0;
					assign node1481 = (inp[1]) ? node1483 : 1'b1;
						assign node1483 = (inp[8]) ? 1'b1 : node1484;
							assign node1484 = (inp[13]) ? node1490 : node1485;
								assign node1485 = (inp[2]) ? 1'b0 : node1486;
									assign node1486 = (inp[14]) ? 1'b1 : 1'b0;
								assign node1490 = (inp[11]) ? node1496 : node1491;
									assign node1491 = (inp[14]) ? node1493 : 1'b1;
										assign node1493 = (inp[2]) ? 1'b1 : 1'b0;
									assign node1496 = (inp[14]) ? node1498 : 1'b0;
										assign node1498 = (inp[2]) ? 1'b0 : 1'b1;
				assign node1502 = (inp[15]) ? node1780 : node1503;
					assign node1503 = (inp[7]) ? node1655 : node1504;
						assign node1504 = (inp[3]) ? node1582 : node1505;
							assign node1505 = (inp[1]) ? node1521 : node1506;
								assign node1506 = (inp[9]) ? node1512 : node1507;
									assign node1507 = (inp[4]) ? 1'b0 : node1508;
										assign node1508 = (inp[14]) ? 1'b0 : 1'b1;
									assign node1512 = (inp[10]) ? 1'b0 : node1513;
										assign node1513 = (inp[0]) ? node1515 : 1'b1;
											assign node1515 = (inp[11]) ? node1517 : 1'b1;
												assign node1517 = (inp[4]) ? 1'b1 : 1'b0;
								assign node1521 = (inp[14]) ? node1561 : node1522;
									assign node1522 = (inp[13]) ? node1546 : node1523;
										assign node1523 = (inp[8]) ? node1533 : node1524;
											assign node1524 = (inp[9]) ? node1526 : 1'b1;
												assign node1526 = (inp[2]) ? 1'b1 : node1527;
													assign node1527 = (inp[11]) ? 1'b0 : node1528;
														assign node1528 = (inp[0]) ? 1'b0 : 1'b1;
											assign node1533 = (inp[0]) ? node1539 : node1534;
												assign node1534 = (inp[10]) ? 1'b0 : node1535;
													assign node1535 = (inp[9]) ? 1'b1 : 1'b0;
												assign node1539 = (inp[4]) ? node1541 : 1'b1;
													assign node1541 = (inp[10]) ? 1'b0 : node1542;
														assign node1542 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1546 = (inp[11]) ? node1552 : node1547;
											assign node1547 = (inp[9]) ? node1549 : 1'b0;
												assign node1549 = (inp[0]) ? 1'b0 : 1'b1;
											assign node1552 = (inp[8]) ? node1556 : node1553;
												assign node1553 = (inp[4]) ? 1'b1 : 1'b0;
												assign node1556 = (inp[10]) ? node1558 : 1'b0;
													assign node1558 = (inp[4]) ? 1'b0 : 1'b1;
									assign node1561 = (inp[4]) ? node1575 : node1562;
										assign node1562 = (inp[2]) ? node1566 : node1563;
											assign node1563 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1566 = (inp[11]) ? node1570 : node1567;
												assign node1567 = (inp[8]) ? 1'b1 : 1'b0;
												assign node1570 = (inp[8]) ? node1572 : 1'b1;
													assign node1572 = (inp[13]) ? 1'b1 : 1'b0;
										assign node1575 = (inp[11]) ? 1'b0 : node1576;
											assign node1576 = (inp[13]) ? 1'b0 : node1577;
												assign node1577 = (inp[8]) ? 1'b0 : 1'b1;
							assign node1582 = (inp[9]) ? node1614 : node1583;
								assign node1583 = (inp[8]) ? node1603 : node1584;
									assign node1584 = (inp[1]) ? node1592 : node1585;
										assign node1585 = (inp[4]) ? 1'b1 : node1586;
											assign node1586 = (inp[0]) ? node1588 : 1'b1;
												assign node1588 = (inp[14]) ? 1'b1 : 1'b0;
										assign node1592 = (inp[0]) ? node1600 : node1593;
											assign node1593 = (inp[13]) ? node1595 : 1'b0;
												assign node1595 = (inp[10]) ? 1'b0 : node1596;
													assign node1596 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1600 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1603 = (inp[0]) ? node1605 : 1'b1;
										assign node1605 = (inp[2]) ? node1607 : 1'b1;
											assign node1607 = (inp[1]) ? 1'b0 : node1608;
												assign node1608 = (inp[13]) ? 1'b1 : node1609;
													assign node1609 = (inp[4]) ? 1'b1 : 1'b0;
								assign node1614 = (inp[10]) ? node1640 : node1615;
									assign node1615 = (inp[0]) ? node1625 : node1616;
										assign node1616 = (inp[8]) ? 1'b0 : node1617;
											assign node1617 = (inp[4]) ? 1'b1 : node1618;
												assign node1618 = (inp[13]) ? node1620 : 1'b0;
													assign node1620 = (inp[11]) ? 1'b1 : 1'b0;
										assign node1625 = (inp[4]) ? 1'b0 : node1626;
											assign node1626 = (inp[1]) ? node1634 : node1627;
												assign node1627 = (inp[11]) ? node1631 : node1628;
													assign node1628 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1631 = (inp[8]) ? 1'b1 : 1'b0;
												assign node1634 = (inp[11]) ? node1636 : 1'b0;
													assign node1636 = (inp[8]) ? 1'b1 : 1'b0;
									assign node1640 = (inp[4]) ? 1'b1 : node1641;
										assign node1641 = (inp[0]) ? node1647 : node1642;
											assign node1642 = (inp[8]) ? 1'b1 : node1643;
												assign node1643 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1647 = (inp[14]) ? node1649 : 1'b0;
												assign node1649 = (inp[8]) ? node1651 : 1'b1;
													assign node1651 = (inp[1]) ? 1'b0 : 1'b1;
						assign node1655 = (inp[9]) ? node1733 : node1656;
							assign node1656 = (inp[11]) ? node1700 : node1657;
								assign node1657 = (inp[4]) ? node1685 : node1658;
									assign node1658 = (inp[0]) ? node1670 : node1659;
										assign node1659 = (inp[1]) ? node1661 : 1'b0;
											assign node1661 = (inp[8]) ? 1'b0 : node1662;
												assign node1662 = (inp[14]) ? node1664 : 1'b0;
													assign node1664 = (inp[13]) ? 1'b1 : node1665;
														assign node1665 = (inp[2]) ? 1'b1 : 1'b0;
										assign node1670 = (inp[8]) ? node1676 : node1671;
											assign node1671 = (inp[1]) ? 1'b0 : node1672;
												assign node1672 = (inp[2]) ? 1'b1 : 1'b0;
											assign node1676 = (inp[2]) ? node1682 : node1677;
												assign node1677 = (inp[1]) ? 1'b1 : node1678;
													assign node1678 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1682 = (inp[13]) ? 1'b0 : 1'b1;
									assign node1685 = (inp[8]) ? 1'b0 : node1686;
										assign node1686 = (inp[0]) ? 1'b0 : node1687;
											assign node1687 = (inp[1]) ? node1689 : 1'b0;
												assign node1689 = (inp[14]) ? node1693 : node1690;
													assign node1690 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1693 = (inp[2]) ? 1'b1 : node1694;
														assign node1694 = (inp[10]) ? 1'b1 : 1'b0;
								assign node1700 = (inp[14]) ? node1714 : node1701;
									assign node1701 = (inp[0]) ? node1707 : node1702;
										assign node1702 = (inp[8]) ? 1'b0 : node1703;
											assign node1703 = (inp[1]) ? 1'b1 : 1'b0;
										assign node1707 = (inp[4]) ? node1709 : 1'b1;
											assign node1709 = (inp[1]) ? node1711 : 1'b0;
												assign node1711 = (inp[8]) ? 1'b0 : 1'b1;
									assign node1714 = (inp[10]) ? 1'b0 : node1715;
										assign node1715 = (inp[4]) ? node1725 : node1716;
											assign node1716 = (inp[0]) ? node1720 : node1717;
												assign node1717 = (inp[1]) ? 1'b1 : 1'b0;
												assign node1720 = (inp[3]) ? node1722 : 1'b1;
													assign node1722 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1725 = (inp[0]) ? 1'b0 : node1726;
												assign node1726 = (inp[8]) ? 1'b0 : node1727;
													assign node1727 = (inp[1]) ? 1'b1 : 1'b0;
							assign node1733 = (inp[10]) ? node1763 : node1734;
								assign node1734 = (inp[13]) ? node1750 : node1735;
									assign node1735 = (inp[14]) ? node1745 : node1736;
										assign node1736 = (inp[8]) ? node1742 : node1737;
											assign node1737 = (inp[11]) ? 1'b0 : node1738;
												assign node1738 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1742 = (inp[4]) ? 1'b1 : 1'b0;
										assign node1745 = (inp[1]) ? node1747 : 1'b1;
											assign node1747 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1750 = (inp[0]) ? node1752 : 1'b1;
										assign node1752 = (inp[11]) ? node1754 : 1'b1;
											assign node1754 = (inp[8]) ? node1760 : node1755;
												assign node1755 = (inp[2]) ? node1757 : 1'b1;
													assign node1757 = (inp[1]) ? 1'b0 : 1'b1;
												assign node1760 = (inp[4]) ? 1'b1 : 1'b0;
								assign node1763 = (inp[1]) ? node1771 : node1764;
									assign node1764 = (inp[14]) ? 1'b0 : node1765;
										assign node1765 = (inp[4]) ? 1'b0 : node1766;
											assign node1766 = (inp[0]) ? 1'b1 : 1'b0;
									assign node1771 = (inp[8]) ? node1773 : 1'b1;
										assign node1773 = (inp[0]) ? node1775 : 1'b0;
											assign node1775 = (inp[3]) ? 1'b0 : node1776;
												assign node1776 = (inp[14]) ? 1'b0 : 1'b1;
					assign node1780 = (inp[8]) ? node1838 : node1781;
						assign node1781 = (inp[1]) ? node1803 : node1782;
							assign node1782 = (inp[0]) ? node1784 : 1'b1;
								assign node1784 = (inp[4]) ? 1'b1 : node1785;
									assign node1785 = (inp[13]) ? node1791 : node1786;
										assign node1786 = (inp[14]) ? node1788 : 1'b0;
											assign node1788 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1791 = (inp[11]) ? node1797 : node1792;
											assign node1792 = (inp[2]) ? 1'b1 : node1793;
												assign node1793 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1797 = (inp[2]) ? 1'b0 : node1798;
												assign node1798 = (inp[14]) ? 1'b1 : 1'b0;
							assign node1803 = (inp[0]) ? node1821 : node1804;
								assign node1804 = (inp[14]) ? node1810 : node1805;
									assign node1805 = (inp[13]) ? node1807 : 1'b0;
										assign node1807 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1810 = (inp[2]) ? node1816 : node1811;
										assign node1811 = (inp[11]) ? 1'b1 : node1812;
											assign node1812 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1816 = (inp[11]) ? 1'b0 : node1817;
											assign node1817 = (inp[13]) ? 1'b1 : 1'b0;
								assign node1821 = (inp[4]) ? node1823 : 1'b1;
									assign node1823 = (inp[2]) ? node1833 : node1824;
										assign node1824 = (inp[3]) ? node1826 : 1'b1;
											assign node1826 = (inp[13]) ? node1828 : 1'b1;
												assign node1828 = (inp[11]) ? node1830 : 1'b0;
													assign node1830 = (inp[14]) ? 1'b1 : 1'b0;
										assign node1833 = (inp[11]) ? 1'b0 : node1834;
											assign node1834 = (inp[13]) ? 1'b1 : 1'b0;
						assign node1838 = (inp[0]) ? node1840 : 1'b1;
							assign node1840 = (inp[4]) ? 1'b1 : node1841;
								assign node1841 = (inp[13]) ? node1847 : node1842;
									assign node1842 = (inp[14]) ? node1844 : 1'b0;
										assign node1844 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1847 = (inp[9]) ? node1853 : node1848;
										assign node1848 = (inp[11]) ? node1850 : 1'b1;
											assign node1850 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1853 = (inp[7]) ? node1869 : node1854;
											assign node1854 = (inp[1]) ? node1864 : node1855;
												assign node1855 = (inp[14]) ? node1857 : 1'b0;
													assign node1857 = (inp[3]) ? node1861 : node1858;
														assign node1858 = (inp[2]) ? 1'b0 : 1'b1;
														assign node1861 = (inp[2]) ? 1'b1 : 1'b0;
												assign node1864 = (inp[2]) ? node1866 : 1'b1;
													assign node1866 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1869 = (inp[11]) ? 1'b0 : node1870;
												assign node1870 = (inp[3]) ? 1'b0 : 1'b1;

endmodule