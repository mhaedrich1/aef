module dtc_split33_bm98 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node114;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node126;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node227;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node254;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node269;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node282;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node290;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node307;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node326;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node360;
	wire [3-1:0] node363;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node373;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node392;
	wire [3-1:0] node395;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node404;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node411;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node430;

	assign outp = (inp[0]) ? node158 : node1;
		assign node1 = (inp[6]) ? node3 : 3'b111;
			assign node3 = (inp[9]) ? node47 : node4;
				assign node4 = (inp[3]) ? node36 : node5;
					assign node5 = (inp[4]) ? node7 : 3'b100;
						assign node7 = (inp[1]) ? node23 : node8;
							assign node8 = (inp[10]) ? node16 : node9;
								assign node9 = (inp[2]) ? 3'b100 : node10;
									assign node10 = (inp[5]) ? 3'b100 : node11;
										assign node11 = (inp[7]) ? 3'b000 : 3'b100;
								assign node16 = (inp[7]) ? node18 : 3'b100;
									assign node18 = (inp[8]) ? 3'b000 : node19;
										assign node19 = (inp[11]) ? 3'b000 : 3'b000;
							assign node23 = (inp[7]) ? node25 : 3'b000;
								assign node25 = (inp[2]) ? node31 : node26;
									assign node26 = (inp[8]) ? 3'b101 : node27;
										assign node27 = (inp[10]) ? 3'b100 : 3'b101;
									assign node31 = (inp[10]) ? 3'b100 : node32;
										assign node32 = (inp[5]) ? 3'b101 : 3'b100;
					assign node36 = (inp[4]) ? node38 : 3'b010;
						assign node38 = (inp[1]) ? node40 : 3'b010;
							assign node40 = (inp[7]) ? node42 : 3'b010;
								assign node42 = (inp[2]) ? node44 : 3'b110;
									assign node44 = (inp[10]) ? 3'b110 : 3'b010;
				assign node47 = (inp[3]) ? node119 : node48;
					assign node48 = (inp[1]) ? node80 : node49;
						assign node49 = (inp[2]) ? node61 : node50;
							assign node50 = (inp[4]) ? node52 : 3'b001;
								assign node52 = (inp[7]) ? node56 : node53;
									assign node53 = (inp[10]) ? 3'b111 : 3'b101;
									assign node56 = (inp[8]) ? 3'b011 : node57;
										assign node57 = (inp[11]) ? 3'b111 : 3'b011;
							assign node61 = (inp[10]) ? node71 : node62;
								assign node62 = (inp[7]) ? node66 : node63;
									assign node63 = (inp[4]) ? 3'b111 : 3'b101;
									assign node66 = (inp[4]) ? node68 : 3'b101;
										assign node68 = (inp[5]) ? 3'b001 : 3'b101;
								assign node71 = (inp[7]) ? node75 : node72;
									assign node72 = (inp[4]) ? 3'b101 : 3'b001;
									assign node75 = (inp[4]) ? node77 : 3'b101;
										assign node77 = (inp[11]) ? 3'b101 : 3'b001;
						assign node80 = (inp[4]) ? node96 : node81;
							assign node81 = (inp[2]) ? node89 : node82;
								assign node82 = (inp[7]) ? 3'b001 : node83;
									assign node83 = (inp[8]) ? node85 : 3'b100;
										assign node85 = (inp[11]) ? 3'b001 : 3'b100;
								assign node89 = (inp[7]) ? 3'b100 : node90;
									assign node90 = (inp[11]) ? node92 : 3'b100;
										assign node92 = (inp[5]) ? 3'b001 : 3'b100;
							assign node96 = (inp[2]) ? node106 : node97;
								assign node97 = (inp[7]) ? node101 : node98;
									assign node98 = (inp[5]) ? 3'b110 : 3'b100;
									assign node101 = (inp[11]) ? node103 : 3'b110;
										assign node103 = (inp[8]) ? 3'b110 : 3'b001;
								assign node106 = (inp[7]) ? node114 : node107;
									assign node107 = (inp[5]) ? node111 : node108;
										assign node108 = (inp[10]) ? 3'b000 : 3'b110;
										assign node111 = (inp[10]) ? 3'b000 : 3'b000;
									assign node114 = (inp[5]) ? node116 : 3'b001;
										assign node116 = (inp[8]) ? 3'b001 : 3'b110;
					assign node119 = (inp[1]) ? node121 : 3'b111;
						assign node121 = (inp[7]) ? node141 : node122;
							assign node122 = (inp[2]) ? node130 : node123;
								assign node123 = (inp[4]) ? 3'b001 : node124;
									assign node124 = (inp[5]) ? node126 : 3'b111;
										assign node126 = (inp[11]) ? 3'b111 : 3'b011;
								assign node130 = (inp[10]) ? node136 : node131;
									assign node131 = (inp[8]) ? node133 : 3'b111;
										assign node133 = (inp[4]) ? 3'b011 : 3'b111;
									assign node136 = (inp[4]) ? 3'b111 : node137;
										assign node137 = (inp[11]) ? 3'b011 : 3'b011;
							assign node141 = (inp[4]) ? node145 : node142;
								assign node142 = (inp[2]) ? 3'b001 : 3'b101;
								assign node145 = (inp[2]) ? node153 : node146;
									assign node146 = (inp[8]) ? node150 : node147;
										assign node147 = (inp[5]) ? 3'b111 : 3'b011;
										assign node150 = (inp[10]) ? 3'b011 : 3'b011;
									assign node153 = (inp[8]) ? 3'b101 : node154;
										assign node154 = (inp[11]) ? 3'b011 : 3'b101;
		assign node158 = (inp[3]) ? node258 : node159;
			assign node159 = (inp[6]) ? node227 : node160;
				assign node160 = (inp[9]) ? node180 : node161;
					assign node161 = (inp[4]) ? node163 : 3'b010;
						assign node163 = (inp[1]) ? node177 : node164;
							assign node164 = (inp[7]) ? node166 : 3'b010;
								assign node166 = (inp[5]) ? node170 : node167;
									assign node167 = (inp[11]) ? 3'b010 : 3'b000;
									assign node170 = (inp[8]) ? node174 : node171;
										assign node171 = (inp[11]) ? 3'b010 : 3'b000;
										assign node174 = (inp[11]) ? 3'b000 : 3'b010;
							assign node177 = (inp[7]) ? 3'b010 : 3'b000;
					assign node180 = (inp[2]) ? node200 : node181;
						assign node181 = (inp[7]) ? node191 : node182;
							assign node182 = (inp[4]) ? 3'b010 : node183;
								assign node183 = (inp[5]) ? node187 : node184;
									assign node184 = (inp[11]) ? 3'b010 : 3'b000;
									assign node187 = (inp[11]) ? 3'b000 : 3'b010;
							assign node191 = (inp[4]) ? node193 : 3'b000;
								assign node193 = (inp[5]) ? node197 : node194;
									assign node194 = (inp[11]) ? 3'b010 : 3'b000;
									assign node197 = (inp[11]) ? 3'b000 : 3'b010;
						assign node200 = (inp[7]) ? node220 : node201;
							assign node201 = (inp[5]) ? node209 : node202;
								assign node202 = (inp[1]) ? node204 : 3'b010;
									assign node204 = (inp[8]) ? 3'b000 : node205;
										assign node205 = (inp[10]) ? 3'b010 : 3'b000;
								assign node209 = (inp[4]) ? node213 : node210;
									assign node210 = (inp[11]) ? 3'b000 : 3'b010;
									assign node213 = (inp[11]) ? node217 : node214;
										assign node214 = (inp[10]) ? 3'b000 : 3'b000;
										assign node217 = (inp[1]) ? 3'b000 : 3'b000;
							assign node220 = (inp[4]) ? node222 : 3'b010;
								assign node222 = (inp[11]) ? 3'b010 : node223;
									assign node223 = (inp[5]) ? 3'b100 : 3'b010;
				assign node227 = (inp[9]) ? node229 : 3'b000;
					assign node229 = (inp[4]) ? node231 : 3'b000;
						assign node231 = (inp[7]) ? node243 : node232;
							assign node232 = (inp[1]) ? 3'b100 : node233;
								assign node233 = (inp[11]) ? node237 : node234;
									assign node234 = (inp[8]) ? 3'b110 : 3'b010;
									assign node237 = (inp[8]) ? 3'b000 : node238;
										assign node238 = (inp[2]) ? 3'b100 : 3'b110;
							assign node243 = (inp[1]) ? 3'b000 : node244;
								assign node244 = (inp[11]) ? node252 : node245;
									assign node245 = (inp[5]) ? node249 : node246;
										assign node246 = (inp[2]) ? 3'b010 : 3'b010;
										assign node249 = (inp[8]) ? 3'b110 : 3'b000;
									assign node252 = (inp[8]) ? node254 : 3'b100;
										assign node254 = (inp[2]) ? 3'b000 : 3'b000;
			assign node258 = (inp[6]) ? node348 : node259;
				assign node259 = (inp[9]) ? node307 : node260;
					assign node260 = (inp[1]) ? node282 : node261;
						assign node261 = (inp[4]) ? node263 : 3'b001;
							assign node263 = (inp[7]) ? node279 : node264;
								assign node264 = (inp[2]) ? node272 : node265;
									assign node265 = (inp[5]) ? node269 : node266;
										assign node266 = (inp[11]) ? 3'b011 : 3'b011;
										assign node269 = (inp[11]) ? 3'b011 : 3'b111;
									assign node272 = (inp[10]) ? node276 : node273;
										assign node273 = (inp[5]) ? 3'b001 : 3'b101;
										assign node276 = (inp[5]) ? 3'b101 : 3'b001;
								assign node279 = (inp[2]) ? 3'b001 : 3'b101;
						assign node282 = (inp[4]) ? node284 : 3'b000;
							assign node284 = (inp[7]) ? node298 : node285;
								assign node285 = (inp[2]) ? node293 : node286;
									assign node286 = (inp[11]) ? node290 : node287;
										assign node287 = (inp[8]) ? 3'b001 : 3'b101;
										assign node290 = (inp[10]) ? 3'b001 : 3'b101;
									assign node293 = (inp[11]) ? 3'b110 : node294;
										assign node294 = (inp[8]) ? 3'b110 : 3'b001;
								assign node298 = (inp[11]) ? node300 : 3'b010;
									assign node300 = (inp[5]) ? node304 : node301;
										assign node301 = (inp[10]) ? 3'b100 : 3'b110;
										assign node304 = (inp[2]) ? 3'b000 : 3'b010;
					assign node307 = (inp[1]) ? node309 : 3'b111;
						assign node309 = (inp[4]) ? node331 : node310;
							assign node310 = (inp[11]) ? node320 : node311;
								assign node311 = (inp[8]) ? node315 : node312;
									assign node312 = (inp[5]) ? 3'b010 : 3'b110;
									assign node315 = (inp[10]) ? 3'b010 : node316;
										assign node316 = (inp[5]) ? 3'b001 : 3'b101;
								assign node320 = (inp[8]) ? node326 : node321;
									assign node321 = (inp[2]) ? 3'b001 : node322;
										assign node322 = (inp[5]) ? 3'b101 : 3'b001;
									assign node326 = (inp[7]) ? node328 : 3'b010;
										assign node328 = (inp[10]) ? 3'b010 : 3'b001;
							assign node331 = (inp[7]) ? node343 : node332;
								assign node332 = (inp[10]) ? node338 : node333;
									assign node333 = (inp[5]) ? node335 : 3'b111;
										assign node335 = (inp[11]) ? 3'b111 : 3'b011;
									assign node338 = (inp[8]) ? 3'b011 : node339;
										assign node339 = (inp[11]) ? 3'b111 : 3'b011;
								assign node343 = (inp[5]) ? 3'b011 : node344;
									assign node344 = (inp[2]) ? 3'b101 : 3'b001;
				assign node348 = (inp[9]) ? node366 : node349;
					assign node349 = (inp[4]) ? node351 : 3'b000;
						assign node351 = (inp[1]) ? node363 : node352;
							assign node352 = (inp[7]) ? node354 : 3'b001;
								assign node354 = (inp[11]) ? node358 : node355;
									assign node355 = (inp[10]) ? 3'b100 : 3'b000;
									assign node358 = (inp[2]) ? node360 : 3'b010;
										assign node360 = (inp[10]) ? 3'b010 : 3'b010;
							assign node363 = (inp[7]) ? 3'b000 : 3'b100;
					assign node366 = (inp[1]) ? node398 : node367;
						assign node367 = (inp[7]) ? node383 : node368;
							assign node368 = (inp[4]) ? node376 : node369;
								assign node369 = (inp[5]) ? node373 : node370;
									assign node370 = (inp[11]) ? 3'b001 : 3'b101;
									assign node373 = (inp[11]) ? 3'b101 : 3'b001;
								assign node376 = (inp[11]) ? 3'b101 : node377;
									assign node377 = (inp[10]) ? 3'b010 : node378;
										assign node378 = (inp[2]) ? 3'b001 : 3'b010;
							assign node383 = (inp[4]) ? node387 : node384;
								assign node384 = (inp[2]) ? 3'b010 : 3'b110;
								assign node387 = (inp[2]) ? node395 : node388;
									assign node388 = (inp[8]) ? node392 : node389;
										assign node389 = (inp[10]) ? 3'b101 : 3'b001;
										assign node392 = (inp[10]) ? 3'b001 : 3'b001;
									assign node395 = (inp[8]) ? 3'b010 : 3'b001;
						assign node398 = (inp[7]) ? node416 : node399;
							assign node399 = (inp[4]) ? node407 : node400;
								assign node400 = (inp[5]) ? node404 : node401;
									assign node401 = (inp[11]) ? 3'b010 : 3'b110;
									assign node404 = (inp[11]) ? 3'b110 : 3'b010;
								assign node407 = (inp[5]) ? node411 : node408;
									assign node408 = (inp[10]) ? 3'b001 : 3'b000;
									assign node411 = (inp[8]) ? node413 : 3'b000;
										assign node413 = (inp[10]) ? 3'b110 : 3'b010;
							assign node416 = (inp[4]) ? node420 : node417;
								assign node417 = (inp[2]) ? 3'b000 : 3'b100;
								assign node420 = (inp[2]) ? node426 : node421;
									assign node421 = (inp[11]) ? 3'b110 : node422;
										assign node422 = (inp[5]) ? 3'b010 : 3'b110;
									assign node426 = (inp[8]) ? node430 : node427;
										assign node427 = (inp[11]) ? 3'b010 : 3'b100;
										assign node430 = (inp[11]) ? 3'b100 : 3'b000;

endmodule