module dtc_split875_bm9 (
	input  wire [8-1:0] inp,
	output wire [8-1:0] outp
);

	wire [8-1:0] node1;
	wire [8-1:0] node2;
	wire [8-1:0] node3;
	wire [8-1:0] node4;
	wire [8-1:0] node5;
	wire [8-1:0] node6;
	wire [8-1:0] node7;
	wire [8-1:0] node10;
	wire [8-1:0] node13;
	wire [8-1:0] node16;
	wire [8-1:0] node17;
	wire [8-1:0] node18;
	wire [8-1:0] node21;
	wire [8-1:0] node24;
	wire [8-1:0] node25;
	wire [8-1:0] node28;
	wire [8-1:0] node31;
	wire [8-1:0] node32;
	wire [8-1:0] node33;
	wire [8-1:0] node34;
	wire [8-1:0] node37;
	wire [8-1:0] node40;
	wire [8-1:0] node41;
	wire [8-1:0] node44;
	wire [8-1:0] node47;
	wire [8-1:0] node48;
	wire [8-1:0] node49;
	wire [8-1:0] node52;
	wire [8-1:0] node55;
	wire [8-1:0] node57;
	wire [8-1:0] node60;
	wire [8-1:0] node61;
	wire [8-1:0] node62;
	wire [8-1:0] node63;
	wire [8-1:0] node64;
	wire [8-1:0] node67;
	wire [8-1:0] node70;
	wire [8-1:0] node73;
	wire [8-1:0] node74;
	wire [8-1:0] node76;
	wire [8-1:0] node79;
	wire [8-1:0] node80;
	wire [8-1:0] node84;
	wire [8-1:0] node85;
	wire [8-1:0] node86;
	wire [8-1:0] node89;
	wire [8-1:0] node92;
	wire [8-1:0] node93;
	wire [8-1:0] node94;
	wire [8-1:0] node97;
	wire [8-1:0] node100;
	wire [8-1:0] node101;
	wire [8-1:0] node105;
	wire [8-1:0] node106;
	wire [8-1:0] node107;
	wire [8-1:0] node108;
	wire [8-1:0] node109;
	wire [8-1:0] node112;
	wire [8-1:0] node114;
	wire [8-1:0] node117;
	wire [8-1:0] node118;
	wire [8-1:0] node119;
	wire [8-1:0] node122;
	wire [8-1:0] node125;
	wire [8-1:0] node127;
	wire [8-1:0] node130;
	wire [8-1:0] node131;
	wire [8-1:0] node132;
	wire [8-1:0] node133;
	wire [8-1:0] node136;
	wire [8-1:0] node139;
	wire [8-1:0] node140;
	wire [8-1:0] node143;
	wire [8-1:0] node146;
	wire [8-1:0] node147;
	wire [8-1:0] node148;
	wire [8-1:0] node151;
	wire [8-1:0] node154;
	wire [8-1:0] node155;
	wire [8-1:0] node158;
	wire [8-1:0] node161;
	wire [8-1:0] node162;
	wire [8-1:0] node163;
	wire [8-1:0] node164;
	wire [8-1:0] node165;
	wire [8-1:0] node168;
	wire [8-1:0] node171;
	wire [8-1:0] node172;
	wire [8-1:0] node175;
	wire [8-1:0] node178;
	wire [8-1:0] node179;
	wire [8-1:0] node180;
	wire [8-1:0] node183;
	wire [8-1:0] node186;
	wire [8-1:0] node188;
	wire [8-1:0] node191;
	wire [8-1:0] node192;
	wire [8-1:0] node193;
	wire [8-1:0] node194;
	wire [8-1:0] node197;
	wire [8-1:0] node200;
	wire [8-1:0] node201;
	wire [8-1:0] node204;
	wire [8-1:0] node207;
	wire [8-1:0] node208;
	wire [8-1:0] node211;
	wire [8-1:0] node214;
	wire [8-1:0] node215;
	wire [8-1:0] node216;
	wire [8-1:0] node217;
	wire [8-1:0] node218;
	wire [8-1:0] node219;
	wire [8-1:0] node221;
	wire [8-1:0] node224;
	wire [8-1:0] node225;
	wire [8-1:0] node228;
	wire [8-1:0] node231;
	wire [8-1:0] node232;
	wire [8-1:0] node233;
	wire [8-1:0] node236;
	wire [8-1:0] node239;
	wire [8-1:0] node240;
	wire [8-1:0] node243;
	wire [8-1:0] node246;
	wire [8-1:0] node247;
	wire [8-1:0] node248;
	wire [8-1:0] node249;
	wire [8-1:0] node252;
	wire [8-1:0] node255;
	wire [8-1:0] node257;
	wire [8-1:0] node260;
	wire [8-1:0] node261;
	wire [8-1:0] node262;
	wire [8-1:0] node265;
	wire [8-1:0] node268;
	wire [8-1:0] node269;
	wire [8-1:0] node272;
	wire [8-1:0] node275;
	wire [8-1:0] node276;
	wire [8-1:0] node277;
	wire [8-1:0] node278;
	wire [8-1:0] node279;
	wire [8-1:0] node282;
	wire [8-1:0] node285;
	wire [8-1:0] node286;
	wire [8-1:0] node289;
	wire [8-1:0] node292;
	wire [8-1:0] node293;
	wire [8-1:0] node295;
	wire [8-1:0] node298;
	wire [8-1:0] node299;
	wire [8-1:0] node302;
	wire [8-1:0] node305;
	wire [8-1:0] node306;
	wire [8-1:0] node307;
	wire [8-1:0] node308;
	wire [8-1:0] node311;
	wire [8-1:0] node314;
	wire [8-1:0] node316;
	wire [8-1:0] node319;
	wire [8-1:0] node320;
	wire [8-1:0] node321;
	wire [8-1:0] node324;
	wire [8-1:0] node327;
	wire [8-1:0] node329;
	wire [8-1:0] node332;
	wire [8-1:0] node333;
	wire [8-1:0] node334;
	wire [8-1:0] node335;
	wire [8-1:0] node336;
	wire [8-1:0] node337;
	wire [8-1:0] node340;
	wire [8-1:0] node343;
	wire [8-1:0] node345;
	wire [8-1:0] node348;
	wire [8-1:0] node349;
	wire [8-1:0] node350;
	wire [8-1:0] node353;
	wire [8-1:0] node356;
	wire [8-1:0] node357;
	wire [8-1:0] node360;
	wire [8-1:0] node363;
	wire [8-1:0] node364;
	wire [8-1:0] node365;
	wire [8-1:0] node366;
	wire [8-1:0] node369;
	wire [8-1:0] node372;
	wire [8-1:0] node374;
	wire [8-1:0] node377;
	wire [8-1:0] node378;
	wire [8-1:0] node380;
	wire [8-1:0] node383;
	wire [8-1:0] node384;
	wire [8-1:0] node388;
	wire [8-1:0] node389;
	wire [8-1:0] node390;
	wire [8-1:0] node391;
	wire [8-1:0] node392;
	wire [8-1:0] node395;
	wire [8-1:0] node398;
	wire [8-1:0] node399;
	wire [8-1:0] node402;
	wire [8-1:0] node405;
	wire [8-1:0] node406;
	wire [8-1:0] node407;
	wire [8-1:0] node410;
	wire [8-1:0] node413;
	wire [8-1:0] node414;
	wire [8-1:0] node417;
	wire [8-1:0] node420;
	wire [8-1:0] node421;
	wire [8-1:0] node422;
	wire [8-1:0] node423;
	wire [8-1:0] node427;
	wire [8-1:0] node428;
	wire [8-1:0] node431;
	wire [8-1:0] node434;
	wire [8-1:0] node435;
	wire [8-1:0] node437;
	wire [8-1:0] node440;
	wire [8-1:0] node441;
	wire [8-1:0] node444;

	assign outp = (inp[5]) ? node214 : node1;
		assign node1 = (inp[2]) ? node105 : node2;
			assign node2 = (inp[4]) ? node60 : node3;
				assign node3 = (inp[1]) ? node31 : node4;
					assign node4 = (inp[7]) ? node16 : node5;
						assign node5 = (inp[0]) ? node13 : node6;
							assign node6 = (inp[6]) ? node10 : node7;
								assign node7 = (inp[3]) ? 8'b10000110 : 8'b10111110;
								assign node10 = (inp[3]) ? 8'b11001010 : 8'b10000100;
							assign node13 = (inp[6]) ? 8'b11001000 : 8'b01100000;
						assign node16 = (inp[3]) ? node24 : node17;
							assign node17 = (inp[6]) ? node21 : node18;
								assign node18 = (inp[0]) ? 8'b01010001 : 8'b00110000;
								assign node21 = (inp[0]) ? 8'b10000000 : 8'b10101010;
							assign node24 = (inp[0]) ? node28 : node25;
								assign node25 = (inp[6]) ? 8'b11000001 : 8'b10011001;
								assign node28 = (inp[6]) ? 8'b00011101 : 8'b10100010;
					assign node31 = (inp[3]) ? node47 : node32;
						assign node32 = (inp[7]) ? node40 : node33;
							assign node33 = (inp[6]) ? node37 : node34;
								assign node34 = (inp[0]) ? 8'b10100100 : 8'b00101111;
								assign node37 = (inp[0]) ? 8'b11010001 : 8'b10110011;
							assign node40 = (inp[6]) ? node44 : node41;
								assign node41 = (inp[0]) ? 8'b10001011 : 8'b01011010;
								assign node44 = (inp[0]) ? 8'b10110110 : 8'b00011110;
						assign node47 = (inp[0]) ? node55 : node48;
							assign node48 = (inp[7]) ? node52 : node49;
								assign node49 = (inp[6]) ? 8'b00011000 : 8'b11011000;
								assign node52 = (inp[6]) ? 8'b01010101 : 8'b01111101;
							assign node55 = (inp[6]) ? node57 : 8'b01110010;
								assign node57 = (inp[7]) ? 8'b01000010 : 8'b01011111;
				assign node60 = (inp[3]) ? node84 : node61;
					assign node61 = (inp[6]) ? node73 : node62;
						assign node62 = (inp[7]) ? node70 : node63;
							assign node63 = (inp[1]) ? node67 : node64;
								assign node64 = (inp[0]) ? 8'b01000000 : 8'b01100100;
								assign node67 = (inp[0]) ? 8'b01001101 : 8'b00000100;
							assign node70 = (inp[0]) ? 8'b11110000 : 8'b01101011;
						assign node73 = (inp[1]) ? node79 : node74;
							assign node74 = (inp[7]) ? node76 : 8'b11111100;
								assign node76 = (inp[0]) ? 8'b01010011 : 8'b01011101;
							assign node79 = (inp[0]) ? 8'b10011011 : node80;
								assign node80 = (inp[7]) ? 8'b01100011 : 8'b01001011;
					assign node84 = (inp[1]) ? node92 : node85;
						assign node85 = (inp[6]) ? node89 : node86;
							assign node86 = (inp[0]) ? 8'b11001011 : 8'b00001101;
							assign node89 = (inp[0]) ? 8'b00111101 : 8'b01110101;
						assign node92 = (inp[0]) ? node100 : node93;
							assign node93 = (inp[7]) ? node97 : node94;
								assign node94 = (inp[6]) ? 8'b10010100 : 8'b10010001;
								assign node97 = (inp[6]) ? 8'b10111000 : 8'b10100011;
							assign node100 = (inp[6]) ? 8'b01000011 : node101;
								assign node101 = (inp[7]) ? 8'b11000100 : 8'b10111100;
			assign node105 = (inp[3]) ? node161 : node106;
				assign node106 = (inp[7]) ? node130 : node107;
					assign node107 = (inp[4]) ? node117 : node108;
						assign node108 = (inp[0]) ? node112 : node109;
							assign node109 = (inp[1]) ? 8'b01110110 : 8'b11110111;
							assign node112 = (inp[1]) ? node114 : 8'b00100001;
								assign node114 = (inp[6]) ? 8'b01111011 : 8'b11010011;
						assign node117 = (inp[6]) ? node125 : node118;
							assign node118 = (inp[0]) ? node122 : node119;
								assign node119 = (inp[1]) ? 8'b10100001 : 8'b10110000;
								assign node122 = (inp[1]) ? 8'b11100001 : 8'b01011011;
							assign node125 = (inp[0]) ? node127 : 8'b10101101;
								assign node127 = (inp[1]) ? 8'b11110100 : 8'b10110111;
					assign node130 = (inp[0]) ? node146 : node131;
						assign node131 = (inp[1]) ? node139 : node132;
							assign node132 = (inp[6]) ? node136 : node133;
								assign node133 = (inp[4]) ? 8'b01010010 : 8'b00111001;
								assign node136 = (inp[4]) ? 8'b10011000 : 8'b11001001;
							assign node139 = (inp[4]) ? node143 : node140;
								assign node140 = (inp[6]) ? 8'b00111000 : 8'b11111011;
								assign node143 = (inp[6]) ? 8'b11100111 : 8'b10101100;
						assign node146 = (inp[4]) ? node154 : node147;
							assign node147 = (inp[1]) ? node151 : node148;
								assign node148 = (inp[6]) ? 8'b11100101 : 8'b10111001;
								assign node151 = (inp[6]) ? 8'b00100011 : 8'b10010111;
							assign node154 = (inp[1]) ? node158 : node155;
								assign node155 = (inp[6]) ? 8'b10111111 : 8'b10011101;
								assign node158 = (inp[6]) ? 8'b11011001 : 8'b11111111;
				assign node161 = (inp[1]) ? node191 : node162;
					assign node162 = (inp[6]) ? node178 : node163;
						assign node163 = (inp[0]) ? node171 : node164;
							assign node164 = (inp[7]) ? node168 : node165;
								assign node165 = (inp[4]) ? 8'b10001100 : 8'b11111010;
								assign node168 = (inp[4]) ? 8'b11100011 : 8'b00110111;
							assign node171 = (inp[4]) ? node175 : node172;
								assign node172 = (inp[7]) ? 8'b01101101 : 8'b01001001;
								assign node175 = (inp[7]) ? 8'b00011001 : 8'b01101000;
						assign node178 = (inp[4]) ? node186 : node179;
							assign node179 = (inp[0]) ? node183 : node180;
								assign node180 = (inp[7]) ? 8'b11100100 : 8'b00000001;
								assign node183 = (inp[7]) ? 8'b10111010 : 8'b10100110;
							assign node186 = (inp[7]) ? node188 : 8'b11100000;
								assign node188 = (inp[0]) ? 8'b01100001 : 8'b00010001;
					assign node191 = (inp[4]) ? node207 : node192;
						assign node192 = (inp[6]) ? node200 : node193;
							assign node193 = (inp[7]) ? node197 : node194;
								assign node194 = (inp[0]) ? 8'b11011111 : 8'b11001110;
								assign node197 = (inp[0]) ? 8'b11101011 : 8'b01100111;
							assign node200 = (inp[0]) ? node204 : node201;
								assign node201 = (inp[7]) ? 8'b00001111 : 8'b00101101;
								assign node204 = (inp[7]) ? 8'b10000001 : 8'b11001111;
						assign node207 = (inp[0]) ? node211 : node208;
							assign node208 = (inp[7]) ? 8'b11110010 : 8'b11100110;
							assign node211 = (inp[6]) ? 8'b00001100 : 8'b10100101;
		assign node214 = (inp[4]) ? node332 : node215;
			assign node215 = (inp[0]) ? node275 : node216;
				assign node216 = (inp[1]) ? node246 : node217;
					assign node217 = (inp[6]) ? node231 : node218;
						assign node218 = (inp[7]) ? node224 : node219;
							assign node219 = (inp[2]) ? node221 : 8'b11000110;
								assign node221 = (inp[3]) ? 8'b10011010 : 8'b11111001;
							assign node224 = (inp[2]) ? node228 : node225;
								assign node225 = (inp[3]) ? 8'b11011101 : 8'b00101000;
								assign node228 = (inp[3]) ? 8'b00001000 : 8'b01011110;
						assign node231 = (inp[3]) ? node239 : node232;
							assign node232 = (inp[2]) ? node236 : node233;
								assign node233 = (inp[7]) ? 8'b10000111 : 8'b10010110;
								assign node236 = (inp[7]) ? 8'b10110100 : 8'b10100111;
							assign node239 = (inp[2]) ? node243 : node240;
								assign node240 = (inp[7]) ? 8'b00010011 : 8'b11010111;
								assign node243 = (inp[7]) ? 8'b10001101 : 8'b01001000;
					assign node246 = (inp[3]) ? node260 : node247;
						assign node247 = (inp[7]) ? node255 : node248;
							assign node248 = (inp[2]) ? node252 : node249;
								assign node249 = (inp[6]) ? 8'b11011011 : 8'b01111111;
								assign node252 = (inp[6]) ? 8'b10011111 : 8'b00010111;
							assign node255 = (inp[6]) ? node257 : 8'b00000011;
								assign node257 = (inp[2]) ? 8'b01000111 : 8'b01011001;
						assign node260 = (inp[6]) ? node268 : node261;
							assign node261 = (inp[2]) ? node265 : node262;
								assign node262 = (inp[7]) ? 8'b01000110 : 8'b01110000;
								assign node265 = (inp[7]) ? 8'b11110011 : 8'b01110011;
							assign node268 = (inp[7]) ? node272 : node269;
								assign node269 = (inp[2]) ? 8'b01001111 : 8'b11101101;
								assign node272 = (inp[2]) ? 8'b11101001 : 8'b11110110;
				assign node275 = (inp[7]) ? node305 : node276;
					assign node276 = (inp[1]) ? node292 : node277;
						assign node277 = (inp[3]) ? node285 : node278;
							assign node278 = (inp[2]) ? node282 : node279;
								assign node279 = (inp[6]) ? 8'b11110101 : 8'b11000000;
								assign node282 = (inp[6]) ? 8'b10101000 : 8'b11101010;
							assign node285 = (inp[6]) ? node289 : node286;
								assign node286 = (inp[2]) ? 8'b00110011 : 8'b10100000;
								assign node289 = (inp[2]) ? 8'b00100101 : 8'b00100111;
						assign node292 = (inp[2]) ? node298 : node293;
							assign node293 = (inp[6]) ? node295 : 8'b11010000;
								assign node295 = (inp[3]) ? 8'b00110010 : 8'b11011010;
							assign node298 = (inp[6]) ? node302 : node299;
								assign node299 = (inp[3]) ? 8'b01111001 : 8'b00100010;
								assign node302 = (inp[3]) ? 8'b00000010 : 8'b01110001;
					assign node305 = (inp[1]) ? node319 : node306;
						assign node306 = (inp[6]) ? node314 : node307;
							assign node307 = (inp[3]) ? node311 : node308;
								assign node308 = (inp[2]) ? 8'b01100010 : 8'b10111101;
								assign node311 = (inp[2]) ? 8'b00111010 : 8'b00011010;
							assign node314 = (inp[3]) ? node316 : 8'b10000011;
								assign node316 = (inp[2]) ? 8'b00101011 : 8'b11101111;
						assign node319 = (inp[6]) ? node327 : node320;
							assign node320 = (inp[3]) ? node324 : node321;
								assign node321 = (inp[2]) ? 8'b11000010 : 8'b01000101;
								assign node324 = (inp[2]) ? 8'b11000101 : 8'b10101001;
							assign node327 = (inp[3]) ? node329 : 8'b00101100;
								assign node329 = (inp[2]) ? 8'b11111101 : 8'b01110111;
			assign node332 = (inp[3]) ? node388 : node333;
				assign node333 = (inp[2]) ? node363 : node334;
					assign node334 = (inp[7]) ? node348 : node335;
						assign node335 = (inp[1]) ? node343 : node336;
							assign node336 = (inp[0]) ? node340 : node337;
								assign node337 = (inp[6]) ? 8'b11010100 : 8'b01111110;
								assign node340 = (inp[6]) ? 8'b00110100 : 8'b11110001;
							assign node343 = (inp[0]) ? node345 : 8'b01101010;
								assign node345 = (inp[6]) ? 8'b01110100 : 8'b01100110;
						assign node348 = (inp[1]) ? node356 : node349;
							assign node349 = (inp[6]) ? node353 : node350;
								assign node350 = (inp[0]) ? 8'b01111000 : 8'b00100000;
								assign node353 = (inp[0]) ? 8'b00001011 : 8'b11101000;
							assign node356 = (inp[0]) ? node360 : node357;
								assign node357 = (inp[6]) ? 8'b00111111 : 8'b01111100;
								assign node360 = (inp[6]) ? 8'b00010000 : 8'b10000101;
					assign node363 = (inp[7]) ? node377 : node364;
						assign node364 = (inp[1]) ? node372 : node365;
							assign node365 = (inp[0]) ? node369 : node366;
								assign node366 = (inp[6]) ? 8'b10001010 : 8'b10010101;
								assign node369 = (inp[6]) ? 8'b00001110 : 8'b00001010;
							assign node372 = (inp[0]) ? node374 : 8'b00110101;
								assign node374 = (inp[6]) ? 8'b11000111 : 8'b01000001;
						assign node377 = (inp[1]) ? node383 : node378;
							assign node378 = (inp[6]) ? node380 : 8'b11111110;
								assign node380 = (inp[0]) ? 8'b00110110 : 8'b00000110;
							assign node383 = (inp[0]) ? 8'b00111110 : node384;
								assign node384 = (inp[6]) ? 8'b01101001 : 8'b00101110;
				assign node388 = (inp[7]) ? node420 : node389;
					assign node389 = (inp[6]) ? node405 : node390;
						assign node390 = (inp[0]) ? node398 : node391;
							assign node391 = (inp[1]) ? node395 : node392;
								assign node392 = (inp[2]) ? 8'b11001100 : 8'b10110010;
								assign node395 = (inp[2]) ? 8'b10000010 : 8'b10001110;
							assign node398 = (inp[2]) ? node402 : node399;
								assign node399 = (inp[1]) ? 8'b01001100 : 8'b00000000;
								assign node402 = (inp[1]) ? 8'b10101011 : 8'b00100110;
						assign node405 = (inp[1]) ? node413 : node406;
							assign node406 = (inp[2]) ? node410 : node407;
								assign node407 = (inp[0]) ? 8'b00011011 : 8'b00000111;
								assign node410 = (inp[0]) ? 8'b00011111 : 8'b10111011;
							assign node413 = (inp[2]) ? node417 : node414;
								assign node414 = (inp[0]) ? 8'b11011110 : 8'b10001111;
								assign node417 = (inp[0]) ? 8'b10010000 : 8'b10001001;
					assign node420 = (inp[1]) ? node434 : node421;
						assign node421 = (inp[6]) ? node427 : node422;
							assign node422 = (inp[2]) ? 8'b00010101 : node423;
								assign node423 = (inp[0]) ? 8'b11010101 : 8'b11011100;
							assign node427 = (inp[2]) ? node431 : node428;
								assign node428 = (inp[0]) ? 8'b00001001 : 8'b00000101;
								assign node431 = (inp[0]) ? 8'b01001110 : 8'b11111000;
						assign node434 = (inp[2]) ? node440 : node435;
							assign node435 = (inp[0]) ? node437 : 8'b11100010;
								assign node437 = (inp[6]) ? 8'b00101010 : 8'b00101001;
							assign node440 = (inp[0]) ? node444 : node441;
								assign node441 = (inp[6]) ? 8'b01011100 : 8'b10001000;
								assign node444 = (inp[6]) ? 8'b01001010 : 8'b01010110;

endmodule