module dtc_split33_bm24 (
	input  wire [13-1:0] inp,
	output wire [13-1:0] outp
);

	wire [13-1:0] node1;
	wire [13-1:0] node2;
	wire [13-1:0] node3;
	wire [13-1:0] node4;
	wire [13-1:0] node5;
	wire [13-1:0] node6;
	wire [13-1:0] node7;
	wire [13-1:0] node8;
	wire [13-1:0] node9;
	wire [13-1:0] node11;
	wire [13-1:0] node14;
	wire [13-1:0] node15;
	wire [13-1:0] node18;
	wire [13-1:0] node21;
	wire [13-1:0] node22;
	wire [13-1:0] node23;
	wire [13-1:0] node27;
	wire [13-1:0] node29;
	wire [13-1:0] node32;
	wire [13-1:0] node33;
	wire [13-1:0] node34;
	wire [13-1:0] node38;
	wire [13-1:0] node39;
	wire [13-1:0] node41;
	wire [13-1:0] node44;
	wire [13-1:0] node45;
	wire [13-1:0] node48;
	wire [13-1:0] node51;
	wire [13-1:0] node52;
	wire [13-1:0] node53;
	wire [13-1:0] node54;
	wire [13-1:0] node56;
	wire [13-1:0] node59;
	wire [13-1:0] node60;
	wire [13-1:0] node63;
	wire [13-1:0] node66;
	wire [13-1:0] node67;
	wire [13-1:0] node70;
	wire [13-1:0] node71;
	wire [13-1:0] node75;
	wire [13-1:0] node76;
	wire [13-1:0] node77;
	wire [13-1:0] node80;
	wire [13-1:0] node82;
	wire [13-1:0] node85;
	wire [13-1:0] node86;
	wire [13-1:0] node89;
	wire [13-1:0] node90;
	wire [13-1:0] node93;
	wire [13-1:0] node96;
	wire [13-1:0] node97;
	wire [13-1:0] node98;
	wire [13-1:0] node99;
	wire [13-1:0] node100;
	wire [13-1:0] node102;
	wire [13-1:0] node105;
	wire [13-1:0] node106;
	wire [13-1:0] node110;
	wire [13-1:0] node111;
	wire [13-1:0] node113;
	wire [13-1:0] node116;
	wire [13-1:0] node117;
	wire [13-1:0] node120;
	wire [13-1:0] node123;
	wire [13-1:0] node124;
	wire [13-1:0] node125;
	wire [13-1:0] node126;
	wire [13-1:0] node129;
	wire [13-1:0] node132;
	wire [13-1:0] node133;
	wire [13-1:0] node137;
	wire [13-1:0] node138;
	wire [13-1:0] node139;
	wire [13-1:0] node143;
	wire [13-1:0] node144;
	wire [13-1:0] node148;
	wire [13-1:0] node149;
	wire [13-1:0] node150;
	wire [13-1:0] node151;
	wire [13-1:0] node154;
	wire [13-1:0] node155;
	wire [13-1:0] node159;
	wire [13-1:0] node160;
	wire [13-1:0] node161;
	wire [13-1:0] node164;
	wire [13-1:0] node167;
	wire [13-1:0] node170;
	wire [13-1:0] node171;
	wire [13-1:0] node172;
	wire [13-1:0] node173;
	wire [13-1:0] node176;
	wire [13-1:0] node179;
	wire [13-1:0] node180;
	wire [13-1:0] node183;
	wire [13-1:0] node186;
	wire [13-1:0] node187;
	wire [13-1:0] node188;
	wire [13-1:0] node191;
	wire [13-1:0] node194;
	wire [13-1:0] node195;
	wire [13-1:0] node198;
	wire [13-1:0] node201;
	wire [13-1:0] node202;
	wire [13-1:0] node203;
	wire [13-1:0] node204;
	wire [13-1:0] node205;
	wire [13-1:0] node206;
	wire [13-1:0] node208;
	wire [13-1:0] node211;
	wire [13-1:0] node213;
	wire [13-1:0] node216;
	wire [13-1:0] node217;
	wire [13-1:0] node218;
	wire [13-1:0] node221;
	wire [13-1:0] node224;
	wire [13-1:0] node225;
	wire [13-1:0] node229;
	wire [13-1:0] node230;
	wire [13-1:0] node231;
	wire [13-1:0] node232;
	wire [13-1:0] node236;
	wire [13-1:0] node237;
	wire [13-1:0] node241;
	wire [13-1:0] node242;
	wire [13-1:0] node243;
	wire [13-1:0] node247;
	wire [13-1:0] node249;
	wire [13-1:0] node252;
	wire [13-1:0] node253;
	wire [13-1:0] node254;
	wire [13-1:0] node255;
	wire [13-1:0] node256;
	wire [13-1:0] node259;
	wire [13-1:0] node262;
	wire [13-1:0] node265;
	wire [13-1:0] node266;
	wire [13-1:0] node267;
	wire [13-1:0] node270;
	wire [13-1:0] node273;
	wire [13-1:0] node274;
	wire [13-1:0] node278;
	wire [13-1:0] node279;
	wire [13-1:0] node281;
	wire [13-1:0] node282;
	wire [13-1:0] node285;
	wire [13-1:0] node288;
	wire [13-1:0] node289;
	wire [13-1:0] node290;
	wire [13-1:0] node293;
	wire [13-1:0] node296;
	wire [13-1:0] node298;
	wire [13-1:0] node301;
	wire [13-1:0] node302;
	wire [13-1:0] node303;
	wire [13-1:0] node304;
	wire [13-1:0] node305;
	wire [13-1:0] node306;
	wire [13-1:0] node309;
	wire [13-1:0] node312;
	wire [13-1:0] node313;
	wire [13-1:0] node317;
	wire [13-1:0] node318;
	wire [13-1:0] node319;
	wire [13-1:0] node322;
	wire [13-1:0] node325;
	wire [13-1:0] node326;
	wire [13-1:0] node329;
	wire [13-1:0] node332;
	wire [13-1:0] node333;
	wire [13-1:0] node334;
	wire [13-1:0] node335;
	wire [13-1:0] node338;
	wire [13-1:0] node342;
	wire [13-1:0] node343;
	wire [13-1:0] node345;
	wire [13-1:0] node348;
	wire [13-1:0] node349;
	wire [13-1:0] node352;
	wire [13-1:0] node355;
	wire [13-1:0] node356;
	wire [13-1:0] node357;
	wire [13-1:0] node358;
	wire [13-1:0] node359;
	wire [13-1:0] node362;
	wire [13-1:0] node365;
	wire [13-1:0] node366;
	wire [13-1:0] node370;
	wire [13-1:0] node372;
	wire [13-1:0] node373;
	wire [13-1:0] node377;
	wire [13-1:0] node378;
	wire [13-1:0] node379;
	wire [13-1:0] node380;
	wire [13-1:0] node383;
	wire [13-1:0] node386;
	wire [13-1:0] node387;
	wire [13-1:0] node390;
	wire [13-1:0] node393;
	wire [13-1:0] node394;
	wire [13-1:0] node395;
	wire [13-1:0] node399;
	wire [13-1:0] node400;
	wire [13-1:0] node403;
	wire [13-1:0] node406;
	wire [13-1:0] node407;
	wire [13-1:0] node408;
	wire [13-1:0] node409;
	wire [13-1:0] node410;
	wire [13-1:0] node411;
	wire [13-1:0] node412;
	wire [13-1:0] node414;
	wire [13-1:0] node417;
	wire [13-1:0] node418;
	wire [13-1:0] node421;
	wire [13-1:0] node424;
	wire [13-1:0] node425;
	wire [13-1:0] node426;
	wire [13-1:0] node429;
	wire [13-1:0] node432;
	wire [13-1:0] node433;
	wire [13-1:0] node437;
	wire [13-1:0] node438;
	wire [13-1:0] node439;
	wire [13-1:0] node440;
	wire [13-1:0] node444;
	wire [13-1:0] node446;
	wire [13-1:0] node449;
	wire [13-1:0] node451;
	wire [13-1:0] node452;
	wire [13-1:0] node455;
	wire [13-1:0] node458;
	wire [13-1:0] node459;
	wire [13-1:0] node460;
	wire [13-1:0] node461;
	wire [13-1:0] node462;
	wire [13-1:0] node465;
	wire [13-1:0] node468;
	wire [13-1:0] node469;
	wire [13-1:0] node472;
	wire [13-1:0] node475;
	wire [13-1:0] node476;
	wire [13-1:0] node477;
	wire [13-1:0] node480;
	wire [13-1:0] node483;
	wire [13-1:0] node484;
	wire [13-1:0] node487;
	wire [13-1:0] node490;
	wire [13-1:0] node491;
	wire [13-1:0] node492;
	wire [13-1:0] node493;
	wire [13-1:0] node496;
	wire [13-1:0] node500;
	wire [13-1:0] node501;
	wire [13-1:0] node502;
	wire [13-1:0] node505;
	wire [13-1:0] node509;
	wire [13-1:0] node510;
	wire [13-1:0] node511;
	wire [13-1:0] node512;
	wire [13-1:0] node513;
	wire [13-1:0] node515;
	wire [13-1:0] node519;
	wire [13-1:0] node520;
	wire [13-1:0] node521;
	wire [13-1:0] node524;
	wire [13-1:0] node527;
	wire [13-1:0] node528;
	wire [13-1:0] node532;
	wire [13-1:0] node533;
	wire [13-1:0] node534;
	wire [13-1:0] node535;
	wire [13-1:0] node538;
	wire [13-1:0] node541;
	wire [13-1:0] node542;
	wire [13-1:0] node545;
	wire [13-1:0] node548;
	wire [13-1:0] node549;
	wire [13-1:0] node550;
	wire [13-1:0] node554;
	wire [13-1:0] node555;
	wire [13-1:0] node559;
	wire [13-1:0] node560;
	wire [13-1:0] node561;
	wire [13-1:0] node562;
	wire [13-1:0] node563;
	wire [13-1:0] node566;
	wire [13-1:0] node569;
	wire [13-1:0] node570;
	wire [13-1:0] node574;
	wire [13-1:0] node575;
	wire [13-1:0] node577;
	wire [13-1:0] node580;
	wire [13-1:0] node581;
	wire [13-1:0] node585;
	wire [13-1:0] node586;
	wire [13-1:0] node587;
	wire [13-1:0] node588;
	wire [13-1:0] node592;
	wire [13-1:0] node593;
	wire [13-1:0] node596;
	wire [13-1:0] node599;
	wire [13-1:0] node600;
	wire [13-1:0] node601;
	wire [13-1:0] node604;
	wire [13-1:0] node607;
	wire [13-1:0] node608;
	wire [13-1:0] node612;
	wire [13-1:0] node613;
	wire [13-1:0] node614;
	wire [13-1:0] node615;
	wire [13-1:0] node616;
	wire [13-1:0] node617;
	wire [13-1:0] node621;
	wire [13-1:0] node622;
	wire [13-1:0] node623;
	wire [13-1:0] node626;
	wire [13-1:0] node629;
	wire [13-1:0] node630;
	wire [13-1:0] node634;
	wire [13-1:0] node635;
	wire [13-1:0] node636;
	wire [13-1:0] node637;
	wire [13-1:0] node640;
	wire [13-1:0] node643;
	wire [13-1:0] node645;
	wire [13-1:0] node648;
	wire [13-1:0] node650;
	wire [13-1:0] node651;
	wire [13-1:0] node654;
	wire [13-1:0] node657;
	wire [13-1:0] node658;
	wire [13-1:0] node659;
	wire [13-1:0] node660;
	wire [13-1:0] node661;
	wire [13-1:0] node664;
	wire [13-1:0] node667;
	wire [13-1:0] node668;
	wire [13-1:0] node671;
	wire [13-1:0] node674;
	wire [13-1:0] node675;
	wire [13-1:0] node676;
	wire [13-1:0] node679;
	wire [13-1:0] node682;
	wire [13-1:0] node683;
	wire [13-1:0] node686;
	wire [13-1:0] node689;
	wire [13-1:0] node690;
	wire [13-1:0] node691;
	wire [13-1:0] node692;
	wire [13-1:0] node695;
	wire [13-1:0] node698;
	wire [13-1:0] node700;
	wire [13-1:0] node703;
	wire [13-1:0] node704;
	wire [13-1:0] node705;
	wire [13-1:0] node708;
	wire [13-1:0] node711;
	wire [13-1:0] node714;
	wire [13-1:0] node715;
	wire [13-1:0] node716;
	wire [13-1:0] node717;
	wire [13-1:0] node718;
	wire [13-1:0] node719;
	wire [13-1:0] node722;
	wire [13-1:0] node726;
	wire [13-1:0] node727;
	wire [13-1:0] node728;
	wire [13-1:0] node732;
	wire [13-1:0] node734;
	wire [13-1:0] node737;
	wire [13-1:0] node738;
	wire [13-1:0] node739;
	wire [13-1:0] node741;
	wire [13-1:0] node744;
	wire [13-1:0] node745;
	wire [13-1:0] node748;
	wire [13-1:0] node751;
	wire [13-1:0] node752;
	wire [13-1:0] node755;
	wire [13-1:0] node758;
	wire [13-1:0] node759;
	wire [13-1:0] node760;
	wire [13-1:0] node761;
	wire [13-1:0] node762;
	wire [13-1:0] node765;
	wire [13-1:0] node769;
	wire [13-1:0] node770;
	wire [13-1:0] node771;
	wire [13-1:0] node774;
	wire [13-1:0] node777;
	wire [13-1:0] node779;
	wire [13-1:0] node782;
	wire [13-1:0] node783;
	wire [13-1:0] node784;
	wire [13-1:0] node785;
	wire [13-1:0] node788;
	wire [13-1:0] node791;
	wire [13-1:0] node793;
	wire [13-1:0] node796;
	wire [13-1:0] node797;
	wire [13-1:0] node798;
	wire [13-1:0] node801;
	wire [13-1:0] node804;
	wire [13-1:0] node806;
	wire [13-1:0] node809;
	wire [13-1:0] node810;
	wire [13-1:0] node811;
	wire [13-1:0] node812;
	wire [13-1:0] node813;
	wire [13-1:0] node814;
	wire [13-1:0] node815;
	wire [13-1:0] node816;
	wire [13-1:0] node818;
	wire [13-1:0] node821;
	wire [13-1:0] node822;
	wire [13-1:0] node826;
	wire [13-1:0] node827;
	wire [13-1:0] node828;
	wire [13-1:0] node831;
	wire [13-1:0] node834;
	wire [13-1:0] node835;
	wire [13-1:0] node838;
	wire [13-1:0] node841;
	wire [13-1:0] node842;
	wire [13-1:0] node844;
	wire [13-1:0] node845;
	wire [13-1:0] node848;
	wire [13-1:0] node851;
	wire [13-1:0] node852;
	wire [13-1:0] node853;
	wire [13-1:0] node856;
	wire [13-1:0] node859;
	wire [13-1:0] node861;
	wire [13-1:0] node864;
	wire [13-1:0] node865;
	wire [13-1:0] node866;
	wire [13-1:0] node867;
	wire [13-1:0] node868;
	wire [13-1:0] node871;
	wire [13-1:0] node874;
	wire [13-1:0] node875;
	wire [13-1:0] node879;
	wire [13-1:0] node880;
	wire [13-1:0] node881;
	wire [13-1:0] node884;
	wire [13-1:0] node887;
	wire [13-1:0] node889;
	wire [13-1:0] node892;
	wire [13-1:0] node893;
	wire [13-1:0] node894;
	wire [13-1:0] node895;
	wire [13-1:0] node898;
	wire [13-1:0] node901;
	wire [13-1:0] node902;
	wire [13-1:0] node906;
	wire [13-1:0] node908;
	wire [13-1:0] node909;
	wire [13-1:0] node913;
	wire [13-1:0] node914;
	wire [13-1:0] node915;
	wire [13-1:0] node916;
	wire [13-1:0] node917;
	wire [13-1:0] node918;
	wire [13-1:0] node921;
	wire [13-1:0] node924;
	wire [13-1:0] node926;
	wire [13-1:0] node929;
	wire [13-1:0] node930;
	wire [13-1:0] node932;
	wire [13-1:0] node935;
	wire [13-1:0] node936;
	wire [13-1:0] node939;
	wire [13-1:0] node942;
	wire [13-1:0] node943;
	wire [13-1:0] node944;
	wire [13-1:0] node945;
	wire [13-1:0] node948;
	wire [13-1:0] node951;
	wire [13-1:0] node952;
	wire [13-1:0] node955;
	wire [13-1:0] node958;
	wire [13-1:0] node959;
	wire [13-1:0] node961;
	wire [13-1:0] node965;
	wire [13-1:0] node966;
	wire [13-1:0] node967;
	wire [13-1:0] node968;
	wire [13-1:0] node970;
	wire [13-1:0] node973;
	wire [13-1:0] node974;
	wire [13-1:0] node977;
	wire [13-1:0] node980;
	wire [13-1:0] node981;
	wire [13-1:0] node983;
	wire [13-1:0] node986;
	wire [13-1:0] node987;
	wire [13-1:0] node991;
	wire [13-1:0] node992;
	wire [13-1:0] node993;
	wire [13-1:0] node996;
	wire [13-1:0] node997;
	wire [13-1:0] node1001;
	wire [13-1:0] node1002;
	wire [13-1:0] node1003;
	wire [13-1:0] node1007;
	wire [13-1:0] node1008;
	wire [13-1:0] node1011;
	wire [13-1:0] node1014;
	wire [13-1:0] node1015;
	wire [13-1:0] node1016;
	wire [13-1:0] node1017;
	wire [13-1:0] node1018;
	wire [13-1:0] node1019;
	wire [13-1:0] node1020;
	wire [13-1:0] node1024;
	wire [13-1:0] node1025;
	wire [13-1:0] node1028;
	wire [13-1:0] node1031;
	wire [13-1:0] node1032;
	wire [13-1:0] node1033;
	wire [13-1:0] node1036;
	wire [13-1:0] node1039;
	wire [13-1:0] node1040;
	wire [13-1:0] node1044;
	wire [13-1:0] node1045;
	wire [13-1:0] node1046;
	wire [13-1:0] node1047;
	wire [13-1:0] node1050;
	wire [13-1:0] node1053;
	wire [13-1:0] node1054;
	wire [13-1:0] node1057;
	wire [13-1:0] node1060;
	wire [13-1:0] node1061;
	wire [13-1:0] node1062;
	wire [13-1:0] node1065;
	wire [13-1:0] node1068;
	wire [13-1:0] node1069;
	wire [13-1:0] node1073;
	wire [13-1:0] node1074;
	wire [13-1:0] node1075;
	wire [13-1:0] node1076;
	wire [13-1:0] node1078;
	wire [13-1:0] node1081;
	wire [13-1:0] node1082;
	wire [13-1:0] node1085;
	wire [13-1:0] node1088;
	wire [13-1:0] node1089;
	wire [13-1:0] node1091;
	wire [13-1:0] node1094;
	wire [13-1:0] node1095;
	wire [13-1:0] node1099;
	wire [13-1:0] node1100;
	wire [13-1:0] node1101;
	wire [13-1:0] node1102;
	wire [13-1:0] node1106;
	wire [13-1:0] node1108;
	wire [13-1:0] node1111;
	wire [13-1:0] node1112;
	wire [13-1:0] node1114;
	wire [13-1:0] node1117;
	wire [13-1:0] node1118;
	wire [13-1:0] node1121;
	wire [13-1:0] node1124;
	wire [13-1:0] node1125;
	wire [13-1:0] node1126;
	wire [13-1:0] node1127;
	wire [13-1:0] node1129;
	wire [13-1:0] node1130;
	wire [13-1:0] node1134;
	wire [13-1:0] node1135;
	wire [13-1:0] node1137;
	wire [13-1:0] node1140;
	wire [13-1:0] node1143;
	wire [13-1:0] node1144;
	wire [13-1:0] node1146;
	wire [13-1:0] node1147;
	wire [13-1:0] node1150;
	wire [13-1:0] node1153;
	wire [13-1:0] node1154;
	wire [13-1:0] node1155;
	wire [13-1:0] node1159;
	wire [13-1:0] node1160;
	wire [13-1:0] node1163;
	wire [13-1:0] node1166;
	wire [13-1:0] node1167;
	wire [13-1:0] node1168;
	wire [13-1:0] node1169;
	wire [13-1:0] node1170;
	wire [13-1:0] node1173;
	wire [13-1:0] node1176;
	wire [13-1:0] node1177;
	wire [13-1:0] node1181;
	wire [13-1:0] node1182;
	wire [13-1:0] node1184;
	wire [13-1:0] node1187;
	wire [13-1:0] node1188;
	wire [13-1:0] node1191;
	wire [13-1:0] node1194;
	wire [13-1:0] node1195;
	wire [13-1:0] node1196;
	wire [13-1:0] node1198;
	wire [13-1:0] node1201;
	wire [13-1:0] node1202;
	wire [13-1:0] node1205;
	wire [13-1:0] node1208;
	wire [13-1:0] node1209;
	wire [13-1:0] node1211;
	wire [13-1:0] node1214;
	wire [13-1:0] node1216;
	wire [13-1:0] node1219;
	wire [13-1:0] node1220;
	wire [13-1:0] node1221;
	wire [13-1:0] node1222;
	wire [13-1:0] node1223;
	wire [13-1:0] node1224;
	wire [13-1:0] node1225;
	wire [13-1:0] node1227;
	wire [13-1:0] node1230;
	wire [13-1:0] node1231;
	wire [13-1:0] node1234;
	wire [13-1:0] node1237;
	wire [13-1:0] node1238;
	wire [13-1:0] node1239;
	wire [13-1:0] node1243;
	wire [13-1:0] node1246;
	wire [13-1:0] node1247;
	wire [13-1:0] node1248;
	wire [13-1:0] node1249;
	wire [13-1:0] node1252;
	wire [13-1:0] node1255;
	wire [13-1:0] node1256;
	wire [13-1:0] node1259;
	wire [13-1:0] node1262;
	wire [13-1:0] node1263;
	wire [13-1:0] node1264;
	wire [13-1:0] node1268;
	wire [13-1:0] node1270;
	wire [13-1:0] node1273;
	wire [13-1:0] node1274;
	wire [13-1:0] node1275;
	wire [13-1:0] node1276;
	wire [13-1:0] node1277;
	wire [13-1:0] node1281;
	wire [13-1:0] node1282;
	wire [13-1:0] node1286;
	wire [13-1:0] node1287;
	wire [13-1:0] node1288;
	wire [13-1:0] node1292;
	wire [13-1:0] node1293;
	wire [13-1:0] node1296;
	wire [13-1:0] node1299;
	wire [13-1:0] node1300;
	wire [13-1:0] node1301;
	wire [13-1:0] node1302;
	wire [13-1:0] node1306;
	wire [13-1:0] node1307;
	wire [13-1:0] node1311;
	wire [13-1:0] node1312;
	wire [13-1:0] node1313;
	wire [13-1:0] node1316;
	wire [13-1:0] node1319;
	wire [13-1:0] node1320;
	wire [13-1:0] node1323;
	wire [13-1:0] node1326;
	wire [13-1:0] node1327;
	wire [13-1:0] node1328;
	wire [13-1:0] node1329;
	wire [13-1:0] node1330;
	wire [13-1:0] node1332;
	wire [13-1:0] node1335;
	wire [13-1:0] node1336;
	wire [13-1:0] node1339;
	wire [13-1:0] node1342;
	wire [13-1:0] node1343;
	wire [13-1:0] node1344;
	wire [13-1:0] node1347;
	wire [13-1:0] node1350;
	wire [13-1:0] node1351;
	wire [13-1:0] node1354;
	wire [13-1:0] node1357;
	wire [13-1:0] node1358;
	wire [13-1:0] node1359;
	wire [13-1:0] node1360;
	wire [13-1:0] node1363;
	wire [13-1:0] node1366;
	wire [13-1:0] node1367;
	wire [13-1:0] node1370;
	wire [13-1:0] node1373;
	wire [13-1:0] node1374;
	wire [13-1:0] node1377;
	wire [13-1:0] node1379;
	wire [13-1:0] node1382;
	wire [13-1:0] node1383;
	wire [13-1:0] node1384;
	wire [13-1:0] node1385;
	wire [13-1:0] node1387;
	wire [13-1:0] node1390;
	wire [13-1:0] node1392;
	wire [13-1:0] node1395;
	wire [13-1:0] node1396;
	wire [13-1:0] node1397;
	wire [13-1:0] node1400;
	wire [13-1:0] node1403;
	wire [13-1:0] node1405;
	wire [13-1:0] node1408;
	wire [13-1:0] node1409;
	wire [13-1:0] node1410;
	wire [13-1:0] node1412;
	wire [13-1:0] node1415;
	wire [13-1:0] node1417;
	wire [13-1:0] node1420;
	wire [13-1:0] node1421;
	wire [13-1:0] node1422;
	wire [13-1:0] node1425;
	wire [13-1:0] node1428;
	wire [13-1:0] node1429;
	wire [13-1:0] node1432;
	wire [13-1:0] node1435;
	wire [13-1:0] node1436;
	wire [13-1:0] node1437;
	wire [13-1:0] node1438;
	wire [13-1:0] node1439;
	wire [13-1:0] node1440;
	wire [13-1:0] node1443;
	wire [13-1:0] node1444;
	wire [13-1:0] node1447;
	wire [13-1:0] node1450;
	wire [13-1:0] node1451;
	wire [13-1:0] node1452;
	wire [13-1:0] node1455;
	wire [13-1:0] node1458;
	wire [13-1:0] node1459;
	wire [13-1:0] node1462;
	wire [13-1:0] node1465;
	wire [13-1:0] node1466;
	wire [13-1:0] node1467;
	wire [13-1:0] node1468;
	wire [13-1:0] node1472;
	wire [13-1:0] node1473;
	wire [13-1:0] node1476;
	wire [13-1:0] node1479;
	wire [13-1:0] node1480;
	wire [13-1:0] node1482;
	wire [13-1:0] node1485;
	wire [13-1:0] node1486;
	wire [13-1:0] node1489;
	wire [13-1:0] node1492;
	wire [13-1:0] node1493;
	wire [13-1:0] node1494;
	wire [13-1:0] node1495;
	wire [13-1:0] node1497;
	wire [13-1:0] node1500;
	wire [13-1:0] node1502;
	wire [13-1:0] node1505;
	wire [13-1:0] node1506;
	wire [13-1:0] node1507;
	wire [13-1:0] node1510;
	wire [13-1:0] node1513;
	wire [13-1:0] node1514;
	wire [13-1:0] node1518;
	wire [13-1:0] node1519;
	wire [13-1:0] node1520;
	wire [13-1:0] node1522;
	wire [13-1:0] node1525;
	wire [13-1:0] node1526;
	wire [13-1:0] node1529;
	wire [13-1:0] node1532;
	wire [13-1:0] node1533;
	wire [13-1:0] node1534;
	wire [13-1:0] node1537;
	wire [13-1:0] node1540;
	wire [13-1:0] node1542;
	wire [13-1:0] node1545;
	wire [13-1:0] node1546;
	wire [13-1:0] node1547;
	wire [13-1:0] node1548;
	wire [13-1:0] node1549;
	wire [13-1:0] node1550;
	wire [13-1:0] node1554;
	wire [13-1:0] node1555;
	wire [13-1:0] node1559;
	wire [13-1:0] node1560;
	wire [13-1:0] node1562;
	wire [13-1:0] node1565;
	wire [13-1:0] node1566;
	wire [13-1:0] node1569;
	wire [13-1:0] node1572;
	wire [13-1:0] node1573;
	wire [13-1:0] node1575;
	wire [13-1:0] node1576;
	wire [13-1:0] node1579;
	wire [13-1:0] node1582;
	wire [13-1:0] node1583;
	wire [13-1:0] node1584;
	wire [13-1:0] node1587;
	wire [13-1:0] node1590;
	wire [13-1:0] node1591;
	wire [13-1:0] node1595;
	wire [13-1:0] node1596;
	wire [13-1:0] node1597;
	wire [13-1:0] node1598;
	wire [13-1:0] node1600;
	wire [13-1:0] node1603;
	wire [13-1:0] node1604;
	wire [13-1:0] node1607;
	wire [13-1:0] node1610;
	wire [13-1:0] node1611;
	wire [13-1:0] node1612;
	wire [13-1:0] node1615;
	wire [13-1:0] node1618;
	wire [13-1:0] node1619;
	wire [13-1:0] node1622;
	wire [13-1:0] node1625;
	wire [13-1:0] node1626;
	wire [13-1:0] node1627;
	wire [13-1:0] node1628;
	wire [13-1:0] node1631;
	wire [13-1:0] node1634;
	wire [13-1:0] node1635;
	wire [13-1:0] node1639;
	wire [13-1:0] node1640;
	wire [13-1:0] node1641;
	wire [13-1:0] node1645;
	wire [13-1:0] node1646;
	wire [13-1:0] node1649;
	wire [13-1:0] node1652;
	wire [13-1:0] node1653;
	wire [13-1:0] node1654;
	wire [13-1:0] node1655;
	wire [13-1:0] node1656;
	wire [13-1:0] node1657;
	wire [13-1:0] node1658;
	wire [13-1:0] node1659;
	wire [13-1:0] node1660;
	wire [13-1:0] node1662;
	wire [13-1:0] node1666;
	wire [13-1:0] node1668;
	wire [13-1:0] node1670;
	wire [13-1:0] node1673;
	wire [13-1:0] node1674;
	wire [13-1:0] node1675;
	wire [13-1:0] node1678;
	wire [13-1:0] node1679;
	wire [13-1:0] node1683;
	wire [13-1:0] node1684;
	wire [13-1:0] node1685;
	wire [13-1:0] node1688;
	wire [13-1:0] node1691;
	wire [13-1:0] node1694;
	wire [13-1:0] node1695;
	wire [13-1:0] node1696;
	wire [13-1:0] node1697;
	wire [13-1:0] node1699;
	wire [13-1:0] node1702;
	wire [13-1:0] node1703;
	wire [13-1:0] node1706;
	wire [13-1:0] node1709;
	wire [13-1:0] node1710;
	wire [13-1:0] node1711;
	wire [13-1:0] node1715;
	wire [13-1:0] node1716;
	wire [13-1:0] node1720;
	wire [13-1:0] node1721;
	wire [13-1:0] node1722;
	wire [13-1:0] node1723;
	wire [13-1:0] node1727;
	wire [13-1:0] node1728;
	wire [13-1:0] node1731;
	wire [13-1:0] node1734;
	wire [13-1:0] node1735;
	wire [13-1:0] node1737;
	wire [13-1:0] node1741;
	wire [13-1:0] node1742;
	wire [13-1:0] node1743;
	wire [13-1:0] node1744;
	wire [13-1:0] node1745;
	wire [13-1:0] node1746;
	wire [13-1:0] node1749;
	wire [13-1:0] node1752;
	wire [13-1:0] node1755;
	wire [13-1:0] node1756;
	wire [13-1:0] node1758;
	wire [13-1:0] node1761;
	wire [13-1:0] node1762;
	wire [13-1:0] node1766;
	wire [13-1:0] node1767;
	wire [13-1:0] node1768;
	wire [13-1:0] node1771;
	wire [13-1:0] node1774;
	wire [13-1:0] node1776;
	wire [13-1:0] node1777;
	wire [13-1:0] node1781;
	wire [13-1:0] node1782;
	wire [13-1:0] node1783;
	wire [13-1:0] node1784;
	wire [13-1:0] node1785;
	wire [13-1:0] node1789;
	wire [13-1:0] node1790;
	wire [13-1:0] node1793;
	wire [13-1:0] node1796;
	wire [13-1:0] node1797;
	wire [13-1:0] node1798;
	wire [13-1:0] node1801;
	wire [13-1:0] node1804;
	wire [13-1:0] node1807;
	wire [13-1:0] node1808;
	wire [13-1:0] node1809;
	wire [13-1:0] node1812;
	wire [13-1:0] node1814;
	wire [13-1:0] node1817;
	wire [13-1:0] node1818;
	wire [13-1:0] node1820;
	wire [13-1:0] node1824;
	wire [13-1:0] node1825;
	wire [13-1:0] node1826;
	wire [13-1:0] node1827;
	wire [13-1:0] node1828;
	wire [13-1:0] node1829;
	wire [13-1:0] node1830;
	wire [13-1:0] node1833;
	wire [13-1:0] node1836;
	wire [13-1:0] node1839;
	wire [13-1:0] node1840;
	wire [13-1:0] node1841;
	wire [13-1:0] node1844;
	wire [13-1:0] node1847;
	wire [13-1:0] node1848;
	wire [13-1:0] node1851;
	wire [13-1:0] node1854;
	wire [13-1:0] node1855;
	wire [13-1:0] node1856;
	wire [13-1:0] node1857;
	wire [13-1:0] node1860;
	wire [13-1:0] node1863;
	wire [13-1:0] node1864;
	wire [13-1:0] node1867;
	wire [13-1:0] node1870;
	wire [13-1:0] node1871;
	wire [13-1:0] node1872;
	wire [13-1:0] node1875;
	wire [13-1:0] node1878;
	wire [13-1:0] node1879;
	wire [13-1:0] node1882;
	wire [13-1:0] node1885;
	wire [13-1:0] node1886;
	wire [13-1:0] node1887;
	wire [13-1:0] node1888;
	wire [13-1:0] node1890;
	wire [13-1:0] node1894;
	wire [13-1:0] node1895;
	wire [13-1:0] node1896;
	wire [13-1:0] node1899;
	wire [13-1:0] node1902;
	wire [13-1:0] node1905;
	wire [13-1:0] node1906;
	wire [13-1:0] node1907;
	wire [13-1:0] node1908;
	wire [13-1:0] node1912;
	wire [13-1:0] node1914;
	wire [13-1:0] node1917;
	wire [13-1:0] node1918;
	wire [13-1:0] node1919;
	wire [13-1:0] node1922;
	wire [13-1:0] node1925;
	wire [13-1:0] node1926;
	wire [13-1:0] node1929;
	wire [13-1:0] node1932;
	wire [13-1:0] node1933;
	wire [13-1:0] node1934;
	wire [13-1:0] node1935;
	wire [13-1:0] node1936;
	wire [13-1:0] node1937;
	wire [13-1:0] node1941;
	wire [13-1:0] node1942;
	wire [13-1:0] node1945;
	wire [13-1:0] node1948;
	wire [13-1:0] node1949;
	wire [13-1:0] node1951;
	wire [13-1:0] node1954;
	wire [13-1:0] node1956;
	wire [13-1:0] node1959;
	wire [13-1:0] node1960;
	wire [13-1:0] node1961;
	wire [13-1:0] node1963;
	wire [13-1:0] node1966;
	wire [13-1:0] node1967;
	wire [13-1:0] node1971;
	wire [13-1:0] node1972;
	wire [13-1:0] node1973;
	wire [13-1:0] node1976;
	wire [13-1:0] node1979;
	wire [13-1:0] node1980;
	wire [13-1:0] node1983;
	wire [13-1:0] node1986;
	wire [13-1:0] node1987;
	wire [13-1:0] node1988;
	wire [13-1:0] node1989;
	wire [13-1:0] node1992;
	wire [13-1:0] node1993;
	wire [13-1:0] node1996;
	wire [13-1:0] node1999;
	wire [13-1:0] node2000;
	wire [13-1:0] node2003;
	wire [13-1:0] node2004;
	wire [13-1:0] node2008;
	wire [13-1:0] node2009;
	wire [13-1:0] node2010;
	wire [13-1:0] node2012;
	wire [13-1:0] node2015;
	wire [13-1:0] node2017;
	wire [13-1:0] node2020;
	wire [13-1:0] node2021;
	wire [13-1:0] node2024;
	wire [13-1:0] node2026;
	wire [13-1:0] node2029;
	wire [13-1:0] node2030;
	wire [13-1:0] node2031;
	wire [13-1:0] node2032;
	wire [13-1:0] node2033;
	wire [13-1:0] node2034;
	wire [13-1:0] node2035;
	wire [13-1:0] node2036;
	wire [13-1:0] node2039;
	wire [13-1:0] node2042;
	wire [13-1:0] node2044;
	wire [13-1:0] node2047;
	wire [13-1:0] node2048;
	wire [13-1:0] node2049;
	wire [13-1:0] node2052;
	wire [13-1:0] node2055;
	wire [13-1:0] node2057;
	wire [13-1:0] node2060;
	wire [13-1:0] node2061;
	wire [13-1:0] node2062;
	wire [13-1:0] node2065;
	wire [13-1:0] node2066;
	wire [13-1:0] node2070;
	wire [13-1:0] node2071;
	wire [13-1:0] node2072;
	wire [13-1:0] node2075;
	wire [13-1:0] node2078;
	wire [13-1:0] node2079;
	wire [13-1:0] node2082;
	wire [13-1:0] node2085;
	wire [13-1:0] node2086;
	wire [13-1:0] node2087;
	wire [13-1:0] node2088;
	wire [13-1:0] node2089;
	wire [13-1:0] node2092;
	wire [13-1:0] node2095;
	wire [13-1:0] node2098;
	wire [13-1:0] node2099;
	wire [13-1:0] node2100;
	wire [13-1:0] node2103;
	wire [13-1:0] node2107;
	wire [13-1:0] node2108;
	wire [13-1:0] node2109;
	wire [13-1:0] node2111;
	wire [13-1:0] node2114;
	wire [13-1:0] node2115;
	wire [13-1:0] node2119;
	wire [13-1:0] node2120;
	wire [13-1:0] node2123;
	wire [13-1:0] node2124;
	wire [13-1:0] node2127;
	wire [13-1:0] node2130;
	wire [13-1:0] node2131;
	wire [13-1:0] node2132;
	wire [13-1:0] node2133;
	wire [13-1:0] node2134;
	wire [13-1:0] node2136;
	wire [13-1:0] node2139;
	wire [13-1:0] node2140;
	wire [13-1:0] node2143;
	wire [13-1:0] node2146;
	wire [13-1:0] node2147;
	wire [13-1:0] node2148;
	wire [13-1:0] node2151;
	wire [13-1:0] node2154;
	wire [13-1:0] node2155;
	wire [13-1:0] node2159;
	wire [13-1:0] node2160;
	wire [13-1:0] node2161;
	wire [13-1:0] node2164;
	wire [13-1:0] node2165;
	wire [13-1:0] node2168;
	wire [13-1:0] node2171;
	wire [13-1:0] node2172;
	wire [13-1:0] node2174;
	wire [13-1:0] node2177;
	wire [13-1:0] node2179;
	wire [13-1:0] node2182;
	wire [13-1:0] node2183;
	wire [13-1:0] node2184;
	wire [13-1:0] node2185;
	wire [13-1:0] node2186;
	wire [13-1:0] node2189;
	wire [13-1:0] node2192;
	wire [13-1:0] node2195;
	wire [13-1:0] node2196;
	wire [13-1:0] node2198;
	wire [13-1:0] node2201;
	wire [13-1:0] node2202;
	wire [13-1:0] node2205;
	wire [13-1:0] node2208;
	wire [13-1:0] node2209;
	wire [13-1:0] node2210;
	wire [13-1:0] node2211;
	wire [13-1:0] node2214;
	wire [13-1:0] node2217;
	wire [13-1:0] node2218;
	wire [13-1:0] node2221;
	wire [13-1:0] node2224;
	wire [13-1:0] node2225;
	wire [13-1:0] node2227;
	wire [13-1:0] node2230;
	wire [13-1:0] node2232;
	wire [13-1:0] node2235;
	wire [13-1:0] node2236;
	wire [13-1:0] node2237;
	wire [13-1:0] node2238;
	wire [13-1:0] node2239;
	wire [13-1:0] node2240;
	wire [13-1:0] node2241;
	wire [13-1:0] node2244;
	wire [13-1:0] node2247;
	wire [13-1:0] node2249;
	wire [13-1:0] node2252;
	wire [13-1:0] node2253;
	wire [13-1:0] node2254;
	wire [13-1:0] node2257;
	wire [13-1:0] node2260;
	wire [13-1:0] node2261;
	wire [13-1:0] node2264;
	wire [13-1:0] node2267;
	wire [13-1:0] node2268;
	wire [13-1:0] node2269;
	wire [13-1:0] node2271;
	wire [13-1:0] node2274;
	wire [13-1:0] node2275;
	wire [13-1:0] node2278;
	wire [13-1:0] node2281;
	wire [13-1:0] node2282;
	wire [13-1:0] node2284;
	wire [13-1:0] node2287;
	wire [13-1:0] node2289;
	wire [13-1:0] node2292;
	wire [13-1:0] node2293;
	wire [13-1:0] node2294;
	wire [13-1:0] node2295;
	wire [13-1:0] node2297;
	wire [13-1:0] node2300;
	wire [13-1:0] node2302;
	wire [13-1:0] node2305;
	wire [13-1:0] node2306;
	wire [13-1:0] node2307;
	wire [13-1:0] node2310;
	wire [13-1:0] node2313;
	wire [13-1:0] node2314;
	wire [13-1:0] node2318;
	wire [13-1:0] node2319;
	wire [13-1:0] node2320;
	wire [13-1:0] node2321;
	wire [13-1:0] node2324;
	wire [13-1:0] node2327;
	wire [13-1:0] node2328;
	wire [13-1:0] node2331;
	wire [13-1:0] node2334;
	wire [13-1:0] node2335;
	wire [13-1:0] node2337;
	wire [13-1:0] node2340;
	wire [13-1:0] node2343;
	wire [13-1:0] node2344;
	wire [13-1:0] node2345;
	wire [13-1:0] node2346;
	wire [13-1:0] node2347;
	wire [13-1:0] node2348;
	wire [13-1:0] node2352;
	wire [13-1:0] node2355;
	wire [13-1:0] node2356;
	wire [13-1:0] node2357;
	wire [13-1:0] node2360;
	wire [13-1:0] node2363;
	wire [13-1:0] node2365;
	wire [13-1:0] node2368;
	wire [13-1:0] node2369;
	wire [13-1:0] node2370;
	wire [13-1:0] node2372;
	wire [13-1:0] node2375;
	wire [13-1:0] node2377;
	wire [13-1:0] node2380;
	wire [13-1:0] node2381;
	wire [13-1:0] node2382;
	wire [13-1:0] node2385;
	wire [13-1:0] node2388;
	wire [13-1:0] node2391;
	wire [13-1:0] node2392;
	wire [13-1:0] node2393;
	wire [13-1:0] node2394;
	wire [13-1:0] node2395;
	wire [13-1:0] node2398;
	wire [13-1:0] node2401;
	wire [13-1:0] node2402;
	wire [13-1:0] node2405;
	wire [13-1:0] node2408;
	wire [13-1:0] node2409;
	wire [13-1:0] node2411;
	wire [13-1:0] node2414;
	wire [13-1:0] node2415;
	wire [13-1:0] node2419;
	wire [13-1:0] node2420;
	wire [13-1:0] node2421;
	wire [13-1:0] node2422;
	wire [13-1:0] node2425;
	wire [13-1:0] node2428;
	wire [13-1:0] node2429;
	wire [13-1:0] node2432;
	wire [13-1:0] node2435;
	wire [13-1:0] node2436;
	wire [13-1:0] node2437;
	wire [13-1:0] node2441;
	wire [13-1:0] node2442;
	wire [13-1:0] node2445;
	wire [13-1:0] node2448;
	wire [13-1:0] node2449;
	wire [13-1:0] node2450;
	wire [13-1:0] node2451;
	wire [13-1:0] node2452;
	wire [13-1:0] node2453;
	wire [13-1:0] node2454;
	wire [13-1:0] node2455;
	wire [13-1:0] node2456;
	wire [13-1:0] node2459;
	wire [13-1:0] node2462;
	wire [13-1:0] node2465;
	wire [13-1:0] node2466;
	wire [13-1:0] node2468;
	wire [13-1:0] node2471;
	wire [13-1:0] node2472;
	wire [13-1:0] node2476;
	wire [13-1:0] node2477;
	wire [13-1:0] node2479;
	wire [13-1:0] node2480;
	wire [13-1:0] node2484;
	wire [13-1:0] node2486;
	wire [13-1:0] node2487;
	wire [13-1:0] node2490;
	wire [13-1:0] node2493;
	wire [13-1:0] node2494;
	wire [13-1:0] node2495;
	wire [13-1:0] node2496;
	wire [13-1:0] node2497;
	wire [13-1:0] node2501;
	wire [13-1:0] node2502;
	wire [13-1:0] node2505;
	wire [13-1:0] node2508;
	wire [13-1:0] node2509;
	wire [13-1:0] node2510;
	wire [13-1:0] node2513;
	wire [13-1:0] node2516;
	wire [13-1:0] node2517;
	wire [13-1:0] node2520;
	wire [13-1:0] node2523;
	wire [13-1:0] node2524;
	wire [13-1:0] node2525;
	wire [13-1:0] node2526;
	wire [13-1:0] node2529;
	wire [13-1:0] node2532;
	wire [13-1:0] node2534;
	wire [13-1:0] node2537;
	wire [13-1:0] node2538;
	wire [13-1:0] node2540;
	wire [13-1:0] node2543;
	wire [13-1:0] node2545;
	wire [13-1:0] node2548;
	wire [13-1:0] node2549;
	wire [13-1:0] node2550;
	wire [13-1:0] node2551;
	wire [13-1:0] node2552;
	wire [13-1:0] node2554;
	wire [13-1:0] node2557;
	wire [13-1:0] node2558;
	wire [13-1:0] node2562;
	wire [13-1:0] node2563;
	wire [13-1:0] node2566;
	wire [13-1:0] node2568;
	wire [13-1:0] node2571;
	wire [13-1:0] node2572;
	wire [13-1:0] node2573;
	wire [13-1:0] node2575;
	wire [13-1:0] node2578;
	wire [13-1:0] node2579;
	wire [13-1:0] node2582;
	wire [13-1:0] node2585;
	wire [13-1:0] node2586;
	wire [13-1:0] node2587;
	wire [13-1:0] node2590;
	wire [13-1:0] node2593;
	wire [13-1:0] node2594;
	wire [13-1:0] node2597;
	wire [13-1:0] node2600;
	wire [13-1:0] node2601;
	wire [13-1:0] node2602;
	wire [13-1:0] node2604;
	wire [13-1:0] node2605;
	wire [13-1:0] node2608;
	wire [13-1:0] node2611;
	wire [13-1:0] node2612;
	wire [13-1:0] node2613;
	wire [13-1:0] node2616;
	wire [13-1:0] node2619;
	wire [13-1:0] node2621;
	wire [13-1:0] node2624;
	wire [13-1:0] node2625;
	wire [13-1:0] node2626;
	wire [13-1:0] node2628;
	wire [13-1:0] node2632;
	wire [13-1:0] node2633;
	wire [13-1:0] node2635;
	wire [13-1:0] node2638;
	wire [13-1:0] node2640;
	wire [13-1:0] node2643;
	wire [13-1:0] node2644;
	wire [13-1:0] node2645;
	wire [13-1:0] node2646;
	wire [13-1:0] node2647;
	wire [13-1:0] node2649;
	wire [13-1:0] node2650;
	wire [13-1:0] node2654;
	wire [13-1:0] node2655;
	wire [13-1:0] node2658;
	wire [13-1:0] node2659;
	wire [13-1:0] node2662;
	wire [13-1:0] node2665;
	wire [13-1:0] node2666;
	wire [13-1:0] node2667;
	wire [13-1:0] node2668;
	wire [13-1:0] node2671;
	wire [13-1:0] node2674;
	wire [13-1:0] node2677;
	wire [13-1:0] node2678;
	wire [13-1:0] node2680;
	wire [13-1:0] node2683;
	wire [13-1:0] node2685;
	wire [13-1:0] node2688;
	wire [13-1:0] node2689;
	wire [13-1:0] node2690;
	wire [13-1:0] node2691;
	wire [13-1:0] node2694;
	wire [13-1:0] node2697;
	wire [13-1:0] node2698;
	wire [13-1:0] node2699;
	wire [13-1:0] node2702;
	wire [13-1:0] node2705;
	wire [13-1:0] node2706;
	wire [13-1:0] node2710;
	wire [13-1:0] node2711;
	wire [13-1:0] node2712;
	wire [13-1:0] node2714;
	wire [13-1:0] node2717;
	wire [13-1:0] node2719;
	wire [13-1:0] node2722;
	wire [13-1:0] node2723;
	wire [13-1:0] node2726;
	wire [13-1:0] node2728;
	wire [13-1:0] node2731;
	wire [13-1:0] node2732;
	wire [13-1:0] node2733;
	wire [13-1:0] node2734;
	wire [13-1:0] node2735;
	wire [13-1:0] node2737;
	wire [13-1:0] node2740;
	wire [13-1:0] node2743;
	wire [13-1:0] node2744;
	wire [13-1:0] node2746;
	wire [13-1:0] node2749;
	wire [13-1:0] node2751;
	wire [13-1:0] node2754;
	wire [13-1:0] node2755;
	wire [13-1:0] node2756;
	wire [13-1:0] node2758;
	wire [13-1:0] node2761;
	wire [13-1:0] node2762;
	wire [13-1:0] node2766;
	wire [13-1:0] node2768;
	wire [13-1:0] node2769;
	wire [13-1:0] node2772;
	wire [13-1:0] node2775;
	wire [13-1:0] node2776;
	wire [13-1:0] node2777;
	wire [13-1:0] node2778;
	wire [13-1:0] node2779;
	wire [13-1:0] node2782;
	wire [13-1:0] node2785;
	wire [13-1:0] node2786;
	wire [13-1:0] node2789;
	wire [13-1:0] node2792;
	wire [13-1:0] node2793;
	wire [13-1:0] node2794;
	wire [13-1:0] node2798;
	wire [13-1:0] node2799;
	wire [13-1:0] node2803;
	wire [13-1:0] node2804;
	wire [13-1:0] node2805;
	wire [13-1:0] node2806;
	wire [13-1:0] node2809;
	wire [13-1:0] node2812;
	wire [13-1:0] node2813;
	wire [13-1:0] node2817;
	wire [13-1:0] node2818;
	wire [13-1:0] node2819;
	wire [13-1:0] node2822;
	wire [13-1:0] node2825;
	wire [13-1:0] node2826;
	wire [13-1:0] node2829;
	wire [13-1:0] node2832;
	wire [13-1:0] node2833;
	wire [13-1:0] node2834;
	wire [13-1:0] node2835;
	wire [13-1:0] node2836;
	wire [13-1:0] node2837;
	wire [13-1:0] node2838;
	wire [13-1:0] node2840;
	wire [13-1:0] node2843;
	wire [13-1:0] node2844;
	wire [13-1:0] node2848;
	wire [13-1:0] node2849;
	wire [13-1:0] node2852;
	wire [13-1:0] node2853;
	wire [13-1:0] node2857;
	wire [13-1:0] node2858;
	wire [13-1:0] node2859;
	wire [13-1:0] node2860;
	wire [13-1:0] node2863;
	wire [13-1:0] node2866;
	wire [13-1:0] node2868;
	wire [13-1:0] node2871;
	wire [13-1:0] node2872;
	wire [13-1:0] node2873;
	wire [13-1:0] node2877;
	wire [13-1:0] node2879;
	wire [13-1:0] node2882;
	wire [13-1:0] node2883;
	wire [13-1:0] node2884;
	wire [13-1:0] node2885;
	wire [13-1:0] node2886;
	wire [13-1:0] node2890;
	wire [13-1:0] node2892;
	wire [13-1:0] node2895;
	wire [13-1:0] node2896;
	wire [13-1:0] node2897;
	wire [13-1:0] node2900;
	wire [13-1:0] node2904;
	wire [13-1:0] node2905;
	wire [13-1:0] node2907;
	wire [13-1:0] node2908;
	wire [13-1:0] node2911;
	wire [13-1:0] node2914;
	wire [13-1:0] node2915;
	wire [13-1:0] node2916;
	wire [13-1:0] node2919;
	wire [13-1:0] node2922;
	wire [13-1:0] node2923;
	wire [13-1:0] node2926;
	wire [13-1:0] node2929;
	wire [13-1:0] node2930;
	wire [13-1:0] node2931;
	wire [13-1:0] node2932;
	wire [13-1:0] node2933;
	wire [13-1:0] node2934;
	wire [13-1:0] node2937;
	wire [13-1:0] node2940;
	wire [13-1:0] node2941;
	wire [13-1:0] node2945;
	wire [13-1:0] node2946;
	wire [13-1:0] node2947;
	wire [13-1:0] node2950;
	wire [13-1:0] node2953;
	wire [13-1:0] node2954;
	wire [13-1:0] node2957;
	wire [13-1:0] node2960;
	wire [13-1:0] node2961;
	wire [13-1:0] node2962;
	wire [13-1:0] node2964;
	wire [13-1:0] node2967;
	wire [13-1:0] node2968;
	wire [13-1:0] node2972;
	wire [13-1:0] node2973;
	wire [13-1:0] node2974;
	wire [13-1:0] node2977;
	wire [13-1:0] node2980;
	wire [13-1:0] node2981;
	wire [13-1:0] node2984;
	wire [13-1:0] node2987;
	wire [13-1:0] node2988;
	wire [13-1:0] node2989;
	wire [13-1:0] node2991;
	wire [13-1:0] node2993;
	wire [13-1:0] node2996;
	wire [13-1:0] node2997;
	wire [13-1:0] node2998;
	wire [13-1:0] node3001;
	wire [13-1:0] node3004;
	wire [13-1:0] node3005;
	wire [13-1:0] node3008;
	wire [13-1:0] node3011;
	wire [13-1:0] node3012;
	wire [13-1:0] node3013;
	wire [13-1:0] node3014;
	wire [13-1:0] node3018;
	wire [13-1:0] node3020;
	wire [13-1:0] node3023;
	wire [13-1:0] node3024;
	wire [13-1:0] node3027;
	wire [13-1:0] node3029;
	wire [13-1:0] node3032;
	wire [13-1:0] node3033;
	wire [13-1:0] node3034;
	wire [13-1:0] node3035;
	wire [13-1:0] node3036;
	wire [13-1:0] node3037;
	wire [13-1:0] node3038;
	wire [13-1:0] node3041;
	wire [13-1:0] node3044;
	wire [13-1:0] node3045;
	wire [13-1:0] node3048;
	wire [13-1:0] node3051;
	wire [13-1:0] node3052;
	wire [13-1:0] node3054;
	wire [13-1:0] node3057;
	wire [13-1:0] node3058;
	wire [13-1:0] node3061;
	wire [13-1:0] node3064;
	wire [13-1:0] node3065;
	wire [13-1:0] node3066;
	wire [13-1:0] node3067;
	wire [13-1:0] node3071;
	wire [13-1:0] node3072;
	wire [13-1:0] node3075;
	wire [13-1:0] node3078;
	wire [13-1:0] node3079;
	wire [13-1:0] node3080;
	wire [13-1:0] node3083;
	wire [13-1:0] node3086;
	wire [13-1:0] node3087;
	wire [13-1:0] node3091;
	wire [13-1:0] node3092;
	wire [13-1:0] node3093;
	wire [13-1:0] node3094;
	wire [13-1:0] node3095;
	wire [13-1:0] node3098;
	wire [13-1:0] node3101;
	wire [13-1:0] node3103;
	wire [13-1:0] node3106;
	wire [13-1:0] node3107;
	wire [13-1:0] node3109;
	wire [13-1:0] node3112;
	wire [13-1:0] node3113;
	wire [13-1:0] node3116;
	wire [13-1:0] node3119;
	wire [13-1:0] node3120;
	wire [13-1:0] node3121;
	wire [13-1:0] node3125;
	wire [13-1:0] node3126;
	wire [13-1:0] node3128;
	wire [13-1:0] node3131;
	wire [13-1:0] node3134;
	wire [13-1:0] node3135;
	wire [13-1:0] node3136;
	wire [13-1:0] node3137;
	wire [13-1:0] node3138;
	wire [13-1:0] node3139;
	wire [13-1:0] node3142;
	wire [13-1:0] node3145;
	wire [13-1:0] node3147;
	wire [13-1:0] node3150;
	wire [13-1:0] node3151;
	wire [13-1:0] node3152;
	wire [13-1:0] node3155;
	wire [13-1:0] node3158;
	wire [13-1:0] node3159;
	wire [13-1:0] node3163;
	wire [13-1:0] node3164;
	wire [13-1:0] node3165;
	wire [13-1:0] node3166;
	wire [13-1:0] node3169;
	wire [13-1:0] node3172;
	wire [13-1:0] node3173;
	wire [13-1:0] node3176;
	wire [13-1:0] node3179;
	wire [13-1:0] node3180;
	wire [13-1:0] node3181;
	wire [13-1:0] node3184;
	wire [13-1:0] node3187;
	wire [13-1:0] node3189;
	wire [13-1:0] node3192;
	wire [13-1:0] node3193;
	wire [13-1:0] node3194;
	wire [13-1:0] node3195;
	wire [13-1:0] node3197;
	wire [13-1:0] node3201;
	wire [13-1:0] node3202;
	wire [13-1:0] node3203;
	wire [13-1:0] node3207;
	wire [13-1:0] node3208;
	wire [13-1:0] node3211;
	wire [13-1:0] node3214;
	wire [13-1:0] node3215;
	wire [13-1:0] node3216;
	wire [13-1:0] node3217;
	wire [13-1:0] node3220;
	wire [13-1:0] node3223;
	wire [13-1:0] node3224;
	wire [13-1:0] node3227;
	wire [13-1:0] node3230;
	wire [13-1:0] node3231;
	wire [13-1:0] node3233;
	wire [13-1:0] node3236;
	wire [13-1:0] node3237;
	wire [13-1:0] node3240;

	assign outp = (inp[5]) ? node1652 : node1;
		assign node1 = (inp[2]) ? node809 : node2;
			assign node2 = (inp[3]) ? node406 : node3;
				assign node3 = (inp[10]) ? node201 : node4;
					assign node4 = (inp[7]) ? node96 : node5;
						assign node5 = (inp[9]) ? node51 : node6;
							assign node6 = (inp[1]) ? node32 : node7;
								assign node7 = (inp[4]) ? node21 : node8;
									assign node8 = (inp[6]) ? node14 : node9;
										assign node9 = (inp[11]) ? node11 : 13'b0111111111111;
											assign node11 = (inp[12]) ? 13'b0001111111111 : 13'b0011111111111;
										assign node14 = (inp[8]) ? node18 : node15;
											assign node15 = (inp[11]) ? 13'b0001111111111 : 13'b0011111111111;
											assign node18 = (inp[11]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node21 = (inp[12]) ? node27 : node22;
										assign node22 = (inp[0]) ? 13'b0000011111111 : node23;
											assign node23 = (inp[11]) ? 13'b0001111111111 : 13'b0011111111111;
										assign node27 = (inp[8]) ? node29 : 13'b0000111111111;
											assign node29 = (inp[0]) ? 13'b0000111111111 : 13'b0000111111111;
								assign node32 = (inp[12]) ? node38 : node33;
									assign node33 = (inp[6]) ? 13'b0000111111111 : node34;
										assign node34 = (inp[11]) ? 13'b0001111111111 : 13'b0011111111111;
									assign node38 = (inp[0]) ? node44 : node39;
										assign node39 = (inp[8]) ? node41 : 13'b0000111111111;
											assign node41 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node44 = (inp[6]) ? node48 : node45;
											assign node45 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node48 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node51 = (inp[12]) ? node75 : node52;
								assign node52 = (inp[4]) ? node66 : node53;
									assign node53 = (inp[1]) ? node59 : node54;
										assign node54 = (inp[8]) ? node56 : 13'b0000111111111;
											assign node56 = (inp[0]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node59 = (inp[8]) ? node63 : node60;
											assign node60 = (inp[0]) ? 13'b0000111111111 : 13'b0000111111111;
											assign node63 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node66 = (inp[6]) ? node70 : node67;
										assign node67 = (inp[8]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node70 = (inp[8]) ? 13'b0000011111111 : node71;
											assign node71 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node75 = (inp[11]) ? node85 : node76;
									assign node76 = (inp[8]) ? node80 : node77;
										assign node77 = (inp[4]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node80 = (inp[4]) ? node82 : 13'b0000011111111;
											assign node82 = (inp[6]) ? 13'b0000011111111 : 13'b0000011111111;
									assign node85 = (inp[0]) ? node89 : node86;
										assign node86 = (inp[4]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node89 = (inp[8]) ? node93 : node90;
											assign node90 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node93 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node96 = (inp[8]) ? node148 : node97;
							assign node97 = (inp[0]) ? node123 : node98;
								assign node98 = (inp[4]) ? node110 : node99;
									assign node99 = (inp[9]) ? node105 : node100;
										assign node100 = (inp[1]) ? node102 : 13'b0011111111111;
											assign node102 = (inp[11]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node105 = (inp[12]) ? 13'b0000111111111 : node106;
											assign node106 = (inp[1]) ? 13'b0000111111111 : 13'b0000111111111;
									assign node110 = (inp[1]) ? node116 : node111;
										assign node111 = (inp[9]) ? node113 : 13'b0000111111111;
											assign node113 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node116 = (inp[11]) ? node120 : node117;
											assign node117 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node120 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node123 = (inp[12]) ? node137 : node124;
									assign node124 = (inp[6]) ? node132 : node125;
										assign node125 = (inp[11]) ? node129 : node126;
											assign node126 = (inp[4]) ? 13'b0000111111111 : 13'b0000111111111;
											assign node129 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node132 = (inp[9]) ? 13'b0000001111111 : node133;
											assign node133 = (inp[4]) ? 13'b0000011111111 : 13'b0000011111111;
									assign node137 = (inp[1]) ? node143 : node138;
										assign node138 = (inp[9]) ? 13'b0000011111111 : node139;
											assign node139 = (inp[4]) ? 13'b0000011111111 : 13'b0000011111111;
										assign node143 = (inp[11]) ? 13'b0000001111111 : node144;
											assign node144 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node148 = (inp[11]) ? node170 : node149;
								assign node149 = (inp[6]) ? node159 : node150;
									assign node150 = (inp[1]) ? node154 : node151;
										assign node151 = (inp[0]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node154 = (inp[0]) ? 13'b0000011111111 : node155;
											assign node155 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node159 = (inp[1]) ? node167 : node160;
										assign node160 = (inp[9]) ? node164 : node161;
											assign node161 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node164 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node167 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node170 = (inp[12]) ? node186 : node171;
									assign node171 = (inp[9]) ? node179 : node172;
										assign node172 = (inp[6]) ? node176 : node173;
											assign node173 = (inp[1]) ? 13'b0000111111111 : 13'b0000111111111;
											assign node176 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node179 = (inp[1]) ? node183 : node180;
											assign node180 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node183 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node186 = (inp[0]) ? node194 : node187;
										assign node187 = (inp[1]) ? node191 : node188;
											assign node188 = (inp[4]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node191 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node194 = (inp[4]) ? node198 : node195;
											assign node195 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node198 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
					assign node201 = (inp[8]) ? node301 : node202;
						assign node202 = (inp[11]) ? node252 : node203;
							assign node203 = (inp[1]) ? node229 : node204;
								assign node204 = (inp[7]) ? node216 : node205;
									assign node205 = (inp[6]) ? node211 : node206;
										assign node206 = (inp[4]) ? node208 : 13'b0011111111111;
											assign node208 = (inp[12]) ? 13'b0001111111111 : 13'b0001111111111;
										assign node211 = (inp[0]) ? node213 : 13'b0001111111111;
											assign node213 = (inp[4]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node216 = (inp[12]) ? node224 : node217;
										assign node217 = (inp[9]) ? node221 : node218;
											assign node218 = (inp[0]) ? 13'b0001111111111 : 13'b0011111111111;
											assign node221 = (inp[4]) ? 13'b0000111111111 : 13'b0000111111111;
										assign node224 = (inp[0]) ? 13'b0000011111111 : node225;
											assign node225 = (inp[4]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node229 = (inp[6]) ? node241 : node230;
									assign node230 = (inp[12]) ? node236 : node231;
										assign node231 = (inp[9]) ? 13'b0000111111111 : node232;
											assign node232 = (inp[0]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node236 = (inp[4]) ? 13'b0000011111111 : node237;
											assign node237 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node241 = (inp[7]) ? node247 : node242;
										assign node242 = (inp[0]) ? 13'b0000011111111 : node243;
											assign node243 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node247 = (inp[12]) ? node249 : 13'b0000011111111;
											assign node249 = (inp[0]) ? 13'b0000000111111 : 13'b0000011111111;
							assign node252 = (inp[7]) ? node278 : node253;
								assign node253 = (inp[12]) ? node265 : node254;
									assign node254 = (inp[4]) ? node262 : node255;
										assign node255 = (inp[6]) ? node259 : node256;
											assign node256 = (inp[1]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node259 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node262 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node265 = (inp[0]) ? node273 : node266;
										assign node266 = (inp[9]) ? node270 : node267;
											assign node267 = (inp[1]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node270 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node273 = (inp[9]) ? 13'b0000001111111 : node274;
											assign node274 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node278 = (inp[9]) ? node288 : node279;
									assign node279 = (inp[1]) ? node281 : 13'b0000011111111;
										assign node281 = (inp[6]) ? node285 : node282;
											assign node282 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node285 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node288 = (inp[0]) ? node296 : node289;
										assign node289 = (inp[1]) ? node293 : node290;
											assign node290 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node293 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node296 = (inp[12]) ? node298 : 13'b0000000111111;
											assign node298 = (inp[4]) ? 13'b0000000001111 : 13'b0000000111111;
						assign node301 = (inp[0]) ? node355 : node302;
							assign node302 = (inp[7]) ? node332 : node303;
								assign node303 = (inp[11]) ? node317 : node304;
									assign node304 = (inp[4]) ? node312 : node305;
										assign node305 = (inp[6]) ? node309 : node306;
											assign node306 = (inp[12]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node309 = (inp[9]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node312 = (inp[6]) ? 13'b0000001111111 : node313;
											assign node313 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node317 = (inp[12]) ? node325 : node318;
										assign node318 = (inp[9]) ? node322 : node319;
											assign node319 = (inp[4]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node322 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node325 = (inp[1]) ? node329 : node326;
											assign node326 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node329 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node332 = (inp[1]) ? node342 : node333;
									assign node333 = (inp[9]) ? 13'b0000001111111 : node334;
										assign node334 = (inp[6]) ? node338 : node335;
											assign node335 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node338 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node342 = (inp[6]) ? node348 : node343;
										assign node343 = (inp[11]) ? node345 : 13'b0000011111111;
											assign node345 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node348 = (inp[11]) ? node352 : node349;
											assign node349 = (inp[9]) ? 13'b0000000011111 : 13'b0000001111111;
											assign node352 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node355 = (inp[6]) ? node377 : node356;
								assign node356 = (inp[12]) ? node370 : node357;
									assign node357 = (inp[7]) ? node365 : node358;
										assign node358 = (inp[11]) ? node362 : node359;
											assign node359 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node362 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node365 = (inp[4]) ? 13'b0000000011111 : node366;
											assign node366 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node370 = (inp[9]) ? node372 : 13'b0000001111111;
										assign node372 = (inp[1]) ? 13'b0000000111111 : node373;
											assign node373 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node377 = (inp[9]) ? node393 : node378;
									assign node378 = (inp[1]) ? node386 : node379;
										assign node379 = (inp[4]) ? node383 : node380;
											assign node380 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node383 = (inp[12]) ? 13'b0000000011111 : 13'b0000001111111;
										assign node386 = (inp[7]) ? node390 : node387;
											assign node387 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node390 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node393 = (inp[4]) ? node399 : node394;
										assign node394 = (inp[12]) ? 13'b0000000111111 : node395;
											assign node395 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node399 = (inp[11]) ? node403 : node400;
											assign node400 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node403 = (inp[1]) ? 13'b0000000001111 : 13'b0000000001111;
				assign node406 = (inp[1]) ? node612 : node407;
					assign node407 = (inp[8]) ? node509 : node408;
						assign node408 = (inp[10]) ? node458 : node409;
							assign node409 = (inp[11]) ? node437 : node410;
								assign node410 = (inp[0]) ? node424 : node411;
									assign node411 = (inp[6]) ? node417 : node412;
										assign node412 = (inp[7]) ? node414 : 13'b0011111111111;
											assign node414 = (inp[9]) ? 13'b0001111111111 : 13'b0001111111111;
										assign node417 = (inp[9]) ? node421 : node418;
											assign node418 = (inp[4]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node421 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node424 = (inp[7]) ? node432 : node425;
										assign node425 = (inp[9]) ? node429 : node426;
											assign node426 = (inp[12]) ? 13'b0000111111111 : 13'b0000111111111;
											assign node429 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node432 = (inp[4]) ? 13'b0000011111111 : node433;
											assign node433 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node437 = (inp[7]) ? node449 : node438;
									assign node438 = (inp[12]) ? node444 : node439;
										assign node439 = (inp[6]) ? 13'b0000111111111 : node440;
											assign node440 = (inp[9]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node444 = (inp[4]) ? node446 : 13'b0000111111111;
											assign node446 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node449 = (inp[6]) ? node451 : 13'b0000011111111;
										assign node451 = (inp[9]) ? node455 : node452;
											assign node452 = (inp[4]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node455 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node458 = (inp[6]) ? node490 : node459;
								assign node459 = (inp[11]) ? node475 : node460;
									assign node460 = (inp[7]) ? node468 : node461;
										assign node461 = (inp[0]) ? node465 : node462;
											assign node462 = (inp[4]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node465 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node468 = (inp[12]) ? node472 : node469;
											assign node469 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node472 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node475 = (inp[7]) ? node483 : node476;
										assign node476 = (inp[0]) ? node480 : node477;
											assign node477 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node480 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node483 = (inp[9]) ? node487 : node484;
											assign node484 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node487 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node490 = (inp[0]) ? node500 : node491;
									assign node491 = (inp[12]) ? 13'b0000001111111 : node492;
										assign node492 = (inp[9]) ? node496 : node493;
											assign node493 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node496 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node500 = (inp[12]) ? 13'b0000000111111 : node501;
										assign node501 = (inp[11]) ? node505 : node502;
											assign node502 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node505 = (inp[7]) ? 13'b0000000111111 : 13'b0000000111111;
						assign node509 = (inp[11]) ? node559 : node510;
							assign node510 = (inp[4]) ? node532 : node511;
								assign node511 = (inp[6]) ? node519 : node512;
									assign node512 = (inp[10]) ? 13'b0000011111111 : node513;
										assign node513 = (inp[7]) ? node515 : 13'b0001111111111;
											assign node515 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node519 = (inp[9]) ? node527 : node520;
										assign node520 = (inp[12]) ? node524 : node521;
											assign node521 = (inp[0]) ? 13'b0000011111111 : 13'b0000011111111;
											assign node524 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node527 = (inp[10]) ? 13'b0000001111111 : node528;
											assign node528 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node532 = (inp[0]) ? node548 : node533;
									assign node533 = (inp[6]) ? node541 : node534;
										assign node534 = (inp[10]) ? node538 : node535;
											assign node535 = (inp[9]) ? 13'b0000011111111 : 13'b0000011111111;
											assign node538 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node541 = (inp[9]) ? node545 : node542;
											assign node542 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node545 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node548 = (inp[7]) ? node554 : node549;
										assign node549 = (inp[10]) ? 13'b0000001111111 : node550;
											assign node550 = (inp[12]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node554 = (inp[10]) ? 13'b0000000111111 : node555;
											assign node555 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node559 = (inp[7]) ? node585 : node560;
								assign node560 = (inp[0]) ? node574 : node561;
									assign node561 = (inp[10]) ? node569 : node562;
										assign node562 = (inp[9]) ? node566 : node563;
											assign node563 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node566 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node569 = (inp[4]) ? 13'b0000001111111 : node570;
											assign node570 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node574 = (inp[4]) ? node580 : node575;
										assign node575 = (inp[9]) ? node577 : 13'b0000011111111;
											assign node577 = (inp[6]) ? 13'b0000000011111 : 13'b0000001111111;
										assign node580 = (inp[6]) ? 13'b0000000111111 : node581;
											assign node581 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node585 = (inp[9]) ? node599 : node586;
									assign node586 = (inp[12]) ? node592 : node587;
										assign node587 = (inp[10]) ? 13'b0000001111111 : node588;
											assign node588 = (inp[0]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node592 = (inp[0]) ? node596 : node593;
											assign node593 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node596 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node599 = (inp[0]) ? node607 : node600;
										assign node600 = (inp[6]) ? node604 : node601;
											assign node601 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node604 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node607 = (inp[12]) ? 13'b0000000001111 : node608;
											assign node608 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
					assign node612 = (inp[4]) ? node714 : node613;
						assign node613 = (inp[7]) ? node657 : node614;
							assign node614 = (inp[8]) ? node634 : node615;
								assign node615 = (inp[12]) ? node621 : node616;
									assign node616 = (inp[6]) ? 13'b0000011111111 : node617;
										assign node617 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node621 = (inp[9]) ? node629 : node622;
										assign node622 = (inp[11]) ? node626 : node623;
											assign node623 = (inp[10]) ? 13'b0000011111111 : 13'b0000011111111;
											assign node626 = (inp[0]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node629 = (inp[6]) ? 13'b0000001111111 : node630;
											assign node630 = (inp[10]) ? 13'b0000001111111 : 13'b0000001111111;
								assign node634 = (inp[12]) ? node648 : node635;
									assign node635 = (inp[11]) ? node643 : node636;
										assign node636 = (inp[6]) ? node640 : node637;
											assign node637 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node640 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node643 = (inp[9]) ? node645 : 13'b0000001111111;
											assign node645 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node648 = (inp[0]) ? node650 : 13'b0000001111111;
										assign node650 = (inp[10]) ? node654 : node651;
											assign node651 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node654 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node657 = (inp[6]) ? node689 : node658;
								assign node658 = (inp[12]) ? node674 : node659;
									assign node659 = (inp[11]) ? node667 : node660;
										assign node660 = (inp[9]) ? node664 : node661;
											assign node661 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node664 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node667 = (inp[8]) ? node671 : node668;
											assign node668 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node671 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node674 = (inp[11]) ? node682 : node675;
										assign node675 = (inp[10]) ? node679 : node676;
											assign node676 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node679 = (inp[9]) ? 13'b0000000111111 : 13'b0000011111111;
										assign node682 = (inp[9]) ? node686 : node683;
											assign node683 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node686 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node689 = (inp[0]) ? node703 : node690;
									assign node690 = (inp[8]) ? node698 : node691;
										assign node691 = (inp[10]) ? node695 : node692;
											assign node692 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node695 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node698 = (inp[12]) ? node700 : 13'b0000000111111;
											assign node700 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node703 = (inp[12]) ? node711 : node704;
										assign node704 = (inp[11]) ? node708 : node705;
											assign node705 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node708 = (inp[10]) ? 13'b0000000001111 : 13'b0000000111111;
										assign node711 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node714 = (inp[8]) ? node758 : node715;
							assign node715 = (inp[0]) ? node737 : node716;
								assign node716 = (inp[7]) ? node726 : node717;
									assign node717 = (inp[11]) ? 13'b0000001111111 : node718;
										assign node718 = (inp[6]) ? node722 : node719;
											assign node719 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node722 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node726 = (inp[10]) ? node732 : node727;
										assign node727 = (inp[9]) ? 13'b0000000111111 : node728;
											assign node728 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node732 = (inp[12]) ? node734 : 13'b0000001111111;
											assign node734 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node737 = (inp[11]) ? node751 : node738;
									assign node738 = (inp[12]) ? node744 : node739;
										assign node739 = (inp[7]) ? node741 : 13'b0000011111111;
											assign node741 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node744 = (inp[9]) ? node748 : node745;
											assign node745 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node748 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node751 = (inp[6]) ? node755 : node752;
										assign node752 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node755 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node758 = (inp[7]) ? node782 : node759;
								assign node759 = (inp[10]) ? node769 : node760;
									assign node760 = (inp[12]) ? 13'b0000000111111 : node761;
										assign node761 = (inp[9]) ? node765 : node762;
											assign node762 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node765 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node769 = (inp[9]) ? node777 : node770;
										assign node770 = (inp[6]) ? node774 : node771;
											assign node771 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node774 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node777 = (inp[11]) ? node779 : 13'b0000000011111;
											assign node779 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node782 = (inp[0]) ? node796 : node783;
									assign node783 = (inp[10]) ? node791 : node784;
										assign node784 = (inp[6]) ? node788 : node785;
											assign node785 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node788 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node791 = (inp[11]) ? node793 : 13'b0000000011111;
											assign node793 = (inp[12]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node796 = (inp[10]) ? node804 : node797;
										assign node797 = (inp[11]) ? node801 : node798;
											assign node798 = (inp[6]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node801 = (inp[9]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node804 = (inp[6]) ? node806 : 13'b0000000001111;
											assign node806 = (inp[12]) ? 13'b0000000000111 : 13'b0000000001111;
			assign node809 = (inp[0]) ? node1219 : node810;
				assign node810 = (inp[8]) ? node1014 : node811;
					assign node811 = (inp[7]) ? node913 : node812;
						assign node812 = (inp[6]) ? node864 : node813;
							assign node813 = (inp[1]) ? node841 : node814;
								assign node814 = (inp[10]) ? node826 : node815;
									assign node815 = (inp[12]) ? node821 : node816;
										assign node816 = (inp[9]) ? node818 : 13'b0011111111111;
											assign node818 = (inp[11]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node821 = (inp[3]) ? 13'b0000111111111 : node822;
											assign node822 = (inp[4]) ? 13'b0000111111111 : 13'b0000111111111;
									assign node826 = (inp[9]) ? node834 : node827;
										assign node827 = (inp[3]) ? node831 : node828;
											assign node828 = (inp[11]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node831 = (inp[4]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node834 = (inp[3]) ? node838 : node835;
											assign node835 = (inp[4]) ? 13'b0000011111111 : 13'b0000011111111;
											assign node838 = (inp[11]) ? 13'b0000001111111 : 13'b0000111111111;
								assign node841 = (inp[4]) ? node851 : node842;
									assign node842 = (inp[9]) ? node844 : 13'b0000111111111;
										assign node844 = (inp[3]) ? node848 : node845;
											assign node845 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node848 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node851 = (inp[3]) ? node859 : node852;
										assign node852 = (inp[11]) ? node856 : node853;
											assign node853 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node856 = (inp[12]) ? 13'b0000001111111 : 13'b0000001111111;
										assign node859 = (inp[11]) ? node861 : 13'b0000001111111;
											assign node861 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node864 = (inp[12]) ? node892 : node865;
								assign node865 = (inp[9]) ? node879 : node866;
									assign node866 = (inp[11]) ? node874 : node867;
										assign node867 = (inp[4]) ? node871 : node868;
											assign node868 = (inp[3]) ? 13'b0001111111111 : 13'b0011111111111;
											assign node871 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node874 = (inp[10]) ? 13'b0000011111111 : node875;
											assign node875 = (inp[1]) ? 13'b0000011111111 : 13'b0000011111111;
									assign node879 = (inp[1]) ? node887 : node880;
										assign node880 = (inp[10]) ? node884 : node881;
											assign node881 = (inp[4]) ? 13'b0000011111111 : 13'b0000011111111;
											assign node884 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node887 = (inp[4]) ? node889 : 13'b0000011111111;
											assign node889 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node892 = (inp[3]) ? node906 : node893;
									assign node893 = (inp[4]) ? node901 : node894;
										assign node894 = (inp[11]) ? node898 : node895;
											assign node895 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node898 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node901 = (inp[1]) ? 13'b0000000111111 : node902;
											assign node902 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node906 = (inp[10]) ? node908 : 13'b0000001111111;
										assign node908 = (inp[1]) ? 13'b0000000111111 : node909;
											assign node909 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node913 = (inp[12]) ? node965 : node914;
							assign node914 = (inp[9]) ? node942 : node915;
								assign node915 = (inp[11]) ? node929 : node916;
									assign node916 = (inp[6]) ? node924 : node917;
										assign node917 = (inp[10]) ? node921 : node918;
											assign node918 = (inp[4]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node921 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node924 = (inp[4]) ? node926 : 13'b0000011111111;
											assign node926 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node929 = (inp[6]) ? node935 : node930;
										assign node930 = (inp[10]) ? node932 : 13'b0000011111111;
											assign node932 = (inp[1]) ? 13'b0000011111111 : 13'b0000011111111;
										assign node935 = (inp[10]) ? node939 : node936;
											assign node936 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node939 = (inp[4]) ? 13'b0000000011111 : 13'b0000001111111;
								assign node942 = (inp[4]) ? node958 : node943;
									assign node943 = (inp[3]) ? node951 : node944;
										assign node944 = (inp[10]) ? node948 : node945;
											assign node945 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node948 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node951 = (inp[6]) ? node955 : node952;
											assign node952 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node955 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node958 = (inp[11]) ? 13'b0000000111111 : node959;
										assign node959 = (inp[1]) ? node961 : 13'b0000001111111;
											assign node961 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node965 = (inp[1]) ? node991 : node966;
								assign node966 = (inp[10]) ? node980 : node967;
									assign node967 = (inp[3]) ? node973 : node968;
										assign node968 = (inp[11]) ? node970 : 13'b0000011111111;
											assign node970 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node973 = (inp[4]) ? node977 : node974;
											assign node974 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node977 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node980 = (inp[6]) ? node986 : node981;
										assign node981 = (inp[3]) ? node983 : 13'b0000001111111;
											assign node983 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node986 = (inp[9]) ? 13'b0000000111111 : node987;
											assign node987 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node991 = (inp[3]) ? node1001 : node992;
									assign node992 = (inp[9]) ? node996 : node993;
										assign node993 = (inp[4]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node996 = (inp[10]) ? 13'b0000000111111 : node997;
											assign node997 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1001 = (inp[11]) ? node1007 : node1002;
										assign node1002 = (inp[4]) ? 13'b0000000111111 : node1003;
											assign node1003 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1007 = (inp[9]) ? node1011 : node1008;
											assign node1008 = (inp[4]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node1011 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
					assign node1014 = (inp[7]) ? node1124 : node1015;
						assign node1015 = (inp[10]) ? node1073 : node1016;
							assign node1016 = (inp[6]) ? node1044 : node1017;
								assign node1017 = (inp[9]) ? node1031 : node1018;
									assign node1018 = (inp[1]) ? node1024 : node1019;
										assign node1019 = (inp[3]) ? 13'b0000111111111 : node1020;
											assign node1020 = (inp[12]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node1024 = (inp[3]) ? node1028 : node1025;
											assign node1025 = (inp[11]) ? 13'b0000011111111 : 13'b0000011111111;
											assign node1028 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1031 = (inp[3]) ? node1039 : node1032;
										assign node1032 = (inp[4]) ? node1036 : node1033;
											assign node1033 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1036 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1039 = (inp[4]) ? 13'b0000000111111 : node1040;
											assign node1040 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node1044 = (inp[4]) ? node1060 : node1045;
									assign node1045 = (inp[11]) ? node1053 : node1046;
										assign node1046 = (inp[12]) ? node1050 : node1047;
											assign node1047 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1050 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1053 = (inp[12]) ? node1057 : node1054;
											assign node1054 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1057 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1060 = (inp[1]) ? node1068 : node1061;
										assign node1061 = (inp[12]) ? node1065 : node1062;
											assign node1062 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1065 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1068 = (inp[3]) ? 13'b0000000111111 : node1069;
											assign node1069 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node1073 = (inp[1]) ? node1099 : node1074;
								assign node1074 = (inp[3]) ? node1088 : node1075;
									assign node1075 = (inp[11]) ? node1081 : node1076;
										assign node1076 = (inp[4]) ? node1078 : 13'b0000111111111;
											assign node1078 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1081 = (inp[6]) ? node1085 : node1082;
											assign node1082 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1085 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1088 = (inp[4]) ? node1094 : node1089;
										assign node1089 = (inp[12]) ? node1091 : 13'b0000001111111;
											assign node1091 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1094 = (inp[9]) ? 13'b0000000011111 : node1095;
											assign node1095 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1099 = (inp[9]) ? node1111 : node1100;
									assign node1100 = (inp[6]) ? node1106 : node1101;
										assign node1101 = (inp[11]) ? 13'b0000001111111 : node1102;
											assign node1102 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1106 = (inp[12]) ? node1108 : 13'b0000001111111;
											assign node1108 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1111 = (inp[11]) ? node1117 : node1112;
										assign node1112 = (inp[6]) ? node1114 : 13'b0000000111111;
											assign node1114 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1117 = (inp[12]) ? node1121 : node1118;
											assign node1118 = (inp[4]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node1121 = (inp[6]) ? 13'b0000000000111 : 13'b0000000011111;
						assign node1124 = (inp[11]) ? node1166 : node1125;
							assign node1125 = (inp[4]) ? node1143 : node1126;
								assign node1126 = (inp[1]) ? node1134 : node1127;
									assign node1127 = (inp[12]) ? node1129 : 13'b0000011111111;
										assign node1129 = (inp[6]) ? 13'b0000000111111 : node1130;
											assign node1130 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1134 = (inp[3]) ? node1140 : node1135;
										assign node1135 = (inp[10]) ? node1137 : 13'b0000001111111;
											assign node1137 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1140 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node1143 = (inp[12]) ? node1153 : node1144;
									assign node1144 = (inp[10]) ? node1146 : 13'b0000000111111;
										assign node1146 = (inp[3]) ? node1150 : node1147;
											assign node1147 = (inp[1]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node1150 = (inp[1]) ? 13'b0000000111111 : 13'b0000000111111;
									assign node1153 = (inp[10]) ? node1159 : node1154;
										assign node1154 = (inp[6]) ? 13'b0000000111111 : node1155;
											assign node1155 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1159 = (inp[6]) ? node1163 : node1160;
											assign node1160 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1163 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node1166 = (inp[1]) ? node1194 : node1167;
								assign node1167 = (inp[3]) ? node1181 : node1168;
									assign node1168 = (inp[12]) ? node1176 : node1169;
										assign node1169 = (inp[10]) ? node1173 : node1170;
											assign node1170 = (inp[4]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node1173 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1176 = (inp[9]) ? 13'b0000000011111 : node1177;
											assign node1177 = (inp[6]) ? 13'b0000000111111 : 13'b0000000111111;
									assign node1181 = (inp[9]) ? node1187 : node1182;
										assign node1182 = (inp[4]) ? node1184 : 13'b0000001111111;
											assign node1184 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1187 = (inp[10]) ? node1191 : node1188;
											assign node1188 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1191 = (inp[6]) ? 13'b0000000000111 : 13'b0000000011111;
								assign node1194 = (inp[9]) ? node1208 : node1195;
									assign node1195 = (inp[10]) ? node1201 : node1196;
										assign node1196 = (inp[4]) ? node1198 : 13'b0000000111111;
											assign node1198 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1201 = (inp[3]) ? node1205 : node1202;
											assign node1202 = (inp[12]) ? 13'b0000000001111 : 13'b0000000111111;
											assign node1205 = (inp[4]) ? 13'b0000000001111 : 13'b0000000001111;
									assign node1208 = (inp[3]) ? node1214 : node1209;
										assign node1209 = (inp[6]) ? node1211 : 13'b0000000011111;
											assign node1211 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1214 = (inp[10]) ? node1216 : 13'b0000000001111;
											assign node1216 = (inp[4]) ? 13'b0000000000011 : 13'b0000000000111;
				assign node1219 = (inp[11]) ? node1435 : node1220;
					assign node1220 = (inp[10]) ? node1326 : node1221;
						assign node1221 = (inp[6]) ? node1273 : node1222;
							assign node1222 = (inp[1]) ? node1246 : node1223;
								assign node1223 = (inp[7]) ? node1237 : node1224;
									assign node1224 = (inp[4]) ? node1230 : node1225;
										assign node1225 = (inp[8]) ? node1227 : 13'b0001111111111;
											assign node1227 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1230 = (inp[8]) ? node1234 : node1231;
											assign node1231 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1234 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1237 = (inp[3]) ? node1243 : node1238;
										assign node1238 = (inp[4]) ? 13'b0000011111111 : node1239;
											assign node1239 = (inp[8]) ? 13'b0000011111111 : 13'b0000011111111;
										assign node1243 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node1246 = (inp[12]) ? node1262 : node1247;
									assign node1247 = (inp[7]) ? node1255 : node1248;
										assign node1248 = (inp[3]) ? node1252 : node1249;
											assign node1249 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1252 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1255 = (inp[9]) ? node1259 : node1256;
											assign node1256 = (inp[8]) ? 13'b0000001111111 : 13'b0000111111111;
											assign node1259 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1262 = (inp[8]) ? node1268 : node1263;
										assign node1263 = (inp[9]) ? 13'b0000001111111 : node1264;
											assign node1264 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1268 = (inp[3]) ? node1270 : 13'b0000001111111;
											assign node1270 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node1273 = (inp[9]) ? node1299 : node1274;
								assign node1274 = (inp[1]) ? node1286 : node1275;
									assign node1275 = (inp[4]) ? node1281 : node1276;
										assign node1276 = (inp[7]) ? 13'b0000011111111 : node1277;
											assign node1277 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1281 = (inp[8]) ? 13'b0000001111111 : node1282;
											assign node1282 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1286 = (inp[12]) ? node1292 : node1287;
										assign node1287 = (inp[4]) ? 13'b0000001111111 : node1288;
											assign node1288 = (inp[7]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node1292 = (inp[4]) ? node1296 : node1293;
											assign node1293 = (inp[8]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node1296 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1299 = (inp[3]) ? node1311 : node1300;
									assign node1300 = (inp[4]) ? node1306 : node1301;
										assign node1301 = (inp[12]) ? 13'b0000001111111 : node1302;
											assign node1302 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1306 = (inp[1]) ? 13'b0000000011111 : node1307;
											assign node1307 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1311 = (inp[8]) ? node1319 : node1312;
										assign node1312 = (inp[7]) ? node1316 : node1313;
											assign node1313 = (inp[12]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node1316 = (inp[4]) ? 13'b0000000011111 : 13'b0000000011111;
										assign node1319 = (inp[12]) ? node1323 : node1320;
											assign node1320 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1323 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node1326 = (inp[1]) ? node1382 : node1327;
							assign node1327 = (inp[9]) ? node1357 : node1328;
								assign node1328 = (inp[4]) ? node1342 : node1329;
									assign node1329 = (inp[7]) ? node1335 : node1330;
										assign node1330 = (inp[6]) ? node1332 : 13'b0000111111111;
											assign node1332 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1335 = (inp[3]) ? node1339 : node1336;
											assign node1336 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1339 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1342 = (inp[8]) ? node1350 : node1343;
										assign node1343 = (inp[6]) ? node1347 : node1344;
											assign node1344 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1347 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1350 = (inp[6]) ? node1354 : node1351;
											assign node1351 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1354 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node1357 = (inp[7]) ? node1373 : node1358;
									assign node1358 = (inp[4]) ? node1366 : node1359;
										assign node1359 = (inp[12]) ? node1363 : node1360;
											assign node1360 = (inp[3]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node1363 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1366 = (inp[6]) ? node1370 : node1367;
											assign node1367 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1370 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1373 = (inp[12]) ? node1377 : node1374;
										assign node1374 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1377 = (inp[4]) ? node1379 : 13'b0000000011111;
											assign node1379 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node1382 = (inp[12]) ? node1408 : node1383;
								assign node1383 = (inp[4]) ? node1395 : node1384;
									assign node1384 = (inp[9]) ? node1390 : node1385;
										assign node1385 = (inp[8]) ? node1387 : 13'b0000001111111;
											assign node1387 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1390 = (inp[6]) ? node1392 : 13'b0000000111111;
											assign node1392 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1395 = (inp[8]) ? node1403 : node1396;
										assign node1396 = (inp[7]) ? node1400 : node1397;
											assign node1397 = (inp[6]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node1400 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1403 = (inp[7]) ? node1405 : 13'b0000000011111;
											assign node1405 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1408 = (inp[9]) ? node1420 : node1409;
									assign node1409 = (inp[8]) ? node1415 : node1410;
										assign node1410 = (inp[6]) ? node1412 : 13'b0000000111111;
											assign node1412 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1415 = (inp[4]) ? node1417 : 13'b0000000011111;
											assign node1417 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1420 = (inp[8]) ? node1428 : node1421;
										assign node1421 = (inp[4]) ? node1425 : node1422;
											assign node1422 = (inp[3]) ? 13'b0000000011111 : 13'b0000001111111;
											assign node1425 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1428 = (inp[6]) ? node1432 : node1429;
											assign node1429 = (inp[3]) ? 13'b0000000001111 : 13'b0000000111111;
											assign node1432 = (inp[4]) ? 13'b0000000000111 : 13'b0000000001111;
					assign node1435 = (inp[4]) ? node1545 : node1436;
						assign node1436 = (inp[8]) ? node1492 : node1437;
							assign node1437 = (inp[9]) ? node1465 : node1438;
								assign node1438 = (inp[12]) ? node1450 : node1439;
									assign node1439 = (inp[3]) ? node1443 : node1440;
										assign node1440 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1443 = (inp[10]) ? node1447 : node1444;
											assign node1444 = (inp[7]) ? 13'b0000001111111 : 13'b0000111111111;
											assign node1447 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1450 = (inp[10]) ? node1458 : node1451;
										assign node1451 = (inp[7]) ? node1455 : node1452;
											assign node1452 = (inp[3]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node1455 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1458 = (inp[6]) ? node1462 : node1459;
											assign node1459 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1462 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node1465 = (inp[3]) ? node1479 : node1466;
									assign node1466 = (inp[7]) ? node1472 : node1467;
										assign node1467 = (inp[1]) ? 13'b0000001111111 : node1468;
											assign node1468 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1472 = (inp[6]) ? node1476 : node1473;
											assign node1473 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1476 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1479 = (inp[10]) ? node1485 : node1480;
										assign node1480 = (inp[12]) ? node1482 : 13'b0000000111111;
											assign node1482 = (inp[1]) ? 13'b0000000011111 : 13'b0000000011111;
										assign node1485 = (inp[12]) ? node1489 : node1486;
											assign node1486 = (inp[7]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node1489 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node1492 = (inp[3]) ? node1518 : node1493;
								assign node1493 = (inp[10]) ? node1505 : node1494;
									assign node1494 = (inp[12]) ? node1500 : node1495;
										assign node1495 = (inp[6]) ? node1497 : 13'b0000001111111;
											assign node1497 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1500 = (inp[7]) ? node1502 : 13'b0000000111111;
											assign node1502 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1505 = (inp[1]) ? node1513 : node1506;
										assign node1506 = (inp[7]) ? node1510 : node1507;
											assign node1507 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1510 = (inp[6]) ? 13'b0000000011111 : 13'b0000000011111;
										assign node1513 = (inp[7]) ? 13'b0000000001111 : node1514;
											assign node1514 = (inp[6]) ? 13'b0000000011111 : 13'b0000000011111;
								assign node1518 = (inp[12]) ? node1532 : node1519;
									assign node1519 = (inp[1]) ? node1525 : node1520;
										assign node1520 = (inp[6]) ? node1522 : 13'b0000001111111;
											assign node1522 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1525 = (inp[9]) ? node1529 : node1526;
											assign node1526 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1529 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1532 = (inp[9]) ? node1540 : node1533;
										assign node1533 = (inp[1]) ? node1537 : node1534;
											assign node1534 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1537 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1540 = (inp[10]) ? node1542 : 13'b0000000001111;
											assign node1542 = (inp[1]) ? 13'b0000000000111 : 13'b0000000001111;
						assign node1545 = (inp[10]) ? node1595 : node1546;
							assign node1546 = (inp[12]) ? node1572 : node1547;
								assign node1547 = (inp[1]) ? node1559 : node1548;
									assign node1548 = (inp[7]) ? node1554 : node1549;
										assign node1549 = (inp[8]) ? 13'b0000001111111 : node1550;
											assign node1550 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1554 = (inp[6]) ? 13'b0000000111111 : node1555;
											assign node1555 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1559 = (inp[3]) ? node1565 : node1560;
										assign node1560 = (inp[7]) ? node1562 : 13'b0000001111111;
											assign node1562 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1565 = (inp[8]) ? node1569 : node1566;
											assign node1566 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1569 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1572 = (inp[3]) ? node1582 : node1573;
									assign node1573 = (inp[1]) ? node1575 : 13'b0000000111111;
										assign node1575 = (inp[7]) ? node1579 : node1576;
											assign node1576 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1579 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1582 = (inp[8]) ? node1590 : node1583;
										assign node1583 = (inp[1]) ? node1587 : node1584;
											assign node1584 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1587 = (inp[7]) ? 13'b0000000000111 : 13'b0000000011111;
										assign node1590 = (inp[1]) ? 13'b0000000000111 : node1591;
											assign node1591 = (inp[6]) ? 13'b0000000001111 : 13'b0000000001111;
							assign node1595 = (inp[8]) ? node1625 : node1596;
								assign node1596 = (inp[1]) ? node1610 : node1597;
									assign node1597 = (inp[12]) ? node1603 : node1598;
										assign node1598 = (inp[3]) ? node1600 : 13'b0000000111111;
											assign node1600 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1603 = (inp[7]) ? node1607 : node1604;
											assign node1604 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1607 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1610 = (inp[3]) ? node1618 : node1611;
										assign node1611 = (inp[7]) ? node1615 : node1612;
											assign node1612 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1615 = (inp[9]) ? 13'b0000000000111 : 13'b0000000011111;
										assign node1618 = (inp[12]) ? node1622 : node1619;
											assign node1619 = (inp[6]) ? 13'b0000000001111 : 13'b0000000001111;
											assign node1622 = (inp[7]) ? 13'b0000000000011 : 13'b0000000000111;
								assign node1625 = (inp[7]) ? node1639 : node1626;
									assign node1626 = (inp[3]) ? node1634 : node1627;
										assign node1627 = (inp[9]) ? node1631 : node1628;
											assign node1628 = (inp[12]) ? 13'b0000000011111 : 13'b0000001111111;
											assign node1631 = (inp[12]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1634 = (inp[12]) ? 13'b0000000000111 : node1635;
											assign node1635 = (inp[1]) ? 13'b0000000001111 : 13'b0000000001111;
									assign node1639 = (inp[9]) ? node1645 : node1640;
										assign node1640 = (inp[12]) ? 13'b0000000001111 : node1641;
											assign node1641 = (inp[3]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node1645 = (inp[12]) ? node1649 : node1646;
											assign node1646 = (inp[3]) ? 13'b0000000000111 : 13'b0000000001111;
											assign node1649 = (inp[1]) ? 13'b0000000000011 : 13'b0000000000011;
		assign node1652 = (inp[6]) ? node2448 : node1653;
			assign node1653 = (inp[8]) ? node2029 : node1654;
				assign node1654 = (inp[10]) ? node1824 : node1655;
					assign node1655 = (inp[0]) ? node1741 : node1656;
						assign node1656 = (inp[7]) ? node1694 : node1657;
							assign node1657 = (inp[4]) ? node1673 : node1658;
								assign node1658 = (inp[11]) ? node1666 : node1659;
									assign node1659 = (inp[2]) ? 13'b0000111111111 : node1660;
										assign node1660 = (inp[1]) ? node1662 : 13'b0011111111111;
											assign node1662 = (inp[12]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node1666 = (inp[9]) ? node1668 : 13'b0000111111111;
										assign node1668 = (inp[3]) ? node1670 : 13'b0000111111111;
											assign node1670 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node1673 = (inp[12]) ? node1683 : node1674;
									assign node1674 = (inp[11]) ? node1678 : node1675;
										assign node1675 = (inp[9]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node1678 = (inp[2]) ? 13'b0000001111111 : node1679;
											assign node1679 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node1683 = (inp[2]) ? node1691 : node1684;
										assign node1684 = (inp[11]) ? node1688 : node1685;
											assign node1685 = (inp[3]) ? 13'b0000011111111 : 13'b0001111111111;
											assign node1688 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1691 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node1694 = (inp[12]) ? node1720 : node1695;
								assign node1695 = (inp[9]) ? node1709 : node1696;
									assign node1696 = (inp[11]) ? node1702 : node1697;
										assign node1697 = (inp[3]) ? node1699 : 13'b0001111111111;
											assign node1699 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1702 = (inp[2]) ? node1706 : node1703;
											assign node1703 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1706 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1709 = (inp[4]) ? node1715 : node1710;
										assign node1710 = (inp[3]) ? 13'b0000001111111 : node1711;
											assign node1711 = (inp[11]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node1715 = (inp[11]) ? 13'b0000001111111 : node1716;
											assign node1716 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node1720 = (inp[3]) ? node1734 : node1721;
									assign node1721 = (inp[1]) ? node1727 : node1722;
										assign node1722 = (inp[9]) ? 13'b0000011111111 : node1723;
											assign node1723 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1727 = (inp[2]) ? node1731 : node1728;
											assign node1728 = (inp[11]) ? 13'b0000001111111 : 13'b0000111111111;
											assign node1731 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1734 = (inp[4]) ? 13'b0000000111111 : node1735;
										assign node1735 = (inp[2]) ? node1737 : 13'b0000011111111;
											assign node1737 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node1741 = (inp[3]) ? node1781 : node1742;
							assign node1742 = (inp[1]) ? node1766 : node1743;
								assign node1743 = (inp[4]) ? node1755 : node1744;
									assign node1744 = (inp[9]) ? node1752 : node1745;
										assign node1745 = (inp[2]) ? node1749 : node1746;
											assign node1746 = (inp[12]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node1749 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1752 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1755 = (inp[11]) ? node1761 : node1756;
										assign node1756 = (inp[9]) ? node1758 : 13'b0000011111111;
											assign node1758 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1761 = (inp[2]) ? 13'b0000001111111 : node1762;
											assign node1762 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node1766 = (inp[11]) ? node1774 : node1767;
									assign node1767 = (inp[7]) ? node1771 : node1768;
										assign node1768 = (inp[4]) ? 13'b0000111111111 : 13'b0000011111111;
										assign node1771 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1774 = (inp[4]) ? node1776 : 13'b0000001111111;
										assign node1776 = (inp[12]) ? 13'b0000000011111 : node1777;
											assign node1777 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node1781 = (inp[9]) ? node1807 : node1782;
								assign node1782 = (inp[2]) ? node1796 : node1783;
									assign node1783 = (inp[12]) ? node1789 : node1784;
										assign node1784 = (inp[11]) ? 13'b0000011111111 : node1785;
											assign node1785 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1789 = (inp[11]) ? node1793 : node1790;
											assign node1790 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1793 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1796 = (inp[12]) ? node1804 : node1797;
										assign node1797 = (inp[1]) ? node1801 : node1798;
											assign node1798 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1801 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1804 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node1807 = (inp[12]) ? node1817 : node1808;
									assign node1808 = (inp[2]) ? node1812 : node1809;
										assign node1809 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1812 = (inp[1]) ? node1814 : 13'b0000000111111;
											assign node1814 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1817 = (inp[4]) ? 13'b0000000001111 : node1818;
										assign node1818 = (inp[1]) ? node1820 : 13'b0000000011111;
											assign node1820 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
					assign node1824 = (inp[1]) ? node1932 : node1825;
						assign node1825 = (inp[2]) ? node1885 : node1826;
							assign node1826 = (inp[4]) ? node1854 : node1827;
								assign node1827 = (inp[3]) ? node1839 : node1828;
									assign node1828 = (inp[12]) ? node1836 : node1829;
										assign node1829 = (inp[7]) ? node1833 : node1830;
											assign node1830 = (inp[11]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node1833 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1836 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node1839 = (inp[7]) ? node1847 : node1840;
										assign node1840 = (inp[11]) ? node1844 : node1841;
											assign node1841 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1844 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1847 = (inp[0]) ? node1851 : node1848;
											assign node1848 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1851 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1854 = (inp[12]) ? node1870 : node1855;
									assign node1855 = (inp[11]) ? node1863 : node1856;
										assign node1856 = (inp[7]) ? node1860 : node1857;
											assign node1857 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node1860 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1863 = (inp[7]) ? node1867 : node1864;
											assign node1864 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1867 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1870 = (inp[7]) ? node1878 : node1871;
										assign node1871 = (inp[11]) ? node1875 : node1872;
											assign node1872 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1875 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1878 = (inp[0]) ? node1882 : node1879;
											assign node1879 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1882 = (inp[11]) ? 13'b0000000011111 : 13'b0000000011111;
							assign node1885 = (inp[12]) ? node1905 : node1886;
								assign node1886 = (inp[4]) ? node1894 : node1887;
									assign node1887 = (inp[3]) ? 13'b0000001111111 : node1888;
										assign node1888 = (inp[9]) ? node1890 : 13'b0000011111111;
											assign node1890 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1894 = (inp[0]) ? node1902 : node1895;
										assign node1895 = (inp[11]) ? node1899 : node1896;
											assign node1896 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1899 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1902 = (inp[7]) ? 13'b0000000011111 : 13'b0000001111111;
								assign node1905 = (inp[11]) ? node1917 : node1906;
									assign node1906 = (inp[7]) ? node1912 : node1907;
										assign node1907 = (inp[4]) ? 13'b0000001111111 : node1908;
											assign node1908 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1912 = (inp[3]) ? node1914 : 13'b0000001111111;
											assign node1914 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1917 = (inp[9]) ? node1925 : node1918;
										assign node1918 = (inp[3]) ? node1922 : node1919;
											assign node1919 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1922 = (inp[0]) ? 13'b0000000011111 : 13'b0000000011111;
										assign node1925 = (inp[7]) ? node1929 : node1926;
											assign node1926 = (inp[4]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node1929 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node1932 = (inp[12]) ? node1986 : node1933;
							assign node1933 = (inp[11]) ? node1959 : node1934;
								assign node1934 = (inp[4]) ? node1948 : node1935;
									assign node1935 = (inp[7]) ? node1941 : node1936;
										assign node1936 = (inp[3]) ? 13'b0000011111111 : node1937;
											assign node1937 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node1941 = (inp[3]) ? node1945 : node1942;
											assign node1942 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node1945 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1948 = (inp[3]) ? node1954 : node1949;
										assign node1949 = (inp[7]) ? node1951 : 13'b0000001111111;
											assign node1951 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1954 = (inp[0]) ? node1956 : 13'b0000001111111;
											assign node1956 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1959 = (inp[2]) ? node1971 : node1960;
									assign node1960 = (inp[0]) ? node1966 : node1961;
										assign node1961 = (inp[4]) ? node1963 : 13'b0000001111111;
											assign node1963 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1966 = (inp[9]) ? 13'b0000000111111 : node1967;
											assign node1967 = (inp[4]) ? 13'b0000001111111 : 13'b0000000111111;
									assign node1971 = (inp[7]) ? node1979 : node1972;
										assign node1972 = (inp[9]) ? node1976 : node1973;
											assign node1973 = (inp[4]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node1976 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1979 = (inp[4]) ? node1983 : node1980;
											assign node1980 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1983 = (inp[3]) ? 13'b0000000001111 : 13'b0000000001111;
							assign node1986 = (inp[3]) ? node2008 : node1987;
								assign node1987 = (inp[7]) ? node1999 : node1988;
									assign node1988 = (inp[9]) ? node1992 : node1989;
										assign node1989 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node1992 = (inp[2]) ? node1996 : node1993;
											assign node1993 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node1996 = (inp[0]) ? 13'b0000000011111 : 13'b0000000011111;
									assign node1999 = (inp[9]) ? node2003 : node2000;
										assign node2000 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2003 = (inp[4]) ? 13'b0000000011111 : node2004;
											assign node2004 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node2008 = (inp[2]) ? node2020 : node2009;
									assign node2009 = (inp[11]) ? node2015 : node2010;
										assign node2010 = (inp[4]) ? node2012 : 13'b0000001111111;
											assign node2012 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2015 = (inp[7]) ? node2017 : 13'b0000000011111;
											assign node2017 = (inp[4]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2020 = (inp[0]) ? node2024 : node2021;
										assign node2021 = (inp[4]) ? 13'b0000000011111 : 13'b0000000001111;
										assign node2024 = (inp[4]) ? node2026 : 13'b0000000001111;
											assign node2026 = (inp[9]) ? 13'b0000000000111 : 13'b0000000001111;
				assign node2029 = (inp[4]) ? node2235 : node2030;
					assign node2030 = (inp[9]) ? node2130 : node2031;
						assign node2031 = (inp[3]) ? node2085 : node2032;
							assign node2032 = (inp[11]) ? node2060 : node2033;
								assign node2033 = (inp[12]) ? node2047 : node2034;
									assign node2034 = (inp[0]) ? node2042 : node2035;
										assign node2035 = (inp[2]) ? node2039 : node2036;
											assign node2036 = (inp[7]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node2039 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node2042 = (inp[1]) ? node2044 : 13'b0000011111111;
											assign node2044 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node2047 = (inp[7]) ? node2055 : node2048;
										assign node2048 = (inp[0]) ? node2052 : node2049;
											assign node2049 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2052 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2055 = (inp[1]) ? node2057 : 13'b0000011111111;
											assign node2057 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node2060 = (inp[7]) ? node2070 : node2061;
									assign node2061 = (inp[1]) ? node2065 : node2062;
										assign node2062 = (inp[12]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node2065 = (inp[0]) ? 13'b0000001111111 : node2066;
											assign node2066 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node2070 = (inp[1]) ? node2078 : node2071;
										assign node2071 = (inp[12]) ? node2075 : node2072;
											assign node2072 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2075 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2078 = (inp[10]) ? node2082 : node2079;
											assign node2079 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2082 = (inp[0]) ? 13'b0000000111111 : 13'b0000000011111;
							assign node2085 = (inp[7]) ? node2107 : node2086;
								assign node2086 = (inp[0]) ? node2098 : node2087;
									assign node2087 = (inp[2]) ? node2095 : node2088;
										assign node2088 = (inp[1]) ? node2092 : node2089;
											assign node2089 = (inp[11]) ? 13'b0000011111111 : 13'b0000011111111;
											assign node2092 = (inp[10]) ? 13'b0000000111111 : 13'b0000011111111;
										assign node2095 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2098 = (inp[2]) ? 13'b0000000111111 : node2099;
										assign node2099 = (inp[1]) ? node2103 : node2100;
											assign node2100 = (inp[11]) ? 13'b0000011111111 : 13'b0000001111111;
											assign node2103 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node2107 = (inp[11]) ? node2119 : node2108;
									assign node2108 = (inp[1]) ? node2114 : node2109;
										assign node2109 = (inp[10]) ? node2111 : 13'b0000001111111;
											assign node2111 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2114 = (inp[10]) ? 13'b0000000111111 : node2115;
											assign node2115 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2119 = (inp[1]) ? node2123 : node2120;
										assign node2120 = (inp[12]) ? 13'b0000000011111 : 13'b0000001111111;
										assign node2123 = (inp[10]) ? node2127 : node2124;
											assign node2124 = (inp[12]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node2127 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node2130 = (inp[11]) ? node2182 : node2131;
							assign node2131 = (inp[12]) ? node2159 : node2132;
								assign node2132 = (inp[0]) ? node2146 : node2133;
									assign node2133 = (inp[2]) ? node2139 : node2134;
										assign node2134 = (inp[3]) ? node2136 : 13'b0000111111111;
											assign node2136 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2139 = (inp[1]) ? node2143 : node2140;
											assign node2140 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2143 = (inp[3]) ? 13'b0000000011111 : 13'b0000001111111;
									assign node2146 = (inp[2]) ? node2154 : node2147;
										assign node2147 = (inp[7]) ? node2151 : node2148;
											assign node2148 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2151 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2154 = (inp[3]) ? 13'b0000000111111 : node2155;
											assign node2155 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node2159 = (inp[3]) ? node2171 : node2160;
									assign node2160 = (inp[10]) ? node2164 : node2161;
										assign node2161 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2164 = (inp[1]) ? node2168 : node2165;
											assign node2165 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2168 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2171 = (inp[1]) ? node2177 : node2172;
										assign node2172 = (inp[0]) ? node2174 : 13'b0000001111111;
											assign node2174 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2177 = (inp[2]) ? node2179 : 13'b0000000111111;
											assign node2179 = (inp[0]) ? 13'b0000000001111 : 13'b0000000001111;
							assign node2182 = (inp[2]) ? node2208 : node2183;
								assign node2183 = (inp[0]) ? node2195 : node2184;
									assign node2184 = (inp[3]) ? node2192 : node2185;
										assign node2185 = (inp[1]) ? node2189 : node2186;
											assign node2186 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2189 = (inp[7]) ? 13'b0000001111111 : 13'b0000000111111;
										assign node2192 = (inp[1]) ? 13'b0000001111111 : 13'b0000000111111;
									assign node2195 = (inp[3]) ? node2201 : node2196;
										assign node2196 = (inp[10]) ? node2198 : 13'b0000000111111;
											assign node2198 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2201 = (inp[10]) ? node2205 : node2202;
											assign node2202 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2205 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node2208 = (inp[12]) ? node2224 : node2209;
									assign node2209 = (inp[0]) ? node2217 : node2210;
										assign node2210 = (inp[1]) ? node2214 : node2211;
											assign node2211 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2214 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2217 = (inp[10]) ? node2221 : node2218;
											assign node2218 = (inp[3]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node2221 = (inp[3]) ? 13'b0000000000111 : 13'b0000000011111;
									assign node2224 = (inp[1]) ? node2230 : node2225;
										assign node2225 = (inp[10]) ? node2227 : 13'b0000000011111;
											assign node2227 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2230 = (inp[7]) ? node2232 : 13'b0000000001111;
											assign node2232 = (inp[10]) ? 13'b0000000000011 : 13'b0000000000111;
					assign node2235 = (inp[1]) ? node2343 : node2236;
						assign node2236 = (inp[10]) ? node2292 : node2237;
							assign node2237 = (inp[3]) ? node2267 : node2238;
								assign node2238 = (inp[0]) ? node2252 : node2239;
									assign node2239 = (inp[12]) ? node2247 : node2240;
										assign node2240 = (inp[7]) ? node2244 : node2241;
											assign node2241 = (inp[11]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node2244 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2247 = (inp[9]) ? node2249 : 13'b0000011111111;
											assign node2249 = (inp[11]) ? 13'b0000001111111 : 13'b0000001111111;
									assign node2252 = (inp[7]) ? node2260 : node2253;
										assign node2253 = (inp[12]) ? node2257 : node2254;
											assign node2254 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2257 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2260 = (inp[9]) ? node2264 : node2261;
											assign node2261 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2264 = (inp[11]) ? 13'b0000000001111 : 13'b0000000111111;
								assign node2267 = (inp[2]) ? node2281 : node2268;
									assign node2268 = (inp[11]) ? node2274 : node2269;
										assign node2269 = (inp[7]) ? node2271 : 13'b0000011111111;
											assign node2271 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2274 = (inp[0]) ? node2278 : node2275;
											assign node2275 = (inp[7]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node2278 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2281 = (inp[9]) ? node2287 : node2282;
										assign node2282 = (inp[7]) ? node2284 : 13'b0000000111111;
											assign node2284 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2287 = (inp[7]) ? node2289 : 13'b0000000011111;
											assign node2289 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node2292 = (inp[7]) ? node2318 : node2293;
								assign node2293 = (inp[12]) ? node2305 : node2294;
									assign node2294 = (inp[11]) ? node2300 : node2295;
										assign node2295 = (inp[0]) ? node2297 : 13'b0000001111111;
											assign node2297 = (inp[9]) ? 13'b0000000111111 : 13'b0000000111111;
										assign node2300 = (inp[9]) ? node2302 : 13'b0000011111111;
											assign node2302 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2305 = (inp[2]) ? node2313 : node2306;
										assign node2306 = (inp[11]) ? node2310 : node2307;
											assign node2307 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2310 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2313 = (inp[3]) ? 13'b0000000001111 : node2314;
											assign node2314 = (inp[11]) ? 13'b0000000001111 : 13'b0000000111111;
								assign node2318 = (inp[12]) ? node2334 : node2319;
									assign node2319 = (inp[2]) ? node2327 : node2320;
										assign node2320 = (inp[3]) ? node2324 : node2321;
											assign node2321 = (inp[0]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node2324 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2327 = (inp[9]) ? node2331 : node2328;
											assign node2328 = (inp[3]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node2331 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2334 = (inp[11]) ? node2340 : node2335;
										assign node2335 = (inp[3]) ? node2337 : 13'b0000000011111;
											assign node2337 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2340 = (inp[3]) ? 13'b0000000000111 : 13'b0000000001111;
						assign node2343 = (inp[11]) ? node2391 : node2344;
							assign node2344 = (inp[0]) ? node2368 : node2345;
								assign node2345 = (inp[12]) ? node2355 : node2346;
									assign node2346 = (inp[3]) ? node2352 : node2347;
										assign node2347 = (inp[10]) ? 13'b0000001111111 : node2348;
											assign node2348 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2352 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2355 = (inp[9]) ? node2363 : node2356;
										assign node2356 = (inp[10]) ? node2360 : node2357;
											assign node2357 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2360 = (inp[3]) ? 13'b0000000001111 : 13'b0000000111111;
										assign node2363 = (inp[2]) ? node2365 : 13'b0000000011111;
											assign node2365 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node2368 = (inp[7]) ? node2380 : node2369;
									assign node2369 = (inp[12]) ? node2375 : node2370;
										assign node2370 = (inp[10]) ? node2372 : 13'b0000001111111;
											assign node2372 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2375 = (inp[3]) ? node2377 : 13'b0000000011111;
											assign node2377 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2380 = (inp[12]) ? node2388 : node2381;
										assign node2381 = (inp[9]) ? node2385 : node2382;
											assign node2382 = (inp[3]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node2385 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2388 = (inp[9]) ? 13'b0000000000111 : 13'b0000000001111;
							assign node2391 = (inp[3]) ? node2419 : node2392;
								assign node2392 = (inp[7]) ? node2408 : node2393;
									assign node2393 = (inp[0]) ? node2401 : node2394;
										assign node2394 = (inp[10]) ? node2398 : node2395;
											assign node2395 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2398 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2401 = (inp[12]) ? node2405 : node2402;
											assign node2402 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node2405 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2408 = (inp[10]) ? node2414 : node2409;
										assign node2409 = (inp[12]) ? node2411 : 13'b0000000011111;
											assign node2411 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2414 = (inp[0]) ? 13'b0000000000111 : node2415;
											assign node2415 = (inp[12]) ? 13'b0000000001111 : 13'b0000000001111;
								assign node2419 = (inp[9]) ? node2435 : node2420;
									assign node2420 = (inp[12]) ? node2428 : node2421;
										assign node2421 = (inp[2]) ? node2425 : node2422;
											assign node2422 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2425 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2428 = (inp[7]) ? node2432 : node2429;
											assign node2429 = (inp[0]) ? 13'b0000000001111 : 13'b0000000001111;
											assign node2432 = (inp[0]) ? 13'b0000000000111 : 13'b0000000000111;
									assign node2435 = (inp[0]) ? node2441 : node2436;
										assign node2436 = (inp[7]) ? 13'b0000000001111 : node2437;
											assign node2437 = (inp[2]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node2441 = (inp[12]) ? node2445 : node2442;
											assign node2442 = (inp[7]) ? 13'b0000000000111 : 13'b0000000000111;
											assign node2445 = (inp[10]) ? 13'b0000000000011 : 13'b0000000000111;
			assign node2448 = (inp[0]) ? node2832 : node2449;
				assign node2449 = (inp[1]) ? node2643 : node2450;
					assign node2450 = (inp[2]) ? node2548 : node2451;
						assign node2451 = (inp[7]) ? node2493 : node2452;
							assign node2452 = (inp[11]) ? node2476 : node2453;
								assign node2453 = (inp[10]) ? node2465 : node2454;
									assign node2454 = (inp[12]) ? node2462 : node2455;
										assign node2455 = (inp[3]) ? node2459 : node2456;
											assign node2456 = (inp[8]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node2459 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node2462 = (inp[4]) ? 13'b0000011111111 : 13'b0000001111111;
									assign node2465 = (inp[3]) ? node2471 : node2466;
										assign node2466 = (inp[4]) ? node2468 : 13'b0000111111111;
											assign node2468 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2471 = (inp[8]) ? 13'b0000001111111 : node2472;
											assign node2472 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node2476 = (inp[9]) ? node2484 : node2477;
									assign node2477 = (inp[8]) ? node2479 : 13'b0000011111111;
										assign node2479 = (inp[4]) ? 13'b0000000011111 : node2480;
											assign node2480 = (inp[3]) ? 13'b0000001111111 : 13'b0000001111111;
									assign node2484 = (inp[3]) ? node2486 : 13'b0000001111111;
										assign node2486 = (inp[4]) ? node2490 : node2487;
											assign node2487 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2490 = (inp[8]) ? 13'b0000000011111 : 13'b0000000011111;
							assign node2493 = (inp[10]) ? node2523 : node2494;
								assign node2494 = (inp[11]) ? node2508 : node2495;
									assign node2495 = (inp[9]) ? node2501 : node2496;
										assign node2496 = (inp[8]) ? 13'b0000011111111 : node2497;
											assign node2497 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node2501 = (inp[8]) ? node2505 : node2502;
											assign node2502 = (inp[4]) ? 13'b0000001111111 : 13'b0000001111111;
											assign node2505 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2508 = (inp[4]) ? node2516 : node2509;
										assign node2509 = (inp[12]) ? node2513 : node2510;
											assign node2510 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2513 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2516 = (inp[9]) ? node2520 : node2517;
											assign node2517 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2520 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node2523 = (inp[3]) ? node2537 : node2524;
									assign node2524 = (inp[9]) ? node2532 : node2525;
										assign node2525 = (inp[8]) ? node2529 : node2526;
											assign node2526 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2529 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2532 = (inp[11]) ? node2534 : 13'b0000000111111;
											assign node2534 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2537 = (inp[9]) ? node2543 : node2538;
										assign node2538 = (inp[4]) ? node2540 : 13'b0000000111111;
											assign node2540 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2543 = (inp[8]) ? node2545 : 13'b0000001111111;
											assign node2545 = (inp[12]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node2548 = (inp[7]) ? node2600 : node2549;
							assign node2549 = (inp[12]) ? node2571 : node2550;
								assign node2550 = (inp[3]) ? node2562 : node2551;
									assign node2551 = (inp[11]) ? node2557 : node2552;
										assign node2552 = (inp[10]) ? node2554 : 13'b0000011111111;
											assign node2554 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2557 = (inp[4]) ? 13'b0000000111111 : node2558;
											assign node2558 = (inp[8]) ? 13'b0000001111111 : 13'b0000001111111;
									assign node2562 = (inp[10]) ? node2566 : node2563;
										assign node2563 = (inp[11]) ? 13'b0000011111111 : 13'b0000001111111;
										assign node2566 = (inp[11]) ? node2568 : 13'b0000000111111;
											assign node2568 = (inp[8]) ? 13'b0000000001111 : 13'b0000000111111;
								assign node2571 = (inp[3]) ? node2585 : node2572;
									assign node2572 = (inp[8]) ? node2578 : node2573;
										assign node2573 = (inp[11]) ? node2575 : 13'b0000001111111;
											assign node2575 = (inp[4]) ? 13'b0000000111111 : 13'b0000000111111;
										assign node2578 = (inp[9]) ? node2582 : node2579;
											assign node2579 = (inp[10]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node2582 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2585 = (inp[11]) ? node2593 : node2586;
										assign node2586 = (inp[9]) ? node2590 : node2587;
											assign node2587 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2590 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2593 = (inp[4]) ? node2597 : node2594;
											assign node2594 = (inp[9]) ? 13'b0000000011111 : 13'b0000000011111;
											assign node2597 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node2600 = (inp[10]) ? node2624 : node2601;
								assign node2601 = (inp[11]) ? node2611 : node2602;
									assign node2602 = (inp[8]) ? node2604 : 13'b0000001111111;
										assign node2604 = (inp[3]) ? node2608 : node2605;
											assign node2605 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2608 = (inp[9]) ? 13'b0000000011111 : 13'b0000000011111;
									assign node2611 = (inp[8]) ? node2619 : node2612;
										assign node2612 = (inp[12]) ? node2616 : node2613;
											assign node2613 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2616 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2619 = (inp[4]) ? node2621 : 13'b0000000111111;
											assign node2621 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node2624 = (inp[8]) ? node2632 : node2625;
									assign node2625 = (inp[3]) ? 13'b0000000011111 : node2626;
										assign node2626 = (inp[11]) ? node2628 : 13'b0000000111111;
											assign node2628 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2632 = (inp[11]) ? node2638 : node2633;
										assign node2633 = (inp[4]) ? node2635 : 13'b0000000011111;
											assign node2635 = (inp[12]) ? 13'b0000000001111 : 13'b0000000001111;
										assign node2638 = (inp[9]) ? node2640 : 13'b0000000011111;
											assign node2640 = (inp[4]) ? 13'b0000000000111 : 13'b0000000001111;
					assign node2643 = (inp[8]) ? node2731 : node2644;
						assign node2644 = (inp[9]) ? node2688 : node2645;
							assign node2645 = (inp[2]) ? node2665 : node2646;
								assign node2646 = (inp[4]) ? node2654 : node2647;
									assign node2647 = (inp[12]) ? node2649 : 13'b0000011111111;
										assign node2649 = (inp[7]) ? 13'b0000001111111 : node2650;
											assign node2650 = (inp[10]) ? 13'b0000001111111 : 13'b0000001111111;
									assign node2654 = (inp[11]) ? node2658 : node2655;
										assign node2655 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2658 = (inp[7]) ? node2662 : node2659;
											assign node2659 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2662 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node2665 = (inp[10]) ? node2677 : node2666;
									assign node2666 = (inp[4]) ? node2674 : node2667;
										assign node2667 = (inp[3]) ? node2671 : node2668;
											assign node2668 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2671 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2674 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2677 = (inp[11]) ? node2683 : node2678;
										assign node2678 = (inp[3]) ? node2680 : 13'b0000001111111;
											assign node2680 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2683 = (inp[4]) ? node2685 : 13'b0000000011111;
											assign node2685 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node2688 = (inp[4]) ? node2710 : node2689;
								assign node2689 = (inp[3]) ? node2697 : node2690;
									assign node2690 = (inp[11]) ? node2694 : node2691;
										assign node2691 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node2694 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node2697 = (inp[11]) ? node2705 : node2698;
										assign node2698 = (inp[12]) ? node2702 : node2699;
											assign node2699 = (inp[2]) ? 13'b0000000111111 : 13'b0000000111111;
											assign node2702 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2705 = (inp[7]) ? 13'b0000000011111 : node2706;
											assign node2706 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node2710 = (inp[2]) ? node2722 : node2711;
									assign node2711 = (inp[12]) ? node2717 : node2712;
										assign node2712 = (inp[7]) ? node2714 : 13'b0000001111111;
											assign node2714 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2717 = (inp[3]) ? node2719 : 13'b0000000011111;
											assign node2719 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2722 = (inp[11]) ? node2726 : node2723;
										assign node2723 = (inp[3]) ? 13'b0000000001111 : 13'b0000000111111;
										assign node2726 = (inp[7]) ? node2728 : 13'b0000000001111;
											assign node2728 = (inp[3]) ? 13'b0000000000011 : 13'b0000000000111;
						assign node2731 = (inp[12]) ? node2775 : node2732;
							assign node2732 = (inp[3]) ? node2754 : node2733;
								assign node2733 = (inp[2]) ? node2743 : node2734;
									assign node2734 = (inp[4]) ? node2740 : node2735;
										assign node2735 = (inp[7]) ? node2737 : 13'b0000001111111;
											assign node2737 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2740 = (inp[7]) ? 13'b0000000011111 : 13'b0000001111111;
									assign node2743 = (inp[10]) ? node2749 : node2744;
										assign node2744 = (inp[4]) ? node2746 : 13'b0000000111111;
											assign node2746 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2749 = (inp[7]) ? node2751 : 13'b0000000011111;
											assign node2751 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node2754 = (inp[10]) ? node2766 : node2755;
									assign node2755 = (inp[4]) ? node2761 : node2756;
										assign node2756 = (inp[9]) ? node2758 : 13'b0000000111111;
											assign node2758 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2761 = (inp[7]) ? 13'b0000000011111 : node2762;
											assign node2762 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2766 = (inp[2]) ? node2768 : 13'b0000000011111;
										assign node2768 = (inp[11]) ? node2772 : node2769;
											assign node2769 = (inp[9]) ? 13'b0000000000111 : 13'b0000000011111;
											assign node2772 = (inp[9]) ? 13'b0000000000111 : 13'b0000000001111;
							assign node2775 = (inp[11]) ? node2803 : node2776;
								assign node2776 = (inp[2]) ? node2792 : node2777;
									assign node2777 = (inp[7]) ? node2785 : node2778;
										assign node2778 = (inp[9]) ? node2782 : node2779;
											assign node2779 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2782 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2785 = (inp[9]) ? node2789 : node2786;
											assign node2786 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2789 = (inp[10]) ? 13'b0000000001111 : 13'b0000000001111;
									assign node2792 = (inp[3]) ? node2798 : node2793;
										assign node2793 = (inp[4]) ? 13'b0000000001111 : node2794;
											assign node2794 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2798 = (inp[7]) ? 13'b0000000001111 : node2799;
											assign node2799 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node2803 = (inp[9]) ? node2817 : node2804;
									assign node2804 = (inp[7]) ? node2812 : node2805;
										assign node2805 = (inp[3]) ? node2809 : node2806;
											assign node2806 = (inp[10]) ? 13'b0000000111111 : 13'b0000000011111;
											assign node2809 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2812 = (inp[4]) ? 13'b0000000000111 : node2813;
											assign node2813 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2817 = (inp[2]) ? node2825 : node2818;
										assign node2818 = (inp[3]) ? node2822 : node2819;
											assign node2819 = (inp[4]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node2822 = (inp[10]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node2825 = (inp[7]) ? node2829 : node2826;
											assign node2826 = (inp[4]) ? 13'b0000000000111 : 13'b0000000001111;
											assign node2829 = (inp[10]) ? 13'b0000000000011 : 13'b0000000000111;
				assign node2832 = (inp[10]) ? node3032 : node2833;
					assign node2833 = (inp[4]) ? node2929 : node2834;
						assign node2834 = (inp[12]) ? node2882 : node2835;
							assign node2835 = (inp[2]) ? node2857 : node2836;
								assign node2836 = (inp[11]) ? node2848 : node2837;
									assign node2837 = (inp[8]) ? node2843 : node2838;
										assign node2838 = (inp[1]) ? node2840 : 13'b0000011111111;
											assign node2840 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node2843 = (inp[9]) ? 13'b0000001111111 : node2844;
											assign node2844 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node2848 = (inp[7]) ? node2852 : node2849;
										assign node2849 = (inp[1]) ? 13'b0000001111111 : 13'b0000111111111;
										assign node2852 = (inp[3]) ? 13'b0000000111111 : node2853;
											assign node2853 = (inp[9]) ? 13'b0000000111111 : 13'b0000011111111;
								assign node2857 = (inp[1]) ? node2871 : node2858;
									assign node2858 = (inp[11]) ? node2866 : node2859;
										assign node2859 = (inp[9]) ? node2863 : node2860;
											assign node2860 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2863 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2866 = (inp[8]) ? node2868 : 13'b0000001111111;
											assign node2868 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2871 = (inp[9]) ? node2877 : node2872;
										assign node2872 = (inp[8]) ? 13'b0000000111111 : node2873;
											assign node2873 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2877 = (inp[3]) ? node2879 : 13'b0000000011111;
											assign node2879 = (inp[8]) ? 13'b0000000011111 : 13'b0000000011111;
							assign node2882 = (inp[7]) ? node2904 : node2883;
								assign node2883 = (inp[11]) ? node2895 : node2884;
									assign node2884 = (inp[3]) ? node2890 : node2885;
										assign node2885 = (inp[2]) ? 13'b0000001111111 : node2886;
											assign node2886 = (inp[8]) ? 13'b0000011111111 : 13'b0000001111111;
										assign node2890 = (inp[8]) ? node2892 : 13'b0000001111111;
											assign node2892 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node2895 = (inp[2]) ? 13'b0000000011111 : node2896;
										assign node2896 = (inp[1]) ? node2900 : node2897;
											assign node2897 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2900 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node2904 = (inp[2]) ? node2914 : node2905;
									assign node2905 = (inp[9]) ? node2907 : 13'b0000000111111;
										assign node2907 = (inp[3]) ? node2911 : node2908;
											assign node2908 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2911 = (inp[8]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node2914 = (inp[8]) ? node2922 : node2915;
										assign node2915 = (inp[3]) ? node2919 : node2916;
											assign node2916 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2919 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2922 = (inp[9]) ? node2926 : node2923;
											assign node2923 = (inp[11]) ? 13'b0000000000111 : 13'b0000000011111;
											assign node2926 = (inp[1]) ? 13'b0000000000111 : 13'b0000000001111;
						assign node2929 = (inp[11]) ? node2987 : node2930;
							assign node2930 = (inp[2]) ? node2960 : node2931;
								assign node2931 = (inp[1]) ? node2945 : node2932;
									assign node2932 = (inp[7]) ? node2940 : node2933;
										assign node2933 = (inp[12]) ? node2937 : node2934;
											assign node2934 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node2937 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node2940 = (inp[9]) ? 13'b0000000011111 : node2941;
											assign node2941 = (inp[3]) ? 13'b0000000111111 : 13'b0000000111111;
									assign node2945 = (inp[7]) ? node2953 : node2946;
										assign node2946 = (inp[9]) ? node2950 : node2947;
											assign node2947 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node2950 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node2953 = (inp[9]) ? node2957 : node2954;
											assign node2954 = (inp[3]) ? 13'b0000000111111 : 13'b0000000011111;
											assign node2957 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node2960 = (inp[3]) ? node2972 : node2961;
									assign node2961 = (inp[7]) ? node2967 : node2962;
										assign node2962 = (inp[12]) ? node2964 : 13'b0000000111111;
											assign node2964 = (inp[9]) ? 13'b0000000011111 : 13'b0000001111111;
										assign node2967 = (inp[1]) ? 13'b0000000011111 : node2968;
											assign node2968 = (inp[9]) ? 13'b0000000001111 : 13'b0000000111111;
									assign node2972 = (inp[7]) ? node2980 : node2973;
										assign node2973 = (inp[9]) ? node2977 : node2974;
											assign node2974 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node2977 = (inp[8]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node2980 = (inp[9]) ? node2984 : node2981;
											assign node2981 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node2984 = (inp[1]) ? 13'b0000000000011 : 13'b0000000001111;
							assign node2987 = (inp[9]) ? node3011 : node2988;
								assign node2988 = (inp[2]) ? node2996 : node2989;
									assign node2989 = (inp[8]) ? node2991 : 13'b0000001111111;
										assign node2991 = (inp[7]) ? node2993 : 13'b0000000111111;
											assign node2993 = (inp[1]) ? 13'b0000000011111 : 13'b0000000011111;
									assign node2996 = (inp[3]) ? node3004 : node2997;
										assign node2997 = (inp[7]) ? node3001 : node2998;
											assign node2998 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3001 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3004 = (inp[12]) ? node3008 : node3005;
											assign node3005 = (inp[8]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3008 = (inp[1]) ? 13'b0000000001111 : 13'b0000000000111;
								assign node3011 = (inp[1]) ? node3023 : node3012;
									assign node3012 = (inp[7]) ? node3018 : node3013;
										assign node3013 = (inp[2]) ? 13'b0000000001111 : node3014;
											assign node3014 = (inp[12]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3018 = (inp[2]) ? node3020 : 13'b0000000001111;
											assign node3020 = (inp[8]) ? 13'b0000000001111 : 13'b0000000000111;
									assign node3023 = (inp[8]) ? node3027 : node3024;
										assign node3024 = (inp[3]) ? 13'b0000000001111 : 13'b0000000111111;
										assign node3027 = (inp[12]) ? node3029 : 13'b0000000000111;
											assign node3029 = (inp[3]) ? 13'b0000000000011 : 13'b0000000000111;
					assign node3032 = (inp[9]) ? node3134 : node3033;
						assign node3033 = (inp[1]) ? node3091 : node3034;
							assign node3034 = (inp[4]) ? node3064 : node3035;
								assign node3035 = (inp[12]) ? node3051 : node3036;
									assign node3036 = (inp[3]) ? node3044 : node3037;
										assign node3037 = (inp[2]) ? node3041 : node3038;
											assign node3038 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
											assign node3041 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node3044 = (inp[7]) ? node3048 : node3045;
											assign node3045 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
											assign node3048 = (inp[11]) ? 13'b0000000111111 : 13'b0000000011111;
									assign node3051 = (inp[3]) ? node3057 : node3052;
										assign node3052 = (inp[8]) ? node3054 : 13'b0000000111111;
											assign node3054 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node3057 = (inp[7]) ? node3061 : node3058;
											assign node3058 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3061 = (inp[11]) ? 13'b0000000000111 : 13'b0000000011111;
								assign node3064 = (inp[2]) ? node3078 : node3065;
									assign node3065 = (inp[8]) ? node3071 : node3066;
										assign node3066 = (inp[7]) ? 13'b0000000011111 : node3067;
											assign node3067 = (inp[12]) ? 13'b0000000111111 : 13'b0000000111111;
										assign node3071 = (inp[11]) ? node3075 : node3072;
											assign node3072 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3075 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3078 = (inp[11]) ? node3086 : node3079;
										assign node3079 = (inp[8]) ? node3083 : node3080;
											assign node3080 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3083 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3086 = (inp[7]) ? 13'b0000000001111 : node3087;
											assign node3087 = (inp[3]) ? 13'b0000000001111 : 13'b0000000111111;
							assign node3091 = (inp[8]) ? node3119 : node3092;
								assign node3092 = (inp[12]) ? node3106 : node3093;
									assign node3093 = (inp[2]) ? node3101 : node3094;
										assign node3094 = (inp[3]) ? node3098 : node3095;
											assign node3095 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3098 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3101 = (inp[11]) ? node3103 : 13'b0000000011111;
											assign node3103 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3106 = (inp[11]) ? node3112 : node3107;
										assign node3107 = (inp[2]) ? node3109 : 13'b0000000111111;
											assign node3109 = (inp[4]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node3112 = (inp[7]) ? node3116 : node3113;
											assign node3113 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3116 = (inp[3]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node3119 = (inp[3]) ? node3125 : node3120;
									assign node3120 = (inp[2]) ? 13'b0000000001111 : node3121;
										assign node3121 = (inp[12]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3125 = (inp[12]) ? node3131 : node3126;
										assign node3126 = (inp[4]) ? node3128 : 13'b0000000001111;
											assign node3128 = (inp[11]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node3131 = (inp[2]) ? 13'b0000000000011 : 13'b0000000000111;
						assign node3134 = (inp[4]) ? node3192 : node3135;
							assign node3135 = (inp[3]) ? node3163 : node3136;
								assign node3136 = (inp[8]) ? node3150 : node3137;
									assign node3137 = (inp[7]) ? node3145 : node3138;
										assign node3138 = (inp[1]) ? node3142 : node3139;
											assign node3139 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3142 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node3145 = (inp[1]) ? node3147 : 13'b0000000111111;
											assign node3147 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3150 = (inp[11]) ? node3158 : node3151;
										assign node3151 = (inp[1]) ? node3155 : node3152;
											assign node3152 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3155 = (inp[7]) ? 13'b0000000001111 : 13'b0000000001111;
										assign node3158 = (inp[7]) ? 13'b0000000001111 : node3159;
											assign node3159 = (inp[12]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node3163 = (inp[7]) ? node3179 : node3164;
									assign node3164 = (inp[1]) ? node3172 : node3165;
										assign node3165 = (inp[2]) ? node3169 : node3166;
											assign node3166 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node3169 = (inp[12]) ? 13'b0000000000111 : 13'b0000000011111;
										assign node3172 = (inp[8]) ? node3176 : node3173;
											assign node3173 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3176 = (inp[12]) ? 13'b0000000000111 : 13'b0000000001111;
									assign node3179 = (inp[11]) ? node3187 : node3180;
										assign node3180 = (inp[12]) ? node3184 : node3181;
											assign node3181 = (inp[8]) ? 13'b0000000000111 : 13'b0000000011111;
											assign node3184 = (inp[8]) ? 13'b0000000000011 : 13'b0000000000111;
										assign node3187 = (inp[12]) ? node3189 : 13'b0000000000111;
											assign node3189 = (inp[8]) ? 13'b0000000000001 : 13'b0000000000011;
							assign node3192 = (inp[8]) ? node3214 : node3193;
								assign node3193 = (inp[7]) ? node3201 : node3194;
									assign node3194 = (inp[11]) ? 13'b0000000001111 : node3195;
										assign node3195 = (inp[12]) ? node3197 : 13'b0000000011111;
											assign node3197 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node3201 = (inp[1]) ? node3207 : node3202;
										assign node3202 = (inp[11]) ? 13'b0000000000111 : node3203;
											assign node3203 = (inp[2]) ? 13'b0000000001111 : 13'b0000000001111;
										assign node3207 = (inp[3]) ? node3211 : node3208;
											assign node3208 = (inp[2]) ? 13'b0000000000111 : 13'b0000000001111;
											assign node3211 = (inp[11]) ? 13'b0000000000011 : 13'b0000000000111;
								assign node3214 = (inp[12]) ? node3230 : node3215;
									assign node3215 = (inp[1]) ? node3223 : node3216;
										assign node3216 = (inp[3]) ? node3220 : node3217;
											assign node3217 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
											assign node3220 = (inp[7]) ? 13'b0000000000111 : 13'b0000000001111;
										assign node3223 = (inp[3]) ? node3227 : node3224;
											assign node3224 = (inp[2]) ? 13'b0000000000111 : 13'b0000000001111;
											assign node3227 = (inp[7]) ? 13'b0000000000011 : 13'b0000000000111;
									assign node3230 = (inp[11]) ? node3236 : node3231;
										assign node3231 = (inp[3]) ? node3233 : 13'b0000000001111;
											assign node3233 = (inp[7]) ? 13'b0000000000011 : 13'b0000000000111;
										assign node3236 = (inp[3]) ? node3240 : node3237;
											assign node3237 = (inp[7]) ? 13'b0000000000011 : 13'b0000000000111;
											assign node3240 = (inp[7]) ? 13'b0000000000000 : 13'b0000000000011;

endmodule