module dtc_split25_bm93 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node100;

	assign outp = (inp[0]) ? node24 : node1;
		assign node1 = (inp[7]) ? 3'b000 : node2;
			assign node2 = (inp[6]) ? 3'b000 : node3;
				assign node3 = (inp[3]) ? node5 : 3'b000;
					assign node5 = (inp[5]) ? node11 : node6;
						assign node6 = (inp[8]) ? 3'b000 : node7;
							assign node7 = (inp[4]) ? 3'b100 : 3'b000;
						assign node11 = (inp[8]) ? node17 : node12;
							assign node12 = (inp[4]) ? node14 : 3'b010;
								assign node14 = (inp[10]) ? 3'b010 : 3'b100;
							assign node17 = (inp[4]) ? node19 : 3'b100;
								assign node19 = (inp[10]) ? 3'b100 : 3'b000;
		assign node24 = (inp[7]) ? node72 : node25;
			assign node25 = (inp[3]) ? node53 : node26;
				assign node26 = (inp[5]) ? node34 : node27;
					assign node27 = (inp[6]) ? 3'b000 : node28;
						assign node28 = (inp[4]) ? node30 : 3'b000;
							assign node30 = (inp[8]) ? 3'b000 : 3'b110;
					assign node34 = (inp[6]) ? 3'b100 : node35;
						assign node35 = (inp[8]) ? node47 : node36;
							assign node36 = (inp[4]) ? node38 : 3'b100;
								assign node38 = (inp[10]) ? node44 : node39;
									assign node39 = (inp[1]) ? 3'b110 : node40;
										assign node40 = (inp[2]) ? 3'b110 : 3'b010;
									assign node44 = (inp[1]) ? 3'b100 : 3'b000;
							assign node47 = (inp[10]) ? 3'b110 : node48;
								assign node48 = (inp[4]) ? 3'b100 : 3'b110;
				assign node53 = (inp[5]) ? node61 : node54;
					assign node54 = (inp[6]) ? 3'b011 : node55;
						assign node55 = (inp[8]) ? 3'b011 : node56;
							assign node56 = (inp[4]) ? 3'b111 : 3'b011;
					assign node61 = (inp[6]) ? 3'b110 : node62;
						assign node62 = (inp[9]) ? node64 : 3'b111;
							assign node64 = (inp[2]) ? 3'b111 : node65;
								assign node65 = (inp[1]) ? 3'b111 : node66;
									assign node66 = (inp[8]) ? 3'b111 : 3'b011;
			assign node72 = (inp[6]) ? 3'b000 : node73;
				assign node73 = (inp[5]) ? node75 : 3'b000;
					assign node75 = (inp[3]) ? node85 : node76;
						assign node76 = (inp[1]) ? node78 : 3'b000;
							assign node78 = (inp[2]) ? node80 : 3'b000;
								assign node80 = (inp[4]) ? node82 : 3'b100;
									assign node82 = (inp[8]) ? 3'b100 : 3'b000;
						assign node85 = (inp[8]) ? node97 : node86;
							assign node86 = (inp[2]) ? node88 : 3'b011;
								assign node88 = (inp[10]) ? 3'b111 : node89;
									assign node89 = (inp[9]) ? node91 : 3'b011;
										assign node91 = (inp[4]) ? node93 : 3'b111;
											assign node93 = (inp[11]) ? 3'b111 : 3'b011;
							assign node97 = (inp[11]) ? 3'b011 : node98;
								assign node98 = (inp[1]) ? node100 : 3'b001;
									assign node100 = (inp[2]) ? 3'b101 : 3'b001;

endmodule