module dtc_split125_bm71 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node201;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node238;
	wire [3-1:0] node240;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node265;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node280;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node297;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node342;
	wire [3-1:0] node347;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node356;

	assign outp = (inp[6]) ? node110 : node1;
		assign node1 = (inp[9]) ? node93 : node2;
			assign node2 = (inp[7]) ? node28 : node3;
				assign node3 = (inp[0]) ? 3'b000 : node4;
					assign node4 = (inp[10]) ? node20 : node5;
						assign node5 = (inp[11]) ? node15 : node6;
							assign node6 = (inp[4]) ? node8 : 3'b100;
								assign node8 = (inp[1]) ? node10 : 3'b110;
									assign node10 = (inp[2]) ? node12 : 3'b010;
										assign node12 = (inp[5]) ? 3'b100 : 3'b010;
							assign node15 = (inp[5]) ? 3'b100 : node16;
								assign node16 = (inp[2]) ? 3'b000 : 3'b100;
						assign node20 = (inp[3]) ? 3'b000 : node21;
							assign node21 = (inp[1]) ? 3'b000 : node22;
								assign node22 = (inp[8]) ? 3'b100 : 3'b000;
				assign node28 = (inp[0]) ? node68 : node29;
					assign node29 = (inp[10]) ? node43 : node30;
						assign node30 = (inp[8]) ? node38 : node31;
							assign node31 = (inp[1]) ? 3'b010 : node32;
								assign node32 = (inp[11]) ? 3'b110 : node33;
									assign node33 = (inp[3]) ? 3'b110 : 3'b001;
							assign node38 = (inp[4]) ? 3'b001 : node39;
								assign node39 = (inp[3]) ? 3'b001 : 3'b101;
						assign node43 = (inp[11]) ? node55 : node44;
							assign node44 = (inp[1]) ? node52 : node45;
								assign node45 = (inp[8]) ? 3'b110 : node46;
									assign node46 = (inp[4]) ? 3'b010 : node47;
										assign node47 = (inp[3]) ? 3'b010 : 3'b110;
								assign node52 = (inp[8]) ? 3'b010 : 3'b100;
							assign node55 = (inp[8]) ? node59 : node56;
								assign node56 = (inp[1]) ? 3'b000 : 3'b100;
								assign node59 = (inp[2]) ? node65 : node60;
									assign node60 = (inp[3]) ? 3'b010 : node61;
										assign node61 = (inp[1]) ? 3'b010 : 3'b110;
									assign node65 = (inp[1]) ? 3'b100 : 3'b010;
					assign node68 = (inp[10]) ? node86 : node69;
						assign node69 = (inp[3]) ? node83 : node70;
							assign node70 = (inp[2]) ? node80 : node71;
								assign node71 = (inp[8]) ? node77 : node72;
									assign node72 = (inp[4]) ? node74 : 3'b010;
										assign node74 = (inp[5]) ? 3'b000 : 3'b100;
									assign node77 = (inp[5]) ? 3'b110 : 3'b010;
								assign node80 = (inp[11]) ? 3'b010 : 3'b100;
							assign node83 = (inp[5]) ? 3'b000 : 3'b100;
						assign node86 = (inp[11]) ? 3'b000 : node87;
							assign node87 = (inp[1]) ? 3'b000 : node88;
								assign node88 = (inp[3]) ? 3'b100 : 3'b000;
			assign node93 = (inp[0]) ? 3'b000 : node94;
				assign node94 = (inp[10]) ? 3'b000 : node95;
					assign node95 = (inp[5]) ? node103 : node96;
						assign node96 = (inp[3]) ? 3'b000 : node97;
							assign node97 = (inp[4]) ? 3'b000 : node98;
								assign node98 = (inp[7]) ? 3'b010 : 3'b000;
						assign node103 = (inp[8]) ? node105 : 3'b000;
							assign node105 = (inp[4]) ? 3'b100 : 3'b000;
		assign node110 = (inp[9]) ? node250 : node111;
			assign node111 = (inp[0]) ? node179 : node112;
				assign node112 = (inp[10]) ? node148 : node113;
					assign node113 = (inp[7]) ? node131 : node114;
						assign node114 = (inp[8]) ? node120 : node115;
							assign node115 = (inp[3]) ? node117 : 3'b101;
								assign node117 = (inp[11]) ? 3'b101 : 3'b011;
							assign node120 = (inp[1]) ? node126 : node121;
								assign node121 = (inp[3]) ? node123 : 3'b111;
									assign node123 = (inp[11]) ? 3'b011 : 3'b111;
								assign node126 = (inp[2]) ? 3'b101 : node127;
									assign node127 = (inp[11]) ? 3'b101 : 3'b011;
						assign node131 = (inp[3]) ? node141 : node132;
							assign node132 = (inp[4]) ? node134 : 3'b111;
								assign node134 = (inp[11]) ? node136 : 3'b111;
									assign node136 = (inp[2]) ? node138 : 3'b111;
										assign node138 = (inp[5]) ? 3'b111 : 3'b011;
							assign node141 = (inp[2]) ? node143 : 3'b011;
								assign node143 = (inp[8]) ? 3'b111 : node144;
									assign node144 = (inp[1]) ? 3'b011 : 3'b111;
					assign node148 = (inp[7]) ? node166 : node149;
						assign node149 = (inp[3]) ? node159 : node150;
							assign node150 = (inp[2]) ? node154 : node151;
								assign node151 = (inp[4]) ? 3'b001 : 3'b011;
								assign node154 = (inp[1]) ? node156 : 3'b001;
									assign node156 = (inp[8]) ? 3'b110 : 3'b010;
							assign node159 = (inp[11]) ? node163 : node160;
								assign node160 = (inp[5]) ? 3'b001 : 3'b110;
								assign node163 = (inp[1]) ? 3'b010 : 3'b110;
						assign node166 = (inp[11]) ? node168 : 3'b011;
							assign node168 = (inp[5]) ? node174 : node169;
								assign node169 = (inp[1]) ? 3'b101 : node170;
									assign node170 = (inp[3]) ? 3'b011 : 3'b111;
								assign node174 = (inp[1]) ? node176 : 3'b101;
									assign node176 = (inp[2]) ? 3'b001 : 3'b101;
				assign node179 = (inp[10]) ? node219 : node180;
					assign node180 = (inp[7]) ? node198 : node181;
						assign node181 = (inp[8]) ? node191 : node182;
							assign node182 = (inp[11]) ? node184 : 3'b110;
								assign node184 = (inp[2]) ? node188 : node185;
									assign node185 = (inp[1]) ? 3'b010 : 3'b110;
									assign node188 = (inp[1]) ? 3'b100 : 3'b010;
							assign node191 = (inp[1]) ? node195 : node192;
								assign node192 = (inp[11]) ? 3'b001 : 3'b101;
								assign node195 = (inp[2]) ? 3'b110 : 3'b001;
						assign node198 = (inp[1]) ? node204 : node199;
							assign node199 = (inp[8]) ? node201 : 3'b011;
								assign node201 = (inp[2]) ? 3'b011 : 3'b111;
							assign node204 = (inp[5]) ? node212 : node205;
								assign node205 = (inp[3]) ? 3'b110 : node206;
									assign node206 = (inp[11]) ? node208 : 3'b101;
										assign node208 = (inp[8]) ? 3'b101 : 3'b001;
								assign node212 = (inp[8]) ? node214 : 3'b001;
									assign node214 = (inp[3]) ? 3'b101 : node215;
										assign node215 = (inp[2]) ? 3'b001 : 3'b011;
					assign node219 = (inp[1]) ? node235 : node220;
						assign node220 = (inp[7]) ? node228 : node221;
							assign node221 = (inp[11]) ? 3'b100 : node222;
								assign node222 = (inp[2]) ? 3'b100 : node223;
									assign node223 = (inp[8]) ? 3'b110 : 3'b010;
							assign node228 = (inp[5]) ? 3'b001 : node229;
								assign node229 = (inp[8]) ? node231 : 3'b110;
									assign node231 = (inp[11]) ? 3'b101 : 3'b001;
						assign node235 = (inp[7]) ? node243 : node236;
							assign node236 = (inp[8]) ? node238 : 3'b000;
								assign node238 = (inp[2]) ? node240 : 3'b010;
									assign node240 = (inp[11]) ? 3'b000 : 3'b100;
							assign node243 = (inp[8]) ? 3'b110 : node244;
								assign node244 = (inp[5]) ? 3'b010 : node245;
									assign node245 = (inp[2]) ? 3'b100 : 3'b010;
			assign node250 = (inp[0]) ? node326 : node251;
				assign node251 = (inp[10]) ? node293 : node252;
					assign node252 = (inp[7]) ? node270 : node253;
						assign node253 = (inp[5]) ? node261 : node254;
							assign node254 = (inp[3]) ? node258 : node255;
								assign node255 = (inp[2]) ? 3'b010 : 3'b110;
								assign node258 = (inp[11]) ? 3'b100 : 3'b110;
							assign node261 = (inp[1]) ? 3'b100 : node262;
								assign node262 = (inp[4]) ? 3'b010 : node263;
									assign node263 = (inp[11]) ? node265 : 3'b010;
										assign node265 = (inp[8]) ? 3'b010 : 3'b100;
						assign node270 = (inp[1]) ? node284 : node271;
							assign node271 = (inp[2]) ? node275 : node272;
								assign node272 = (inp[3]) ? 3'b001 : 3'b101;
								assign node275 = (inp[8]) ? node277 : 3'b110;
									assign node277 = (inp[4]) ? 3'b101 : node278;
										assign node278 = (inp[5]) ? node280 : 3'b101;
											assign node280 = (inp[11]) ? 3'b101 : 3'b011;
							assign node284 = (inp[8]) ? node288 : node285;
								assign node285 = (inp[11]) ? 3'b010 : 3'b110;
								assign node288 = (inp[11]) ? 3'b110 : node289;
									assign node289 = (inp[2]) ? 3'b001 : 3'b101;
					assign node293 = (inp[7]) ? node301 : node294;
						assign node294 = (inp[11]) ? 3'b000 : node295;
							assign node295 = (inp[4]) ? node297 : 3'b100;
								assign node297 = (inp[3]) ? 3'b100 : 3'b000;
						assign node301 = (inp[8]) ? node313 : node302;
							assign node302 = (inp[2]) ? node310 : node303;
								assign node303 = (inp[11]) ? node307 : node304;
									assign node304 = (inp[1]) ? 3'b010 : 3'b110;
									assign node307 = (inp[1]) ? 3'b100 : 3'b010;
								assign node310 = (inp[1]) ? 3'b000 : 3'b010;
							assign node313 = (inp[3]) ? node321 : node314;
								assign node314 = (inp[11]) ? node318 : node315;
									assign node315 = (inp[1]) ? 3'b010 : 3'b001;
									assign node318 = (inp[2]) ? 3'b100 : 3'b110;
								assign node321 = (inp[5]) ? 3'b110 : node322;
									assign node322 = (inp[4]) ? 3'b010 : 3'b110;
				assign node326 = (inp[7]) ? node336 : node327;
					assign node327 = (inp[2]) ? 3'b000 : node328;
						assign node328 = (inp[1]) ? 3'b000 : node329;
							assign node329 = (inp[3]) ? 3'b000 : node330;
								assign node330 = (inp[11]) ? 3'b000 : 3'b010;
					assign node336 = (inp[5]) ? node350 : node337;
						assign node337 = (inp[1]) ? node347 : node338;
							assign node338 = (inp[2]) ? 3'b100 : node339;
								assign node339 = (inp[11]) ? 3'b110 : node340;
									assign node340 = (inp[3]) ? node342 : 3'b010;
										assign node342 = (inp[10]) ? 3'b100 : 3'b010;
							assign node347 = (inp[11]) ? 3'b000 : 3'b010;
						assign node350 = (inp[3]) ? node356 : node351;
							assign node351 = (inp[8]) ? 3'b100 : node352;
								assign node352 = (inp[10]) ? 3'b000 : 3'b100;
							assign node356 = (inp[11]) ? 3'b000 : 3'b100;

endmodule