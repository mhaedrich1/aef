module dtc_split5_bm80 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node44;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node71;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node106;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node131;
	wire [3-1:0] node135;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node140;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node185;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node205;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node255;
	wire [3-1:0] node257;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node285;
	wire [3-1:0] node287;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node352;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node365;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node383;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node404;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node425;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node433;
	wire [3-1:0] node435;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node445;
	wire [3-1:0] node448;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node466;
	wire [3-1:0] node468;
	wire [3-1:0] node472;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node498;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node509;
	wire [3-1:0] node512;
	wire [3-1:0] node514;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node520;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node543;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node550;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node558;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node571;
	wire [3-1:0] node574;
	wire [3-1:0] node576;
	wire [3-1:0] node579;
	wire [3-1:0] node581;
	wire [3-1:0] node583;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node605;
	wire [3-1:0] node608;
	wire [3-1:0] node611;
	wire [3-1:0] node612;
	wire [3-1:0] node613;
	wire [3-1:0] node617;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node648;
	wire [3-1:0] node650;
	wire [3-1:0] node654;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node660;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node683;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node703;
	wire [3-1:0] node706;
	wire [3-1:0] node708;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node738;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node754;
	wire [3-1:0] node756;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node767;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node782;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node789;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node796;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node804;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node812;
	wire [3-1:0] node814;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node835;
	wire [3-1:0] node837;
	wire [3-1:0] node839;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node855;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node866;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node874;
	wire [3-1:0] node877;
	wire [3-1:0] node880;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node884;
	wire [3-1:0] node889;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node894;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node900;
	wire [3-1:0] node903;
	wire [3-1:0] node905;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node918;
	wire [3-1:0] node919;
	wire [3-1:0] node921;
	wire [3-1:0] node925;
	wire [3-1:0] node927;
	wire [3-1:0] node930;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node939;
	wire [3-1:0] node942;
	wire [3-1:0] node944;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node950;
	wire [3-1:0] node952;
	wire [3-1:0] node953;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node962;
	wire [3-1:0] node965;
	wire [3-1:0] node967;
	wire [3-1:0] node969;
	wire [3-1:0] node970;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node981;
	wire [3-1:0] node984;
	wire [3-1:0] node986;
	wire [3-1:0] node989;
	wire [3-1:0] node990;
	wire [3-1:0] node991;
	wire [3-1:0] node993;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node999;
	wire [3-1:0] node1002;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1013;
	wire [3-1:0] node1015;
	wire [3-1:0] node1018;
	wire [3-1:0] node1019;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1026;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1033;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1040;
	wire [3-1:0] node1043;
	wire [3-1:0] node1045;
	wire [3-1:0] node1048;
	wire [3-1:0] node1049;
	wire [3-1:0] node1050;
	wire [3-1:0] node1055;
	wire [3-1:0] node1056;
	wire [3-1:0] node1057;
	wire [3-1:0] node1058;
	wire [3-1:0] node1059;
	wire [3-1:0] node1060;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1063;
	wire [3-1:0] node1066;
	wire [3-1:0] node1070;
	wire [3-1:0] node1072;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1079;
	wire [3-1:0] node1081;
	wire [3-1:0] node1082;
	wire [3-1:0] node1086;
	wire [3-1:0] node1087;
	wire [3-1:0] node1088;
	wire [3-1:0] node1092;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1095;
	wire [3-1:0] node1100;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1107;
	wire [3-1:0] node1108;
	wire [3-1:0] node1109;
	wire [3-1:0] node1110;
	wire [3-1:0] node1112;
	wire [3-1:0] node1115;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1121;
	wire [3-1:0] node1124;
	wire [3-1:0] node1125;
	wire [3-1:0] node1129;
	wire [3-1:0] node1131;
	wire [3-1:0] node1132;
	wire [3-1:0] node1134;
	wire [3-1:0] node1137;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1142;
	wire [3-1:0] node1143;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1154;
	wire [3-1:0] node1157;
	wire [3-1:0] node1158;
	wire [3-1:0] node1159;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1166;
	wire [3-1:0] node1167;
	wire [3-1:0] node1171;
	wire [3-1:0] node1172;
	wire [3-1:0] node1174;
	wire [3-1:0] node1177;
	wire [3-1:0] node1180;
	wire [3-1:0] node1181;
	wire [3-1:0] node1182;
	wire [3-1:0] node1184;
	wire [3-1:0] node1185;
	wire [3-1:0] node1188;
	wire [3-1:0] node1191;
	wire [3-1:0] node1192;
	wire [3-1:0] node1195;
	wire [3-1:0] node1197;
	wire [3-1:0] node1200;
	wire [3-1:0] node1201;
	wire [3-1:0] node1203;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1210;
	wire [3-1:0] node1211;
	wire [3-1:0] node1212;
	wire [3-1:0] node1215;
	wire [3-1:0] node1218;
	wire [3-1:0] node1220;
	wire [3-1:0] node1223;
	wire [3-1:0] node1224;
	wire [3-1:0] node1225;
	wire [3-1:0] node1226;
	wire [3-1:0] node1227;
	wire [3-1:0] node1228;
	wire [3-1:0] node1229;
	wire [3-1:0] node1234;
	wire [3-1:0] node1235;
	wire [3-1:0] node1236;
	wire [3-1:0] node1239;
	wire [3-1:0] node1241;
	wire [3-1:0] node1244;
	wire [3-1:0] node1245;
	wire [3-1:0] node1248;
	wire [3-1:0] node1251;
	wire [3-1:0] node1252;
	wire [3-1:0] node1253;
	wire [3-1:0] node1255;
	wire [3-1:0] node1256;
	wire [3-1:0] node1259;
	wire [3-1:0] node1263;
	wire [3-1:0] node1264;
	wire [3-1:0] node1266;
	wire [3-1:0] node1269;
	wire [3-1:0] node1270;
	wire [3-1:0] node1271;
	wire [3-1:0] node1276;
	wire [3-1:0] node1277;
	wire [3-1:0] node1278;
	wire [3-1:0] node1279;
	wire [3-1:0] node1281;
	wire [3-1:0] node1285;
	wire [3-1:0] node1286;
	wire [3-1:0] node1288;
	wire [3-1:0] node1291;
	wire [3-1:0] node1292;
	wire [3-1:0] node1296;
	wire [3-1:0] node1297;
	wire [3-1:0] node1298;
	wire [3-1:0] node1301;
	wire [3-1:0] node1303;
	wire [3-1:0] node1306;
	wire [3-1:0] node1307;
	wire [3-1:0] node1309;
	wire [3-1:0] node1312;
	wire [3-1:0] node1314;
	wire [3-1:0] node1315;
	wire [3-1:0] node1319;
	wire [3-1:0] node1320;
	wire [3-1:0] node1321;
	wire [3-1:0] node1322;
	wire [3-1:0] node1324;
	wire [3-1:0] node1326;
	wire [3-1:0] node1328;
	wire [3-1:0] node1331;
	wire [3-1:0] node1332;
	wire [3-1:0] node1334;
	wire [3-1:0] node1335;
	wire [3-1:0] node1339;
	wire [3-1:0] node1340;
	wire [3-1:0] node1342;
	wire [3-1:0] node1345;
	wire [3-1:0] node1348;
	wire [3-1:0] node1349;
	wire [3-1:0] node1350;
	wire [3-1:0] node1353;
	wire [3-1:0] node1354;
	wire [3-1:0] node1358;
	wire [3-1:0] node1359;
	wire [3-1:0] node1361;
	wire [3-1:0] node1364;
	wire [3-1:0] node1365;
	wire [3-1:0] node1368;
	wire [3-1:0] node1369;
	wire [3-1:0] node1373;
	wire [3-1:0] node1374;
	wire [3-1:0] node1375;
	wire [3-1:0] node1376;
	wire [3-1:0] node1378;
	wire [3-1:0] node1381;
	wire [3-1:0] node1384;
	wire [3-1:0] node1385;
	wire [3-1:0] node1386;
	wire [3-1:0] node1391;
	wire [3-1:0] node1392;
	wire [3-1:0] node1394;
	wire [3-1:0] node1395;
	wire [3-1:0] node1398;
	wire [3-1:0] node1399;
	wire [3-1:0] node1403;
	wire [3-1:0] node1404;
	wire [3-1:0] node1405;
	wire [3-1:0] node1408;
	wire [3-1:0] node1409;
	wire [3-1:0] node1413;
	wire [3-1:0] node1414;
	wire [3-1:0] node1418;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1421;
	wire [3-1:0] node1422;
	wire [3-1:0] node1423;
	wire [3-1:0] node1424;
	wire [3-1:0] node1426;
	wire [3-1:0] node1427;
	wire [3-1:0] node1431;
	wire [3-1:0] node1432;
	wire [3-1:0] node1433;
	wire [3-1:0] node1437;
	wire [3-1:0] node1438;
	wire [3-1:0] node1439;
	wire [3-1:0] node1443;
	wire [3-1:0] node1446;
	wire [3-1:0] node1447;
	wire [3-1:0] node1449;
	wire [3-1:0] node1451;
	wire [3-1:0] node1452;
	wire [3-1:0] node1455;
	wire [3-1:0] node1458;
	wire [3-1:0] node1459;
	wire [3-1:0] node1462;
	wire [3-1:0] node1463;
	wire [3-1:0] node1466;
	wire [3-1:0] node1469;
	wire [3-1:0] node1470;
	wire [3-1:0] node1471;
	wire [3-1:0] node1472;
	wire [3-1:0] node1473;
	wire [3-1:0] node1477;
	wire [3-1:0] node1480;
	wire [3-1:0] node1482;
	wire [3-1:0] node1485;
	wire [3-1:0] node1486;
	wire [3-1:0] node1487;
	wire [3-1:0] node1491;
	wire [3-1:0] node1494;
	wire [3-1:0] node1495;
	wire [3-1:0] node1496;
	wire [3-1:0] node1497;
	wire [3-1:0] node1498;
	wire [3-1:0] node1499;
	wire [3-1:0] node1502;
	wire [3-1:0] node1503;
	wire [3-1:0] node1506;
	wire [3-1:0] node1509;
	wire [3-1:0] node1510;
	wire [3-1:0] node1514;
	wire [3-1:0] node1515;
	wire [3-1:0] node1518;
	wire [3-1:0] node1520;
	wire [3-1:0] node1522;
	wire [3-1:0] node1525;
	wire [3-1:0] node1526;
	wire [3-1:0] node1527;
	wire [3-1:0] node1530;
	wire [3-1:0] node1533;
	wire [3-1:0] node1534;
	wire [3-1:0] node1536;
	wire [3-1:0] node1537;
	wire [3-1:0] node1541;
	wire [3-1:0] node1544;
	wire [3-1:0] node1545;
	wire [3-1:0] node1546;
	wire [3-1:0] node1547;
	wire [3-1:0] node1548;
	wire [3-1:0] node1549;
	wire [3-1:0] node1555;
	wire [3-1:0] node1556;
	wire [3-1:0] node1557;
	wire [3-1:0] node1558;
	wire [3-1:0] node1562;
	wire [3-1:0] node1566;
	wire [3-1:0] node1567;
	wire [3-1:0] node1568;
	wire [3-1:0] node1569;
	wire [3-1:0] node1572;
	wire [3-1:0] node1575;
	wire [3-1:0] node1576;
	wire [3-1:0] node1581;
	wire [3-1:0] node1582;
	wire [3-1:0] node1583;
	wire [3-1:0] node1584;
	wire [3-1:0] node1586;
	wire [3-1:0] node1587;
	wire [3-1:0] node1591;
	wire [3-1:0] node1592;
	wire [3-1:0] node1593;
	wire [3-1:0] node1594;
	wire [3-1:0] node1599;
	wire [3-1:0] node1600;
	wire [3-1:0] node1603;
	wire [3-1:0] node1605;
	wire [3-1:0] node1608;
	wire [3-1:0] node1609;
	wire [3-1:0] node1610;
	wire [3-1:0] node1611;
	wire [3-1:0] node1612;
	wire [3-1:0] node1617;
	wire [3-1:0] node1618;
	wire [3-1:0] node1621;
	wire [3-1:0] node1623;
	wire [3-1:0] node1626;
	wire [3-1:0] node1627;
	wire [3-1:0] node1628;
	wire [3-1:0] node1629;
	wire [3-1:0] node1633;
	wire [3-1:0] node1635;
	wire [3-1:0] node1638;
	wire [3-1:0] node1639;
	wire [3-1:0] node1641;
	wire [3-1:0] node1645;
	wire [3-1:0] node1646;
	wire [3-1:0] node1647;
	wire [3-1:0] node1648;
	wire [3-1:0] node1650;
	wire [3-1:0] node1651;
	wire [3-1:0] node1652;
	wire [3-1:0] node1656;
	wire [3-1:0] node1659;
	wire [3-1:0] node1662;
	wire [3-1:0] node1663;
	wire [3-1:0] node1664;
	wire [3-1:0] node1665;
	wire [3-1:0] node1666;
	wire [3-1:0] node1670;
	wire [3-1:0] node1673;
	wire [3-1:0] node1674;
	wire [3-1:0] node1677;
	wire [3-1:0] node1678;
	wire [3-1:0] node1682;
	wire [3-1:0] node1683;
	wire [3-1:0] node1684;
	wire [3-1:0] node1686;
	wire [3-1:0] node1689;
	wire [3-1:0] node1691;
	wire [3-1:0] node1694;
	wire [3-1:0] node1695;
	wire [3-1:0] node1699;
	wire [3-1:0] node1700;
	wire [3-1:0] node1701;
	wire [3-1:0] node1703;
	wire [3-1:0] node1705;
	wire [3-1:0] node1708;
	wire [3-1:0] node1710;
	wire [3-1:0] node1712;
	wire [3-1:0] node1715;
	wire [3-1:0] node1716;
	wire [3-1:0] node1718;
	wire [3-1:0] node1721;
	wire [3-1:0] node1722;
	wire [3-1:0] node1724;
	wire [3-1:0] node1727;
	wire [3-1:0] node1728;
	wire [3-1:0] node1731;
	wire [3-1:0] node1732;
	wire [3-1:0] node1736;
	wire [3-1:0] node1737;
	wire [3-1:0] node1738;
	wire [3-1:0] node1739;
	wire [3-1:0] node1740;
	wire [3-1:0] node1741;
	wire [3-1:0] node1742;
	wire [3-1:0] node1744;
	wire [3-1:0] node1747;
	wire [3-1:0] node1748;
	wire [3-1:0] node1752;
	wire [3-1:0] node1753;
	wire [3-1:0] node1755;
	wire [3-1:0] node1758;
	wire [3-1:0] node1759;
	wire [3-1:0] node1763;
	wire [3-1:0] node1764;
	wire [3-1:0] node1765;
	wire [3-1:0] node1766;
	wire [3-1:0] node1767;
	wire [3-1:0] node1772;
	wire [3-1:0] node1773;
	wire [3-1:0] node1777;
	wire [3-1:0] node1779;
	wire [3-1:0] node1782;
	wire [3-1:0] node1783;
	wire [3-1:0] node1784;
	wire [3-1:0] node1785;
	wire [3-1:0] node1786;
	wire [3-1:0] node1790;
	wire [3-1:0] node1793;
	wire [3-1:0] node1794;
	wire [3-1:0] node1797;
	wire [3-1:0] node1800;
	wire [3-1:0] node1801;
	wire [3-1:0] node1802;
	wire [3-1:0] node1803;
	wire [3-1:0] node1807;
	wire [3-1:0] node1810;
	wire [3-1:0] node1811;
	wire [3-1:0] node1812;
	wire [3-1:0] node1814;
	wire [3-1:0] node1819;
	wire [3-1:0] node1820;
	wire [3-1:0] node1821;
	wire [3-1:0] node1822;
	wire [3-1:0] node1824;
	wire [3-1:0] node1826;
	wire [3-1:0] node1827;
	wire [3-1:0] node1830;
	wire [3-1:0] node1833;
	wire [3-1:0] node1834;
	wire [3-1:0] node1836;
	wire [3-1:0] node1839;
	wire [3-1:0] node1842;
	wire [3-1:0] node1843;
	wire [3-1:0] node1844;
	wire [3-1:0] node1845;
	wire [3-1:0] node1848;
	wire [3-1:0] node1851;
	wire [3-1:0] node1852;
	wire [3-1:0] node1854;
	wire [3-1:0] node1858;
	wire [3-1:0] node1859;
	wire [3-1:0] node1860;
	wire [3-1:0] node1862;
	wire [3-1:0] node1867;
	wire [3-1:0] node1868;
	wire [3-1:0] node1869;
	wire [3-1:0] node1870;
	wire [3-1:0] node1872;
	wire [3-1:0] node1874;
	wire [3-1:0] node1877;
	wire [3-1:0] node1878;
	wire [3-1:0] node1882;
	wire [3-1:0] node1883;
	wire [3-1:0] node1885;
	wire [3-1:0] node1888;
	wire [3-1:0] node1890;
	wire [3-1:0] node1892;
	wire [3-1:0] node1895;
	wire [3-1:0] node1896;
	wire [3-1:0] node1897;
	wire [3-1:0] node1898;
	wire [3-1:0] node1899;
	wire [3-1:0] node1905;
	wire [3-1:0] node1906;
	wire [3-1:0] node1908;
	wire [3-1:0] node1911;
	wire [3-1:0] node1912;
	wire [3-1:0] node1916;
	wire [3-1:0] node1917;
	wire [3-1:0] node1918;
	wire [3-1:0] node1919;
	wire [3-1:0] node1920;
	wire [3-1:0] node1921;
	wire [3-1:0] node1922;
	wire [3-1:0] node1924;
	wire [3-1:0] node1928;
	wire [3-1:0] node1931;
	wire [3-1:0] node1933;
	wire [3-1:0] node1934;
	wire [3-1:0] node1938;
	wire [3-1:0] node1939;
	wire [3-1:0] node1940;
	wire [3-1:0] node1941;
	wire [3-1:0] node1944;
	wire [3-1:0] node1949;
	wire [3-1:0] node1950;
	wire [3-1:0] node1951;
	wire [3-1:0] node1952;
	wire [3-1:0] node1953;
	wire [3-1:0] node1957;
	wire [3-1:0] node1958;
	wire [3-1:0] node1962;
	wire [3-1:0] node1963;
	wire [3-1:0] node1965;
	wire [3-1:0] node1969;
	wire [3-1:0] node1970;
	wire [3-1:0] node1972;
	wire [3-1:0] node1975;
	wire [3-1:0] node1976;
	wire [3-1:0] node1979;
	wire [3-1:0] node1980;
	wire [3-1:0] node1984;
	wire [3-1:0] node1986;
	wire [3-1:0] node1987;
	wire [3-1:0] node1988;
	wire [3-1:0] node1989;
	wire [3-1:0] node1991;
	wire [3-1:0] node1994;
	wire [3-1:0] node1995;
	wire [3-1:0] node1999;
	wire [3-1:0] node2000;
	wire [3-1:0] node2001;
	wire [3-1:0] node2006;
	wire [3-1:0] node2007;
	wire [3-1:0] node2008;
	wire [3-1:0] node2009;

	assign outp = (inp[6]) ? node824 : node1;
		assign node1 = (inp[3]) ? node627 : node2;
			assign node2 = (inp[9]) ? node326 : node3;
				assign node3 = (inp[7]) ? node173 : node4;
					assign node4 = (inp[4]) ? node98 : node5;
						assign node5 = (inp[0]) ? node47 : node6;
							assign node6 = (inp[8]) ? node24 : node7;
								assign node7 = (inp[11]) ? node19 : node8;
									assign node8 = (inp[5]) ? node12 : node9;
										assign node9 = (inp[10]) ? 3'b110 : 3'b011;
										assign node12 = (inp[1]) ? node16 : node13;
											assign node13 = (inp[10]) ? 3'b001 : 3'b101;
											assign node16 = (inp[10]) ? 3'b110 : 3'b001;
									assign node19 = (inp[10]) ? 3'b110 : node20;
										assign node20 = (inp[2]) ? 3'b001 : 3'b110;
								assign node24 = (inp[10]) ? node36 : node25;
									assign node25 = (inp[1]) ? node29 : node26;
										assign node26 = (inp[2]) ? 3'b001 : 3'b011;
										assign node29 = (inp[11]) ? node33 : node30;
											assign node30 = (inp[5]) ? 3'b101 : 3'b011;
											assign node33 = (inp[5]) ? 3'b001 : 3'b101;
									assign node36 = (inp[1]) ? node38 : 3'b101;
										assign node38 = (inp[2]) ? node44 : node39;
											assign node39 = (inp[11]) ? 3'b001 : node40;
												assign node40 = (inp[5]) ? 3'b001 : 3'b101;
											assign node44 = (inp[5]) ? 3'b110 : 3'b001;
							assign node47 = (inp[10]) ? node75 : node48;
								assign node48 = (inp[8]) ? node64 : node49;
									assign node49 = (inp[2]) ? node57 : node50;
										assign node50 = (inp[5]) ? 3'b110 : node51;
											assign node51 = (inp[11]) ? node53 : 3'b001;
												assign node53 = (inp[1]) ? 3'b000 : 3'b010;
										assign node57 = (inp[11]) ? node59 : 3'b110;
											assign node59 = (inp[1]) ? 3'b010 : node60;
												assign node60 = (inp[5]) ? 3'b010 : 3'b110;
									assign node64 = (inp[1]) ? 3'b110 : node65;
										assign node65 = (inp[11]) ? node71 : node66;
											assign node66 = (inp[5]) ? 3'b001 : node67;
												assign node67 = (inp[2]) ? 3'b001 : 3'b101;
											assign node71 = (inp[2]) ? 3'b001 : 3'b000;
								assign node75 = (inp[11]) ? node89 : node76;
									assign node76 = (inp[2]) ? node84 : node77;
										assign node77 = (inp[8]) ? node79 : 3'b110;
											assign node79 = (inp[5]) ? 3'b110 : node80;
												assign node80 = (inp[1]) ? 3'b110 : 3'b010;
										assign node84 = (inp[1]) ? 3'b010 : node85;
											assign node85 = (inp[5]) ? 3'b010 : 3'b110;
									assign node89 = (inp[1]) ? 3'b100 : node90;
										assign node90 = (inp[5]) ? node92 : 3'b110;
											assign node92 = (inp[2]) ? 3'b100 : node93;
												assign node93 = (inp[8]) ? 3'b010 : 3'b000;
						assign node98 = (inp[0]) ? node144 : node99;
							assign node99 = (inp[8]) ? node121 : node100;
								assign node100 = (inp[2]) ? node116 : node101;
									assign node101 = (inp[1]) ? node109 : node102;
										assign node102 = (inp[11]) ? node106 : node103;
											assign node103 = (inp[5]) ? 3'b110 : 3'b100;
											assign node106 = (inp[10]) ? 3'b110 : 3'b010;
										assign node109 = (inp[10]) ? node111 : 3'b010;
											assign node111 = (inp[11]) ? 3'b100 : node112;
												assign node112 = (inp[5]) ? 3'b000 : 3'b010;
									assign node116 = (inp[1]) ? 3'b010 : node117;
										assign node117 = (inp[11]) ? 3'b010 : 3'b000;
								assign node121 = (inp[1]) ? node135 : node122;
									assign node122 = (inp[10]) ? node128 : node123;
										assign node123 = (inp[2]) ? 3'b010 : node124;
											assign node124 = (inp[5]) ? 3'b000 : 3'b100;
										assign node128 = (inp[5]) ? 3'b110 : node129;
											assign node129 = (inp[2]) ? node131 : 3'b000;
												assign node131 = (inp[11]) ? 3'b110 : 3'b000;
									assign node135 = (inp[10]) ? node137 : 3'b110;
										assign node137 = (inp[5]) ? 3'b010 : node138;
											assign node138 = (inp[2]) ? node140 : 3'b110;
												assign node140 = (inp[11]) ? 3'b010 : 3'b110;
							assign node144 = (inp[1]) ? node162 : node145;
								assign node145 = (inp[10]) ? node151 : node146;
									assign node146 = (inp[5]) ? 3'b010 : node147;
										assign node147 = (inp[8]) ? 3'b110 : 3'b010;
									assign node151 = (inp[8]) ? node157 : node152;
										assign node152 = (inp[2]) ? node154 : 3'b100;
											assign node154 = (inp[5]) ? 3'b000 : 3'b100;
										assign node157 = (inp[11]) ? node159 : 3'b010;
											assign node159 = (inp[5]) ? 3'b100 : 3'b000;
								assign node162 = (inp[10]) ? 3'b000 : node163;
									assign node163 = (inp[5]) ? node165 : 3'b100;
										assign node165 = (inp[11]) ? 3'b000 : node166;
											assign node166 = (inp[2]) ? 3'b100 : node167;
												assign node167 = (inp[8]) ? 3'b000 : 3'b100;
					assign node173 = (inp[0]) ? node249 : node174;
						assign node174 = (inp[4]) ? node208 : node175;
							assign node175 = (inp[1]) ? node189 : node176;
								assign node176 = (inp[2]) ? 3'b001 : node177;
									assign node177 = (inp[5]) ? node183 : node178;
										assign node178 = (inp[8]) ? node180 : 3'b001;
											assign node180 = (inp[10]) ? 3'b001 : 3'b000;
										assign node183 = (inp[10]) ? node185 : 3'b001;
											assign node185 = (inp[8]) ? 3'b001 : 3'b000;
								assign node189 = (inp[10]) ? node201 : node190;
									assign node190 = (inp[8]) ? node198 : node191;
										assign node191 = (inp[5]) ? 3'b101 : node192;
											assign node192 = (inp[11]) ? 3'b001 : node193;
												assign node193 = (inp[2]) ? 3'b011 : 3'b111;
										assign node198 = (inp[5]) ? 3'b011 : 3'b111;
									assign node201 = (inp[5]) ? node203 : 3'b001;
										assign node203 = (inp[2]) ? node205 : 3'b101;
											assign node205 = (inp[8]) ? 3'b101 : 3'b001;
							assign node208 = (inp[1]) ? node234 : node209;
								assign node209 = (inp[10]) ? node223 : node210;
									assign node210 = (inp[11]) ? node218 : node211;
										assign node211 = (inp[5]) ? node215 : node212;
											assign node212 = (inp[8]) ? 3'b011 : 3'b111;
											assign node215 = (inp[2]) ? 3'b101 : 3'b111;
										assign node218 = (inp[2]) ? 3'b101 : node219;
											assign node219 = (inp[8]) ? 3'b011 : 3'b001;
									assign node223 = (inp[11]) ? node229 : node224;
										assign node224 = (inp[8]) ? node226 : 3'b001;
											assign node226 = (inp[2]) ? 3'b101 : 3'b001;
										assign node229 = (inp[5]) ? 3'b110 : node230;
											assign node230 = (inp[8]) ? 3'b101 : 3'b001;
								assign node234 = (inp[10]) ? node240 : node235;
									assign node235 = (inp[2]) ? node237 : 3'b001;
										assign node237 = (inp[8]) ? 3'b101 : 3'b001;
									assign node240 = (inp[8]) ? node244 : node241;
										assign node241 = (inp[5]) ? 3'b010 : 3'b110;
										assign node244 = (inp[5]) ? 3'b110 : node245;
											assign node245 = (inp[2]) ? 3'b001 : 3'b101;
						assign node249 = (inp[10]) ? node295 : node250;
							assign node250 = (inp[4]) ? node280 : node251;
								assign node251 = (inp[11]) ? node267 : node252;
									assign node252 = (inp[1]) ? node260 : node253;
										assign node253 = (inp[2]) ? node255 : 3'b001;
											assign node255 = (inp[8]) ? node257 : 3'b101;
												assign node257 = (inp[5]) ? 3'b101 : 3'b011;
										assign node260 = (inp[8]) ? node264 : node261;
											assign node261 = (inp[5]) ? 3'b110 : 3'b101;
											assign node264 = (inp[5]) ? 3'b001 : 3'b101;
									assign node267 = (inp[8]) ? node269 : 3'b001;
										assign node269 = (inp[1]) ? node275 : node270;
											assign node270 = (inp[5]) ? 3'b101 : node271;
												assign node271 = (inp[2]) ? 3'b101 : 3'b010;
											assign node275 = (inp[2]) ? 3'b001 : node276;
												assign node276 = (inp[5]) ? 3'b001 : 3'b101;
								assign node280 = (inp[11]) ? node290 : node281;
									assign node281 = (inp[1]) ? node285 : node282;
										assign node282 = (inp[2]) ? 3'b001 : 3'b101;
										assign node285 = (inp[5]) ? node287 : 3'b111;
											assign node287 = (inp[8]) ? 3'b110 : 3'b010;
									assign node290 = (inp[5]) ? 3'b010 : node291;
										assign node291 = (inp[2]) ? 3'b010 : 3'b100;
							assign node295 = (inp[4]) ? node311 : node296;
								assign node296 = (inp[1]) ? node306 : node297;
									assign node297 = (inp[8]) ? node301 : node298;
										assign node298 = (inp[5]) ? 3'b110 : 3'b001;
										assign node301 = (inp[11]) ? 3'b001 : node302;
											assign node302 = (inp[5]) ? 3'b001 : 3'b101;
									assign node306 = (inp[5]) ? 3'b110 : node307;
										assign node307 = (inp[11]) ? 3'b110 : 3'b001;
								assign node311 = (inp[11]) ? node315 : node312;
									assign node312 = (inp[5]) ? 3'b010 : 3'b110;
									assign node315 = (inp[5]) ? node321 : node316;
										assign node316 = (inp[2]) ? node318 : 3'b010;
											assign node318 = (inp[8]) ? 3'b010 : 3'b100;
										assign node321 = (inp[1]) ? node323 : 3'b000;
											assign node323 = (inp[2]) ? 3'b000 : 3'b100;
				assign node326 = (inp[4]) ? node502 : node327;
					assign node327 = (inp[7]) ? node409 : node328;
						assign node328 = (inp[11]) ? node356 : node329;
							assign node329 = (inp[10]) ? node341 : node330;
								assign node330 = (inp[1]) ? node336 : node331;
									assign node331 = (inp[8]) ? 3'b010 : node332;
										assign node332 = (inp[5]) ? 3'b100 : 3'b010;
									assign node336 = (inp[0]) ? 3'b100 : node337;
										assign node337 = (inp[5]) ? 3'b010 : 3'b111;
								assign node341 = (inp[1]) ? node349 : node342;
									assign node342 = (inp[8]) ? node346 : node343;
										assign node343 = (inp[5]) ? 3'b000 : 3'b100;
										assign node346 = (inp[5]) ? 3'b100 : 3'b000;
									assign node349 = (inp[0]) ? 3'b000 : node350;
										assign node350 = (inp[5]) ? node352 : 3'b010;
											assign node352 = (inp[2]) ? 3'b100 : 3'b110;
							assign node356 = (inp[0]) ? node386 : node357;
								assign node357 = (inp[10]) ? node379 : node358;
									assign node358 = (inp[8]) ? node370 : node359;
										assign node359 = (inp[5]) ? node365 : node360;
											assign node360 = (inp[1]) ? 3'b010 : node361;
												assign node361 = (inp[2]) ? 3'b100 : 3'b000;
											assign node365 = (inp[2]) ? node367 : 3'b100;
												assign node367 = (inp[1]) ? 3'b100 : 3'b000;
										assign node370 = (inp[2]) ? node372 : 3'b000;
											assign node372 = (inp[1]) ? node376 : node373;
												assign node373 = (inp[5]) ? 3'b100 : 3'b010;
												assign node376 = (inp[5]) ? 3'b010 : 3'b110;
									assign node379 = (inp[2]) ? node381 : 3'b100;
										assign node381 = (inp[5]) ? node383 : 3'b100;
											assign node383 = (inp[1]) ? 3'b100 : 3'b000;
								assign node386 = (inp[1]) ? node400 : node387;
									assign node387 = (inp[5]) ? node389 : 3'b100;
										assign node389 = (inp[8]) ? node395 : node390;
											assign node390 = (inp[2]) ? 3'b000 : node391;
												assign node391 = (inp[10]) ? 3'b000 : 3'b100;
											assign node395 = (inp[10]) ? 3'b100 : node396;
												assign node396 = (inp[2]) ? 3'b100 : 3'b000;
									assign node400 = (inp[5]) ? 3'b000 : node401;
										assign node401 = (inp[10]) ? 3'b000 : node402;
											assign node402 = (inp[2]) ? node404 : 3'b000;
												assign node404 = (inp[8]) ? 3'b100 : 3'b000;
						assign node409 = (inp[0]) ? node461 : node410;
							assign node410 = (inp[1]) ? node438 : node411;
								assign node411 = (inp[8]) ? node425 : node412;
									assign node412 = (inp[10]) ? node420 : node413;
										assign node413 = (inp[5]) ? 3'b000 : node414;
											assign node414 = (inp[11]) ? 3'b000 : node415;
												assign node415 = (inp[2]) ? 3'b101 : 3'b001;
										assign node420 = (inp[11]) ? 3'b100 : node421;
											assign node421 = (inp[5]) ? 3'b100 : 3'b000;
									assign node425 = (inp[11]) ? node427 : 3'b101;
										assign node427 = (inp[10]) ? node433 : node428;
											assign node428 = (inp[2]) ? 3'b101 : node429;
												assign node429 = (inp[5]) ? 3'b101 : 3'b100;
											assign node433 = (inp[5]) ? node435 : 3'b001;
												assign node435 = (inp[2]) ? 3'b100 : 3'b000;
								assign node438 = (inp[10]) ? node448 : node439;
									assign node439 = (inp[8]) ? node445 : node440;
										assign node440 = (inp[11]) ? 3'b110 : node441;
											assign node441 = (inp[2]) ? 3'b110 : 3'b101;
										assign node445 = (inp[2]) ? 3'b001 : 3'b101;
									assign node448 = (inp[11]) ? node450 : 3'b110;
										assign node450 = (inp[8]) ? node456 : node451;
											assign node451 = (inp[5]) ? 3'b010 : node452;
												assign node452 = (inp[2]) ? 3'b010 : 3'b110;
											assign node456 = (inp[5]) ? 3'b110 : node457;
												assign node457 = (inp[2]) ? 3'b110 : 3'b001;
							assign node461 = (inp[10]) ? node481 : node462;
								assign node462 = (inp[2]) ? node472 : node463;
									assign node463 = (inp[11]) ? 3'b010 : node464;
										assign node464 = (inp[8]) ? node466 : 3'b100;
											assign node466 = (inp[1]) ? node468 : 3'b000;
												assign node468 = (inp[5]) ? 3'b010 : 3'b110;
									assign node472 = (inp[1]) ? node474 : 3'b110;
										assign node474 = (inp[5]) ? node478 : node475;
											assign node475 = (inp[8]) ? 3'b110 : 3'b010;
											assign node478 = (inp[8]) ? 3'b010 : 3'b100;
								assign node481 = (inp[1]) ? node491 : node482;
									assign node482 = (inp[11]) ? node486 : node483;
										assign node483 = (inp[2]) ? 3'b100 : 3'b000;
										assign node486 = (inp[5]) ? 3'b010 : node487;
											assign node487 = (inp[8]) ? 3'b110 : 3'b010;
									assign node491 = (inp[11]) ? node495 : node492;
										assign node492 = (inp[5]) ? 3'b100 : 3'b010;
										assign node495 = (inp[5]) ? 3'b000 : node496;
											assign node496 = (inp[8]) ? node498 : 3'b100;
												assign node498 = (inp[2]) ? 3'b100 : 3'b000;
					assign node502 = (inp[0]) ? node586 : node503;
						assign node503 = (inp[10]) ? node553 : node504;
							assign node504 = (inp[11]) ? node528 : node505;
								assign node505 = (inp[5]) ? node517 : node506;
									assign node506 = (inp[2]) ? node512 : node507;
										assign node507 = (inp[1]) ? node509 : 3'b010;
											assign node509 = (inp[8]) ? 3'b001 : 3'b011;
										assign node512 = (inp[8]) ? node514 : 3'b010;
											assign node514 = (inp[7]) ? 3'b110 : 3'b010;
									assign node517 = (inp[7]) ? node523 : node518;
										assign node518 = (inp[1]) ? node520 : 3'b010;
											assign node520 = (inp[8]) ? 3'b100 : 3'b000;
										assign node523 = (inp[1]) ? 3'b010 : node524;
											assign node524 = (inp[8]) ? 3'b010 : 3'b100;
								assign node528 = (inp[1]) ? node538 : node529;
									assign node529 = (inp[7]) ? node531 : 3'b010;
										assign node531 = (inp[8]) ? node535 : node532;
											assign node532 = (inp[5]) ? 3'b000 : 3'b100;
											assign node535 = (inp[5]) ? 3'b100 : 3'b010;
									assign node538 = (inp[7]) ? node546 : node539;
										assign node539 = (inp[5]) ? node543 : node540;
											assign node540 = (inp[8]) ? 3'b000 : 3'b100;
											assign node543 = (inp[8]) ? 3'b100 : 3'b000;
										assign node546 = (inp[8]) ? node550 : node547;
											assign node547 = (inp[5]) ? 3'b100 : 3'b110;
											assign node550 = (inp[5]) ? 3'b010 : 3'b110;
							assign node553 = (inp[1]) ? node565 : node554;
								assign node554 = (inp[5]) ? node558 : node555;
									assign node555 = (inp[7]) ? 3'b000 : 3'b010;
									assign node558 = (inp[8]) ? node560 : 3'b000;
										assign node560 = (inp[11]) ? 3'b000 : node561;
											assign node561 = (inp[7]) ? 3'b100 : 3'b000;
								assign node565 = (inp[5]) ? node579 : node566;
									assign node566 = (inp[2]) ? node574 : node567;
										assign node567 = (inp[8]) ? node571 : node568;
											assign node568 = (inp[11]) ? 3'b000 : 3'b100;
											assign node571 = (inp[7]) ? 3'b110 : 3'b100;
										assign node574 = (inp[8]) ? node576 : 3'b100;
											assign node576 = (inp[7]) ? 3'b000 : 3'b100;
									assign node579 = (inp[7]) ? node581 : 3'b000;
										assign node581 = (inp[11]) ? node583 : 3'b010;
											assign node583 = (inp[2]) ? 3'b000 : 3'b100;
						assign node586 = (inp[7]) ? node598 : node587;
							assign node587 = (inp[2]) ? node589 : 3'b000;
								assign node589 = (inp[10]) ? 3'b000 : node590;
									assign node590 = (inp[8]) ? node592 : 3'b000;
										assign node592 = (inp[5]) ? 3'b000 : node593;
											assign node593 = (inp[11]) ? 3'b000 : 3'b100;
							assign node598 = (inp[10]) ? node622 : node599;
								assign node599 = (inp[1]) ? node611 : node600;
									assign node600 = (inp[2]) ? node608 : node601;
										assign node601 = (inp[11]) ? node605 : node602;
											assign node602 = (inp[5]) ? 3'b100 : 3'b010;
											assign node605 = (inp[5]) ? 3'b000 : 3'b100;
										assign node608 = (inp[5]) ? 3'b110 : 3'b010;
									assign node611 = (inp[8]) ? node617 : node612;
										assign node612 = (inp[11]) ? 3'b000 : node613;
											assign node613 = (inp[5]) ? 3'b000 : 3'b100;
										assign node617 = (inp[5]) ? node619 : 3'b100;
											assign node619 = (inp[11]) ? 3'b000 : 3'b100;
								assign node622 = (inp[1]) ? 3'b000 : node623;
									assign node623 = (inp[11]) ? 3'b000 : 3'b100;
			assign node627 = (inp[9]) ? node789 : node628;
				assign node628 = (inp[4]) ? node748 : node629;
					assign node629 = (inp[7]) ? node669 : node630;
						assign node630 = (inp[11]) ? node654 : node631;
							assign node631 = (inp[10]) ? node645 : node632;
								assign node632 = (inp[1]) ? node638 : node633;
									assign node633 = (inp[8]) ? 3'b100 : node634;
										assign node634 = (inp[5]) ? 3'b000 : 3'b100;
									assign node638 = (inp[0]) ? 3'b000 : node639;
										assign node639 = (inp[5]) ? 3'b100 : node640;
											assign node640 = (inp[8]) ? 3'b110 : 3'b010;
								assign node645 = (inp[0]) ? 3'b000 : node646;
									assign node646 = (inp[1]) ? node648 : 3'b000;
										assign node648 = (inp[5]) ? node650 : 3'b100;
											assign node650 = (inp[8]) ? 3'b100 : 3'b000;
							assign node654 = (inp[1]) ? node656 : 3'b000;
								assign node656 = (inp[0]) ? 3'b000 : node657;
									assign node657 = (inp[5]) ? node663 : node658;
										assign node658 = (inp[10]) ? node660 : 3'b100;
											assign node660 = (inp[8]) ? 3'b100 : 3'b000;
										assign node663 = (inp[10]) ? 3'b000 : node664;
											assign node664 = (inp[2]) ? 3'b100 : 3'b000;
						assign node669 = (inp[0]) ? node711 : node670;
							assign node670 = (inp[5]) ? node692 : node671;
								assign node671 = (inp[11]) ? node681 : node672;
									assign node672 = (inp[1]) ? node678 : node673;
										assign node673 = (inp[10]) ? node675 : 3'b100;
											assign node675 = (inp[2]) ? 3'b110 : 3'b000;
										assign node678 = (inp[8]) ? 3'b001 : 3'b010;
									assign node681 = (inp[10]) ? node687 : node682;
										assign node682 = (inp[8]) ? 3'b110 : node683;
											assign node683 = (inp[2]) ? 3'b010 : 3'b000;
										assign node687 = (inp[8]) ? 3'b010 : node688;
											assign node688 = (inp[2]) ? 3'b100 : 3'b110;
								assign node692 = (inp[8]) ? node698 : node693;
									assign node693 = (inp[10]) ? 3'b010 : node694;
										assign node694 = (inp[1]) ? 3'b010 : 3'b110;
									assign node698 = (inp[11]) ? node706 : node699;
										assign node699 = (inp[1]) ? node703 : node700;
											assign node700 = (inp[10]) ? 3'b110 : 3'b000;
											assign node703 = (inp[10]) ? 3'b010 : 3'b110;
										assign node706 = (inp[10]) ? node708 : 3'b110;
											assign node708 = (inp[1]) ? 3'b100 : 3'b110;
							assign node711 = (inp[10]) ? node735 : node712;
								assign node712 = (inp[1]) ? node718 : node713;
									assign node713 = (inp[8]) ? 3'b010 : node714;
										assign node714 = (inp[2]) ? 3'b010 : 3'b110;
									assign node718 = (inp[8]) ? node730 : node719;
										assign node719 = (inp[5]) ? node725 : node720;
											assign node720 = (inp[11]) ? 3'b100 : node721;
												assign node721 = (inp[2]) ? 3'b100 : 3'b000;
											assign node725 = (inp[11]) ? 3'b000 : node726;
												assign node726 = (inp[2]) ? 3'b000 : 3'b100;
										assign node730 = (inp[2]) ? 3'b100 : node731;
											assign node731 = (inp[11]) ? 3'b100 : 3'b010;
								assign node735 = (inp[5]) ? node741 : node736;
									assign node736 = (inp[11]) ? node738 : 3'b100;
										assign node738 = (inp[2]) ? 3'b100 : 3'b000;
									assign node741 = (inp[8]) ? 3'b100 : node742;
										assign node742 = (inp[2]) ? 3'b000 : node743;
											assign node743 = (inp[1]) ? 3'b000 : 3'b100;
					assign node748 = (inp[7]) ? node762 : node749;
						assign node749 = (inp[0]) ? 3'b000 : node750;
							assign node750 = (inp[5]) ? 3'b000 : node751;
								assign node751 = (inp[10]) ? 3'b000 : node752;
									assign node752 = (inp[1]) ? node754 : 3'b000;
										assign node754 = (inp[8]) ? node756 : 3'b000;
											assign node756 = (inp[2]) ? 3'b100 : 3'b000;
						assign node762 = (inp[10]) ? node782 : node763;
							assign node763 = (inp[1]) ? node771 : node764;
								assign node764 = (inp[8]) ? 3'b100 : node765;
									assign node765 = (inp[2]) ? node767 : 3'b000;
										assign node767 = (inp[0]) ? 3'b100 : 3'b000;
								assign node771 = (inp[0]) ? 3'b000 : node772;
									assign node772 = (inp[11]) ? node776 : node773;
										assign node773 = (inp[2]) ? 3'b010 : 3'b110;
										assign node776 = (inp[5]) ? 3'b000 : node777;
											assign node777 = (inp[2]) ? 3'b010 : 3'b000;
							assign node782 = (inp[1]) ? node784 : 3'b000;
								assign node784 = (inp[0]) ? 3'b000 : node785;
									assign node785 = (inp[8]) ? 3'b100 : 3'b000;
				assign node789 = (inp[7]) ? node791 : 3'b000;
					assign node791 = (inp[0]) ? 3'b000 : node792;
						assign node792 = (inp[4]) ? 3'b000 : node793;
							assign node793 = (inp[1]) ? node799 : node794;
								assign node794 = (inp[10]) ? node796 : 3'b010;
									assign node796 = (inp[5]) ? 3'b000 : 3'b010;
								assign node799 = (inp[10]) ? node817 : node800;
									assign node800 = (inp[2]) ? node808 : node801;
										assign node801 = (inp[11]) ? 3'b100 : node802;
											assign node802 = (inp[8]) ? node804 : 3'b100;
												assign node804 = (inp[5]) ? 3'b100 : 3'b000;
										assign node808 = (inp[5]) ? node812 : node809;
											assign node809 = (inp[11]) ? 3'b100 : 3'b010;
											assign node812 = (inp[8]) ? node814 : 3'b000;
												assign node814 = (inp[11]) ? 3'b000 : 3'b100;
									assign node817 = (inp[11]) ? 3'b000 : node818;
										assign node818 = (inp[8]) ? 3'b100 : 3'b000;
		assign node824 = (inp[3]) ? node1418 : node825;
			assign node825 = (inp[9]) ? node1055 : node826;
				assign node826 = (inp[0]) ? node908 : node827;
					assign node827 = (inp[1]) ? node843 : node828;
						assign node828 = (inp[7]) ? 3'b111 : node829;
							assign node829 = (inp[4]) ? node831 : 3'b111;
								assign node831 = (inp[2]) ? node835 : node832;
									assign node832 = (inp[10]) ? 3'b011 : 3'b111;
									assign node835 = (inp[8]) ? node837 : 3'b111;
										assign node837 = (inp[5]) ? node839 : 3'b111;
											assign node839 = (inp[11]) ? 3'b011 : 3'b111;
						assign node843 = (inp[7]) ? node889 : node844;
							assign node844 = (inp[4]) ? node870 : node845;
								assign node845 = (inp[10]) ? node859 : node846;
									assign node846 = (inp[5]) ? node852 : node847;
										assign node847 = (inp[11]) ? 3'b011 : node848;
											assign node848 = (inp[8]) ? 3'b011 : 3'b111;
										assign node852 = (inp[11]) ? 3'b111 : node853;
											assign node853 = (inp[8]) ? node855 : 3'b111;
												assign node855 = (inp[2]) ? 3'b111 : 3'b011;
									assign node859 = (inp[5]) ? node863 : node860;
										assign node860 = (inp[8]) ? 3'b111 : 3'b011;
										assign node863 = (inp[8]) ? 3'b011 : node864;
											assign node864 = (inp[11]) ? node866 : 3'b011;
												assign node866 = (inp[2]) ? 3'b110 : 3'b010;
								assign node870 = (inp[10]) ? node880 : node871;
									assign node871 = (inp[5]) ? node877 : node872;
										assign node872 = (inp[8]) ? node874 : 3'b011;
											assign node874 = (inp[2]) ? 3'b111 : 3'b011;
										assign node877 = (inp[8]) ? 3'b011 : 3'b101;
									assign node880 = (inp[8]) ? 3'b101 : node881;
										assign node881 = (inp[11]) ? 3'b001 : node882;
											assign node882 = (inp[2]) ? node884 : 3'b101;
												assign node884 = (inp[5]) ? 3'b001 : 3'b101;
							assign node889 = (inp[4]) ? node891 : 3'b111;
								assign node891 = (inp[10]) ? node897 : node892;
									assign node892 = (inp[11]) ? node894 : 3'b111;
										assign node894 = (inp[8]) ? 3'b111 : 3'b101;
									assign node897 = (inp[8]) ? node903 : node898;
										assign node898 = (inp[11]) ? node900 : 3'b011;
											assign node900 = (inp[5]) ? 3'b101 : 3'b011;
										assign node903 = (inp[5]) ? node905 : 3'b111;
											assign node905 = (inp[2]) ? 3'b011 : 3'b111;
					assign node908 = (inp[4]) ? node974 : node909;
						assign node909 = (inp[7]) ? node947 : node910;
							assign node910 = (inp[5]) ? node930 : node911;
								assign node911 = (inp[11]) ? node925 : node912;
									assign node912 = (inp[10]) ? node918 : node913;
										assign node913 = (inp[2]) ? 3'b011 : node914;
											assign node914 = (inp[8]) ? 3'b111 : 3'b011;
										assign node918 = (inp[1]) ? 3'b101 : node919;
											assign node919 = (inp[8]) ? node921 : 3'b111;
												assign node921 = (inp[2]) ? 3'b011 : 3'b111;
									assign node925 = (inp[8]) ? node927 : 3'b101;
										assign node927 = (inp[2]) ? 3'b011 : 3'b111;
								assign node930 = (inp[2]) ? node932 : 3'b101;
									assign node932 = (inp[8]) ? node942 : node933;
										assign node933 = (inp[1]) ? node935 : 3'b011;
											assign node935 = (inp[10]) ? node939 : node936;
												assign node936 = (inp[11]) ? 3'b001 : 3'b101;
												assign node939 = (inp[11]) ? 3'b110 : 3'b001;
										assign node942 = (inp[1]) ? node944 : 3'b101;
											assign node944 = (inp[10]) ? 3'b001 : 3'b101;
							assign node947 = (inp[10]) ? node957 : node948;
								assign node948 = (inp[1]) ? node950 : 3'b111;
									assign node950 = (inp[5]) ? node952 : 3'b111;
										assign node952 = (inp[11]) ? 3'b011 : node953;
											assign node953 = (inp[8]) ? 3'b111 : 3'b011;
								assign node957 = (inp[8]) ? node965 : node958;
									assign node958 = (inp[1]) ? node962 : node959;
										assign node959 = (inp[11]) ? 3'b011 : 3'b111;
										assign node962 = (inp[11]) ? 3'b111 : 3'b011;
									assign node965 = (inp[1]) ? node967 : 3'b111;
										assign node967 = (inp[2]) ? node969 : 3'b111;
											assign node969 = (inp[5]) ? 3'b011 : node970;
												assign node970 = (inp[11]) ? 3'b011 : 3'b111;
						assign node974 = (inp[7]) ? node1006 : node975;
							assign node975 = (inp[8]) ? node989 : node976;
								assign node976 = (inp[5]) ? node984 : node977;
									assign node977 = (inp[1]) ? node981 : node978;
										assign node978 = (inp[11]) ? 3'b000 : 3'b001;
										assign node981 = (inp[10]) ? 3'b110 : 3'b001;
									assign node984 = (inp[11]) ? node986 : 3'b110;
										assign node986 = (inp[1]) ? 3'b010 : 3'b110;
								assign node989 = (inp[1]) ? 3'b001 : node990;
									assign node990 = (inp[11]) ? node996 : node991;
										assign node991 = (inp[5]) ? node993 : 3'b011;
											assign node993 = (inp[10]) ? 3'b001 : 3'b101;
										assign node996 = (inp[5]) ? node1002 : node997;
											assign node997 = (inp[10]) ? node999 : 3'b101;
												assign node999 = (inp[2]) ? 3'b001 : 3'b101;
											assign node1002 = (inp[10]) ? 3'b110 : 3'b101;
							assign node1006 = (inp[1]) ? node1036 : node1007;
								assign node1007 = (inp[10]) ? node1023 : node1008;
									assign node1008 = (inp[2]) ? node1018 : node1009;
										assign node1009 = (inp[8]) ? node1013 : node1010;
											assign node1010 = (inp[5]) ? 3'b101 : 3'b111;
											assign node1013 = (inp[5]) ? node1015 : 3'b111;
												assign node1015 = (inp[11]) ? 3'b011 : 3'b111;
										assign node1018 = (inp[5]) ? 3'b011 : node1019;
											assign node1019 = (inp[8]) ? 3'b111 : 3'b011;
									assign node1023 = (inp[11]) ? node1029 : node1024;
										assign node1024 = (inp[8]) ? node1026 : 3'b111;
											assign node1026 = (inp[2]) ? 3'b101 : 3'b011;
										assign node1029 = (inp[8]) ? node1033 : node1030;
											assign node1030 = (inp[5]) ? 3'b001 : 3'b101;
											assign node1033 = (inp[5]) ? 3'b101 : 3'b011;
								assign node1036 = (inp[8]) ? node1048 : node1037;
									assign node1037 = (inp[5]) ? node1043 : node1038;
										assign node1038 = (inp[11]) ? node1040 : 3'b101;
											assign node1040 = (inp[2]) ? 3'b101 : 3'b001;
										assign node1043 = (inp[10]) ? node1045 : 3'b001;
											assign node1045 = (inp[11]) ? 3'b010 : 3'b001;
									assign node1048 = (inp[5]) ? 3'b101 : node1049;
										assign node1049 = (inp[10]) ? 3'b101 : node1050;
											assign node1050 = (inp[11]) ? 3'b011 : 3'b001;
				assign node1055 = (inp[0]) ? node1223 : node1056;
					assign node1056 = (inp[4]) ? node1140 : node1057;
						assign node1057 = (inp[7]) ? node1107 : node1058;
							assign node1058 = (inp[1]) ? node1086 : node1059;
								assign node1059 = (inp[8]) ? node1075 : node1060;
									assign node1060 = (inp[5]) ? node1070 : node1061;
										assign node1061 = (inp[11]) ? 3'b011 : node1062;
											assign node1062 = (inp[2]) ? node1066 : node1063;
												assign node1063 = (inp[10]) ? 3'b011 : 3'b101;
												assign node1066 = (inp[10]) ? 3'b101 : 3'b011;
										assign node1070 = (inp[11]) ? node1072 : 3'b011;
											assign node1072 = (inp[10]) ? 3'b001 : 3'b101;
									assign node1075 = (inp[10]) ? node1079 : node1076;
										assign node1076 = (inp[2]) ? 3'b011 : 3'b111;
										assign node1079 = (inp[11]) ? node1081 : 3'b011;
											assign node1081 = (inp[5]) ? 3'b101 : node1082;
												assign node1082 = (inp[2]) ? 3'b111 : 3'b011;
								assign node1086 = (inp[2]) ? node1092 : node1087;
									assign node1087 = (inp[11]) ? 3'b001 : node1088;
										assign node1088 = (inp[8]) ? 3'b101 : 3'b001;
									assign node1092 = (inp[8]) ? node1100 : node1093;
										assign node1093 = (inp[10]) ? 3'b111 : node1094;
											assign node1094 = (inp[5]) ? 3'b101 : node1095;
												assign node1095 = (inp[11]) ? 3'b101 : 3'b111;
										assign node1100 = (inp[11]) ? 3'b101 : node1101;
											assign node1101 = (inp[5]) ? 3'b101 : node1102;
												assign node1102 = (inp[10]) ? 3'b101 : 3'b011;
							assign node1107 = (inp[8]) ? node1129 : node1108;
								assign node1108 = (inp[10]) ? node1118 : node1109;
									assign node1109 = (inp[5]) ? node1115 : node1110;
										assign node1110 = (inp[2]) ? node1112 : 3'b111;
											assign node1112 = (inp[11]) ? 3'b011 : 3'b111;
										assign node1115 = (inp[1]) ? 3'b011 : 3'b111;
									assign node1118 = (inp[1]) ? node1124 : node1119;
										assign node1119 = (inp[11]) ? node1121 : 3'b011;
											assign node1121 = (inp[5]) ? 3'b011 : 3'b111;
										assign node1124 = (inp[5]) ? 3'b101 : node1125;
											assign node1125 = (inp[11]) ? 3'b011 : 3'b001;
								assign node1129 = (inp[10]) ? node1131 : 3'b111;
									assign node1131 = (inp[1]) ? node1137 : node1132;
										assign node1132 = (inp[5]) ? node1134 : 3'b111;
											assign node1134 = (inp[11]) ? 3'b111 : 3'b011;
										assign node1137 = (inp[5]) ? 3'b111 : 3'b011;
						assign node1140 = (inp[7]) ? node1180 : node1141;
							assign node1141 = (inp[10]) ? node1157 : node1142;
								assign node1142 = (inp[1]) ? node1150 : node1143;
									assign node1143 = (inp[5]) ? 3'b001 : node1144;
										assign node1144 = (inp[11]) ? 3'b101 : node1145;
											assign node1145 = (inp[8]) ? 3'b101 : 3'b001;
									assign node1150 = (inp[8]) ? node1154 : node1151;
										assign node1151 = (inp[2]) ? 3'b110 : 3'b010;
										assign node1154 = (inp[11]) ? 3'b001 : 3'b101;
								assign node1157 = (inp[1]) ? node1163 : node1158;
									assign node1158 = (inp[11]) ? 3'b000 : node1159;
										assign node1159 = (inp[5]) ? 3'b001 : 3'b110;
									assign node1163 = (inp[11]) ? node1171 : node1164;
										assign node1164 = (inp[2]) ? node1166 : 3'b110;
											assign node1166 = (inp[5]) ? 3'b001 : node1167;
												assign node1167 = (inp[8]) ? 3'b001 : 3'b110;
										assign node1171 = (inp[5]) ? node1177 : node1172;
											assign node1172 = (inp[8]) ? node1174 : 3'b110;
												assign node1174 = (inp[2]) ? 3'b110 : 3'b001;
											assign node1177 = (inp[8]) ? 3'b110 : 3'b010;
							assign node1180 = (inp[8]) ? node1200 : node1181;
								assign node1181 = (inp[1]) ? node1191 : node1182;
									assign node1182 = (inp[2]) ? node1184 : 3'b101;
										assign node1184 = (inp[10]) ? node1188 : node1185;
											assign node1185 = (inp[5]) ? 3'b101 : 3'b011;
											assign node1188 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1191 = (inp[11]) ? node1195 : node1192;
										assign node1192 = (inp[10]) ? 3'b001 : 3'b111;
										assign node1195 = (inp[2]) ? node1197 : 3'b001;
											assign node1197 = (inp[10]) ? 3'b001 : 3'b101;
								assign node1200 = (inp[10]) ? node1210 : node1201;
									assign node1201 = (inp[5]) ? node1203 : 3'b011;
										assign node1203 = (inp[1]) ? node1205 : 3'b011;
											assign node1205 = (inp[2]) ? 3'b101 : node1206;
												assign node1206 = (inp[11]) ? 3'b101 : 3'b011;
									assign node1210 = (inp[1]) ? node1218 : node1211;
										assign node1211 = (inp[11]) ? node1215 : node1212;
											assign node1212 = (inp[2]) ? 3'b111 : 3'b011;
											assign node1215 = (inp[5]) ? 3'b101 : 3'b111;
										assign node1218 = (inp[5]) ? node1220 : 3'b101;
											assign node1220 = (inp[11]) ? 3'b001 : 3'b101;
					assign node1223 = (inp[7]) ? node1319 : node1224;
						assign node1224 = (inp[10]) ? node1276 : node1225;
							assign node1225 = (inp[4]) ? node1251 : node1226;
								assign node1226 = (inp[5]) ? node1234 : node1227;
									assign node1227 = (inp[8]) ? 3'b101 : node1228;
										assign node1228 = (inp[2]) ? 3'b001 : node1229;
											assign node1229 = (inp[1]) ? 3'b001 : 3'b101;
									assign node1234 = (inp[8]) ? node1244 : node1235;
										assign node1235 = (inp[11]) ? node1239 : node1236;
											assign node1236 = (inp[1]) ? 3'b110 : 3'b001;
											assign node1239 = (inp[2]) ? node1241 : 3'b110;
												assign node1241 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1244 = (inp[1]) ? node1248 : node1245;
											assign node1245 = (inp[11]) ? 3'b001 : 3'b101;
											assign node1248 = (inp[2]) ? 3'b110 : 3'b001;
								assign node1251 = (inp[5]) ? node1263 : node1252;
									assign node1252 = (inp[1]) ? 3'b010 : node1253;
										assign node1253 = (inp[2]) ? node1255 : 3'b101;
											assign node1255 = (inp[8]) ? node1259 : node1256;
												assign node1256 = (inp[11]) ? 3'b010 : 3'b110;
												assign node1259 = (inp[11]) ? 3'b110 : 3'b001;
									assign node1263 = (inp[2]) ? node1269 : node1264;
										assign node1264 = (inp[8]) ? node1266 : 3'b010;
											assign node1266 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1269 = (inp[11]) ? 3'b100 : node1270;
											assign node1270 = (inp[8]) ? 3'b010 : node1271;
												assign node1271 = (inp[1]) ? 3'b100 : 3'b010;
							assign node1276 = (inp[4]) ? node1296 : node1277;
								assign node1277 = (inp[1]) ? node1285 : node1278;
									assign node1278 = (inp[2]) ? 3'b110 : node1279;
										assign node1279 = (inp[8]) ? node1281 : 3'b110;
											assign node1281 = (inp[5]) ? 3'b110 : 3'b001;
									assign node1285 = (inp[5]) ? node1291 : node1286;
										assign node1286 = (inp[11]) ? node1288 : 3'b110;
											assign node1288 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1291 = (inp[8]) ? 3'b010 : node1292;
											assign node1292 = (inp[11]) ? 3'b100 : 3'b010;
								assign node1296 = (inp[1]) ? node1306 : node1297;
									assign node1297 = (inp[5]) ? node1301 : node1298;
										assign node1298 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1301 = (inp[8]) ? node1303 : 3'b100;
											assign node1303 = (inp[2]) ? 3'b100 : 3'b010;
									assign node1306 = (inp[8]) ? node1312 : node1307;
										assign node1307 = (inp[2]) ? node1309 : 3'b100;
											assign node1309 = (inp[5]) ? 3'b000 : 3'b100;
										assign node1312 = (inp[11]) ? node1314 : 3'b010;
											assign node1314 = (inp[2]) ? 3'b100 : node1315;
												assign node1315 = (inp[5]) ? 3'b100 : 3'b000;
						assign node1319 = (inp[4]) ? node1373 : node1320;
							assign node1320 = (inp[5]) ? node1348 : node1321;
								assign node1321 = (inp[8]) ? node1331 : node1322;
									assign node1322 = (inp[1]) ? node1324 : 3'b101;
										assign node1324 = (inp[2]) ? node1326 : 3'b011;
											assign node1326 = (inp[11]) ? node1328 : 3'b001;
												assign node1328 = (inp[10]) ? 3'b110 : 3'b001;
									assign node1331 = (inp[10]) ? node1339 : node1332;
										assign node1332 = (inp[2]) ? node1334 : 3'b111;
											assign node1334 = (inp[1]) ? 3'b011 : node1335;
												assign node1335 = (inp[11]) ? 3'b011 : 3'b111;
										assign node1339 = (inp[1]) ? node1345 : node1340;
											assign node1340 = (inp[2]) ? node1342 : 3'b011;
												assign node1342 = (inp[11]) ? 3'b101 : 3'b011;
											assign node1345 = (inp[2]) ? 3'b101 : 3'b001;
								assign node1348 = (inp[8]) ? node1358 : node1349;
									assign node1349 = (inp[10]) ? node1353 : node1350;
										assign node1350 = (inp[1]) ? 3'b001 : 3'b101;
										assign node1353 = (inp[1]) ? 3'b110 : node1354;
											assign node1354 = (inp[11]) ? 3'b001 : 3'b011;
									assign node1358 = (inp[2]) ? node1364 : node1359;
										assign node1359 = (inp[1]) ? node1361 : 3'b101;
											assign node1361 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1364 = (inp[1]) ? node1368 : node1365;
											assign node1365 = (inp[11]) ? 3'b001 : 3'b011;
											assign node1368 = (inp[10]) ? 3'b001 : node1369;
												assign node1369 = (inp[11]) ? 3'b001 : 3'b101;
							assign node1373 = (inp[10]) ? node1391 : node1374;
								assign node1374 = (inp[5]) ? node1384 : node1375;
									assign node1375 = (inp[8]) ? node1381 : node1376;
										assign node1376 = (inp[1]) ? node1378 : 3'b001;
											assign node1378 = (inp[11]) ? 3'b010 : 3'b001;
										assign node1381 = (inp[1]) ? 3'b001 : 3'b101;
									assign node1384 = (inp[11]) ? 3'b110 : node1385;
										assign node1385 = (inp[8]) ? 3'b001 : node1386;
											assign node1386 = (inp[1]) ? 3'b110 : 3'b001;
								assign node1391 = (inp[1]) ? node1403 : node1392;
									assign node1392 = (inp[8]) ? node1394 : 3'b110;
										assign node1394 = (inp[5]) ? node1398 : node1395;
											assign node1395 = (inp[2]) ? 3'b001 : 3'b101;
											assign node1398 = (inp[2]) ? 3'b110 : node1399;
												assign node1399 = (inp[11]) ? 3'b110 : 3'b001;
									assign node1403 = (inp[5]) ? node1413 : node1404;
										assign node1404 = (inp[2]) ? node1408 : node1405;
											assign node1405 = (inp[11]) ? 3'b110 : 3'b010;
											assign node1408 = (inp[8]) ? 3'b110 : node1409;
												assign node1409 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1413 = (inp[2]) ? 3'b010 : node1414;
											assign node1414 = (inp[8]) ? 3'b010 : 3'b000;
			assign node1418 = (inp[0]) ? node1736 : node1419;
				assign node1419 = (inp[7]) ? node1581 : node1420;
					assign node1420 = (inp[4]) ? node1494 : node1421;
						assign node1421 = (inp[5]) ? node1469 : node1422;
							assign node1422 = (inp[10]) ? node1446 : node1423;
								assign node1423 = (inp[2]) ? node1431 : node1424;
									assign node1424 = (inp[1]) ? node1426 : 3'b111;
										assign node1426 = (inp[11]) ? 3'b110 : node1427;
											assign node1427 = (inp[8]) ? 3'b011 : 3'b001;
									assign node1431 = (inp[9]) ? node1437 : node1432;
										assign node1432 = (inp[8]) ? 3'b101 : node1433;
											assign node1433 = (inp[1]) ? 3'b001 : 3'b101;
										assign node1437 = (inp[1]) ? node1443 : node1438;
											assign node1438 = (inp[11]) ? 3'b001 : node1439;
												assign node1439 = (inp[8]) ? 3'b000 : 3'b001;
											assign node1443 = (inp[11]) ? 3'b010 : 3'b100;
								assign node1446 = (inp[8]) ? node1458 : node1447;
									assign node1447 = (inp[9]) ? node1449 : 3'b110;
										assign node1449 = (inp[2]) ? node1451 : 3'b100;
											assign node1451 = (inp[1]) ? node1455 : node1452;
												assign node1452 = (inp[11]) ? 3'b010 : 3'b110;
												assign node1455 = (inp[11]) ? 3'b100 : 3'b010;
									assign node1458 = (inp[9]) ? node1462 : node1459;
										assign node1459 = (inp[1]) ? 3'b001 : 3'b100;
										assign node1462 = (inp[11]) ? node1466 : node1463;
											assign node1463 = (inp[2]) ? 3'b111 : 3'b011;
											assign node1466 = (inp[1]) ? 3'b010 : 3'b110;
							assign node1469 = (inp[10]) ? node1485 : node1470;
								assign node1470 = (inp[11]) ? node1480 : node1471;
									assign node1471 = (inp[1]) ? node1477 : node1472;
										assign node1472 = (inp[2]) ? 3'b110 : node1473;
											assign node1473 = (inp[9]) ? 3'b001 : 3'b100;
										assign node1477 = (inp[9]) ? 3'b010 : 3'b001;
									assign node1480 = (inp[1]) ? node1482 : 3'b110;
										assign node1482 = (inp[8]) ? 3'b010 : 3'b110;
								assign node1485 = (inp[9]) ? node1491 : node1486;
									assign node1486 = (inp[8]) ? 3'b110 : node1487;
										assign node1487 = (inp[1]) ? 3'b110 : 3'b100;
									assign node1491 = (inp[1]) ? 3'b100 : 3'b010;
						assign node1494 = (inp[1]) ? node1544 : node1495;
							assign node1495 = (inp[11]) ? node1525 : node1496;
								assign node1496 = (inp[9]) ? node1514 : node1497;
									assign node1497 = (inp[2]) ? node1509 : node1498;
										assign node1498 = (inp[5]) ? node1502 : node1499;
											assign node1499 = (inp[10]) ? 3'b000 : 3'b100;
											assign node1502 = (inp[8]) ? node1506 : node1503;
												assign node1503 = (inp[10]) ? 3'b100 : 3'b110;
												assign node1506 = (inp[10]) ? 3'b110 : 3'b000;
										assign node1509 = (inp[10]) ? 3'b000 : node1510;
											assign node1510 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1514 = (inp[10]) ? node1518 : node1515;
										assign node1515 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1518 = (inp[5]) ? node1520 : 3'b010;
											assign node1520 = (inp[2]) ? node1522 : 3'b100;
												assign node1522 = (inp[8]) ? 3'b100 : 3'b000;
								assign node1525 = (inp[5]) ? node1533 : node1526;
									assign node1526 = (inp[10]) ? node1530 : node1527;
										assign node1527 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1530 = (inp[2]) ? 3'b110 : 3'b010;
									assign node1533 = (inp[10]) ? node1541 : node1534;
										assign node1534 = (inp[8]) ? node1536 : 3'b110;
											assign node1536 = (inp[2]) ? 3'b110 : node1537;
												assign node1537 = (inp[9]) ? 3'b010 : 3'b000;
										assign node1541 = (inp[8]) ? 3'b100 : 3'b000;
							assign node1544 = (inp[9]) ? node1566 : node1545;
								assign node1545 = (inp[10]) ? node1555 : node1546;
									assign node1546 = (inp[5]) ? 3'b010 : node1547;
										assign node1547 = (inp[8]) ? 3'b001 : node1548;
											assign node1548 = (inp[2]) ? 3'b010 : node1549;
												assign node1549 = (inp[11]) ? 3'b000 : 3'b010;
									assign node1555 = (inp[2]) ? 3'b100 : node1556;
										assign node1556 = (inp[5]) ? node1562 : node1557;
											assign node1557 = (inp[11]) ? 3'b010 : node1558;
												assign node1558 = (inp[8]) ? 3'b110 : 3'b010;
											assign node1562 = (inp[11]) ? 3'b100 : 3'b000;
								assign node1566 = (inp[5]) ? 3'b000 : node1567;
									assign node1567 = (inp[10]) ? node1575 : node1568;
										assign node1568 = (inp[8]) ? node1572 : node1569;
											assign node1569 = (inp[11]) ? 3'b000 : 3'b100;
											assign node1572 = (inp[11]) ? 3'b100 : 3'b000;
										assign node1575 = (inp[2]) ? 3'b000 : node1576;
											assign node1576 = (inp[8]) ? 3'b100 : 3'b000;
					assign node1581 = (inp[9]) ? node1645 : node1582;
						assign node1582 = (inp[1]) ? node1608 : node1583;
							assign node1583 = (inp[4]) ? node1591 : node1584;
								assign node1584 = (inp[10]) ? node1586 : 3'b111;
									assign node1586 = (inp[11]) ? 3'b011 : node1587;
										assign node1587 = (inp[5]) ? 3'b011 : 3'b111;
								assign node1591 = (inp[10]) ? node1599 : node1592;
									assign node1592 = (inp[8]) ? 3'b011 : node1593;
										assign node1593 = (inp[11]) ? 3'b100 : node1594;
											assign node1594 = (inp[5]) ? 3'b111 : 3'b011;
									assign node1599 = (inp[11]) ? node1603 : node1600;
										assign node1600 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1603 = (inp[5]) ? node1605 : 3'b001;
											assign node1605 = (inp[8]) ? 3'b001 : 3'b110;
							assign node1608 = (inp[4]) ? node1626 : node1609;
								assign node1609 = (inp[11]) ? node1617 : node1610;
									assign node1610 = (inp[5]) ? 3'b101 : node1611;
										assign node1611 = (inp[8]) ? 3'b011 : node1612;
											assign node1612 = (inp[2]) ? 3'b101 : 3'b111;
									assign node1617 = (inp[10]) ? node1621 : node1618;
										assign node1618 = (inp[5]) ? 3'b101 : 3'b011;
										assign node1621 = (inp[8]) ? node1623 : 3'b001;
											assign node1623 = (inp[5]) ? 3'b001 : 3'b101;
								assign node1626 = (inp[8]) ? node1638 : node1627;
									assign node1627 = (inp[10]) ? node1633 : node1628;
										assign node1628 = (inp[5]) ? 3'b110 : node1629;
											assign node1629 = (inp[11]) ? 3'b101 : 3'b001;
										assign node1633 = (inp[2]) ? node1635 : 3'b110;
											assign node1635 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1638 = (inp[5]) ? 3'b001 : node1639;
										assign node1639 = (inp[2]) ? node1641 : 3'b101;
											assign node1641 = (inp[10]) ? 3'b001 : 3'b101;
						assign node1645 = (inp[4]) ? node1699 : node1646;
							assign node1646 = (inp[1]) ? node1662 : node1647;
								assign node1647 = (inp[11]) ? node1659 : node1648;
									assign node1648 = (inp[8]) ? node1650 : 3'b001;
										assign node1650 = (inp[5]) ? node1656 : node1651;
											assign node1651 = (inp[2]) ? 3'b011 : node1652;
												assign node1652 = (inp[10]) ? 3'b101 : 3'b011;
											assign node1656 = (inp[10]) ? 3'b110 : 3'b101;
									assign node1659 = (inp[10]) ? 3'b001 : 3'b101;
								assign node1662 = (inp[11]) ? node1682 : node1663;
									assign node1663 = (inp[8]) ? node1673 : node1664;
										assign node1664 = (inp[10]) ? node1670 : node1665;
											assign node1665 = (inp[5]) ? 3'b110 : node1666;
												assign node1666 = (inp[2]) ? 3'b001 : 3'b101;
											assign node1670 = (inp[5]) ? 3'b101 : 3'b110;
										assign node1673 = (inp[2]) ? node1677 : node1674;
											assign node1674 = (inp[5]) ? 3'b110 : 3'b001;
											assign node1677 = (inp[10]) ? 3'b001 : node1678;
												assign node1678 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1682 = (inp[5]) ? node1694 : node1683;
										assign node1683 = (inp[8]) ? node1689 : node1684;
											assign node1684 = (inp[2]) ? node1686 : 3'b010;
												assign node1686 = (inp[10]) ? 3'b010 : 3'b110;
											assign node1689 = (inp[10]) ? node1691 : 3'b001;
												assign node1691 = (inp[2]) ? 3'b110 : 3'b001;
										assign node1694 = (inp[8]) ? 3'b110 : node1695;
											assign node1695 = (inp[10]) ? 3'b010 : 3'b110;
							assign node1699 = (inp[1]) ? node1715 : node1700;
								assign node1700 = (inp[10]) ? node1708 : node1701;
									assign node1701 = (inp[8]) ? node1703 : 3'b110;
										assign node1703 = (inp[5]) ? node1705 : 3'b001;
											assign node1705 = (inp[11]) ? 3'b110 : 3'b001;
									assign node1708 = (inp[11]) ? node1710 : 3'b110;
										assign node1710 = (inp[2]) ? node1712 : 3'b010;
											assign node1712 = (inp[8]) ? 3'b110 : 3'b010;
								assign node1715 = (inp[10]) ? node1721 : node1716;
									assign node1716 = (inp[2]) ? node1718 : 3'b110;
										assign node1718 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1721 = (inp[8]) ? node1727 : node1722;
										assign node1722 = (inp[5]) ? node1724 : 3'b100;
											assign node1724 = (inp[2]) ? 3'b000 : 3'b100;
										assign node1727 = (inp[5]) ? node1731 : node1728;
											assign node1728 = (inp[2]) ? 3'b010 : 3'b110;
											assign node1731 = (inp[2]) ? 3'b100 : node1732;
												assign node1732 = (inp[11]) ? 3'b100 : 3'b010;
				assign node1736 = (inp[9]) ? node1916 : node1737;
					assign node1737 = (inp[4]) ? node1819 : node1738;
						assign node1738 = (inp[7]) ? node1782 : node1739;
							assign node1739 = (inp[8]) ? node1763 : node1740;
								assign node1740 = (inp[5]) ? node1752 : node1741;
									assign node1741 = (inp[1]) ? node1747 : node1742;
										assign node1742 = (inp[10]) ? node1744 : 3'b001;
											assign node1744 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1747 = (inp[10]) ? 3'b010 : node1748;
											assign node1748 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1752 = (inp[10]) ? node1758 : node1753;
										assign node1753 = (inp[1]) ? node1755 : 3'b010;
											assign node1755 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1758 = (inp[1]) ? 3'b100 : node1759;
											assign node1759 = (inp[2]) ? 3'b100 : 3'b000;
								assign node1763 = (inp[2]) ? node1777 : node1764;
									assign node1764 = (inp[5]) ? node1772 : node1765;
										assign node1765 = (inp[10]) ? 3'b100 : node1766;
											assign node1766 = (inp[11]) ? 3'b110 : node1767;
												assign node1767 = (inp[1]) ? 3'b001 : 3'b011;
										assign node1772 = (inp[10]) ? 3'b010 : node1773;
											assign node1773 = (inp[1]) ? 3'b110 : 3'b100;
									assign node1777 = (inp[1]) ? node1779 : 3'b110;
										assign node1779 = (inp[10]) ? 3'b010 : 3'b110;
							assign node1782 = (inp[10]) ? node1800 : node1783;
								assign node1783 = (inp[8]) ? node1793 : node1784;
									assign node1784 = (inp[5]) ? node1790 : node1785;
										assign node1785 = (inp[1]) ? 3'b001 : node1786;
											assign node1786 = (inp[2]) ? 3'b101 : 3'b111;
										assign node1790 = (inp[1]) ? 3'b110 : 3'b001;
									assign node1793 = (inp[1]) ? node1797 : node1794;
										assign node1794 = (inp[5]) ? 3'b101 : 3'b011;
										assign node1797 = (inp[5]) ? 3'b001 : 3'b101;
								assign node1800 = (inp[1]) ? node1810 : node1801;
									assign node1801 = (inp[8]) ? node1807 : node1802;
										assign node1802 = (inp[11]) ? 3'b110 : node1803;
											assign node1803 = (inp[5]) ? 3'b010 : 3'b001;
										assign node1807 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1810 = (inp[2]) ? 3'b110 : node1811;
										assign node1811 = (inp[8]) ? 3'b110 : node1812;
											assign node1812 = (inp[11]) ? node1814 : 3'b110;
												assign node1814 = (inp[5]) ? 3'b010 : 3'b110;
						assign node1819 = (inp[7]) ? node1867 : node1820;
							assign node1820 = (inp[10]) ? node1842 : node1821;
								assign node1821 = (inp[11]) ? node1833 : node1822;
									assign node1822 = (inp[8]) ? node1824 : 3'b100;
										assign node1824 = (inp[2]) ? node1826 : 3'b010;
											assign node1826 = (inp[5]) ? node1830 : node1827;
												assign node1827 = (inp[1]) ? 3'b010 : 3'b110;
												assign node1830 = (inp[1]) ? 3'b100 : 3'b010;
									assign node1833 = (inp[8]) ? node1839 : node1834;
										assign node1834 = (inp[1]) ? node1836 : 3'b100;
											assign node1836 = (inp[5]) ? 3'b000 : 3'b100;
										assign node1839 = (inp[1]) ? 3'b100 : 3'b110;
								assign node1842 = (inp[1]) ? node1858 : node1843;
									assign node1843 = (inp[2]) ? node1851 : node1844;
										assign node1844 = (inp[5]) ? node1848 : node1845;
											assign node1845 = (inp[11]) ? 3'b000 : 3'b010;
											assign node1848 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1851 = (inp[11]) ? 3'b100 : node1852;
											assign node1852 = (inp[5]) ? node1854 : 3'b100;
												assign node1854 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1858 = (inp[11]) ? 3'b000 : node1859;
										assign node1859 = (inp[2]) ? 3'b000 : node1860;
											assign node1860 = (inp[5]) ? node1862 : 3'b100;
												assign node1862 = (inp[8]) ? 3'b100 : 3'b000;
							assign node1867 = (inp[8]) ? node1895 : node1868;
								assign node1868 = (inp[10]) ? node1882 : node1869;
									assign node1869 = (inp[5]) ? node1877 : node1870;
										assign node1870 = (inp[2]) ? node1872 : 3'b100;
											assign node1872 = (inp[1]) ? node1874 : 3'b110;
												assign node1874 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1877 = (inp[1]) ? 3'b010 : node1878;
											assign node1878 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1882 = (inp[1]) ? node1888 : node1883;
										assign node1883 = (inp[2]) ? node1885 : 3'b010;
											assign node1885 = (inp[5]) ? 3'b100 : 3'b000;
										assign node1888 = (inp[5]) ? node1890 : 3'b100;
											assign node1890 = (inp[2]) ? node1892 : 3'b100;
												assign node1892 = (inp[11]) ? 3'b000 : 3'b100;
								assign node1895 = (inp[10]) ? node1905 : node1896;
									assign node1896 = (inp[5]) ? 3'b110 : node1897;
										assign node1897 = (inp[1]) ? 3'b110 : node1898;
											assign node1898 = (inp[2]) ? 3'b001 : node1899;
												assign node1899 = (inp[11]) ? 3'b001 : 3'b101;
									assign node1905 = (inp[5]) ? node1911 : node1906;
										assign node1906 = (inp[2]) ? node1908 : 3'b110;
											assign node1908 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1911 = (inp[2]) ? 3'b010 : node1912;
											assign node1912 = (inp[11]) ? 3'b010 : 3'b110;
					assign node1916 = (inp[4]) ? node1984 : node1917;
						assign node1917 = (inp[7]) ? node1949 : node1918;
							assign node1918 = (inp[11]) ? node1938 : node1919;
								assign node1919 = (inp[5]) ? node1931 : node1920;
									assign node1920 = (inp[1]) ? node1928 : node1921;
										assign node1921 = (inp[10]) ? 3'b100 : node1922;
											assign node1922 = (inp[8]) ? node1924 : 3'b010;
												assign node1924 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1928 = (inp[10]) ? 3'b000 : 3'b100;
									assign node1931 = (inp[10]) ? node1933 : 3'b100;
										assign node1933 = (inp[1]) ? 3'b000 : node1934;
											assign node1934 = (inp[8]) ? 3'b100 : 3'b000;
								assign node1938 = (inp[10]) ? 3'b000 : node1939;
									assign node1939 = (inp[1]) ? 3'b000 : node1940;
										assign node1940 = (inp[8]) ? node1944 : node1941;
											assign node1941 = (inp[5]) ? 3'b000 : 3'b100;
											assign node1944 = (inp[5]) ? 3'b100 : 3'b010;
							assign node1949 = (inp[10]) ? node1969 : node1950;
								assign node1950 = (inp[2]) ? node1962 : node1951;
									assign node1951 = (inp[5]) ? node1957 : node1952;
										assign node1952 = (inp[1]) ? 3'b010 : node1953;
											assign node1953 = (inp[11]) ? 3'b101 : 3'b010;
										assign node1957 = (inp[1]) ? 3'b100 : node1958;
											assign node1958 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1962 = (inp[11]) ? 3'b010 : node1963;
										assign node1963 = (inp[5]) ? node1965 : 3'b110;
											assign node1965 = (inp[8]) ? 3'b110 : 3'b010;
								assign node1969 = (inp[8]) ? node1975 : node1970;
									assign node1970 = (inp[1]) ? node1972 : 3'b100;
										assign node1972 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1975 = (inp[11]) ? node1979 : node1976;
										assign node1976 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1979 = (inp[2]) ? 3'b100 : node1980;
											assign node1980 = (inp[5]) ? 3'b010 : 3'b000;
						assign node1984 = (inp[7]) ? node1986 : 3'b000;
							assign node1986 = (inp[10]) ? node2006 : node1987;
								assign node1987 = (inp[1]) ? node1999 : node1988;
									assign node1988 = (inp[8]) ? node1994 : node1989;
										assign node1989 = (inp[5]) ? node1991 : 3'b010;
											assign node1991 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1994 = (inp[2]) ? 3'b010 : node1995;
											assign node1995 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1999 = (inp[8]) ? 3'b100 : node2000;
										assign node2000 = (inp[5]) ? 3'b000 : node2001;
											assign node2001 = (inp[2]) ? 3'b000 : 3'b100;
								assign node2006 = (inp[5]) ? 3'b000 : node2007;
									assign node2007 = (inp[1]) ? 3'b000 : node2008;
										assign node2008 = (inp[2]) ? 3'b100 : node2009;
											assign node2009 = (inp[11]) ? 3'b000 : 3'b010;

endmodule