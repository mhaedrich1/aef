module dtc_split33_bm64 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node14;
	wire [4-1:0] node15;
	wire [4-1:0] node20;
	wire [4-1:0] node22;
	wire [4-1:0] node24;
	wire [4-1:0] node28;
	wire [4-1:0] node30;
	wire [4-1:0] node31;
	wire [4-1:0] node32;
	wire [4-1:0] node33;
	wire [4-1:0] node38;
	wire [4-1:0] node40;
	wire [4-1:0] node41;
	wire [4-1:0] node42;
	wire [4-1:0] node48;
	wire [4-1:0] node50;
	wire [4-1:0] node51;
	wire [4-1:0] node52;
	wire [4-1:0] node53;
	wire [4-1:0] node54;
	wire [4-1:0] node55;
	wire [4-1:0] node57;
	wire [4-1:0] node60;
	wire [4-1:0] node62;
	wire [4-1:0] node64;
	wire [4-1:0] node68;
	wire [4-1:0] node70;
	wire [4-1:0] node72;
	wire [4-1:0] node73;
	wire [4-1:0] node78;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node82;
	wire [4-1:0] node83;
	wire [4-1:0] node85;
	wire [4-1:0] node88;
	wire [4-1:0] node90;
	wire [4-1:0] node94;
	wire [4-1:0] node96;
	wire [4-1:0] node97;
	wire [4-1:0] node98;
	wire [4-1:0] node104;
	wire [4-1:0] node105;
	wire [4-1:0] node106;
	wire [4-1:0] node107;
	wire [4-1:0] node108;
	wire [4-1:0] node109;
	wire [4-1:0] node110;
	wire [4-1:0] node111;
	wire [4-1:0] node112;
	wire [4-1:0] node114;
	wire [4-1:0] node118;
	wire [4-1:0] node119;
	wire [4-1:0] node124;
	wire [4-1:0] node126;
	wire [4-1:0] node127;
	wire [4-1:0] node128;
	wire [4-1:0] node129;
	wire [4-1:0] node136;
	wire [4-1:0] node138;
	wire [4-1:0] node139;
	wire [4-1:0] node140;
	wire [4-1:0] node141;
	wire [4-1:0] node142;
	wire [4-1:0] node146;
	wire [4-1:0] node148;
	wire [4-1:0] node152;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node156;
	wire [4-1:0] node160;
	wire [4-1:0] node162;
	wire [4-1:0] node164;
	wire [4-1:0] node166;
	wire [4-1:0] node170;
	wire [4-1:0] node171;
	wire [4-1:0] node172;
	wire [4-1:0] node173;
	wire [4-1:0] node174;
	wire [4-1:0] node176;
	wire [4-1:0] node177;
	wire [4-1:0] node178;
	wire [4-1:0] node179;
	wire [4-1:0] node184;
	wire [4-1:0] node185;
	wire [4-1:0] node187;
	wire [4-1:0] node188;
	wire [4-1:0] node195;
	wire [4-1:0] node196;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node200;
	wire [4-1:0] node205;
	wire [4-1:0] node206;
	wire [4-1:0] node208;
	wire [4-1:0] node209;
	wire [4-1:0] node210;
	wire [4-1:0] node215;
	wire [4-1:0] node216;
	wire [4-1:0] node217;
	wire [4-1:0] node219;
	wire [4-1:0] node223;
	wire [4-1:0] node224;
	wire [4-1:0] node225;
	wire [4-1:0] node226;
	wire [4-1:0] node231;
	wire [4-1:0] node232;
	wire [4-1:0] node236;
	wire [4-1:0] node237;
	wire [4-1:0] node238;
	wire [4-1:0] node239;
	wire [4-1:0] node240;
	wire [4-1:0] node241;
	wire [4-1:0] node242;
	wire [4-1:0] node248;
	wire [4-1:0] node250;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node256;
	wire [4-1:0] node258;
	wire [4-1:0] node260;
	wire [4-1:0] node264;
	wire [4-1:0] node266;
	wire [4-1:0] node267;
	wire [4-1:0] node268;
	wire [4-1:0] node270;
	wire [4-1:0] node272;
	wire [4-1:0] node274;
	wire [4-1:0] node278;
	wire [4-1:0] node279;
	wire [4-1:0] node281;
	wire [4-1:0] node282;
	wire [4-1:0] node284;
	wire [4-1:0] node289;
	wire [4-1:0] node290;
	wire [4-1:0] node292;
	wire [4-1:0] node293;
	wire [4-1:0] node294;
	wire [4-1:0] node295;
	wire [4-1:0] node296;
	wire [4-1:0] node297;
	wire [4-1:0] node298;
	wire [4-1:0] node299;
	wire [4-1:0] node300;
	wire [4-1:0] node305;
	wire [4-1:0] node306;
	wire [4-1:0] node310;
	wire [4-1:0] node312;
	wire [4-1:0] node314;
	wire [4-1:0] node318;
	wire [4-1:0] node320;
	wire [4-1:0] node321;
	wire [4-1:0] node322;
	wire [4-1:0] node323;
	wire [4-1:0] node324;
	wire [4-1:0] node330;
	wire [4-1:0] node332;
	wire [4-1:0] node334;
	wire [4-1:0] node338;
	wire [4-1:0] node340;
	wire [4-1:0] node341;
	wire [4-1:0] node342;
	wire [4-1:0] node343;
	wire [4-1:0] node344;
	wire [4-1:0] node345;
	wire [4-1:0] node350;
	wire [4-1:0] node352;
	wire [4-1:0] node354;
	wire [4-1:0] node356;
	wire [4-1:0] node360;
	wire [4-1:0] node362;
	wire [4-1:0] node363;
	wire [4-1:0] node364;
	wire [4-1:0] node366;
	wire [4-1:0] node370;
	wire [4-1:0] node372;
	wire [4-1:0] node375;
	wire [4-1:0] node376;
	wire [4-1:0] node377;
	wire [4-1:0] node378;
	wire [4-1:0] node379;
	wire [4-1:0] node380;
	wire [4-1:0] node381;
	wire [4-1:0] node382;
	wire [4-1:0] node384;
	wire [4-1:0] node388;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node396;
	wire [4-1:0] node397;
	wire [4-1:0] node398;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node408;
	wire [4-1:0] node409;
	wire [4-1:0] node410;
	wire [4-1:0] node411;
	wire [4-1:0] node415;
	wire [4-1:0] node418;
	wire [4-1:0] node419;
	wire [4-1:0] node421;
	wire [4-1:0] node425;
	wire [4-1:0] node426;
	wire [4-1:0] node427;
	wire [4-1:0] node428;
	wire [4-1:0] node429;
	wire [4-1:0] node430;
	wire [4-1:0] node431;
	wire [4-1:0] node437;
	wire [4-1:0] node439;
	wire [4-1:0] node440;
	wire [4-1:0] node441;
	wire [4-1:0] node447;
	wire [4-1:0] node449;
	wire [4-1:0] node451;
	wire [4-1:0] node452;
	wire [4-1:0] node456;
	wire [4-1:0] node457;
	wire [4-1:0] node458;
	wire [4-1:0] node459;
	wire [4-1:0] node460;
	wire [4-1:0] node461;
	wire [4-1:0] node463;
	wire [4-1:0] node464;
	wire [4-1:0] node468;
	wire [4-1:0] node471;
	wire [4-1:0] node472;
	wire [4-1:0] node473;
	wire [4-1:0] node475;
	wire [4-1:0] node477;
	wire [4-1:0] node482;
	wire [4-1:0] node483;
	wire [4-1:0] node484;
	wire [4-1:0] node487;
	wire [4-1:0] node490;
	wire [4-1:0] node491;
	wire [4-1:0] node492;
	wire [4-1:0] node493;
	wire [4-1:0] node496;
	wire [4-1:0] node497;
	wire [4-1:0] node502;
	wire [4-1:0] node503;
	wire [4-1:0] node504;
	wire [4-1:0] node507;
	wire [4-1:0] node510;
	wire [4-1:0] node511;
	wire [4-1:0] node512;
	wire [4-1:0] node514;
	wire [4-1:0] node518;
	wire [4-1:0] node520;
	wire [4-1:0] node523;
	wire [4-1:0] node524;
	wire [4-1:0] node525;
	wire [4-1:0] node526;
	wire [4-1:0] node527;
	wire [4-1:0] node528;
	wire [4-1:0] node532;
	wire [4-1:0] node534;
	wire [4-1:0] node537;
	wire [4-1:0] node538;
	wire [4-1:0] node542;
	wire [4-1:0] node543;
	wire [4-1:0] node544;
	wire [4-1:0] node546;
	wire [4-1:0] node550;
	wire [4-1:0] node551;
	wire [4-1:0] node555;
	wire [4-1:0] node556;
	wire [4-1:0] node557;
	wire [4-1:0] node560;
	wire [4-1:0] node561;
	wire [4-1:0] node565;
	wire [4-1:0] node566;
	wire [4-1:0] node567;
	wire [4-1:0] node568;
	wire [4-1:0] node570;
	wire [4-1:0] node575;
	wire [4-1:0] node576;
	wire [4-1:0] node579;
	wire [4-1:0] node581;
	wire [4-1:0] node582;
	wire [4-1:0] node586;
	wire [4-1:0] node587;
	wire [4-1:0] node588;
	wire [4-1:0] node589;
	wire [4-1:0] node590;
	wire [4-1:0] node591;
	wire [4-1:0] node593;
	wire [4-1:0] node597;
	wire [4-1:0] node600;
	wire [4-1:0] node601;
	wire [4-1:0] node602;
	wire [4-1:0] node603;
	wire [4-1:0] node608;
	wire [4-1:0] node609;
	wire [4-1:0] node610;
	wire [4-1:0] node615;
	wire [4-1:0] node616;
	wire [4-1:0] node618;
	wire [4-1:0] node621;
	wire [4-1:0] node622;
	wire [4-1:0] node624;
	wire [4-1:0] node628;
	wire [4-1:0] node629;
	wire [4-1:0] node630;
	wire [4-1:0] node631;
	wire [4-1:0] node633;
	wire [4-1:0] node635;
	wire [4-1:0] node638;
	wire [4-1:0] node639;
	wire [4-1:0] node640;
	wire [4-1:0] node643;
	wire [4-1:0] node646;
	wire [4-1:0] node648;
	wire [4-1:0] node651;
	wire [4-1:0] node652;
	wire [4-1:0] node654;
	wire [4-1:0] node657;
	wire [4-1:0] node660;
	wire [4-1:0] node661;
	wire [4-1:0] node662;
	wire [4-1:0] node663;
	wire [4-1:0] node664;
	wire [4-1:0] node666;
	wire [4-1:0] node671;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node676;
	wire [4-1:0] node677;
	wire [4-1:0] node682;
	wire [4-1:0] node683;
	wire [4-1:0] node686;
	wire [4-1:0] node689;
	wire [4-1:0] node690;
	wire [4-1:0] node691;
	wire [4-1:0] node692;
	wire [4-1:0] node693;
	wire [4-1:0] node694;
	wire [4-1:0] node696;
	wire [4-1:0] node697;
	wire [4-1:0] node701;
	wire [4-1:0] node702;
	wire [4-1:0] node703;
	wire [4-1:0] node708;
	wire [4-1:0] node709;
	wire [4-1:0] node711;
	wire [4-1:0] node712;
	wire [4-1:0] node714;
	wire [4-1:0] node718;
	wire [4-1:0] node720;
	wire [4-1:0] node723;
	wire [4-1:0] node724;
	wire [4-1:0] node725;
	wire [4-1:0] node727;
	wire [4-1:0] node729;
	wire [4-1:0] node732;
	wire [4-1:0] node733;
	wire [4-1:0] node734;
	wire [4-1:0] node739;
	wire [4-1:0] node740;
	wire [4-1:0] node742;
	wire [4-1:0] node745;
	wire [4-1:0] node747;
	wire [4-1:0] node748;
	wire [4-1:0] node752;
	wire [4-1:0] node753;
	wire [4-1:0] node754;
	wire [4-1:0] node755;
	wire [4-1:0] node756;
	wire [4-1:0] node758;
	wire [4-1:0] node762;
	wire [4-1:0] node763;
	wire [4-1:0] node764;
	wire [4-1:0] node766;
	wire [4-1:0] node771;
	wire [4-1:0] node773;
	wire [4-1:0] node774;
	wire [4-1:0] node776;
	wire [4-1:0] node777;
	wire [4-1:0] node782;
	wire [4-1:0] node783;
	wire [4-1:0] node784;
	wire [4-1:0] node786;
	wire [4-1:0] node789;
	wire [4-1:0] node790;
	wire [4-1:0] node792;
	wire [4-1:0] node796;
	wire [4-1:0] node797;
	wire [4-1:0] node799;
	wire [4-1:0] node801;
	wire [4-1:0] node802;
	wire [4-1:0] node806;
	wire [4-1:0] node808;
	wire [4-1:0] node810;
	wire [4-1:0] node813;
	wire [4-1:0] node814;
	wire [4-1:0] node815;
	wire [4-1:0] node816;
	wire [4-1:0] node817;
	wire [4-1:0] node818;
	wire [4-1:0] node819;
	wire [4-1:0] node823;
	wire [4-1:0] node824;
	wire [4-1:0] node826;
	wire [4-1:0] node830;
	wire [4-1:0] node831;
	wire [4-1:0] node832;
	wire [4-1:0] node835;
	wire [4-1:0] node837;
	wire [4-1:0] node840;
	wire [4-1:0] node841;
	wire [4-1:0] node844;
	wire [4-1:0] node845;
	wire [4-1:0] node849;
	wire [4-1:0] node850;
	wire [4-1:0] node851;
	wire [4-1:0] node852;
	wire [4-1:0] node855;
	wire [4-1:0] node858;
	wire [4-1:0] node860;
	wire [4-1:0] node861;
	wire [4-1:0] node863;
	wire [4-1:0] node867;
	wire [4-1:0] node868;
	wire [4-1:0] node869;
	wire [4-1:0] node870;
	wire [4-1:0] node874;
	wire [4-1:0] node877;
	wire [4-1:0] node878;
	wire [4-1:0] node882;
	wire [4-1:0] node883;
	wire [4-1:0] node884;
	wire [4-1:0] node885;
	wire [4-1:0] node886;
	wire [4-1:0] node889;
	wire [4-1:0] node891;
	wire [4-1:0] node893;
	wire [4-1:0] node896;
	wire [4-1:0] node899;
	wire [4-1:0] node902;
	wire [4-1:0] node903;
	wire [4-1:0] node904;
	wire [4-1:0] node905;
	wire [4-1:0] node908;
	wire [4-1:0] node910;
	wire [4-1:0] node913;
	wire [4-1:0] node914;
	wire [4-1:0] node917;
	wire [4-1:0] node918;
	wire [4-1:0] node922;
	wire [4-1:0] node925;
	wire [4-1:0] node926;
	wire [4-1:0] node927;
	wire [4-1:0] node928;
	wire [4-1:0] node929;
	wire [4-1:0] node930;
	wire [4-1:0] node931;
	wire [4-1:0] node932;
	wire [4-1:0] node935;
	wire [4-1:0] node939;
	wire [4-1:0] node940;
	wire [4-1:0] node941;
	wire [4-1:0] node946;
	wire [4-1:0] node947;
	wire [4-1:0] node950;
	wire [4-1:0] node951;
	wire [4-1:0] node952;
	wire [4-1:0] node954;
	wire [4-1:0] node958;
	wire [4-1:0] node961;
	wire [4-1:0] node962;
	wire [4-1:0] node965;
	wire [4-1:0] node968;
	wire [4-1:0] node969;
	wire [4-1:0] node970;
	wire [4-1:0] node971;
	wire [4-1:0] node972;
	wire [4-1:0] node976;
	wire [4-1:0] node979;
	wire [4-1:0] node981;
	wire [4-1:0] node982;
	wire [4-1:0] node983;
	wire [4-1:0] node987;
	wire [4-1:0] node990;
	wire [4-1:0] node991;
	wire [4-1:0] node994;
	wire [4-1:0] node997;
	wire [4-1:0] node998;
	wire [4-1:0] node999;
	wire [4-1:0] node1000;
	wire [4-1:0] node1003;
	wire [4-1:0] node1006;
	wire [4-1:0] node1007;
	wire [4-1:0] node1010;
	wire [4-1:0] node1014;
	wire [4-1:0] node1016;
	wire [4-1:0] node1017;
	wire [4-1:0] node1018;
	wire [4-1:0] node1019;
	wire [4-1:0] node1020;
	wire [4-1:0] node1021;
	wire [4-1:0] node1022;
	wire [4-1:0] node1023;
	wire [4-1:0] node1025;
	wire [4-1:0] node1026;
	wire [4-1:0] node1028;
	wire [4-1:0] node1030;
	wire [4-1:0] node1034;
	wire [4-1:0] node1036;
	wire [4-1:0] node1037;
	wire [4-1:0] node1038;
	wire [4-1:0] node1042;
	wire [4-1:0] node1044;
	wire [4-1:0] node1048;
	wire [4-1:0] node1050;
	wire [4-1:0] node1051;
	wire [4-1:0] node1052;
	wire [4-1:0] node1053;
	wire [4-1:0] node1054;
	wire [4-1:0] node1056;
	wire [4-1:0] node1062;
	wire [4-1:0] node1064;
	wire [4-1:0] node1065;
	wire [4-1:0] node1066;
	wire [4-1:0] node1070;
	wire [4-1:0] node1071;
	wire [4-1:0] node1076;
	wire [4-1:0] node1077;
	wire [4-1:0] node1078;
	wire [4-1:0] node1079;
	wire [4-1:0] node1080;
	wire [4-1:0] node1082;
	wire [4-1:0] node1084;
	wire [4-1:0] node1087;
	wire [4-1:0] node1089;
	wire [4-1:0] node1091;
	wire [4-1:0] node1094;
	wire [4-1:0] node1095;
	wire [4-1:0] node1096;
	wire [4-1:0] node1097;
	wire [4-1:0] node1101;
	wire [4-1:0] node1102;
	wire [4-1:0] node1104;
	wire [4-1:0] node1107;
	wire [4-1:0] node1110;
	wire [4-1:0] node1111;
	wire [4-1:0] node1112;
	wire [4-1:0] node1113;
	wire [4-1:0] node1114;
	wire [4-1:0] node1120;
	wire [4-1:0] node1121;
	wire [4-1:0] node1122;
	wire [4-1:0] node1126;
	wire [4-1:0] node1128;
	wire [4-1:0] node1131;
	wire [4-1:0] node1132;
	wire [4-1:0] node1133;
	wire [4-1:0] node1134;
	wire [4-1:0] node1138;
	wire [4-1:0] node1139;
	wire [4-1:0] node1140;
	wire [4-1:0] node1141;
	wire [4-1:0] node1147;
	wire [4-1:0] node1149;
	wire [4-1:0] node1151;
	wire [4-1:0] node1153;
	wire [4-1:0] node1155;
	wire [4-1:0] node1158;
	wire [4-1:0] node1160;
	wire [4-1:0] node1161;
	wire [4-1:0] node1162;
	wire [4-1:0] node1164;
	wire [4-1:0] node1166;
	wire [4-1:0] node1167;
	wire [4-1:0] node1172;
	wire [4-1:0] node1174;
	wire [4-1:0] node1175;
	wire [4-1:0] node1176;
	wire [4-1:0] node1181;
	wire [4-1:0] node1182;
	wire [4-1:0] node1184;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1187;
	wire [4-1:0] node1188;
	wire [4-1:0] node1190;
	wire [4-1:0] node1192;
	wire [4-1:0] node1196;
	wire [4-1:0] node1198;
	wire [4-1:0] node1199;
	wire [4-1:0] node1201;
	wire [4-1:0] node1206;
	wire [4-1:0] node1208;
	wire [4-1:0] node1209;
	wire [4-1:0] node1211;
	wire [4-1:0] node1212;
	wire [4-1:0] node1214;
	wire [4-1:0] node1215;
	wire [4-1:0] node1220;
	wire [4-1:0] node1222;
	wire [4-1:0] node1223;
	wire [4-1:0] node1224;
	wire [4-1:0] node1226;
	wire [4-1:0] node1230;
	wire [4-1:0] node1232;
	wire [4-1:0] node1235;
	wire [4-1:0] node1236;
	wire [4-1:0] node1237;
	wire [4-1:0] node1238;
	wire [4-1:0] node1239;
	wire [4-1:0] node1240;
	wire [4-1:0] node1241;
	wire [4-1:0] node1242;
	wire [4-1:0] node1246;
	wire [4-1:0] node1249;
	wire [4-1:0] node1250;
	wire [4-1:0] node1253;
	wire [4-1:0] node1254;
	wire [4-1:0] node1256;
	wire [4-1:0] node1259;
	wire [4-1:0] node1262;
	wire [4-1:0] node1263;
	wire [4-1:0] node1265;
	wire [4-1:0] node1266;
	wire [4-1:0] node1270;
	wire [4-1:0] node1271;
	wire [4-1:0] node1272;
	wire [4-1:0] node1277;
	wire [4-1:0] node1278;
	wire [4-1:0] node1279;
	wire [4-1:0] node1280;
	wire [4-1:0] node1283;
	wire [4-1:0] node1286;
	wire [4-1:0] node1287;
	wire [4-1:0] node1290;
	wire [4-1:0] node1293;
	wire [4-1:0] node1294;
	wire [4-1:0] node1295;
	wire [4-1:0] node1300;
	wire [4-1:0] node1301;
	wire [4-1:0] node1302;
	wire [4-1:0] node1303;
	wire [4-1:0] node1304;
	wire [4-1:0] node1308;
	wire [4-1:0] node1309;
	wire [4-1:0] node1312;
	wire [4-1:0] node1313;
	wire [4-1:0] node1315;
	wire [4-1:0] node1319;
	wire [4-1:0] node1320;
	wire [4-1:0] node1321;
	wire [4-1:0] node1326;
	wire [4-1:0] node1327;
	wire [4-1:0] node1328;
	wire [4-1:0] node1329;
	wire [4-1:0] node1334;
	wire [4-1:0] node1335;
	wire [4-1:0] node1337;
	wire [4-1:0] node1339;
	wire [4-1:0] node1341;
	wire [4-1:0] node1344;
	wire [4-1:0] node1346;
	wire [4-1:0] node1349;
	wire [4-1:0] node1350;
	wire [4-1:0] node1351;
	wire [4-1:0] node1352;
	wire [4-1:0] node1353;
	wire [4-1:0] node1355;
	wire [4-1:0] node1358;
	wire [4-1:0] node1359;
	wire [4-1:0] node1363;
	wire [4-1:0] node1364;
	wire [4-1:0] node1366;
	wire [4-1:0] node1368;
	wire [4-1:0] node1369;
	wire [4-1:0] node1370;
	wire [4-1:0] node1373;
	wire [4-1:0] node1377;
	wire [4-1:0] node1379;
	wire [4-1:0] node1380;
	wire [4-1:0] node1384;
	wire [4-1:0] node1385;
	wire [4-1:0] node1386;
	wire [4-1:0] node1388;
	wire [4-1:0] node1391;
	wire [4-1:0] node1393;
	wire [4-1:0] node1395;
	wire [4-1:0] node1397;
	wire [4-1:0] node1400;
	wire [4-1:0] node1401;
	wire [4-1:0] node1402;
	wire [4-1:0] node1406;
	wire [4-1:0] node1407;
	wire [4-1:0] node1411;
	wire [4-1:0] node1412;
	wire [4-1:0] node1413;
	wire [4-1:0] node1414;
	wire [4-1:0] node1415;
	wire [4-1:0] node1416;
	wire [4-1:0] node1421;
	wire [4-1:0] node1422;
	wire [4-1:0] node1423;
	wire [4-1:0] node1428;
	wire [4-1:0] node1429;
	wire [4-1:0] node1430;
	wire [4-1:0] node1431;
	wire [4-1:0] node1435;
	wire [4-1:0] node1436;
	wire [4-1:0] node1437;
	wire [4-1:0] node1440;
	wire [4-1:0] node1442;
	wire [4-1:0] node1446;
	wire [4-1:0] node1447;
	wire [4-1:0] node1449;
	wire [4-1:0] node1452;
	wire [4-1:0] node1455;
	wire [4-1:0] node1456;
	wire [4-1:0] node1457;
	wire [4-1:0] node1458;
	wire [4-1:0] node1461;
	wire [4-1:0] node1464;
	wire [4-1:0] node1465;
	wire [4-1:0] node1470;
	wire [4-1:0] node1472;
	wire [4-1:0] node1473;
	wire [4-1:0] node1474;
	wire [4-1:0] node1475;
	wire [4-1:0] node1476;
	wire [4-1:0] node1477;
	wire [4-1:0] node1478;
	wire [4-1:0] node1479;
	wire [4-1:0] node1480;
	wire [4-1:0] node1482;
	wire [4-1:0] node1488;
	wire [4-1:0] node1490;
	wire [4-1:0] node1494;
	wire [4-1:0] node1495;
	wire [4-1:0] node1496;
	wire [4-1:0] node1498;
	wire [4-1:0] node1500;
	wire [4-1:0] node1503;
	wire [4-1:0] node1506;
	wire [4-1:0] node1508;
	wire [4-1:0] node1510;
	wire [4-1:0] node1512;
	wire [4-1:0] node1515;
	wire [4-1:0] node1516;
	wire [4-1:0] node1518;
	wire [4-1:0] node1519;
	wire [4-1:0] node1521;
	wire [4-1:0] node1522;
	wire [4-1:0] node1523;
	wire [4-1:0] node1528;
	wire [4-1:0] node1530;
	wire [4-1:0] node1531;
	wire [4-1:0] node1532;
	wire [4-1:0] node1537;
	wire [4-1:0] node1538;
	wire [4-1:0] node1539;
	wire [4-1:0] node1540;
	wire [4-1:0] node1542;
	wire [4-1:0] node1545;
	wire [4-1:0] node1546;
	wire [4-1:0] node1547;
	wire [4-1:0] node1551;
	wire [4-1:0] node1552;
	wire [4-1:0] node1556;
	wire [4-1:0] node1557;
	wire [4-1:0] node1559;
	wire [4-1:0] node1562;
	wire [4-1:0] node1563;
	wire [4-1:0] node1564;
	wire [4-1:0] node1569;
	wire [4-1:0] node1570;
	wire [4-1:0] node1571;
	wire [4-1:0] node1572;
	wire [4-1:0] node1575;
	wire [4-1:0] node1577;
	wire [4-1:0] node1580;
	wire [4-1:0] node1581;
	wire [4-1:0] node1582;
	wire [4-1:0] node1585;
	wire [4-1:0] node1586;
	wire [4-1:0] node1589;
	wire [4-1:0] node1593;
	wire [4-1:0] node1594;
	wire [4-1:0] node1595;
	wire [4-1:0] node1598;
	wire [4-1:0] node1601;
	wire [4-1:0] node1602;
	wire [4-1:0] node1603;
	wire [4-1:0] node1606;
	wire [4-1:0] node1610;
	wire [4-1:0] node1612;
	wire [4-1:0] node1613;
	wire [4-1:0] node1614;
	wire [4-1:0] node1615;
	wire [4-1:0] node1616;
	wire [4-1:0] node1617;
	wire [4-1:0] node1618;
	wire [4-1:0] node1619;
	wire [4-1:0] node1624;
	wire [4-1:0] node1626;
	wire [4-1:0] node1627;
	wire [4-1:0] node1631;
	wire [4-1:0] node1633;
	wire [4-1:0] node1634;
	wire [4-1:0] node1638;
	wire [4-1:0] node1640;
	wire [4-1:0] node1641;
	wire [4-1:0] node1644;
	wire [4-1:0] node1645;
	wire [4-1:0] node1648;
	wire [4-1:0] node1649;
	wire [4-1:0] node1653;
	wire [4-1:0] node1654;
	wire [4-1:0] node1655;
	wire [4-1:0] node1656;
	wire [4-1:0] node1657;
	wire [4-1:0] node1658;
	wire [4-1:0] node1662;
	wire [4-1:0] node1665;
	wire [4-1:0] node1666;
	wire [4-1:0] node1668;
	wire [4-1:0] node1671;
	wire [4-1:0] node1675;
	wire [4-1:0] node1676;
	wire [4-1:0] node1677;
	wire [4-1:0] node1681;
	wire [4-1:0] node1682;
	wire [4-1:0] node1684;
	wire [4-1:0] node1687;
	wire [4-1:0] node1688;
	wire [4-1:0] node1692;
	wire [4-1:0] node1694;
	wire [4-1:0] node1695;
	wire [4-1:0] node1696;
	wire [4-1:0] node1697;
	wire [4-1:0] node1701;
	wire [4-1:0] node1702;
	wire [4-1:0] node1705;
	wire [4-1:0] node1706;
	wire [4-1:0] node1710;
	wire [4-1:0] node1712;
	wire [4-1:0] node1713;
	wire [4-1:0] node1715;
	wire [4-1:0] node1718;
	wire [4-1:0] node1720;

	assign outp = (inp[14]) ? node2 : 4'b0000;
		assign node2 = (inp[12]) ? node1014 : node3;
			assign node3 = (inp[3]) ? node289 : node4;
				assign node4 = (inp[0]) ? node104 : node5;
					assign node5 = (inp[4]) ? 4'b0000 : node6;
						assign node6 = (inp[11]) ? node48 : node7;
							assign node7 = (inp[7]) ? 4'b0010 : node8;
								assign node8 = (inp[9]) ? node28 : node9;
									assign node9 = (inp[5]) ? 4'b0000 : node10;
										assign node10 = (inp[13]) ? node20 : node11;
											assign node11 = (inp[15]) ? 4'b0000 : node12;
												assign node12 = (inp[8]) ? node14 : 4'b0010;
													assign node14 = (inp[10]) ? 4'b0000 : node15;
														assign node15 = (inp[1]) ? 4'b0010 : 4'b0000;
											assign node20 = (inp[15]) ? node22 : 4'b0010;
												assign node22 = (inp[10]) ? node24 : 4'b0010;
													assign node24 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node28 = (inp[5]) ? node30 : 4'b0010;
										assign node30 = (inp[15]) ? node38 : node31;
											assign node31 = (inp[13]) ? 4'b0010 : node32;
												assign node32 = (inp[1]) ? 4'b0010 : node33;
													assign node33 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node38 = (inp[13]) ? node40 : 4'b0000;
												assign node40 = (inp[6]) ? 4'b0010 : node41;
													assign node41 = (inp[8]) ? 4'b0000 : node42;
														assign node42 = (inp[10]) ? 4'b0000 : 4'b0010;
							assign node48 = (inp[7]) ? node50 : 4'b0000;
								assign node50 = (inp[5]) ? node78 : node51;
									assign node51 = (inp[9]) ? 4'b0010 : node52;
										assign node52 = (inp[13]) ? node68 : node53;
											assign node53 = (inp[15]) ? 4'b0000 : node54;
												assign node54 = (inp[8]) ? node60 : node55;
													assign node55 = (inp[10]) ? node57 : 4'b0010;
														assign node57 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node60 = (inp[1]) ? node62 : 4'b0000;
														assign node62 = (inp[10]) ? node64 : 4'b0010;
															assign node64 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node68 = (inp[15]) ? node70 : 4'b0010;
												assign node70 = (inp[8]) ? node72 : 4'b0010;
													assign node72 = (inp[10]) ? 4'b0000 : node73;
														assign node73 = (inp[1]) ? 4'b0010 : 4'b0000;
									assign node78 = (inp[9]) ? node80 : 4'b0000;
										assign node80 = (inp[15]) ? node94 : node81;
											assign node81 = (inp[13]) ? 4'b0010 : node82;
												assign node82 = (inp[8]) ? node88 : node83;
													assign node83 = (inp[10]) ? node85 : 4'b0010;
														assign node85 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node88 = (inp[1]) ? node90 : 4'b0000;
														assign node90 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node94 = (inp[13]) ? node96 : 4'b0000;
												assign node96 = (inp[1]) ? 4'b0010 : node97;
													assign node97 = (inp[8]) ? 4'b0000 : node98;
														assign node98 = (inp[2]) ? 4'b0000 : 4'b0010;
					assign node104 = (inp[7]) ? node170 : node105;
						assign node105 = (inp[4]) ? 4'b0010 : node106;
							assign node106 = (inp[11]) ? node136 : node107;
								assign node107 = (inp[9]) ? 4'b0000 : node108;
									assign node108 = (inp[5]) ? node124 : node109;
										assign node109 = (inp[13]) ? 4'b0000 : node110;
											assign node110 = (inp[15]) ? node118 : node111;
												assign node111 = (inp[6]) ? 4'b0000 : node112;
													assign node112 = (inp[8]) ? node114 : 4'b0000;
														assign node114 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node118 = (inp[10]) ? 4'b0010 : node119;
													assign node119 = (inp[1]) ? 4'b0000 : 4'b0010;
										assign node124 = (inp[13]) ? node126 : 4'b0010;
											assign node126 = (inp[1]) ? 4'b0000 : node127;
												assign node127 = (inp[15]) ? 4'b0010 : node128;
													assign node128 = (inp[6]) ? 4'b0000 : node129;
														assign node129 = (inp[10]) ? 4'b0010 : 4'b0000;
								assign node136 = (inp[9]) ? node138 : 4'b0010;
									assign node138 = (inp[5]) ? node152 : node139;
										assign node139 = (inp[13]) ? 4'b0000 : node140;
											assign node140 = (inp[1]) ? node146 : node141;
												assign node141 = (inp[8]) ? 4'b0010 : node142;
													assign node142 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node146 = (inp[15]) ? node148 : 4'b0000;
													assign node148 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node152 = (inp[13]) ? node154 : 4'b0010;
											assign node154 = (inp[1]) ? node160 : node155;
												assign node155 = (inp[15]) ? 4'b0010 : node156;
													assign node156 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node160 = (inp[8]) ? node162 : 4'b0000;
													assign node162 = (inp[10]) ? node164 : 4'b0010;
														assign node164 = (inp[15]) ? node166 : 4'b0000;
															assign node166 = (inp[6]) ? 4'b0000 : 4'b0010;
						assign node170 = (inp[4]) ? node236 : node171;
							assign node171 = (inp[9]) ? node195 : node172;
								assign node172 = (inp[5]) ? 4'b0000 : node173;
									assign node173 = (inp[11]) ? 4'b0000 : node174;
										assign node174 = (inp[13]) ? node176 : 4'b0000;
											assign node176 = (inp[1]) ? node184 : node177;
												assign node177 = (inp[15]) ? 4'b0000 : node178;
													assign node178 = (inp[8]) ? 4'b0000 : node179;
														assign node179 = (inp[6]) ? 4'b0010 : 4'b0000;
												assign node184 = (inp[6]) ? 4'b0010 : node185;
													assign node185 = (inp[15]) ? node187 : 4'b0010;
														assign node187 = (inp[10]) ? 4'b0000 : node188;
															assign node188 = (inp[8]) ? 4'b0000 : 4'b0010;
								assign node195 = (inp[11]) ? node205 : node196;
									assign node196 = (inp[5]) ? node198 : 4'b0010;
										assign node198 = (inp[13]) ? 4'b0010 : node199;
											assign node199 = (inp[1]) ? 4'b0010 : node200;
												assign node200 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node205 = (inp[13]) ? node215 : node206;
										assign node206 = (inp[1]) ? node208 : 4'b0000;
											assign node208 = (inp[15]) ? 4'b0000 : node209;
												assign node209 = (inp[5]) ? 4'b0000 : node210;
													assign node210 = (inp[6]) ? 4'b0010 : 4'b0000;
										assign node215 = (inp[5]) ? node223 : node216;
											assign node216 = (inp[2]) ? 4'b0010 : node217;
												assign node217 = (inp[8]) ? node219 : 4'b0010;
													assign node219 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node223 = (inp[1]) ? node231 : node224;
												assign node224 = (inp[10]) ? 4'b0000 : node225;
													assign node225 = (inp[15]) ? 4'b0000 : node226;
														assign node226 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node231 = (inp[6]) ? 4'b0010 : node232;
													assign node232 = (inp[8]) ? 4'b0000 : 4'b0010;
							assign node236 = (inp[9]) ? node264 : node237;
								assign node237 = (inp[11]) ? 4'b0010 : node238;
									assign node238 = (inp[13]) ? node248 : node239;
										assign node239 = (inp[5]) ? 4'b0010 : node240;
											assign node240 = (inp[1]) ? 4'b0000 : node241;
												assign node241 = (inp[15]) ? 4'b0010 : node242;
													assign node242 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node248 = (inp[5]) ? node250 : 4'b0000;
											assign node250 = (inp[15]) ? node256 : node251;
												assign node251 = (inp[6]) ? 4'b0000 : node252;
													assign node252 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node256 = (inp[1]) ? node258 : 4'b0010;
													assign node258 = (inp[8]) ? node260 : 4'b0000;
														assign node260 = (inp[6]) ? 4'b0000 : 4'b0010;
								assign node264 = (inp[11]) ? node266 : 4'b0000;
									assign node266 = (inp[13]) ? node278 : node267;
										assign node267 = (inp[5]) ? 4'b0010 : node268;
											assign node268 = (inp[15]) ? node270 : 4'b0000;
												assign node270 = (inp[1]) ? node272 : 4'b0010;
													assign node272 = (inp[8]) ? node274 : 4'b0000;
														assign node274 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node278 = (inp[1]) ? 4'b0000 : node279;
											assign node279 = (inp[5]) ? node281 : 4'b0000;
												assign node281 = (inp[15]) ? 4'b0010 : node282;
													assign node282 = (inp[8]) ? node284 : 4'b0000;
														assign node284 = (inp[6]) ? 4'b0000 : 4'b0010;
				assign node289 = (inp[0]) ? node375 : node290;
					assign node290 = (inp[4]) ? node292 : 4'b0010;
						assign node292 = (inp[11]) ? node338 : node293;
							assign node293 = (inp[7]) ? 4'b0010 : node294;
								assign node294 = (inp[5]) ? node318 : node295;
									assign node295 = (inp[9]) ? 4'b0010 : node296;
										assign node296 = (inp[15]) ? node310 : node297;
											assign node297 = (inp[8]) ? node305 : node298;
												assign node298 = (inp[1]) ? 4'b0010 : node299;
													assign node299 = (inp[2]) ? 4'b0010 : node300;
														assign node300 = (inp[6]) ? 4'b0010 : 4'b0000;
												assign node305 = (inp[6]) ? 4'b0010 : node306;
													assign node306 = (inp[13]) ? 4'b0010 : 4'b0000;
											assign node310 = (inp[13]) ? node312 : 4'b0000;
												assign node312 = (inp[8]) ? node314 : 4'b0010;
													assign node314 = (inp[1]) ? 4'b0010 : 4'b0000;
									assign node318 = (inp[9]) ? node320 : 4'b0000;
										assign node320 = (inp[13]) ? node330 : node321;
											assign node321 = (inp[15]) ? 4'b0000 : node322;
												assign node322 = (inp[1]) ? 4'b0010 : node323;
													assign node323 = (inp[8]) ? 4'b0000 : node324;
														assign node324 = (inp[2]) ? 4'b0000 : 4'b0010;
											assign node330 = (inp[8]) ? node332 : 4'b0010;
												assign node332 = (inp[15]) ? node334 : 4'b0010;
													assign node334 = (inp[2]) ? 4'b0010 : 4'b0000;
							assign node338 = (inp[7]) ? node340 : 4'b0000;
								assign node340 = (inp[9]) ? node360 : node341;
									assign node341 = (inp[5]) ? 4'b0000 : node342;
										assign node342 = (inp[15]) ? node350 : node343;
											assign node343 = (inp[1]) ? 4'b0010 : node344;
												assign node344 = (inp[13]) ? 4'b0010 : node345;
													assign node345 = (inp[2]) ? 4'b0010 : 4'b0000;
											assign node350 = (inp[13]) ? node352 : 4'b0000;
												assign node352 = (inp[8]) ? node354 : 4'b0010;
													assign node354 = (inp[1]) ? node356 : 4'b0000;
														assign node356 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node360 = (inp[5]) ? node362 : 4'b0010;
										assign node362 = (inp[13]) ? node370 : node363;
											assign node363 = (inp[15]) ? 4'b0000 : node364;
												assign node364 = (inp[10]) ? node366 : 4'b0010;
													assign node366 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node370 = (inp[15]) ? node372 : 4'b0010;
												assign node372 = (inp[8]) ? 4'b0000 : 4'b0010;
					assign node375 = (inp[9]) ? node689 : node376;
						assign node376 = (inp[7]) ? node456 : node377;
							assign node377 = (inp[4]) ? node425 : node378;
								assign node378 = (inp[13]) ? node396 : node379;
									assign node379 = (inp[11]) ? 4'b0010 : node380;
										assign node380 = (inp[5]) ? node388 : node381;
											assign node381 = (inp[6]) ? 4'b1000 : node382;
												assign node382 = (inp[8]) ? node384 : 4'b1000;
													assign node384 = (inp[1]) ? 4'b1000 : 4'b0010;
											assign node388 = (inp[1]) ? node390 : 4'b0010;
												assign node390 = (inp[6]) ? 4'b1000 : node391;
													assign node391 = (inp[15]) ? 4'b0010 : 4'b1000;
									assign node396 = (inp[11]) ? node408 : node397;
										assign node397 = (inp[5]) ? 4'b1000 : node398;
											assign node398 = (inp[1]) ? node400 : 4'b1000;
												assign node400 = (inp[6]) ? 4'b1010 : node401;
													assign node401 = (inp[10]) ? 4'b1000 : node402;
														assign node402 = (inp[8]) ? 4'b1010 : 4'b1000;
										assign node408 = (inp[1]) ? node418 : node409;
											assign node409 = (inp[6]) ? node415 : node410;
												assign node410 = (inp[15]) ? 4'b0010 : node411;
													assign node411 = (inp[5]) ? 4'b0010 : 4'b1000;
												assign node415 = (inp[5]) ? 4'b0010 : 4'b1000;
											assign node418 = (inp[6]) ? 4'b1000 : node419;
												assign node419 = (inp[15]) ? node421 : 4'b1000;
													assign node421 = (inp[10]) ? 4'b1000 : 4'b0010;
								assign node425 = (inp[11]) ? node447 : node426;
									assign node426 = (inp[13]) ? 4'b0010 : node427;
										assign node427 = (inp[5]) ? node437 : node428;
											assign node428 = (inp[6]) ? 4'b0010 : node429;
												assign node429 = (inp[1]) ? 4'b0010 : node430;
													assign node430 = (inp[15]) ? 4'b0000 : node431;
														assign node431 = (inp[2]) ? 4'b0000 : 4'b0010;
											assign node437 = (inp[1]) ? node439 : 4'b0000;
												assign node439 = (inp[15]) ? 4'b0000 : node440;
													assign node440 = (inp[10]) ? 4'b0000 : node441;
														assign node441 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node447 = (inp[1]) ? node449 : 4'b0000;
										assign node449 = (inp[13]) ? node451 : 4'b0000;
											assign node451 = (inp[5]) ? 4'b0000 : node452;
												assign node452 = (inp[15]) ? 4'b0000 : 4'b0010;
							assign node456 = (inp[13]) ? node586 : node457;
								assign node457 = (inp[4]) ? node523 : node458;
									assign node458 = (inp[1]) ? node482 : node459;
										assign node459 = (inp[11]) ? node471 : node460;
											assign node460 = (inp[5]) ? node468 : node461;
												assign node461 = (inp[6]) ? node463 : 4'b0000;
													assign node463 = (inp[15]) ? 4'b0000 : node464;
														assign node464 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node468 = (inp[6]) ? 4'b0000 : 4'b1010;
											assign node471 = (inp[6]) ? 4'b1010 : node472;
												assign node472 = (inp[5]) ? 4'b1000 : node473;
													assign node473 = (inp[15]) ? node475 : 4'b1010;
														assign node475 = (inp[8]) ? node477 : 4'b1010;
															assign node477 = (inp[10]) ? 4'b1000 : 4'b1010;
										assign node482 = (inp[6]) ? node490 : node483;
											assign node483 = (inp[5]) ? node487 : node484;
												assign node484 = (inp[11]) ? 4'b0000 : 4'b0010;
												assign node487 = (inp[11]) ? 4'b1010 : 4'b0000;
											assign node490 = (inp[2]) ? node502 : node491;
												assign node491 = (inp[15]) ? 4'b0000 : node492;
													assign node492 = (inp[10]) ? node496 : node493;
														assign node493 = (inp[11]) ? 4'b0010 : 4'b0000;
														assign node496 = (inp[8]) ? 4'b0000 : node497;
															assign node497 = (inp[11]) ? 4'b0000 : 4'b0010;
												assign node502 = (inp[8]) ? node510 : node503;
													assign node503 = (inp[5]) ? node507 : node504;
														assign node504 = (inp[10]) ? 4'b0010 : 4'b0000;
														assign node507 = (inp[11]) ? 4'b0000 : 4'b0010;
													assign node510 = (inp[15]) ? node518 : node511;
														assign node511 = (inp[10]) ? 4'b0010 : node512;
															assign node512 = (inp[11]) ? node514 : 4'b0000;
																assign node514 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node518 = (inp[5]) ? node520 : 4'b0000;
															assign node520 = (inp[11]) ? 4'b0000 : 4'b0010;
									assign node523 = (inp[1]) ? node555 : node524;
										assign node524 = (inp[15]) ? node542 : node525;
											assign node525 = (inp[8]) ? node537 : node526;
												assign node526 = (inp[10]) ? node532 : node527;
													assign node527 = (inp[5]) ? 4'b1010 : node528;
														assign node528 = (inp[11]) ? 4'b1010 : 4'b1000;
													assign node532 = (inp[2]) ? node534 : 4'b1000;
														assign node534 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node537 = (inp[6]) ? 4'b1000 : node538;
													assign node538 = (inp[11]) ? 4'b1000 : 4'b1010;
											assign node542 = (inp[11]) ? node550 : node543;
												assign node543 = (inp[5]) ? 4'b1010 : node544;
													assign node544 = (inp[8]) ? node546 : 4'b1000;
														assign node546 = (inp[6]) ? 4'b1000 : 4'b1010;
												assign node550 = (inp[5]) ? 4'b1000 : node551;
													assign node551 = (inp[10]) ? 4'b1000 : 4'b1010;
										assign node555 = (inp[15]) ? node565 : node556;
											assign node556 = (inp[5]) ? node560 : node557;
												assign node557 = (inp[11]) ? 4'b1000 : 4'b1010;
												assign node560 = (inp[6]) ? 4'b1010 : node561;
													assign node561 = (inp[11]) ? 4'b1010 : 4'b1000;
											assign node565 = (inp[11]) ? node575 : node566;
												assign node566 = (inp[5]) ? 4'b1000 : node567;
													assign node567 = (inp[6]) ? 4'b1010 : node568;
														assign node568 = (inp[2]) ? node570 : 4'b1000;
															assign node570 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node575 = (inp[5]) ? node579 : node576;
													assign node576 = (inp[6]) ? 4'b1000 : 4'b1010;
													assign node579 = (inp[10]) ? node581 : 4'b1010;
														assign node581 = (inp[6]) ? 4'b1010 : node582;
															assign node582 = (inp[8]) ? 4'b1000 : 4'b1010;
								assign node586 = (inp[11]) ? node628 : node587;
									assign node587 = (inp[4]) ? node615 : node588;
										assign node588 = (inp[1]) ? node600 : node589;
											assign node589 = (inp[5]) ? node597 : node590;
												assign node590 = (inp[6]) ? 4'b1000 : node591;
													assign node591 = (inp[10]) ? node593 : 4'b0010;
														assign node593 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node597 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node600 = (inp[5]) ? node608 : node601;
												assign node601 = (inp[15]) ? 4'b1010 : node602;
													assign node602 = (inp[6]) ? 4'b1010 : node603;
														assign node603 = (inp[8]) ? 4'b1010 : 4'b1000;
												assign node608 = (inp[6]) ? 4'b1000 : node609;
													assign node609 = (inp[15]) ? 4'b1000 : node610;
														assign node610 = (inp[8]) ? 4'b1000 : 4'b1010;
										assign node615 = (inp[6]) ? node621 : node616;
											assign node616 = (inp[5]) ? node618 : 4'b0000;
												assign node618 = (inp[1]) ? 4'b0010 : 4'b1010;
											assign node621 = (inp[5]) ? 4'b0000 : node622;
												assign node622 = (inp[15]) ? node624 : 4'b0010;
													assign node624 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node628 = (inp[4]) ? node660 : node629;
										assign node629 = (inp[6]) ? node651 : node630;
											assign node630 = (inp[10]) ? node638 : node631;
												assign node631 = (inp[15]) ? node633 : 4'b0010;
													assign node633 = (inp[5]) ? node635 : 4'b0010;
														assign node635 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node638 = (inp[2]) ? node646 : node639;
													assign node639 = (inp[5]) ? node643 : node640;
														assign node640 = (inp[8]) ? 4'b1000 : 4'b0000;
														assign node643 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node646 = (inp[5]) ? node648 : 4'b0010;
														assign node648 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node651 = (inp[1]) ? node657 : node652;
												assign node652 = (inp[5]) ? node654 : 4'b0000;
													assign node654 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node657 = (inp[5]) ? 4'b1000 : 4'b1010;
										assign node660 = (inp[1]) ? node682 : node661;
											assign node661 = (inp[5]) ? node671 : node662;
												assign node662 = (inp[6]) ? 4'b1010 : node663;
													assign node663 = (inp[15]) ? 4'b1000 : node664;
														assign node664 = (inp[10]) ? node666 : 4'b1010;
															assign node666 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node671 = (inp[2]) ? 4'b1000 : node672;
													assign node672 = (inp[6]) ? node676 : node673;
														assign node673 = (inp[8]) ? 4'b1010 : 4'b1000;
														assign node676 = (inp[15]) ? 4'b1000 : node677;
															assign node677 = (inp[8]) ? 4'b1000 : 4'b1010;
											assign node682 = (inp[6]) ? node686 : node683;
												assign node683 = (inp[5]) ? 4'b1010 : 4'b0000;
												assign node686 = (inp[5]) ? 4'b0000 : 4'b0010;
						assign node689 = (inp[7]) ? node813 : node690;
							assign node690 = (inp[4]) ? node752 : node691;
								assign node691 = (inp[11]) ? node723 : node692;
									assign node692 = (inp[13]) ? node708 : node693;
										assign node693 = (inp[1]) ? node701 : node694;
											assign node694 = (inp[5]) ? node696 : 4'b1010;
												assign node696 = (inp[6]) ? 4'b1010 : node697;
													assign node697 = (inp[8]) ? 4'b1000 : 4'b1010;
											assign node701 = (inp[5]) ? 4'b1010 : node702;
												assign node702 = (inp[6]) ? 4'b1000 : node703;
													assign node703 = (inp[8]) ? 4'b1010 : 4'b1000;
										assign node708 = (inp[1]) ? node718 : node709;
											assign node709 = (inp[5]) ? node711 : 4'b1000;
												assign node711 = (inp[2]) ? 4'b1010 : node712;
													assign node712 = (inp[15]) ? node714 : 4'b1000;
														assign node714 = (inp[6]) ? 4'b1000 : 4'b1010;
											assign node718 = (inp[5]) ? node720 : 4'b1010;
												assign node720 = (inp[6]) ? 4'b1010 : 4'b1000;
									assign node723 = (inp[15]) ? node739 : node724;
										assign node724 = (inp[13]) ? node732 : node725;
											assign node725 = (inp[5]) ? node727 : 4'b1010;
												assign node727 = (inp[1]) ? node729 : 4'b1000;
													assign node729 = (inp[6]) ? 4'b1010 : 4'b1000;
											assign node732 = (inp[1]) ? 4'b1000 : node733;
												assign node733 = (inp[5]) ? 4'b1010 : node734;
													assign node734 = (inp[6]) ? 4'b1000 : 4'b1010;
										assign node739 = (inp[13]) ? node745 : node740;
											assign node740 = (inp[1]) ? node742 : 4'b1000;
												assign node742 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node745 = (inp[1]) ? node747 : 4'b1010;
												assign node747 = (inp[6]) ? 4'b1000 : node748;
													assign node748 = (inp[5]) ? 4'b1010 : 4'b1000;
								assign node752 = (inp[13]) ? node782 : node753;
									assign node753 = (inp[11]) ? node771 : node754;
										assign node754 = (inp[1]) ? node762 : node755;
											assign node755 = (inp[5]) ? 4'b0010 : node756;
												assign node756 = (inp[15]) ? node758 : 4'b1000;
													assign node758 = (inp[6]) ? 4'b1000 : 4'b0010;
											assign node762 = (inp[6]) ? 4'b1000 : node763;
												assign node763 = (inp[10]) ? 4'b1000 : node764;
													assign node764 = (inp[5]) ? node766 : 4'b1000;
														assign node766 = (inp[15]) ? 4'b0010 : 4'b1000;
										assign node771 = (inp[15]) ? node773 : 4'b0010;
											assign node773 = (inp[1]) ? 4'b0010 : node774;
												assign node774 = (inp[5]) ? node776 : 4'b0010;
													assign node776 = (inp[8]) ? 4'b0000 : node777;
														assign node777 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node782 = (inp[11]) ? node796 : node783;
										assign node783 = (inp[1]) ? node789 : node784;
											assign node784 = (inp[6]) ? node786 : 4'b1000;
												assign node786 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node789 = (inp[6]) ? 4'b1010 : node790;
												assign node790 = (inp[15]) ? node792 : 4'b1010;
													assign node792 = (inp[5]) ? 4'b1000 : 4'b1010;
										assign node796 = (inp[5]) ? node806 : node797;
											assign node797 = (inp[2]) ? node799 : 4'b1000;
												assign node799 = (inp[15]) ? node801 : 4'b1000;
													assign node801 = (inp[6]) ? 4'b1000 : node802;
														assign node802 = (inp[1]) ? 4'b1000 : 4'b0010;
											assign node806 = (inp[1]) ? node808 : 4'b0010;
												assign node808 = (inp[15]) ? node810 : 4'b1000;
													assign node810 = (inp[6]) ? 4'b1000 : 4'b0010;
							assign node813 = (inp[13]) ? node925 : node814;
								assign node814 = (inp[1]) ? node882 : node815;
									assign node815 = (inp[4]) ? node849 : node816;
										assign node816 = (inp[6]) ? node830 : node817;
											assign node817 = (inp[11]) ? node823 : node818;
												assign node818 = (inp[5]) ? 4'b0001 : node819;
													assign node819 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node823 = (inp[5]) ? 4'b1000 : node824;
													assign node824 = (inp[10]) ? node826 : 4'b1010;
														assign node826 = (inp[8]) ? 4'b1000 : 4'b1010;
											assign node830 = (inp[11]) ? node840 : node831;
												assign node831 = (inp[5]) ? node835 : node832;
													assign node832 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node835 = (inp[8]) ? node837 : 4'b0011;
														assign node837 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node840 = (inp[5]) ? node844 : node841;
													assign node841 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node844 = (inp[15]) ? 4'b0001 : node845;
														assign node845 = (inp[8]) ? 4'b0001 : 4'b0011;
										assign node849 = (inp[11]) ? node867 : node850;
											assign node850 = (inp[6]) ? node858 : node851;
												assign node851 = (inp[5]) ? node855 : node852;
													assign node852 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node855 = (inp[15]) ? 4'b0010 : 4'b1000;
												assign node858 = (inp[2]) ? node860 : 4'b1010;
													assign node860 = (inp[8]) ? 4'b1000 : node861;
														assign node861 = (inp[5]) ? node863 : 4'b1010;
															assign node863 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node867 = (inp[5]) ? node877 : node868;
												assign node868 = (inp[6]) ? node874 : node869;
													assign node869 = (inp[15]) ? 4'b0000 : node870;
														assign node870 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node874 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node877 = (inp[6]) ? 4'b0010 : node878;
													assign node878 = (inp[15]) ? 4'b0010 : 4'b0000;
									assign node882 = (inp[15]) ? node902 : node883;
										assign node883 = (inp[6]) ? node899 : node884;
											assign node884 = (inp[11]) ? node896 : node885;
												assign node885 = (inp[4]) ? node889 : node886;
													assign node886 = (inp[5]) ? 4'b1011 : 4'b0011;
													assign node889 = (inp[5]) ? node891 : 4'b0001;
														assign node891 = (inp[8]) ? node893 : 4'b0011;
															assign node893 = (inp[10]) ? 4'b0001 : 4'b0011;
												assign node896 = (inp[4]) ? 4'b1010 : 4'b1001;
											assign node899 = (inp[11]) ? 4'b0011 : 4'b1011;
										assign node902 = (inp[6]) ? node922 : node903;
											assign node903 = (inp[11]) ? node913 : node904;
												assign node904 = (inp[4]) ? node908 : node905;
													assign node905 = (inp[5]) ? 4'b1001 : 4'b0001;
													assign node908 = (inp[8]) ? node910 : 4'b0001;
														assign node910 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node913 = (inp[4]) ? node917 : node914;
													assign node914 = (inp[5]) ? 4'b0011 : 4'b1011;
													assign node917 = (inp[5]) ? 4'b1010 : node918;
														assign node918 = (inp[10]) ? 4'b1000 : 4'b1010;
											assign node922 = (inp[11]) ? 4'b0001 : 4'b1001;
								assign node925 = (inp[1]) ? node997 : node926;
									assign node926 = (inp[8]) ? node968 : node927;
										assign node927 = (inp[6]) ? node961 : node928;
											assign node928 = (inp[4]) ? node946 : node929;
												assign node929 = (inp[2]) ? node939 : node930;
													assign node930 = (inp[15]) ? 4'b1000 : node931;
														assign node931 = (inp[11]) ? node935 : node932;
															assign node932 = (inp[5]) ? 4'b1010 : 4'b0000;
															assign node935 = (inp[5]) ? 4'b0000 : 4'b1000;
													assign node939 = (inp[15]) ? 4'b0010 : node940;
														assign node940 = (inp[10]) ? 4'b0000 : node941;
															assign node941 = (inp[5]) ? 4'b1010 : 4'b0000;
												assign node946 = (inp[2]) ? node950 : node947;
													assign node947 = (inp[15]) ? 4'b0011 : 4'b1011;
													assign node950 = (inp[11]) ? node958 : node951;
														assign node951 = (inp[15]) ? 4'b1001 : node952;
															assign node952 = (inp[5]) ? node954 : 4'b1011;
																assign node954 = (inp[10]) ? 4'b1001 : 4'b1011;
														assign node958 = (inp[5]) ? 4'b1001 : 4'b0001;
											assign node961 = (inp[5]) ? node965 : node962;
												assign node962 = (inp[4]) ? 4'b1010 : 4'b1011;
												assign node965 = (inp[4]) ? 4'b0010 : 4'b0011;
										assign node968 = (inp[6]) ? node990 : node969;
											assign node969 = (inp[4]) ? node979 : node970;
												assign node970 = (inp[11]) ? node976 : node971;
													assign node971 = (inp[5]) ? 4'b1010 : node972;
														assign node972 = (inp[10]) ? 4'b0010 : 4'b0000;
													assign node976 = (inp[5]) ? 4'b0000 : 4'b1000;
												assign node979 = (inp[2]) ? node981 : 4'b0001;
													assign node981 = (inp[11]) ? node987 : node982;
														assign node982 = (inp[5]) ? 4'b1001 : node983;
															assign node983 = (inp[10]) ? 4'b1001 : 4'b1011;
														assign node987 = (inp[5]) ? 4'b1011 : 4'b0011;
											assign node990 = (inp[5]) ? node994 : node991;
												assign node991 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node994 = (inp[4]) ? 4'b0000 : 4'b0001;
									assign node997 = (inp[6]) ? 4'b0000 : node998;
										assign node998 = (inp[11]) ? node1006 : node999;
											assign node999 = (inp[10]) ? node1003 : node1000;
												assign node1000 = (inp[15]) ? 4'b0111 : 4'b1111;
												assign node1003 = (inp[15]) ? 4'b0101 : 4'b1101;
											assign node1006 = (inp[10]) ? node1010 : node1007;
												assign node1007 = (inp[15]) ? 4'b0110 : 4'b1110;
												assign node1010 = (inp[15]) ? 4'b0100 : 4'b1100;
			assign node1014 = (inp[0]) ? node1016 : 4'b0000;
				assign node1016 = (inp[4]) ? node1470 : node1017;
					assign node1017 = (inp[7]) ? node1181 : node1018;
						assign node1018 = (inp[3]) ? node1076 : node1019;
							assign node1019 = (inp[11]) ? 4'b0000 : node1020;
								assign node1020 = (inp[9]) ? node1048 : node1021;
									assign node1021 = (inp[5]) ? 4'b0000 : node1022;
										assign node1022 = (inp[15]) ? node1034 : node1023;
											assign node1023 = (inp[8]) ? node1025 : 4'b0010;
												assign node1025 = (inp[13]) ? 4'b0010 : node1026;
													assign node1026 = (inp[10]) ? node1028 : 4'b0010;
														assign node1028 = (inp[6]) ? node1030 : 4'b0000;
															assign node1030 = (inp[1]) ? 4'b0010 : 4'b0000;
											assign node1034 = (inp[13]) ? node1036 : 4'b0000;
												assign node1036 = (inp[8]) ? node1042 : node1037;
													assign node1037 = (inp[1]) ? 4'b0010 : node1038;
														assign node1038 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1042 = (inp[1]) ? node1044 : 4'b0000;
														assign node1044 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node1048 = (inp[5]) ? node1050 : 4'b0010;
										assign node1050 = (inp[15]) ? node1062 : node1051;
											assign node1051 = (inp[13]) ? 4'b0010 : node1052;
												assign node1052 = (inp[1]) ? 4'b0010 : node1053;
													assign node1053 = (inp[8]) ? 4'b0000 : node1054;
														assign node1054 = (inp[10]) ? node1056 : 4'b0010;
															assign node1056 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node1062 = (inp[13]) ? node1064 : 4'b0000;
												assign node1064 = (inp[1]) ? node1070 : node1065;
													assign node1065 = (inp[2]) ? 4'b0000 : node1066;
														assign node1066 = (inp[8]) ? 4'b0000 : 4'b0010;
													assign node1070 = (inp[6]) ? 4'b0010 : node1071;
														assign node1071 = (inp[2]) ? 4'b0000 : 4'b0010;
							assign node1076 = (inp[11]) ? node1158 : node1077;
								assign node1077 = (inp[15]) ? node1131 : node1078;
									assign node1078 = (inp[8]) ? node1094 : node1079;
										assign node1079 = (inp[13]) ? node1087 : node1080;
											assign node1080 = (inp[1]) ? node1082 : 4'b0000;
												assign node1082 = (inp[6]) ? node1084 : 4'b0000;
													assign node1084 = (inp[9]) ? 4'b0000 : 4'b0010;
											assign node1087 = (inp[9]) ? node1089 : 4'b0000;
												assign node1089 = (inp[5]) ? node1091 : 4'b0010;
													assign node1091 = (inp[1]) ? 4'b0010 : 4'b0000;
										assign node1094 = (inp[10]) ? node1110 : node1095;
											assign node1095 = (inp[1]) ? node1101 : node1096;
												assign node1096 = (inp[6]) ? 4'b0000 : node1097;
													assign node1097 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node1101 = (inp[9]) ? node1107 : node1102;
													assign node1102 = (inp[5]) ? node1104 : 4'b0000;
														assign node1104 = (inp[13]) ? 4'b0000 : 4'b0010;
													assign node1107 = (inp[13]) ? 4'b0010 : 4'b0000;
											assign node1110 = (inp[6]) ? node1120 : node1111;
												assign node1111 = (inp[9]) ? 4'b0000 : node1112;
													assign node1112 = (inp[1]) ? 4'b0000 : node1113;
														assign node1113 = (inp[5]) ? 4'b0010 : node1114;
															assign node1114 = (inp[13]) ? 4'b0000 : 4'b0010;
												assign node1120 = (inp[13]) ? node1126 : node1121;
													assign node1121 = (inp[5]) ? 4'b0010 : node1122;
														assign node1122 = (inp[9]) ? 4'b0010 : 4'b0000;
													assign node1126 = (inp[9]) ? node1128 : 4'b0000;
														assign node1128 = (inp[1]) ? 4'b0010 : 4'b0000;
									assign node1131 = (inp[9]) ? node1147 : node1132;
										assign node1132 = (inp[1]) ? node1138 : node1133;
											assign node1133 = (inp[5]) ? 4'b0010 : node1134;
												assign node1134 = (inp[13]) ? 4'b0000 : 4'b0010;
											assign node1138 = (inp[13]) ? 4'b0000 : node1139;
												assign node1139 = (inp[5]) ? 4'b0010 : node1140;
													assign node1140 = (inp[6]) ? 4'b0000 : node1141;
														assign node1141 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node1147 = (inp[13]) ? node1149 : 4'b0000;
											assign node1149 = (inp[5]) ? node1151 : 4'b0010;
												assign node1151 = (inp[1]) ? node1153 : 4'b0000;
													assign node1153 = (inp[10]) ? node1155 : 4'b0010;
														assign node1155 = (inp[6]) ? 4'b0010 : 4'b0000;
								assign node1158 = (inp[9]) ? node1160 : 4'b0010;
									assign node1160 = (inp[5]) ? node1172 : node1161;
										assign node1161 = (inp[13]) ? 4'b0000 : node1162;
											assign node1162 = (inp[15]) ? node1164 : 4'b0000;
												assign node1164 = (inp[1]) ? node1166 : 4'b0010;
													assign node1166 = (inp[6]) ? 4'b0000 : node1167;
														assign node1167 = (inp[8]) ? 4'b0010 : 4'b0000;
										assign node1172 = (inp[13]) ? node1174 : 4'b0010;
											assign node1174 = (inp[1]) ? 4'b0000 : node1175;
												assign node1175 = (inp[15]) ? 4'b0010 : node1176;
													assign node1176 = (inp[6]) ? 4'b0000 : 4'b0010;
						assign node1181 = (inp[3]) ? node1235 : node1182;
							assign node1182 = (inp[11]) ? node1184 : 4'b0010;
								assign node1184 = (inp[5]) ? node1206 : node1185;
									assign node1185 = (inp[9]) ? 4'b0010 : node1186;
										assign node1186 = (inp[13]) ? node1196 : node1187;
											assign node1187 = (inp[15]) ? 4'b0000 : node1188;
												assign node1188 = (inp[8]) ? node1190 : 4'b0010;
													assign node1190 = (inp[6]) ? node1192 : 4'b0000;
														assign node1192 = (inp[2]) ? 4'b0010 : 4'b0000;
											assign node1196 = (inp[15]) ? node1198 : 4'b0010;
												assign node1198 = (inp[6]) ? 4'b0010 : node1199;
													assign node1199 = (inp[1]) ? node1201 : 4'b0000;
														assign node1201 = (inp[2]) ? 4'b0000 : 4'b0010;
									assign node1206 = (inp[9]) ? node1208 : 4'b0000;
										assign node1208 = (inp[15]) ? node1220 : node1209;
											assign node1209 = (inp[8]) ? node1211 : 4'b0010;
												assign node1211 = (inp[13]) ? 4'b0010 : node1212;
													assign node1212 = (inp[1]) ? node1214 : 4'b0000;
														assign node1214 = (inp[6]) ? 4'b0010 : node1215;
															assign node1215 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node1220 = (inp[13]) ? node1222 : 4'b0000;
												assign node1222 = (inp[8]) ? node1230 : node1223;
													assign node1223 = (inp[1]) ? 4'b0010 : node1224;
														assign node1224 = (inp[10]) ? node1226 : 4'b0010;
															assign node1226 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1230 = (inp[6]) ? node1232 : 4'b0000;
														assign node1232 = (inp[1]) ? 4'b0010 : 4'b0000;
							assign node1235 = (inp[13]) ? node1349 : node1236;
								assign node1236 = (inp[15]) ? node1300 : node1237;
									assign node1237 = (inp[6]) ? node1277 : node1238;
										assign node1238 = (inp[10]) ? node1262 : node1239;
											assign node1239 = (inp[9]) ? node1249 : node1240;
												assign node1240 = (inp[11]) ? node1246 : node1241;
													assign node1241 = (inp[1]) ? 4'b1000 : node1242;
														assign node1242 = (inp[5]) ? 4'b0010 : 4'b1000;
													assign node1246 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node1249 = (inp[1]) ? node1253 : node1250;
													assign node1250 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node1253 = (inp[11]) ? node1259 : node1254;
														assign node1254 = (inp[5]) ? node1256 : 4'b1000;
															assign node1256 = (inp[2]) ? 4'b0000 : 4'b0010;
														assign node1259 = (inp[5]) ? 4'b1010 : 4'b0010;
											assign node1262 = (inp[5]) ? node1270 : node1263;
												assign node1263 = (inp[9]) ? node1265 : 4'b1000;
													assign node1265 = (inp[11]) ? 4'b1000 : node1266;
														assign node1266 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node1270 = (inp[9]) ? 4'b1010 : node1271;
													assign node1271 = (inp[1]) ? 4'b1000 : node1272;
														assign node1272 = (inp[11]) ? 4'b0000 : 4'b0010;
										assign node1277 = (inp[1]) ? node1293 : node1278;
											assign node1278 = (inp[9]) ? node1286 : node1279;
												assign node1279 = (inp[11]) ? node1283 : node1280;
													assign node1280 = (inp[5]) ? 4'b0010 : 4'b1000;
													assign node1283 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node1286 = (inp[11]) ? node1290 : node1287;
													assign node1287 = (inp[2]) ? 4'b0010 : 4'b0000;
													assign node1290 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node1293 = (inp[11]) ? 4'b0010 : node1294;
												assign node1294 = (inp[9]) ? 4'b1010 : node1295;
													assign node1295 = (inp[5]) ? 4'b1000 : 4'b1010;
									assign node1300 = (inp[11]) ? node1326 : node1301;
										assign node1301 = (inp[1]) ? node1319 : node1302;
											assign node1302 = (inp[9]) ? node1308 : node1303;
												assign node1303 = (inp[5]) ? 4'b0010 : node1304;
													assign node1304 = (inp[6]) ? 4'b1000 : 4'b0010;
												assign node1308 = (inp[5]) ? node1312 : node1309;
													assign node1309 = (inp[6]) ? 4'b0010 : 4'b0000;
													assign node1312 = (inp[6]) ? 4'b0000 : node1313;
														assign node1313 = (inp[8]) ? node1315 : 4'b1010;
															assign node1315 = (inp[2]) ? 4'b1000 : 4'b1010;
											assign node1319 = (inp[6]) ? 4'b1000 : node1320;
												assign node1320 = (inp[9]) ? 4'b0010 : node1321;
													assign node1321 = (inp[5]) ? 4'b0010 : 4'b1000;
										assign node1326 = (inp[9]) ? node1334 : node1327;
											assign node1327 = (inp[5]) ? 4'b0000 : node1328;
												assign node1328 = (inp[1]) ? 4'b0010 : node1329;
													assign node1329 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node1334 = (inp[1]) ? node1344 : node1335;
												assign node1335 = (inp[10]) ? node1337 : 4'b1000;
													assign node1337 = (inp[8]) ? node1339 : 4'b1010;
														assign node1339 = (inp[6]) ? node1341 : 4'b1010;
															assign node1341 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node1344 = (inp[5]) ? node1346 : 4'b0000;
													assign node1346 = (inp[6]) ? 4'b0000 : 4'b1000;
								assign node1349 = (inp[9]) ? node1411 : node1350;
									assign node1350 = (inp[11]) ? node1384 : node1351;
										assign node1351 = (inp[1]) ? node1363 : node1352;
											assign node1352 = (inp[15]) ? node1358 : node1353;
												assign node1353 = (inp[5]) ? node1355 : 4'b1000;
													assign node1355 = (inp[6]) ? 4'b1010 : 4'b1000;
												assign node1358 = (inp[10]) ? 4'b1010 : node1359;
													assign node1359 = (inp[2]) ? 4'b1000 : 4'b1010;
											assign node1363 = (inp[10]) ? node1377 : node1364;
												assign node1364 = (inp[8]) ? node1366 : 4'b1010;
													assign node1366 = (inp[15]) ? node1368 : 4'b1000;
														assign node1368 = (inp[2]) ? 4'b1010 : node1369;
															assign node1369 = (inp[5]) ? node1373 : node1370;
																assign node1370 = (inp[6]) ? 4'b1010 : 4'b1000;
																assign node1373 = (inp[6]) ? 4'b1000 : 4'b1010;
												assign node1377 = (inp[8]) ? node1379 : 4'b1000;
													assign node1379 = (inp[2]) ? 4'b1000 : node1380;
														assign node1380 = (inp[5]) ? 4'b1010 : 4'b1000;
										assign node1384 = (inp[1]) ? node1400 : node1385;
											assign node1385 = (inp[5]) ? node1391 : node1386;
												assign node1386 = (inp[15]) ? node1388 : 4'b1000;
													assign node1388 = (inp[2]) ? 4'b1000 : 4'b0010;
												assign node1391 = (inp[15]) ? node1393 : 4'b0010;
													assign node1393 = (inp[2]) ? node1395 : 4'b0010;
														assign node1395 = (inp[10]) ? node1397 : 4'b0010;
															assign node1397 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node1400 = (inp[5]) ? node1406 : node1401;
												assign node1401 = (inp[6]) ? 4'b1010 : node1402;
													assign node1402 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node1406 = (inp[6]) ? 4'b1000 : node1407;
													assign node1407 = (inp[15]) ? 4'b0010 : 4'b1000;
									assign node1411 = (inp[1]) ? node1455 : node1412;
										assign node1412 = (inp[5]) ? node1428 : node1413;
											assign node1413 = (inp[8]) ? node1421 : node1414;
												assign node1414 = (inp[6]) ? 4'b1011 : node1415;
													assign node1415 = (inp[11]) ? 4'b1010 : node1416;
														assign node1416 = (inp[15]) ? 4'b0011 : 4'b1011;
												assign node1421 = (inp[6]) ? 4'b1001 : node1422;
													assign node1422 = (inp[11]) ? 4'b1010 : node1423;
														assign node1423 = (inp[15]) ? 4'b0011 : 4'b1001;
											assign node1428 = (inp[11]) ? node1446 : node1429;
												assign node1429 = (inp[10]) ? node1435 : node1430;
													assign node1430 = (inp[8]) ? 4'b0001 : node1431;
														assign node1431 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node1435 = (inp[15]) ? 4'b0001 : node1436;
														assign node1436 = (inp[2]) ? node1440 : node1437;
															assign node1437 = (inp[8]) ? 4'b0011 : 4'b0001;
															assign node1440 = (inp[8]) ? node1442 : 4'b0011;
																assign node1442 = (inp[6]) ? 4'b0001 : 4'b0011;
												assign node1446 = (inp[6]) ? node1452 : node1447;
													assign node1447 = (inp[10]) ? node1449 : 4'b0010;
														assign node1449 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node1452 = (inp[8]) ? 4'b0001 : 4'b0011;
										assign node1455 = (inp[6]) ? 4'b0000 : node1456;
											assign node1456 = (inp[10]) ? node1464 : node1457;
												assign node1457 = (inp[11]) ? node1461 : node1458;
													assign node1458 = (inp[15]) ? 4'b0011 : 4'b1011;
													assign node1461 = (inp[15]) ? 4'b0010 : 4'b1010;
												assign node1464 = (inp[11]) ? 4'b1000 : node1465;
													assign node1465 = (inp[15]) ? 4'b0001 : 4'b1001;
					assign node1470 = (inp[3]) ? node1472 : 4'b0000;
						assign node1472 = (inp[11]) ? node1610 : node1473;
							assign node1473 = (inp[9]) ? node1515 : node1474;
								assign node1474 = (inp[7]) ? node1494 : node1475;
									assign node1475 = (inp[5]) ? 4'b0000 : node1476;
										assign node1476 = (inp[15]) ? node1488 : node1477;
											assign node1477 = (inp[1]) ? 4'b0010 : node1478;
												assign node1478 = (inp[13]) ? 4'b0010 : node1479;
													assign node1479 = (inp[8]) ? 4'b0000 : node1480;
														assign node1480 = (inp[10]) ? node1482 : 4'b0010;
															assign node1482 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node1488 = (inp[13]) ? node1490 : 4'b0000;
												assign node1490 = (inp[1]) ? 4'b0010 : 4'b0000;
									assign node1494 = (inp[5]) ? node1506 : node1495;
										assign node1495 = (inp[13]) ? node1503 : node1496;
											assign node1496 = (inp[15]) ? node1498 : 4'b0000;
												assign node1498 = (inp[1]) ? node1500 : 4'b0010;
													assign node1500 = (inp[6]) ? 4'b0000 : 4'b0010;
											assign node1503 = (inp[1]) ? 4'b0010 : 4'b0000;
										assign node1506 = (inp[13]) ? node1508 : 4'b0010;
											assign node1508 = (inp[1]) ? node1510 : 4'b0010;
												assign node1510 = (inp[8]) ? node1512 : 4'b0000;
													assign node1512 = (inp[6]) ? 4'b0000 : 4'b0010;
								assign node1515 = (inp[7]) ? node1537 : node1516;
									assign node1516 = (inp[5]) ? node1518 : 4'b0010;
										assign node1518 = (inp[15]) ? node1528 : node1519;
											assign node1519 = (inp[2]) ? node1521 : 4'b0010;
												assign node1521 = (inp[13]) ? 4'b0010 : node1522;
													assign node1522 = (inp[6]) ? 4'b0010 : node1523;
														assign node1523 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node1528 = (inp[13]) ? node1530 : 4'b0000;
												assign node1530 = (inp[1]) ? 4'b0010 : node1531;
													assign node1531 = (inp[8]) ? 4'b0000 : node1532;
														assign node1532 = (inp[10]) ? 4'b0000 : 4'b0010;
									assign node1537 = (inp[5]) ? node1569 : node1538;
										assign node1538 = (inp[13]) ? node1556 : node1539;
											assign node1539 = (inp[1]) ? node1545 : node1540;
												assign node1540 = (inp[15]) ? node1542 : 4'b1000;
													assign node1542 = (inp[6]) ? 4'b1000 : 4'b0010;
												assign node1545 = (inp[15]) ? node1551 : node1546;
													assign node1546 = (inp[6]) ? 4'b1010 : node1547;
														assign node1547 = (inp[2]) ? 4'b1000 : 4'b1010;
													assign node1551 = (inp[8]) ? 4'b1000 : node1552;
														assign node1552 = (inp[2]) ? 4'b1010 : 4'b1000;
											assign node1556 = (inp[1]) ? node1562 : node1557;
												assign node1557 = (inp[6]) ? node1559 : 4'b0000;
													assign node1559 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node1562 = (inp[6]) ? 4'b0000 : node1563;
													assign node1563 = (inp[10]) ? 4'b1001 : node1564;
														assign node1564 = (inp[15]) ? 4'b0011 : 4'b1011;
										assign node1569 = (inp[1]) ? node1593 : node1570;
											assign node1570 = (inp[8]) ? node1580 : node1571;
												assign node1571 = (inp[2]) ? node1575 : node1572;
													assign node1572 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node1575 = (inp[13]) ? node1577 : 4'b0010;
														assign node1577 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node1580 = (inp[15]) ? 4'b0000 : node1581;
													assign node1581 = (inp[10]) ? node1585 : node1582;
														assign node1582 = (inp[13]) ? 4'b1010 : 4'b0010;
														assign node1585 = (inp[6]) ? node1589 : node1586;
															assign node1586 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node1589 = (inp[13]) ? 4'b0000 : 4'b0010;
											assign node1593 = (inp[13]) ? node1601 : node1594;
												assign node1594 = (inp[15]) ? node1598 : node1595;
													assign node1595 = (inp[6]) ? 4'b1010 : 4'b1000;
													assign node1598 = (inp[6]) ? 4'b1000 : 4'b0010;
												assign node1601 = (inp[6]) ? 4'b0000 : node1602;
													assign node1602 = (inp[10]) ? node1606 : node1603;
														assign node1603 = (inp[2]) ? 4'b0011 : 4'b1011;
														assign node1606 = (inp[15]) ? 4'b0001 : 4'b1001;
							assign node1610 = (inp[7]) ? node1612 : 4'b0000;
								assign node1612 = (inp[5]) ? node1692 : node1613;
									assign node1613 = (inp[8]) ? node1653 : node1614;
										assign node1614 = (inp[13]) ? node1638 : node1615;
											assign node1615 = (inp[10]) ? node1631 : node1616;
												assign node1616 = (inp[2]) ? node1624 : node1617;
													assign node1617 = (inp[6]) ? 4'b0010 : node1618;
														assign node1618 = (inp[15]) ? 4'b0000 : node1619;
															assign node1619 = (inp[1]) ? 4'b0010 : 4'b0000;
													assign node1624 = (inp[6]) ? node1626 : 4'b0010;
														assign node1626 = (inp[1]) ? 4'b0010 : node1627;
															assign node1627 = (inp[9]) ? 4'b0000 : 4'b0010;
												assign node1631 = (inp[6]) ? node1633 : 4'b0000;
													assign node1633 = (inp[9]) ? 4'b0000 : node1634;
														assign node1634 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node1638 = (inp[9]) ? node1640 : 4'b0010;
												assign node1640 = (inp[1]) ? node1644 : node1641;
													assign node1641 = (inp[6]) ? 4'b1010 : 4'b0010;
													assign node1644 = (inp[15]) ? node1648 : node1645;
														assign node1645 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node1648 = (inp[10]) ? 4'b0000 : node1649;
															assign node1649 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node1653 = (inp[2]) ? node1675 : node1654;
											assign node1654 = (inp[10]) ? 4'b0010 : node1655;
												assign node1655 = (inp[13]) ? node1665 : node1656;
													assign node1656 = (inp[6]) ? node1662 : node1657;
														assign node1657 = (inp[1]) ? 4'b0010 : node1658;
															assign node1658 = (inp[9]) ? 4'b0010 : 4'b0000;
														assign node1662 = (inp[1]) ? 4'b0000 : 4'b0010;
													assign node1665 = (inp[9]) ? node1671 : node1666;
														assign node1666 = (inp[15]) ? node1668 : 4'b0010;
															assign node1668 = (inp[6]) ? 4'b0010 : 4'b0000;
														assign node1671 = (inp[1]) ? 4'b0000 : 4'b1000;
											assign node1675 = (inp[9]) ? node1681 : node1676;
												assign node1676 = (inp[15]) ? 4'b0000 : node1677;
													assign node1677 = (inp[10]) ? 4'b0010 : 4'b0000;
												assign node1681 = (inp[6]) ? node1687 : node1682;
													assign node1682 = (inp[1]) ? node1684 : 4'b0010;
														assign node1684 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node1687 = (inp[1]) ? 4'b0000 : node1688;
														assign node1688 = (inp[15]) ? 4'b0010 : 4'b0000;
									assign node1692 = (inp[9]) ? node1694 : 4'b0000;
										assign node1694 = (inp[15]) ? node1710 : node1695;
											assign node1695 = (inp[13]) ? node1701 : node1696;
												assign node1696 = (inp[1]) ? 4'b0010 : node1697;
													assign node1697 = (inp[8]) ? 4'b0000 : 4'b0010;
												assign node1701 = (inp[6]) ? node1705 : node1702;
													assign node1702 = (inp[1]) ? 4'b1010 : 4'b0010;
													assign node1705 = (inp[8]) ? 4'b0000 : node1706;
														assign node1706 = (inp[1]) ? 4'b0000 : 4'b0010;
											assign node1710 = (inp[13]) ? node1712 : 4'b0000;
												assign node1712 = (inp[8]) ? node1718 : node1713;
													assign node1713 = (inp[1]) ? node1715 : 4'b0010;
														assign node1715 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1718 = (inp[1]) ? node1720 : 4'b0000;
														assign node1720 = (inp[10]) ? 4'b0000 : 4'b0010;

endmodule