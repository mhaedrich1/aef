module dtc_split75_bm85 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node118;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node213;
	wire [3-1:0] node217;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node281;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node289;
	wire [3-1:0] node292;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node310;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node344;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node352;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node360;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node389;
	wire [3-1:0] node392;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node407;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node413;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node422;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node433;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node458;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node477;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node488;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node494;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node500;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node522;
	wire [3-1:0] node524;
	wire [3-1:0] node526;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node569;
	wire [3-1:0] node571;
	wire [3-1:0] node574;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node580;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node598;
	wire [3-1:0] node600;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node607;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node614;

	assign outp = (inp[6]) ? node522 : node1;
		assign node1 = (inp[0]) ? node111 : node2;
			assign node2 = (inp[9]) ? node4 : 3'b000;
				assign node4 = (inp[3]) ? node6 : 3'b000;
					assign node6 = (inp[4]) ? node22 : node7;
						assign node7 = (inp[1]) ? node9 : 3'b000;
							assign node9 = (inp[2]) ? node11 : 3'b000;
								assign node11 = (inp[7]) ? 3'b000 : node12;
									assign node12 = (inp[10]) ? node16 : node13;
										assign node13 = (inp[8]) ? 3'b100 : 3'b000;
										assign node16 = (inp[5]) ? 3'b100 : node17;
											assign node17 = (inp[8]) ? 3'b000 : 3'b100;
						assign node22 = (inp[1]) ? node46 : node23;
							assign node23 = (inp[7]) ? 3'b000 : node24;
								assign node24 = (inp[2]) ? node36 : node25;
									assign node25 = (inp[5]) ? node31 : node26;
										assign node26 = (inp[8]) ? 3'b000 : node27;
											assign node27 = (inp[11]) ? 3'b100 : 3'b000;
										assign node31 = (inp[10]) ? node33 : 3'b100;
											assign node33 = (inp[8]) ? 3'b100 : 3'b010;
									assign node36 = (inp[10]) ? node42 : node37;
										assign node37 = (inp[8]) ? node39 : 3'b010;
											assign node39 = (inp[5]) ? 3'b011 : 3'b010;
										assign node42 = (inp[5]) ? 3'b001 : 3'b000;
							assign node46 = (inp[7]) ? node84 : node47;
								assign node47 = (inp[10]) ? node65 : node48;
									assign node48 = (inp[11]) ? node56 : node49;
										assign node49 = (inp[2]) ? node53 : node50;
											assign node50 = (inp[8]) ? 3'b010 : 3'b110;
											assign node53 = (inp[5]) ? 3'b001 : 3'b010;
										assign node56 = (inp[2]) ? node60 : node57;
											assign node57 = (inp[8]) ? 3'b010 : 3'b001;
											assign node60 = (inp[8]) ? 3'b001 : node61;
												assign node61 = (inp[5]) ? 3'b101 : 3'b110;
									assign node65 = (inp[8]) ? node75 : node66;
										assign node66 = (inp[11]) ? node70 : node67;
											assign node67 = (inp[2]) ? 3'b101 : 3'b001;
											assign node70 = (inp[2]) ? node72 : 3'b101;
												assign node72 = (inp[5]) ? 3'b011 : 3'b001;
										assign node75 = (inp[11]) ? node79 : node76;
											assign node76 = (inp[5]) ? 3'b110 : 3'b010;
											assign node79 = (inp[5]) ? 3'b101 : node80;
												assign node80 = (inp[2]) ? 3'b110 : 3'b101;
								assign node84 = (inp[2]) ? node96 : node85;
									assign node85 = (inp[8]) ? node91 : node86;
										assign node86 = (inp[10]) ? node88 : 3'b100;
											assign node88 = (inp[5]) ? 3'b010 : 3'b110;
										assign node91 = (inp[10]) ? 3'b100 : node92;
											assign node92 = (inp[5]) ? 3'b000 : 3'b100;
									assign node96 = (inp[8]) ? node108 : node97;
										assign node97 = (inp[10]) ? node103 : node98;
											assign node98 = (inp[5]) ? 3'b010 : node99;
												assign node99 = (inp[11]) ? 3'b110 : 3'b010;
											assign node103 = (inp[11]) ? node105 : 3'b110;
												assign node105 = (inp[5]) ? 3'b110 : 3'b010;
										assign node108 = (inp[10]) ? 3'b010 : 3'b100;
			assign node111 = (inp[3]) ? node247 : node112;
				assign node112 = (inp[4]) ? node130 : node113;
					assign node113 = (inp[5]) ? node115 : 3'b000;
						assign node115 = (inp[7]) ? 3'b000 : node116;
							assign node116 = (inp[9]) ? node118 : 3'b000;
								assign node118 = (inp[1]) ? node120 : 3'b000;
									assign node120 = (inp[2]) ? node122 : 3'b000;
										assign node122 = (inp[10]) ? node126 : node123;
											assign node123 = (inp[8]) ? 3'b100 : 3'b000;
											assign node126 = (inp[8]) ? 3'b000 : 3'b100;
					assign node130 = (inp[9]) ? node166 : node131;
						assign node131 = (inp[7]) ? 3'b100 : node132;
							assign node132 = (inp[5]) ? node142 : node133;
								assign node133 = (inp[11]) ? node135 : 3'b100;
									assign node135 = (inp[10]) ? node139 : node136;
										assign node136 = (inp[8]) ? 3'b100 : 3'b000;
										assign node139 = (inp[8]) ? 3'b000 : 3'b100;
								assign node142 = (inp[11]) ? node158 : node143;
									assign node143 = (inp[2]) ? node151 : node144;
										assign node144 = (inp[10]) ? node148 : node145;
											assign node145 = (inp[8]) ? 3'b000 : 3'b100;
											assign node148 = (inp[8]) ? 3'b100 : 3'b000;
										assign node151 = (inp[8]) ? node155 : node152;
											assign node152 = (inp[10]) ? 3'b000 : 3'b100;
											assign node155 = (inp[10]) ? 3'b100 : 3'b000;
									assign node158 = (inp[10]) ? node162 : node159;
										assign node159 = (inp[8]) ? 3'b000 : 3'b100;
										assign node162 = (inp[8]) ? 3'b100 : 3'b000;
						assign node166 = (inp[1]) ? node206 : node167;
							assign node167 = (inp[7]) ? node181 : node168;
								assign node168 = (inp[2]) ? 3'b100 : node169;
									assign node169 = (inp[5]) ? node175 : node170;
										assign node170 = (inp[8]) ? 3'b100 : node171;
											assign node171 = (inp[11]) ? 3'b000 : 3'b100;
										assign node175 = (inp[8]) ? 3'b000 : node176;
											assign node176 = (inp[11]) ? 3'b100 : 3'b000;
								assign node181 = (inp[11]) ? node199 : node182;
									assign node182 = (inp[5]) ? node192 : node183;
										assign node183 = (inp[2]) ? node189 : node184;
											assign node184 = (inp[8]) ? 3'b000 : node185;
												assign node185 = (inp[10]) ? 3'b000 : 3'b100;
											assign node189 = (inp[10]) ? 3'b100 : 3'b000;
										assign node192 = (inp[10]) ? node196 : node193;
											assign node193 = (inp[8]) ? 3'b000 : 3'b100;
											assign node196 = (inp[8]) ? 3'b100 : 3'b000;
									assign node199 = (inp[10]) ? node203 : node200;
										assign node200 = (inp[8]) ? 3'b000 : 3'b100;
										assign node203 = (inp[8]) ? 3'b100 : 3'b000;
							assign node206 = (inp[7]) ? node226 : node207;
								assign node207 = (inp[2]) ? node217 : node208;
									assign node208 = (inp[11]) ? node210 : 3'b000;
										assign node210 = (inp[8]) ? 3'b000 : node211;
											assign node211 = (inp[10]) ? node213 : 3'b100;
												assign node213 = (inp[5]) ? 3'b100 : 3'b000;
									assign node217 = (inp[5]) ? node219 : 3'b010;
										assign node219 = (inp[10]) ? node223 : node220;
											assign node220 = (inp[8]) ? 3'b011 : 3'b110;
											assign node223 = (inp[8]) ? 3'b100 : 3'b001;
								assign node226 = (inp[2]) ? node240 : node227;
									assign node227 = (inp[11]) ? node235 : node228;
										assign node228 = (inp[8]) ? node232 : node229;
											assign node229 = (inp[10]) ? 3'b000 : 3'b100;
											assign node232 = (inp[10]) ? 3'b100 : 3'b000;
										assign node235 = (inp[8]) ? node237 : 3'b100;
											assign node237 = (inp[10]) ? 3'b100 : 3'b000;
									assign node240 = (inp[10]) ? node244 : node241;
										assign node241 = (inp[8]) ? 3'b000 : 3'b100;
										assign node244 = (inp[8]) ? 3'b100 : 3'b000;
				assign node247 = (inp[9]) ? node303 : node248;
					assign node248 = (inp[7]) ? 3'b001 : node249;
						assign node249 = (inp[4]) ? 3'b111 : node250;
							assign node250 = (inp[11]) ? node260 : node251;
								assign node251 = (inp[5]) ? node253 : 3'b001;
									assign node253 = (inp[8]) ? node257 : node254;
										assign node254 = (inp[10]) ? 3'b101 : 3'b001;
										assign node257 = (inp[10]) ? 3'b001 : 3'b101;
								assign node260 = (inp[1]) ? node284 : node261;
									assign node261 = (inp[2]) ? node271 : node262;
										assign node262 = (inp[5]) ? 3'b001 : node263;
											assign node263 = (inp[10]) ? node267 : node264;
												assign node264 = (inp[8]) ? 3'b001 : 3'b101;
												assign node267 = (inp[8]) ? 3'b101 : 3'b001;
										assign node271 = (inp[8]) ? node279 : node272;
											assign node272 = (inp[5]) ? node276 : node273;
												assign node273 = (inp[10]) ? 3'b001 : 3'b101;
												assign node276 = (inp[10]) ? 3'b101 : 3'b001;
											assign node279 = (inp[5]) ? node281 : 3'b001;
												assign node281 = (inp[10]) ? 3'b001 : 3'b101;
									assign node284 = (inp[8]) ? node292 : node285;
										assign node285 = (inp[10]) ? node289 : node286;
											assign node286 = (inp[5]) ? 3'b001 : 3'b101;
											assign node289 = (inp[5]) ? 3'b101 : 3'b001;
										assign node292 = (inp[2]) ? node294 : 3'b101;
											assign node294 = (inp[5]) ? node298 : node295;
												assign node295 = (inp[10]) ? 3'b101 : 3'b001;
												assign node298 = (inp[10]) ? 3'b001 : 3'b101;
					assign node303 = (inp[4]) ? node395 : node304;
						assign node304 = (inp[1]) ? node330 : node305;
							assign node305 = (inp[8]) ? node321 : node306;
								assign node306 = (inp[7]) ? node318 : node307;
									assign node307 = (inp[5]) ? node313 : node308;
										assign node308 = (inp[11]) ? node310 : 3'b010;
											assign node310 = (inp[2]) ? 3'b010 : 3'b110;
										assign node313 = (inp[11]) ? 3'b001 : node314;
											assign node314 = (inp[2]) ? 3'b010 : 3'b110;
									assign node318 = (inp[10]) ? 3'b110 : 3'b010;
								assign node321 = (inp[7]) ? node327 : node322;
									assign node322 = (inp[5]) ? node324 : 3'b010;
										assign node324 = (inp[2]) ? 3'b010 : 3'b110;
									assign node327 = (inp[10]) ? 3'b001 : 3'b101;
							assign node330 = (inp[7]) ? node370 : node331;
								assign node331 = (inp[5]) ? node347 : node332;
									assign node332 = (inp[2]) ? node338 : node333;
										assign node333 = (inp[8]) ? node335 : 3'b101;
											assign node335 = (inp[10]) ? 3'b011 : 3'b101;
										assign node338 = (inp[11]) ? node340 : 3'b001;
											assign node340 = (inp[10]) ? node344 : node341;
												assign node341 = (inp[8]) ? 3'b001 : 3'b101;
												assign node344 = (inp[8]) ? 3'b101 : 3'b011;
									assign node347 = (inp[2]) ? node355 : node348;
										assign node348 = (inp[10]) ? node352 : node349;
											assign node349 = (inp[8]) ? 3'b011 : 3'b101;
											assign node352 = (inp[8]) ? 3'b101 : 3'b011;
										assign node355 = (inp[11]) ? node363 : node356;
											assign node356 = (inp[8]) ? node360 : node357;
												assign node357 = (inp[10]) ? 3'b111 : 3'b011;
												assign node360 = (inp[10]) ? 3'b011 : 3'b111;
											assign node363 = (inp[8]) ? node367 : node364;
												assign node364 = (inp[10]) ? 3'b111 : 3'b011;
												assign node367 = (inp[10]) ? 3'b011 : 3'b111;
								assign node370 = (inp[2]) ? node378 : node371;
									assign node371 = (inp[8]) ? node375 : node372;
										assign node372 = (inp[10]) ? 3'b101 : 3'b010;
										assign node375 = (inp[10]) ? 3'b010 : 3'b101;
									assign node378 = (inp[5]) ? node386 : node379;
										assign node379 = (inp[11]) ? node381 : 3'b110;
											assign node381 = (inp[8]) ? 3'b010 : node382;
												assign node382 = (inp[10]) ? 3'b110 : 3'b010;
										assign node386 = (inp[10]) ? node392 : node387;
											assign node387 = (inp[11]) ? node389 : 3'b001;
												assign node389 = (inp[8]) ? 3'b110 : 3'b010;
											assign node392 = (inp[11]) ? 3'b101 : 3'b110;
						assign node395 = (inp[7]) ? node441 : node396;
							assign node396 = (inp[1]) ? node430 : node397;
								assign node397 = (inp[2]) ? node417 : node398;
									assign node398 = (inp[11]) ? node410 : node399;
										assign node399 = (inp[10]) ? node403 : node400;
											assign node400 = (inp[5]) ? 3'b101 : 3'b110;
											assign node403 = (inp[8]) ? node407 : node404;
												assign node404 = (inp[5]) ? 3'b011 : 3'b101;
												assign node407 = (inp[5]) ? 3'b101 : 3'b001;
										assign node410 = (inp[5]) ? 3'b011 : node411;
											assign node411 = (inp[10]) ? node413 : 3'b001;
												assign node413 = (inp[8]) ? 3'b001 : 3'b101;
									assign node417 = (inp[5]) ? node425 : node418;
										assign node418 = (inp[10]) ? node422 : node419;
											assign node419 = (inp[8]) ? 3'b011 : 3'b101;
											assign node422 = (inp[8]) ? 3'b101 : 3'b111;
										assign node425 = (inp[10]) ? 3'b111 : node426;
											assign node426 = (inp[8]) ? 3'b011 : 3'b111;
								assign node430 = (inp[2]) ? 3'b111 : node431;
									assign node431 = (inp[8]) ? node433 : 3'b111;
										assign node433 = (inp[5]) ? node435 : 3'b111;
											assign node435 = (inp[10]) ? 3'b111 : node436;
												assign node436 = (inp[11]) ? 3'b111 : 3'b011;
							assign node441 = (inp[1]) ? node491 : node442;
								assign node442 = (inp[5]) ? node466 : node443;
									assign node443 = (inp[10]) ? node453 : node444;
										assign node444 = (inp[11]) ? node446 : 3'b110;
											assign node446 = (inp[8]) ? node450 : node447;
												assign node447 = (inp[2]) ? 3'b100 : 3'b000;
												assign node450 = (inp[2]) ? 3'b001 : 3'b101;
										assign node453 = (inp[8]) ? node461 : node454;
											assign node454 = (inp[2]) ? node458 : node455;
												assign node455 = (inp[11]) ? 3'b110 : 3'b100;
												assign node458 = (inp[11]) ? 3'b011 : 3'b001;
											assign node461 = (inp[2]) ? 3'b110 : node462;
												assign node462 = (inp[11]) ? 3'b010 : 3'b110;
									assign node466 = (inp[11]) ? node480 : node467;
										assign node467 = (inp[2]) ? node473 : node468;
											assign node468 = (inp[8]) ? 3'b110 : node469;
												assign node469 = (inp[10]) ? 3'b101 : 3'b110;
											assign node473 = (inp[8]) ? node477 : node474;
												assign node474 = (inp[10]) ? 3'b001 : 3'b111;
												assign node477 = (inp[10]) ? 3'b111 : 3'b001;
										assign node480 = (inp[10]) ? node484 : node481;
											assign node481 = (inp[2]) ? 3'b101 : 3'b001;
											assign node484 = (inp[8]) ? node488 : node485;
												assign node485 = (inp[2]) ? 3'b011 : 3'b111;
												assign node488 = (inp[2]) ? 3'b111 : 3'b011;
								assign node491 = (inp[2]) ? node503 : node492;
									assign node492 = (inp[5]) ? node494 : 3'b001;
										assign node494 = (inp[11]) ? node496 : 3'b101;
											assign node496 = (inp[10]) ? node500 : node497;
												assign node497 = (inp[8]) ? 3'b101 : 3'b011;
												assign node500 = (inp[8]) ? 3'b011 : 3'b111;
									assign node503 = (inp[5]) ? node511 : node504;
										assign node504 = (inp[8]) ? node506 : 3'b111;
											assign node506 = (inp[10]) ? 3'b111 : node507;
												assign node507 = (inp[11]) ? 3'b111 : 3'b101;
										assign node511 = (inp[8]) ? node517 : node512;
											assign node512 = (inp[11]) ? 3'b111 : node513;
												assign node513 = (inp[10]) ? 3'b111 : 3'b011;
											assign node517 = (inp[11]) ? 3'b011 : node518;
												assign node518 = (inp[10]) ? 3'b011 : 3'b101;
		assign node522 = (inp[0]) ? node524 : 3'b000;
			assign node524 = (inp[3]) ? node526 : 3'b000;
				assign node526 = (inp[9]) ? node528 : 3'b000;
					assign node528 = (inp[4]) ? node560 : node529;
						assign node529 = (inp[7]) ? 3'b000 : node530;
							assign node530 = (inp[2]) ? node538 : node531;
								assign node531 = (inp[5]) ? node533 : 3'b000;
									assign node533 = (inp[8]) ? 3'b000 : node534;
										assign node534 = (inp[11]) ? 3'b010 : 3'b000;
								assign node538 = (inp[1]) ? node544 : node539;
									assign node539 = (inp[8]) ? 3'b000 : node540;
										assign node540 = (inp[5]) ? 3'b010 : 3'b000;
									assign node544 = (inp[10]) ? node554 : node545;
										assign node545 = (inp[5]) ? node549 : node546;
											assign node546 = (inp[8]) ? 3'b100 : 3'b000;
											assign node549 = (inp[8]) ? 3'b000 : node550;
												assign node550 = (inp[11]) ? 3'b010 : 3'b000;
										assign node554 = (inp[5]) ? 3'b100 : node555;
											assign node555 = (inp[8]) ? 3'b000 : 3'b100;
						assign node560 = (inp[7]) ? node598 : node561;
							assign node561 = (inp[8]) ? node583 : node562;
								assign node562 = (inp[1]) ? node566 : node563;
									assign node563 = (inp[10]) ? 3'b110 : 3'b100;
									assign node566 = (inp[10]) ? node574 : node567;
										assign node567 = (inp[2]) ? node569 : 3'b110;
											assign node569 = (inp[5]) ? node571 : 3'b110;
												assign node571 = (inp[11]) ? 3'b101 : 3'b001;
										assign node574 = (inp[2]) ? node576 : 3'b001;
											assign node576 = (inp[11]) ? node580 : node577;
												assign node577 = (inp[5]) ? 3'b101 : 3'b111;
												assign node580 = (inp[5]) ? 3'b011 : 3'b111;
								assign node583 = (inp[1]) ? node587 : node584;
									assign node584 = (inp[10]) ? 3'b010 : 3'b000;
									assign node587 = (inp[10]) ? node591 : node588;
										assign node588 = (inp[2]) ? 3'b110 : 3'b010;
										assign node591 = (inp[5]) ? node595 : node592;
											assign node592 = (inp[2]) ? 3'b110 : 3'b101;
											assign node595 = (inp[2]) ? 3'b001 : 3'b101;
							assign node598 = (inp[1]) ? node600 : 3'b000;
								assign node600 = (inp[2]) ? node602 : 3'b000;
									assign node602 = (inp[8]) ? node610 : node603;
										assign node603 = (inp[10]) ? node607 : node604;
											assign node604 = (inp[5]) ? 3'b010 : 3'b100;
											assign node607 = (inp[5]) ? 3'b110 : 3'b010;
										assign node610 = (inp[10]) ? node614 : node611;
											assign node611 = (inp[5]) ? 3'b100 : 3'b000;
											assign node614 = (inp[5]) ? 3'b010 : 3'b000;

endmodule