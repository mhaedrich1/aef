module dtc_split25_bm62 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node14;
	wire [4-1:0] node19;
	wire [4-1:0] node20;
	wire [4-1:0] node24;
	wire [4-1:0] node25;
	wire [4-1:0] node27;
	wire [4-1:0] node30;
	wire [4-1:0] node31;
	wire [4-1:0] node34;
	wire [4-1:0] node35;
	wire [4-1:0] node38;
	wire [4-1:0] node41;
	wire [4-1:0] node42;
	wire [4-1:0] node43;
	wire [4-1:0] node46;
	wire [4-1:0] node47;
	wire [4-1:0] node49;
	wire [4-1:0] node52;
	wire [4-1:0] node55;
	wire [4-1:0] node56;
	wire [4-1:0] node57;
	wire [4-1:0] node59;
	wire [4-1:0] node62;
	wire [4-1:0] node64;
	wire [4-1:0] node67;
	wire [4-1:0] node68;
	wire [4-1:0] node71;
	wire [4-1:0] node74;
	wire [4-1:0] node75;
	wire [4-1:0] node76;
	wire [4-1:0] node77;
	wire [4-1:0] node80;
	wire [4-1:0] node83;
	wire [4-1:0] node84;
	wire [4-1:0] node85;
	wire [4-1:0] node86;
	wire [4-1:0] node90;
	wire [4-1:0] node93;
	wire [4-1:0] node96;
	wire [4-1:0] node97;
	wire [4-1:0] node98;
	wire [4-1:0] node99;
	wire [4-1:0] node103;
	wire [4-1:0] node105;
	wire [4-1:0] node108;
	wire [4-1:0] node109;
	wire [4-1:0] node111;
	wire [4-1:0] node114;
	wire [4-1:0] node115;
	wire [4-1:0] node116;
	wire [4-1:0] node119;
	wire [4-1:0] node123;
	wire [4-1:0] node124;
	wire [4-1:0] node125;
	wire [4-1:0] node126;
	wire [4-1:0] node127;
	wire [4-1:0] node128;
	wire [4-1:0] node131;
	wire [4-1:0] node134;
	wire [4-1:0] node137;
	wire [4-1:0] node138;
	wire [4-1:0] node139;
	wire [4-1:0] node142;
	wire [4-1:0] node145;
	wire [4-1:0] node147;
	wire [4-1:0] node150;
	wire [4-1:0] node151;
	wire [4-1:0] node152;
	wire [4-1:0] node154;
	wire [4-1:0] node156;
	wire [4-1:0] node159;
	wire [4-1:0] node161;
	wire [4-1:0] node162;
	wire [4-1:0] node166;
	wire [4-1:0] node168;
	wire [4-1:0] node169;
	wire [4-1:0] node170;
	wire [4-1:0] node173;
	wire [4-1:0] node177;
	wire [4-1:0] node178;
	wire [4-1:0] node179;
	wire [4-1:0] node180;
	wire [4-1:0] node183;
	wire [4-1:0] node185;
	wire [4-1:0] node186;
	wire [4-1:0] node190;
	wire [4-1:0] node191;
	wire [4-1:0] node193;
	wire [4-1:0] node196;
	wire [4-1:0] node198;
	wire [4-1:0] node201;
	wire [4-1:0] node202;
	wire [4-1:0] node203;
	wire [4-1:0] node206;
	wire [4-1:0] node208;
	wire [4-1:0] node211;
	wire [4-1:0] node212;
	wire [4-1:0] node213;
	wire [4-1:0] node217;
	wire [4-1:0] node219;
	wire [4-1:0] node222;
	wire [4-1:0] node223;
	wire [4-1:0] node224;
	wire [4-1:0] node225;
	wire [4-1:0] node226;
	wire [4-1:0] node227;
	wire [4-1:0] node229;
	wire [4-1:0] node232;
	wire [4-1:0] node233;
	wire [4-1:0] node237;
	wire [4-1:0] node238;
	wire [4-1:0] node239;
	wire [4-1:0] node244;
	wire [4-1:0] node245;
	wire [4-1:0] node246;
	wire [4-1:0] node248;
	wire [4-1:0] node252;
	wire [4-1:0] node253;
	wire [4-1:0] node257;
	wire [4-1:0] node258;
	wire [4-1:0] node259;
	wire [4-1:0] node260;
	wire [4-1:0] node264;
	wire [4-1:0] node265;
	wire [4-1:0] node268;
	wire [4-1:0] node269;
	wire [4-1:0] node271;
	wire [4-1:0] node274;
	wire [4-1:0] node277;
	wire [4-1:0] node278;
	wire [4-1:0] node279;
	wire [4-1:0] node282;
	wire [4-1:0] node283;
	wire [4-1:0] node284;
	wire [4-1:0] node289;
	wire [4-1:0] node290;
	wire [4-1:0] node291;
	wire [4-1:0] node293;
	wire [4-1:0] node297;
	wire [4-1:0] node298;
	wire [4-1:0] node299;
	wire [4-1:0] node302;
	wire [4-1:0] node306;
	wire [4-1:0] node307;
	wire [4-1:0] node308;
	wire [4-1:0] node309;
	wire [4-1:0] node310;
	wire [4-1:0] node312;
	wire [4-1:0] node315;
	wire [4-1:0] node318;
	wire [4-1:0] node319;
	wire [4-1:0] node320;
	wire [4-1:0] node321;
	wire [4-1:0] node324;
	wire [4-1:0] node327;
	wire [4-1:0] node330;
	wire [4-1:0] node331;
	wire [4-1:0] node334;
	wire [4-1:0] node337;
	wire [4-1:0] node338;
	wire [4-1:0] node340;
	wire [4-1:0] node341;
	wire [4-1:0] node343;
	wire [4-1:0] node347;
	wire [4-1:0] node348;
	wire [4-1:0] node349;
	wire [4-1:0] node351;
	wire [4-1:0] node354;
	wire [4-1:0] node357;
	wire [4-1:0] node360;
	wire [4-1:0] node361;
	wire [4-1:0] node362;
	wire [4-1:0] node363;
	wire [4-1:0] node366;
	wire [4-1:0] node368;
	wire [4-1:0] node371;
	wire [4-1:0] node374;
	wire [4-1:0] node375;
	wire [4-1:0] node376;
	wire [4-1:0] node378;
	wire [4-1:0] node380;
	wire [4-1:0] node383;
	wire [4-1:0] node384;
	wire [4-1:0] node387;
	wire [4-1:0] node388;
	wire [4-1:0] node391;
	wire [4-1:0] node394;
	wire [4-1:0] node395;
	wire [4-1:0] node398;
	wire [4-1:0] node399;
	wire [4-1:0] node402;
	wire [4-1:0] node405;
	wire [4-1:0] node406;
	wire [4-1:0] node407;
	wire [4-1:0] node408;
	wire [4-1:0] node409;
	wire [4-1:0] node410;
	wire [4-1:0] node411;
	wire [4-1:0] node412;
	wire [4-1:0] node417;
	wire [4-1:0] node418;
	wire [4-1:0] node419;
	wire [4-1:0] node422;
	wire [4-1:0] node426;
	wire [4-1:0] node427;
	wire [4-1:0] node428;
	wire [4-1:0] node430;
	wire [4-1:0] node432;
	wire [4-1:0] node435;
	wire [4-1:0] node436;
	wire [4-1:0] node438;
	wire [4-1:0] node442;
	wire [4-1:0] node445;
	wire [4-1:0] node446;
	wire [4-1:0] node447;
	wire [4-1:0] node448;
	wire [4-1:0] node451;
	wire [4-1:0] node452;
	wire [4-1:0] node453;
	wire [4-1:0] node457;
	wire [4-1:0] node459;
	wire [4-1:0] node462;
	wire [4-1:0] node463;
	wire [4-1:0] node466;
	wire [4-1:0] node469;
	wire [4-1:0] node470;
	wire [4-1:0] node471;
	wire [4-1:0] node473;
	wire [4-1:0] node476;
	wire [4-1:0] node477;
	wire [4-1:0] node481;
	wire [4-1:0] node482;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node490;
	wire [4-1:0] node491;
	wire [4-1:0] node492;
	wire [4-1:0] node493;
	wire [4-1:0] node494;
	wire [4-1:0] node495;
	wire [4-1:0] node498;
	wire [4-1:0] node500;
	wire [4-1:0] node503;
	wire [4-1:0] node504;
	wire [4-1:0] node505;
	wire [4-1:0] node509;
	wire [4-1:0] node512;
	wire [4-1:0] node514;
	wire [4-1:0] node516;
	wire [4-1:0] node519;
	wire [4-1:0] node520;
	wire [4-1:0] node521;
	wire [4-1:0] node523;
	wire [4-1:0] node526;
	wire [4-1:0] node529;
	wire [4-1:0] node530;
	wire [4-1:0] node531;
	wire [4-1:0] node532;
	wire [4-1:0] node537;
	wire [4-1:0] node539;
	wire [4-1:0] node541;
	wire [4-1:0] node544;
	wire [4-1:0] node545;
	wire [4-1:0] node546;
	wire [4-1:0] node547;
	wire [4-1:0] node549;
	wire [4-1:0] node552;
	wire [4-1:0] node553;
	wire [4-1:0] node557;
	wire [4-1:0] node558;
	wire [4-1:0] node559;
	wire [4-1:0] node561;
	wire [4-1:0] node564;
	wire [4-1:0] node567;
	wire [4-1:0] node568;
	wire [4-1:0] node572;
	wire [4-1:0] node573;
	wire [4-1:0] node574;
	wire [4-1:0] node575;
	wire [4-1:0] node579;
	wire [4-1:0] node581;
	wire [4-1:0] node583;
	wire [4-1:0] node586;
	wire [4-1:0] node587;
	wire [4-1:0] node588;
	wire [4-1:0] node590;
	wire [4-1:0] node595;
	wire [4-1:0] node596;
	wire [4-1:0] node597;
	wire [4-1:0] node598;
	wire [4-1:0] node599;
	wire [4-1:0] node600;
	wire [4-1:0] node602;
	wire [4-1:0] node604;
	wire [4-1:0] node607;
	wire [4-1:0] node608;
	wire [4-1:0] node612;
	wire [4-1:0] node613;
	wire [4-1:0] node615;
	wire [4-1:0] node616;
	wire [4-1:0] node620;
	wire [4-1:0] node621;
	wire [4-1:0] node625;
	wire [4-1:0] node626;
	wire [4-1:0] node628;
	wire [4-1:0] node630;
	wire [4-1:0] node631;
	wire [4-1:0] node634;
	wire [4-1:0] node637;
	wire [4-1:0] node639;
	wire [4-1:0] node640;
	wire [4-1:0] node644;
	wire [4-1:0] node645;
	wire [4-1:0] node646;
	wire [4-1:0] node647;
	wire [4-1:0] node649;
	wire [4-1:0] node652;
	wire [4-1:0] node655;
	wire [4-1:0] node656;
	wire [4-1:0] node657;
	wire [4-1:0] node658;
	wire [4-1:0] node661;
	wire [4-1:0] node665;
	wire [4-1:0] node668;
	wire [4-1:0] node669;
	wire [4-1:0] node670;
	wire [4-1:0] node672;
	wire [4-1:0] node675;
	wire [4-1:0] node677;
	wire [4-1:0] node680;
	wire [4-1:0] node681;
	wire [4-1:0] node683;
	wire [4-1:0] node686;
	wire [4-1:0] node687;
	wire [4-1:0] node691;
	wire [4-1:0] node692;
	wire [4-1:0] node693;
	wire [4-1:0] node694;
	wire [4-1:0] node695;
	wire [4-1:0] node697;
	wire [4-1:0] node701;
	wire [4-1:0] node702;
	wire [4-1:0] node704;
	wire [4-1:0] node706;
	wire [4-1:0] node709;
	wire [4-1:0] node711;
	wire [4-1:0] node713;
	wire [4-1:0] node716;
	wire [4-1:0] node717;
	wire [4-1:0] node718;
	wire [4-1:0] node720;
	wire [4-1:0] node723;
	wire [4-1:0] node725;
	wire [4-1:0] node727;
	wire [4-1:0] node730;
	wire [4-1:0] node731;
	wire [4-1:0] node732;
	wire [4-1:0] node736;
	wire [4-1:0] node737;
	wire [4-1:0] node739;
	wire [4-1:0] node743;
	wire [4-1:0] node744;
	wire [4-1:0] node745;
	wire [4-1:0] node746;
	wire [4-1:0] node748;
	wire [4-1:0] node750;
	wire [4-1:0] node753;
	wire [4-1:0] node754;
	wire [4-1:0] node755;
	wire [4-1:0] node760;
	wire [4-1:0] node761;
	wire [4-1:0] node762;
	wire [4-1:0] node764;
	wire [4-1:0] node768;
	wire [4-1:0] node769;
	wire [4-1:0] node770;
	wire [4-1:0] node775;
	wire [4-1:0] node776;
	wire [4-1:0] node777;
	wire [4-1:0] node780;
	wire [4-1:0] node781;
	wire [4-1:0] node784;
	wire [4-1:0] node787;
	wire [4-1:0] node788;
	wire [4-1:0] node789;
	wire [4-1:0] node790;
	wire [4-1:0] node793;
	wire [4-1:0] node798;
	wire [4-1:0] node799;
	wire [4-1:0] node800;
	wire [4-1:0] node801;
	wire [4-1:0] node802;
	wire [4-1:0] node803;
	wire [4-1:0] node804;
	wire [4-1:0] node805;
	wire [4-1:0] node807;
	wire [4-1:0] node809;
	wire [4-1:0] node812;
	wire [4-1:0] node813;
	wire [4-1:0] node814;
	wire [4-1:0] node819;
	wire [4-1:0] node820;
	wire [4-1:0] node823;
	wire [4-1:0] node824;
	wire [4-1:0] node825;
	wire [4-1:0] node830;
	wire [4-1:0] node831;
	wire [4-1:0] node833;
	wire [4-1:0] node836;
	wire [4-1:0] node837;
	wire [4-1:0] node840;
	wire [4-1:0] node842;
	wire [4-1:0] node845;
	wire [4-1:0] node846;
	wire [4-1:0] node847;
	wire [4-1:0] node848;
	wire [4-1:0] node852;
	wire [4-1:0] node854;
	wire [4-1:0] node856;
	wire [4-1:0] node858;
	wire [4-1:0] node861;
	wire [4-1:0] node862;
	wire [4-1:0] node863;
	wire [4-1:0] node864;
	wire [4-1:0] node868;
	wire [4-1:0] node870;
	wire [4-1:0] node873;
	wire [4-1:0] node874;
	wire [4-1:0] node877;
	wire [4-1:0] node878;
	wire [4-1:0] node879;
	wire [4-1:0] node882;
	wire [4-1:0] node886;
	wire [4-1:0] node887;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node891;
	wire [4-1:0] node894;
	wire [4-1:0] node895;
	wire [4-1:0] node898;
	wire [4-1:0] node900;
	wire [4-1:0] node903;
	wire [4-1:0] node904;
	wire [4-1:0] node905;
	wire [4-1:0] node908;
	wire [4-1:0] node909;
	wire [4-1:0] node913;
	wire [4-1:0] node914;
	wire [4-1:0] node916;
	wire [4-1:0] node918;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node924;
	wire [4-1:0] node925;
	wire [4-1:0] node928;
	wire [4-1:0] node930;
	wire [4-1:0] node933;
	wire [4-1:0] node934;
	wire [4-1:0] node935;
	wire [4-1:0] node938;
	wire [4-1:0] node941;
	wire [4-1:0] node943;
	wire [4-1:0] node946;
	wire [4-1:0] node947;
	wire [4-1:0] node948;
	wire [4-1:0] node951;
	wire [4-1:0] node954;
	wire [4-1:0] node956;
	wire [4-1:0] node958;
	wire [4-1:0] node960;
	wire [4-1:0] node963;
	wire [4-1:0] node964;
	wire [4-1:0] node965;
	wire [4-1:0] node966;
	wire [4-1:0] node967;
	wire [4-1:0] node968;
	wire [4-1:0] node969;
	wire [4-1:0] node974;
	wire [4-1:0] node975;
	wire [4-1:0] node978;
	wire [4-1:0] node980;
	wire [4-1:0] node982;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node987;
	wire [4-1:0] node989;
	wire [4-1:0] node993;
	wire [4-1:0] node994;
	wire [4-1:0] node995;
	wire [4-1:0] node996;
	wire [4-1:0] node1000;
	wire [4-1:0] node1001;
	wire [4-1:0] node1005;
	wire [4-1:0] node1006;
	wire [4-1:0] node1010;
	wire [4-1:0] node1011;
	wire [4-1:0] node1012;
	wire [4-1:0] node1014;
	wire [4-1:0] node1015;
	wire [4-1:0] node1016;
	wire [4-1:0] node1021;
	wire [4-1:0] node1022;
	wire [4-1:0] node1024;
	wire [4-1:0] node1028;
	wire [4-1:0] node1029;
	wire [4-1:0] node1030;
	wire [4-1:0] node1032;
	wire [4-1:0] node1033;
	wire [4-1:0] node1036;
	wire [4-1:0] node1039;
	wire [4-1:0] node1040;
	wire [4-1:0] node1041;
	wire [4-1:0] node1046;
	wire [4-1:0] node1047;
	wire [4-1:0] node1050;
	wire [4-1:0] node1053;
	wire [4-1:0] node1054;
	wire [4-1:0] node1055;
	wire [4-1:0] node1056;
	wire [4-1:0] node1057;
	wire [4-1:0] node1061;
	wire [4-1:0] node1063;
	wire [4-1:0] node1065;
	wire [4-1:0] node1068;
	wire [4-1:0] node1069;
	wire [4-1:0] node1070;
	wire [4-1:0] node1071;
	wire [4-1:0] node1075;
	wire [4-1:0] node1078;
	wire [4-1:0] node1080;
	wire [4-1:0] node1081;
	wire [4-1:0] node1085;
	wire [4-1:0] node1086;
	wire [4-1:0] node1087;
	wire [4-1:0] node1088;
	wire [4-1:0] node1089;
	wire [4-1:0] node1093;
	wire [4-1:0] node1096;
	wire [4-1:0] node1097;
	wire [4-1:0] node1100;
	wire [4-1:0] node1103;
	wire [4-1:0] node1104;
	wire [4-1:0] node1105;
	wire [4-1:0] node1106;
	wire [4-1:0] node1107;
	wire [4-1:0] node1111;
	wire [4-1:0] node1114;
	wire [4-1:0] node1116;
	wire [4-1:0] node1119;
	wire [4-1:0] node1120;
	wire [4-1:0] node1121;
	wire [4-1:0] node1125;
	wire [4-1:0] node1126;
	wire [4-1:0] node1129;
	wire [4-1:0] node1132;
	wire [4-1:0] node1133;
	wire [4-1:0] node1134;
	wire [4-1:0] node1135;
	wire [4-1:0] node1136;
	wire [4-1:0] node1137;
	wire [4-1:0] node1138;
	wire [4-1:0] node1141;
	wire [4-1:0] node1142;
	wire [4-1:0] node1143;
	wire [4-1:0] node1148;
	wire [4-1:0] node1149;
	wire [4-1:0] node1152;
	wire [4-1:0] node1153;
	wire [4-1:0] node1155;
	wire [4-1:0] node1159;
	wire [4-1:0] node1160;
	wire [4-1:0] node1161;
	wire [4-1:0] node1162;
	wire [4-1:0] node1164;
	wire [4-1:0] node1170;
	wire [4-1:0] node1171;
	wire [4-1:0] node1172;
	wire [4-1:0] node1175;
	wire [4-1:0] node1176;
	wire [4-1:0] node1177;
	wire [4-1:0] node1181;
	wire [4-1:0] node1182;
	wire [4-1:0] node1186;
	wire [4-1:0] node1187;
	wire [4-1:0] node1189;
	wire [4-1:0] node1190;
	wire [4-1:0] node1192;
	wire [4-1:0] node1196;
	wire [4-1:0] node1199;
	wire [4-1:0] node1200;
	wire [4-1:0] node1201;
	wire [4-1:0] node1202;
	wire [4-1:0] node1203;
	wire [4-1:0] node1204;
	wire [4-1:0] node1205;
	wire [4-1:0] node1208;
	wire [4-1:0] node1212;
	wire [4-1:0] node1215;
	wire [4-1:0] node1217;
	wire [4-1:0] node1220;
	wire [4-1:0] node1221;
	wire [4-1:0] node1222;
	wire [4-1:0] node1224;
	wire [4-1:0] node1226;
	wire [4-1:0] node1229;
	wire [4-1:0] node1230;
	wire [4-1:0] node1234;
	wire [4-1:0] node1235;
	wire [4-1:0] node1236;
	wire [4-1:0] node1239;
	wire [4-1:0] node1240;
	wire [4-1:0] node1243;
	wire [4-1:0] node1247;
	wire [4-1:0] node1248;
	wire [4-1:0] node1249;
	wire [4-1:0] node1250;
	wire [4-1:0] node1253;
	wire [4-1:0] node1256;
	wire [4-1:0] node1257;
	wire [4-1:0] node1259;
	wire [4-1:0] node1263;
	wire [4-1:0] node1264;
	wire [4-1:0] node1265;
	wire [4-1:0] node1266;
	wire [4-1:0] node1270;
	wire [4-1:0] node1273;
	wire [4-1:0] node1274;
	wire [4-1:0] node1276;
	wire [4-1:0] node1280;
	wire [4-1:0] node1281;
	wire [4-1:0] node1282;
	wire [4-1:0] node1283;
	wire [4-1:0] node1284;
	wire [4-1:0] node1285;
	wire [4-1:0] node1286;
	wire [4-1:0] node1290;
	wire [4-1:0] node1293;
	wire [4-1:0] node1294;
	wire [4-1:0] node1297;
	wire [4-1:0] node1299;
	wire [4-1:0] node1301;
	wire [4-1:0] node1304;
	wire [4-1:0] node1305;
	wire [4-1:0] node1306;
	wire [4-1:0] node1307;
	wire [4-1:0] node1311;
	wire [4-1:0] node1313;
	wire [4-1:0] node1316;
	wire [4-1:0] node1317;
	wire [4-1:0] node1321;
	wire [4-1:0] node1322;
	wire [4-1:0] node1323;
	wire [4-1:0] node1324;
	wire [4-1:0] node1325;
	wire [4-1:0] node1329;
	wire [4-1:0] node1330;
	wire [4-1:0] node1333;
	wire [4-1:0] node1334;
	wire [4-1:0] node1337;
	wire [4-1:0] node1340;
	wire [4-1:0] node1341;
	wire [4-1:0] node1343;
	wire [4-1:0] node1344;
	wire [4-1:0] node1348;
	wire [4-1:0] node1349;
	wire [4-1:0] node1352;
	wire [4-1:0] node1355;
	wire [4-1:0] node1356;
	wire [4-1:0] node1359;
	wire [4-1:0] node1360;
	wire [4-1:0] node1362;
	wire [4-1:0] node1363;
	wire [4-1:0] node1366;
	wire [4-1:0] node1369;
	wire [4-1:0] node1372;
	wire [4-1:0] node1373;
	wire [4-1:0] node1374;
	wire [4-1:0] node1375;
	wire [4-1:0] node1376;
	wire [4-1:0] node1377;
	wire [4-1:0] node1378;
	wire [4-1:0] node1383;
	wire [4-1:0] node1385;
	wire [4-1:0] node1387;
	wire [4-1:0] node1390;
	wire [4-1:0] node1392;
	wire [4-1:0] node1394;
	wire [4-1:0] node1396;
	wire [4-1:0] node1399;
	wire [4-1:0] node1400;
	wire [4-1:0] node1402;
	wire [4-1:0] node1403;
	wire [4-1:0] node1407;
	wire [4-1:0] node1409;
	wire [4-1:0] node1411;
	wire [4-1:0] node1412;
	wire [4-1:0] node1415;
	wire [4-1:0] node1418;
	wire [4-1:0] node1419;
	wire [4-1:0] node1420;
	wire [4-1:0] node1421;
	wire [4-1:0] node1424;
	wire [4-1:0] node1426;
	wire [4-1:0] node1429;
	wire [4-1:0] node1430;
	wire [4-1:0] node1431;
	wire [4-1:0] node1434;
	wire [4-1:0] node1437;
	wire [4-1:0] node1439;
	wire [4-1:0] node1442;
	wire [4-1:0] node1443;
	wire [4-1:0] node1444;
	wire [4-1:0] node1447;
	wire [4-1:0] node1450;
	wire [4-1:0] node1451;
	wire [4-1:0] node1452;
	wire [4-1:0] node1455;
	wire [4-1:0] node1457;
	wire [4-1:0] node1461;
	wire [4-1:0] node1462;
	wire [4-1:0] node1463;
	wire [4-1:0] node1464;
	wire [4-1:0] node1465;
	wire [4-1:0] node1466;
	wire [4-1:0] node1467;
	wire [4-1:0] node1468;
	wire [4-1:0] node1469;
	wire [4-1:0] node1471;
	wire [4-1:0] node1474;
	wire [4-1:0] node1477;
	wire [4-1:0] node1479;
	wire [4-1:0] node1480;
	wire [4-1:0] node1481;
	wire [4-1:0] node1485;
	wire [4-1:0] node1486;
	wire [4-1:0] node1490;
	wire [4-1:0] node1491;
	wire [4-1:0] node1493;
	wire [4-1:0] node1494;
	wire [4-1:0] node1498;
	wire [4-1:0] node1499;
	wire [4-1:0] node1502;
	wire [4-1:0] node1504;
	wire [4-1:0] node1507;
	wire [4-1:0] node1508;
	wire [4-1:0] node1509;
	wire [4-1:0] node1510;
	wire [4-1:0] node1512;
	wire [4-1:0] node1515;
	wire [4-1:0] node1518;
	wire [4-1:0] node1519;
	wire [4-1:0] node1522;
	wire [4-1:0] node1523;
	wire [4-1:0] node1525;
	wire [4-1:0] node1529;
	wire [4-1:0] node1530;
	wire [4-1:0] node1531;
	wire [4-1:0] node1532;
	wire [4-1:0] node1533;
	wire [4-1:0] node1536;
	wire [4-1:0] node1541;
	wire [4-1:0] node1543;
	wire [4-1:0] node1546;
	wire [4-1:0] node1547;
	wire [4-1:0] node1548;
	wire [4-1:0] node1549;
	wire [4-1:0] node1550;
	wire [4-1:0] node1552;
	wire [4-1:0] node1554;
	wire [4-1:0] node1557;
	wire [4-1:0] node1558;
	wire [4-1:0] node1562;
	wire [4-1:0] node1563;
	wire [4-1:0] node1565;
	wire [4-1:0] node1566;
	wire [4-1:0] node1571;
	wire [4-1:0] node1572;
	wire [4-1:0] node1573;
	wire [4-1:0] node1574;
	wire [4-1:0] node1575;
	wire [4-1:0] node1581;
	wire [4-1:0] node1582;
	wire [4-1:0] node1583;
	wire [4-1:0] node1586;
	wire [4-1:0] node1588;
	wire [4-1:0] node1592;
	wire [4-1:0] node1593;
	wire [4-1:0] node1594;
	wire [4-1:0] node1595;
	wire [4-1:0] node1598;
	wire [4-1:0] node1600;
	wire [4-1:0] node1602;
	wire [4-1:0] node1606;
	wire [4-1:0] node1607;
	wire [4-1:0] node1608;
	wire [4-1:0] node1611;
	wire [4-1:0] node1612;
	wire [4-1:0] node1614;
	wire [4-1:0] node1618;
	wire [4-1:0] node1619;
	wire [4-1:0] node1622;
	wire [4-1:0] node1624;
	wire [4-1:0] node1627;
	wire [4-1:0] node1628;
	wire [4-1:0] node1629;
	wire [4-1:0] node1630;
	wire [4-1:0] node1631;
	wire [4-1:0] node1632;
	wire [4-1:0] node1633;
	wire [4-1:0] node1636;
	wire [4-1:0] node1638;
	wire [4-1:0] node1641;
	wire [4-1:0] node1642;
	wire [4-1:0] node1646;
	wire [4-1:0] node1647;
	wire [4-1:0] node1648;
	wire [4-1:0] node1649;
	wire [4-1:0] node1654;
	wire [4-1:0] node1655;
	wire [4-1:0] node1657;
	wire [4-1:0] node1661;
	wire [4-1:0] node1662;
	wire [4-1:0] node1663;
	wire [4-1:0] node1665;
	wire [4-1:0] node1668;
	wire [4-1:0] node1671;
	wire [4-1:0] node1672;
	wire [4-1:0] node1674;
	wire [4-1:0] node1678;
	wire [4-1:0] node1679;
	wire [4-1:0] node1680;
	wire [4-1:0] node1682;
	wire [4-1:0] node1683;
	wire [4-1:0] node1687;
	wire [4-1:0] node1688;
	wire [4-1:0] node1689;
	wire [4-1:0] node1693;
	wire [4-1:0] node1694;
	wire [4-1:0] node1698;
	wire [4-1:0] node1699;
	wire [4-1:0] node1700;
	wire [4-1:0] node1702;
	wire [4-1:0] node1704;
	wire [4-1:0] node1707;
	wire [4-1:0] node1709;
	wire [4-1:0] node1712;
	wire [4-1:0] node1713;
	wire [4-1:0] node1714;
	wire [4-1:0] node1718;
	wire [4-1:0] node1720;
	wire [4-1:0] node1723;
	wire [4-1:0] node1724;
	wire [4-1:0] node1725;
	wire [4-1:0] node1726;
	wire [4-1:0] node1727;
	wire [4-1:0] node1728;
	wire [4-1:0] node1732;
	wire [4-1:0] node1735;
	wire [4-1:0] node1736;
	wire [4-1:0] node1739;
	wire [4-1:0] node1742;
	wire [4-1:0] node1743;
	wire [4-1:0] node1744;
	wire [4-1:0] node1745;
	wire [4-1:0] node1747;
	wire [4-1:0] node1750;
	wire [4-1:0] node1754;
	wire [4-1:0] node1756;
	wire [4-1:0] node1757;
	wire [4-1:0] node1761;
	wire [4-1:0] node1762;
	wire [4-1:0] node1763;
	wire [4-1:0] node1764;
	wire [4-1:0] node1768;
	wire [4-1:0] node1769;
	wire [4-1:0] node1771;
	wire [4-1:0] node1774;
	wire [4-1:0] node1776;
	wire [4-1:0] node1779;
	wire [4-1:0] node1780;
	wire [4-1:0] node1781;
	wire [4-1:0] node1784;
	wire [4-1:0] node1785;
	wire [4-1:0] node1789;
	wire [4-1:0] node1790;
	wire [4-1:0] node1794;
	wire [4-1:0] node1795;
	wire [4-1:0] node1796;
	wire [4-1:0] node1797;
	wire [4-1:0] node1798;
	wire [4-1:0] node1799;
	wire [4-1:0] node1801;
	wire [4-1:0] node1803;
	wire [4-1:0] node1806;
	wire [4-1:0] node1808;
	wire [4-1:0] node1810;
	wire [4-1:0] node1813;
	wire [4-1:0] node1814;
	wire [4-1:0] node1815;
	wire [4-1:0] node1817;
	wire [4-1:0] node1819;
	wire [4-1:0] node1823;
	wire [4-1:0] node1825;
	wire [4-1:0] node1826;
	wire [4-1:0] node1830;
	wire [4-1:0] node1831;
	wire [4-1:0] node1832;
	wire [4-1:0] node1833;
	wire [4-1:0] node1834;
	wire [4-1:0] node1836;
	wire [4-1:0] node1839;
	wire [4-1:0] node1841;
	wire [4-1:0] node1844;
	wire [4-1:0] node1846;
	wire [4-1:0] node1849;
	wire [4-1:0] node1851;
	wire [4-1:0] node1852;
	wire [4-1:0] node1856;
	wire [4-1:0] node1857;
	wire [4-1:0] node1859;
	wire [4-1:0] node1862;
	wire [4-1:0] node1863;
	wire [4-1:0] node1864;
	wire [4-1:0] node1869;
	wire [4-1:0] node1870;
	wire [4-1:0] node1871;
	wire [4-1:0] node1872;
	wire [4-1:0] node1873;
	wire [4-1:0] node1874;
	wire [4-1:0] node1878;
	wire [4-1:0] node1880;
	wire [4-1:0] node1883;
	wire [4-1:0] node1884;
	wire [4-1:0] node1885;
	wire [4-1:0] node1888;
	wire [4-1:0] node1892;
	wire [4-1:0] node1893;
	wire [4-1:0] node1894;
	wire [4-1:0] node1895;
	wire [4-1:0] node1897;
	wire [4-1:0] node1900;
	wire [4-1:0] node1904;
	wire [4-1:0] node1905;
	wire [4-1:0] node1906;
	wire [4-1:0] node1908;
	wire [4-1:0] node1913;
	wire [4-1:0] node1914;
	wire [4-1:0] node1915;
	wire [4-1:0] node1916;
	wire [4-1:0] node1919;
	wire [4-1:0] node1921;
	wire [4-1:0] node1923;
	wire [4-1:0] node1927;
	wire [4-1:0] node1928;
	wire [4-1:0] node1929;
	wire [4-1:0] node1931;
	wire [4-1:0] node1933;
	wire [4-1:0] node1936;
	wire [4-1:0] node1938;
	wire [4-1:0] node1941;
	wire [4-1:0] node1942;
	wire [4-1:0] node1944;
	wire [4-1:0] node1945;
	wire [4-1:0] node1949;
	wire [4-1:0] node1951;
	wire [4-1:0] node1953;
	wire [4-1:0] node1956;
	wire [4-1:0] node1957;
	wire [4-1:0] node1958;
	wire [4-1:0] node1959;
	wire [4-1:0] node1960;
	wire [4-1:0] node1961;
	wire [4-1:0] node1964;
	wire [4-1:0] node1965;
	wire [4-1:0] node1969;
	wire [4-1:0] node1970;
	wire [4-1:0] node1972;
	wire [4-1:0] node1975;
	wire [4-1:0] node1978;
	wire [4-1:0] node1979;
	wire [4-1:0] node1980;
	wire [4-1:0] node1981;
	wire [4-1:0] node1985;
	wire [4-1:0] node1986;
	wire [4-1:0] node1987;
	wire [4-1:0] node1990;
	wire [4-1:0] node1994;
	wire [4-1:0] node1995;
	wire [4-1:0] node1997;
	wire [4-1:0] node1998;
	wire [4-1:0] node2002;
	wire [4-1:0] node2003;
	wire [4-1:0] node2006;
	wire [4-1:0] node2009;
	wire [4-1:0] node2010;
	wire [4-1:0] node2011;
	wire [4-1:0] node2012;
	wire [4-1:0] node2013;
	wire [4-1:0] node2016;
	wire [4-1:0] node2019;
	wire [4-1:0] node2022;
	wire [4-1:0] node2023;
	wire [4-1:0] node2024;
	wire [4-1:0] node2025;
	wire [4-1:0] node2029;
	wire [4-1:0] node2033;
	wire [4-1:0] node2034;
	wire [4-1:0] node2035;
	wire [4-1:0] node2036;
	wire [4-1:0] node2039;
	wire [4-1:0] node2040;
	wire [4-1:0] node2045;
	wire [4-1:0] node2047;
	wire [4-1:0] node2048;
	wire [4-1:0] node2050;
	wire [4-1:0] node2054;
	wire [4-1:0] node2055;
	wire [4-1:0] node2056;
	wire [4-1:0] node2057;
	wire [4-1:0] node2058;
	wire [4-1:0] node2060;
	wire [4-1:0] node2062;
	wire [4-1:0] node2065;
	wire [4-1:0] node2069;
	wire [4-1:0] node2070;
	wire [4-1:0] node2071;
	wire [4-1:0] node2073;
	wire [4-1:0] node2074;
	wire [4-1:0] node2078;
	wire [4-1:0] node2081;
	wire [4-1:0] node2083;
	wire [4-1:0] node2085;
	wire [4-1:0] node2086;
	wire [4-1:0] node2090;
	wire [4-1:0] node2091;
	wire [4-1:0] node2092;
	wire [4-1:0] node2093;
	wire [4-1:0] node2096;
	wire [4-1:0] node2099;
	wire [4-1:0] node2100;
	wire [4-1:0] node2101;
	wire [4-1:0] node2102;
	wire [4-1:0] node2105;
	wire [4-1:0] node2109;
	wire [4-1:0] node2111;
	wire [4-1:0] node2114;
	wire [4-1:0] node2115;
	wire [4-1:0] node2116;
	wire [4-1:0] node2117;
	wire [4-1:0] node2119;
	wire [4-1:0] node2122;
	wire [4-1:0] node2125;
	wire [4-1:0] node2128;
	wire [4-1:0] node2129;
	wire [4-1:0] node2131;
	wire [4-1:0] node2132;
	wire [4-1:0] node2135;
	wire [4-1:0] node2138;
	wire [4-1:0] node2140;
	wire [4-1:0] node2143;
	wire [4-1:0] node2144;
	wire [4-1:0] node2145;
	wire [4-1:0] node2146;
	wire [4-1:0] node2147;
	wire [4-1:0] node2148;
	wire [4-1:0] node2149;
	wire [4-1:0] node2150;
	wire [4-1:0] node2153;
	wire [4-1:0] node2154;
	wire [4-1:0] node2156;
	wire [4-1:0] node2160;
	wire [4-1:0] node2161;
	wire [4-1:0] node2164;
	wire [4-1:0] node2166;
	wire [4-1:0] node2168;
	wire [4-1:0] node2171;
	wire [4-1:0] node2172;
	wire [4-1:0] node2173;
	wire [4-1:0] node2175;
	wire [4-1:0] node2176;
	wire [4-1:0] node2180;
	wire [4-1:0] node2181;
	wire [4-1:0] node2182;
	wire [4-1:0] node2187;
	wire [4-1:0] node2189;
	wire [4-1:0] node2190;
	wire [4-1:0] node2192;
	wire [4-1:0] node2196;
	wire [4-1:0] node2197;
	wire [4-1:0] node2198;
	wire [4-1:0] node2199;
	wire [4-1:0] node2200;
	wire [4-1:0] node2203;
	wire [4-1:0] node2207;
	wire [4-1:0] node2208;
	wire [4-1:0] node2210;
	wire [4-1:0] node2213;
	wire [4-1:0] node2214;
	wire [4-1:0] node2215;
	wire [4-1:0] node2218;
	wire [4-1:0] node2222;
	wire [4-1:0] node2223;
	wire [4-1:0] node2224;
	wire [4-1:0] node2225;
	wire [4-1:0] node2228;
	wire [4-1:0] node2230;
	wire [4-1:0] node2234;
	wire [4-1:0] node2235;
	wire [4-1:0] node2238;
	wire [4-1:0] node2240;
	wire [4-1:0] node2241;
	wire [4-1:0] node2244;
	wire [4-1:0] node2247;
	wire [4-1:0] node2248;
	wire [4-1:0] node2249;
	wire [4-1:0] node2250;
	wire [4-1:0] node2251;
	wire [4-1:0] node2253;
	wire [4-1:0] node2256;
	wire [4-1:0] node2257;
	wire [4-1:0] node2258;
	wire [4-1:0] node2262;
	wire [4-1:0] node2264;
	wire [4-1:0] node2267;
	wire [4-1:0] node2268;
	wire [4-1:0] node2270;
	wire [4-1:0] node2271;
	wire [4-1:0] node2275;
	wire [4-1:0] node2276;
	wire [4-1:0] node2278;
	wire [4-1:0] node2282;
	wire [4-1:0] node2283;
	wire [4-1:0] node2284;
	wire [4-1:0] node2288;
	wire [4-1:0] node2289;
	wire [4-1:0] node2290;
	wire [4-1:0] node2293;
	wire [4-1:0] node2296;
	wire [4-1:0] node2299;
	wire [4-1:0] node2300;
	wire [4-1:0] node2301;
	wire [4-1:0] node2303;
	wire [4-1:0] node2305;
	wire [4-1:0] node2308;
	wire [4-1:0] node2309;
	wire [4-1:0] node2311;
	wire [4-1:0] node2313;
	wire [4-1:0] node2316;
	wire [4-1:0] node2318;
	wire [4-1:0] node2319;
	wire [4-1:0] node2322;
	wire [4-1:0] node2325;
	wire [4-1:0] node2326;
	wire [4-1:0] node2327;
	wire [4-1:0] node2330;
	wire [4-1:0] node2332;
	wire [4-1:0] node2334;
	wire [4-1:0] node2337;
	wire [4-1:0] node2338;
	wire [4-1:0] node2339;
	wire [4-1:0] node2341;
	wire [4-1:0] node2344;
	wire [4-1:0] node2348;
	wire [4-1:0] node2349;
	wire [4-1:0] node2350;
	wire [4-1:0] node2351;
	wire [4-1:0] node2352;
	wire [4-1:0] node2355;
	wire [4-1:0] node2357;
	wire [4-1:0] node2358;
	wire [4-1:0] node2362;
	wire [4-1:0] node2363;
	wire [4-1:0] node2364;
	wire [4-1:0] node2367;
	wire [4-1:0] node2368;
	wire [4-1:0] node2372;
	wire [4-1:0] node2373;
	wire [4-1:0] node2375;
	wire [4-1:0] node2378;
	wire [4-1:0] node2381;
	wire [4-1:0] node2382;
	wire [4-1:0] node2383;
	wire [4-1:0] node2384;
	wire [4-1:0] node2387;
	wire [4-1:0] node2390;
	wire [4-1:0] node2391;
	wire [4-1:0] node2394;
	wire [4-1:0] node2396;
	wire [4-1:0] node2399;
	wire [4-1:0] node2400;
	wire [4-1:0] node2402;
	wire [4-1:0] node2403;
	wire [4-1:0] node2406;
	wire [4-1:0] node2409;
	wire [4-1:0] node2410;
	wire [4-1:0] node2413;
	wire [4-1:0] node2414;
	wire [4-1:0] node2415;
	wire [4-1:0] node2420;
	wire [4-1:0] node2421;
	wire [4-1:0] node2422;
	wire [4-1:0] node2423;
	wire [4-1:0] node2424;
	wire [4-1:0] node2425;
	wire [4-1:0] node2428;
	wire [4-1:0] node2430;
	wire [4-1:0] node2434;
	wire [4-1:0] node2436;
	wire [4-1:0] node2437;
	wire [4-1:0] node2439;
	wire [4-1:0] node2443;
	wire [4-1:0] node2444;
	wire [4-1:0] node2445;
	wire [4-1:0] node2446;
	wire [4-1:0] node2450;
	wire [4-1:0] node2451;
	wire [4-1:0] node2453;
	wire [4-1:0] node2456;
	wire [4-1:0] node2457;
	wire [4-1:0] node2460;
	wire [4-1:0] node2463;
	wire [4-1:0] node2464;
	wire [4-1:0] node2466;
	wire [4-1:0] node2468;
	wire [4-1:0] node2471;
	wire [4-1:0] node2472;
	wire [4-1:0] node2475;
	wire [4-1:0] node2477;
	wire [4-1:0] node2480;
	wire [4-1:0] node2481;
	wire [4-1:0] node2482;
	wire [4-1:0] node2483;
	wire [4-1:0] node2486;
	wire [4-1:0] node2489;
	wire [4-1:0] node2490;
	wire [4-1:0] node2491;
	wire [4-1:0] node2494;
	wire [4-1:0] node2496;
	wire [4-1:0] node2499;
	wire [4-1:0] node2500;
	wire [4-1:0] node2504;
	wire [4-1:0] node2505;
	wire [4-1:0] node2506;
	wire [4-1:0] node2509;
	wire [4-1:0] node2510;
	wire [4-1:0] node2511;
	wire [4-1:0] node2514;
	wire [4-1:0] node2517;
	wire [4-1:0] node2520;
	wire [4-1:0] node2522;
	wire [4-1:0] node2524;
	wire [4-1:0] node2527;
	wire [4-1:0] node2528;
	wire [4-1:0] node2529;
	wire [4-1:0] node2530;
	wire [4-1:0] node2531;
	wire [4-1:0] node2532;
	wire [4-1:0] node2533;
	wire [4-1:0] node2534;
	wire [4-1:0] node2535;
	wire [4-1:0] node2540;
	wire [4-1:0] node2542;
	wire [4-1:0] node2545;
	wire [4-1:0] node2546;
	wire [4-1:0] node2547;
	wire [4-1:0] node2552;
	wire [4-1:0] node2553;
	wire [4-1:0] node2554;
	wire [4-1:0] node2557;
	wire [4-1:0] node2560;
	wire [4-1:0] node2561;
	wire [4-1:0] node2562;
	wire [4-1:0] node2564;
	wire [4-1:0] node2567;
	wire [4-1:0] node2568;
	wire [4-1:0] node2571;
	wire [4-1:0] node2574;
	wire [4-1:0] node2577;
	wire [4-1:0] node2578;
	wire [4-1:0] node2579;
	wire [4-1:0] node2580;
	wire [4-1:0] node2582;
	wire [4-1:0] node2584;
	wire [4-1:0] node2587;
	wire [4-1:0] node2589;
	wire [4-1:0] node2591;
	wire [4-1:0] node2594;
	wire [4-1:0] node2595;
	wire [4-1:0] node2598;
	wire [4-1:0] node2599;
	wire [4-1:0] node2601;
	wire [4-1:0] node2605;
	wire [4-1:0] node2606;
	wire [4-1:0] node2607;
	wire [4-1:0] node2609;
	wire [4-1:0] node2610;
	wire [4-1:0] node2614;
	wire [4-1:0] node2615;
	wire [4-1:0] node2617;
	wire [4-1:0] node2620;
	wire [4-1:0] node2621;
	wire [4-1:0] node2625;
	wire [4-1:0] node2626;
	wire [4-1:0] node2629;
	wire [4-1:0] node2630;
	wire [4-1:0] node2633;
	wire [4-1:0] node2635;
	wire [4-1:0] node2638;
	wire [4-1:0] node2639;
	wire [4-1:0] node2640;
	wire [4-1:0] node2641;
	wire [4-1:0] node2642;
	wire [4-1:0] node2643;
	wire [4-1:0] node2645;
	wire [4-1:0] node2648;
	wire [4-1:0] node2650;
	wire [4-1:0] node2653;
	wire [4-1:0] node2655;
	wire [4-1:0] node2656;
	wire [4-1:0] node2660;
	wire [4-1:0] node2661;
	wire [4-1:0] node2665;
	wire [4-1:0] node2666;
	wire [4-1:0] node2667;
	wire [4-1:0] node2668;
	wire [4-1:0] node2670;
	wire [4-1:0] node2673;
	wire [4-1:0] node2676;
	wire [4-1:0] node2677;
	wire [4-1:0] node2679;
	wire [4-1:0] node2683;
	wire [4-1:0] node2684;
	wire [4-1:0] node2687;
	wire [4-1:0] node2688;
	wire [4-1:0] node2690;
	wire [4-1:0] node2694;
	wire [4-1:0] node2695;
	wire [4-1:0] node2696;
	wire [4-1:0] node2697;
	wire [4-1:0] node2698;
	wire [4-1:0] node2702;
	wire [4-1:0] node2703;
	wire [4-1:0] node2707;
	wire [4-1:0] node2708;
	wire [4-1:0] node2709;
	wire [4-1:0] node2713;
	wire [4-1:0] node2714;
	wire [4-1:0] node2716;
	wire [4-1:0] node2720;
	wire [4-1:0] node2721;
	wire [4-1:0] node2722;
	wire [4-1:0] node2724;
	wire [4-1:0] node2726;
	wire [4-1:0] node2729;
	wire [4-1:0] node2731;
	wire [4-1:0] node2734;
	wire [4-1:0] node2735;
	wire [4-1:0] node2736;
	wire [4-1:0] node2739;
	wire [4-1:0] node2742;
	wire [4-1:0] node2743;
	wire [4-1:0] node2747;
	wire [4-1:0] node2748;
	wire [4-1:0] node2749;
	wire [4-1:0] node2750;
	wire [4-1:0] node2751;
	wire [4-1:0] node2754;
	wire [4-1:0] node2756;
	wire [4-1:0] node2757;
	wire [4-1:0] node2760;
	wire [4-1:0] node2763;
	wire [4-1:0] node2764;
	wire [4-1:0] node2765;
	wire [4-1:0] node2769;
	wire [4-1:0] node2771;
	wire [4-1:0] node2772;
	wire [4-1:0] node2774;
	wire [4-1:0] node2778;
	wire [4-1:0] node2779;
	wire [4-1:0] node2780;
	wire [4-1:0] node2781;
	wire [4-1:0] node2782;
	wire [4-1:0] node2785;
	wire [4-1:0] node2789;
	wire [4-1:0] node2791;
	wire [4-1:0] node2794;
	wire [4-1:0] node2795;
	wire [4-1:0] node2796;
	wire [4-1:0] node2800;
	wire [4-1:0] node2801;
	wire [4-1:0] node2802;
	wire [4-1:0] node2803;
	wire [4-1:0] node2807;
	wire [4-1:0] node2810;
	wire [4-1:0] node2812;
	wire [4-1:0] node2815;
	wire [4-1:0] node2816;
	wire [4-1:0] node2817;
	wire [4-1:0] node2818;
	wire [4-1:0] node2819;
	wire [4-1:0] node2820;
	wire [4-1:0] node2824;
	wire [4-1:0] node2827;
	wire [4-1:0] node2828;
	wire [4-1:0] node2830;
	wire [4-1:0] node2831;
	wire [4-1:0] node2835;
	wire [4-1:0] node2836;
	wire [4-1:0] node2840;
	wire [4-1:0] node2841;
	wire [4-1:0] node2842;
	wire [4-1:0] node2843;
	wire [4-1:0] node2844;
	wire [4-1:0] node2848;
	wire [4-1:0] node2849;
	wire [4-1:0] node2854;
	wire [4-1:0] node2855;
	wire [4-1:0] node2857;
	wire [4-1:0] node2858;
	wire [4-1:0] node2861;
	wire [4-1:0] node2864;
	wire [4-1:0] node2865;
	wire [4-1:0] node2869;
	wire [4-1:0] node2870;
	wire [4-1:0] node2871;
	wire [4-1:0] node2872;
	wire [4-1:0] node2874;
	wire [4-1:0] node2877;
	wire [4-1:0] node2879;
	wire [4-1:0] node2880;
	wire [4-1:0] node2884;
	wire [4-1:0] node2885;
	wire [4-1:0] node2886;
	wire [4-1:0] node2888;
	wire [4-1:0] node2892;
	wire [4-1:0] node2893;
	wire [4-1:0] node2897;
	wire [4-1:0] node2898;
	wire [4-1:0] node2899;
	wire [4-1:0] node2900;
	wire [4-1:0] node2901;
	wire [4-1:0] node2904;
	wire [4-1:0] node2907;
	wire [4-1:0] node2911;
	wire [4-1:0] node2912;
	wire [4-1:0] node2913;
	wire [4-1:0] node2917;
	wire [4-1:0] node2920;
	wire [4-1:0] node2921;
	wire [4-1:0] node2922;
	wire [4-1:0] node2923;
	wire [4-1:0] node2924;
	wire [4-1:0] node2925;
	wire [4-1:0] node2926;
	wire [4-1:0] node2927;
	wire [4-1:0] node2928;
	wire [4-1:0] node2929;
	wire [4-1:0] node2930;
	wire [4-1:0] node2931;
	wire [4-1:0] node2935;
	wire [4-1:0] node2938;
	wire [4-1:0] node2941;
	wire [4-1:0] node2943;
	wire [4-1:0] node2946;
	wire [4-1:0] node2947;
	wire [4-1:0] node2949;
	wire [4-1:0] node2951;
	wire [4-1:0] node2953;
	wire [4-1:0] node2956;
	wire [4-1:0] node2957;
	wire [4-1:0] node2959;
	wire [4-1:0] node2962;
	wire [4-1:0] node2964;
	wire [4-1:0] node2967;
	wire [4-1:0] node2968;
	wire [4-1:0] node2969;
	wire [4-1:0] node2971;
	wire [4-1:0] node2974;
	wire [4-1:0] node2975;
	wire [4-1:0] node2976;
	wire [4-1:0] node2977;
	wire [4-1:0] node2980;
	wire [4-1:0] node2983;
	wire [4-1:0] node2986;
	wire [4-1:0] node2988;
	wire [4-1:0] node2991;
	wire [4-1:0] node2992;
	wire [4-1:0] node2993;
	wire [4-1:0] node2994;
	wire [4-1:0] node2998;
	wire [4-1:0] node2999;
	wire [4-1:0] node3003;
	wire [4-1:0] node3004;
	wire [4-1:0] node3006;
	wire [4-1:0] node3009;
	wire [4-1:0] node3010;
	wire [4-1:0] node3013;
	wire [4-1:0] node3016;
	wire [4-1:0] node3017;
	wire [4-1:0] node3018;
	wire [4-1:0] node3019;
	wire [4-1:0] node3020;
	wire [4-1:0] node3021;
	wire [4-1:0] node3024;
	wire [4-1:0] node3027;
	wire [4-1:0] node3028;
	wire [4-1:0] node3029;
	wire [4-1:0] node3032;
	wire [4-1:0] node3035;
	wire [4-1:0] node3038;
	wire [4-1:0] node3039;
	wire [4-1:0] node3043;
	wire [4-1:0] node3044;
	wire [4-1:0] node3045;
	wire [4-1:0] node3048;
	wire [4-1:0] node3050;
	wire [4-1:0] node3053;
	wire [4-1:0] node3054;
	wire [4-1:0] node3058;
	wire [4-1:0] node3059;
	wire [4-1:0] node3060;
	wire [4-1:0] node3061;
	wire [4-1:0] node3062;
	wire [4-1:0] node3066;
	wire [4-1:0] node3069;
	wire [4-1:0] node3070;
	wire [4-1:0] node3073;
	wire [4-1:0] node3074;
	wire [4-1:0] node3077;
	wire [4-1:0] node3080;
	wire [4-1:0] node3082;
	wire [4-1:0] node3083;
	wire [4-1:0] node3084;
	wire [4-1:0] node3089;
	wire [4-1:0] node3090;
	wire [4-1:0] node3091;
	wire [4-1:0] node3092;
	wire [4-1:0] node3093;
	wire [4-1:0] node3094;
	wire [4-1:0] node3097;
	wire [4-1:0] node3098;
	wire [4-1:0] node3102;
	wire [4-1:0] node3103;
	wire [4-1:0] node3105;
	wire [4-1:0] node3108;
	wire [4-1:0] node3111;
	wire [4-1:0] node3112;
	wire [4-1:0] node3114;
	wire [4-1:0] node3117;
	wire [4-1:0] node3118;
	wire [4-1:0] node3120;
	wire [4-1:0] node3121;
	wire [4-1:0] node3124;
	wire [4-1:0] node3127;
	wire [4-1:0] node3129;
	wire [4-1:0] node3132;
	wire [4-1:0] node3133;
	wire [4-1:0] node3134;
	wire [4-1:0] node3135;
	wire [4-1:0] node3137;
	wire [4-1:0] node3141;
	wire [4-1:0] node3143;
	wire [4-1:0] node3145;
	wire [4-1:0] node3148;
	wire [4-1:0] node3149;
	wire [4-1:0] node3151;
	wire [4-1:0] node3154;
	wire [4-1:0] node3156;
	wire [4-1:0] node3157;
	wire [4-1:0] node3158;
	wire [4-1:0] node3163;
	wire [4-1:0] node3164;
	wire [4-1:0] node3165;
	wire [4-1:0] node3166;
	wire [4-1:0] node3168;
	wire [4-1:0] node3170;
	wire [4-1:0] node3172;
	wire [4-1:0] node3175;
	wire [4-1:0] node3177;
	wire [4-1:0] node3179;
	wire [4-1:0] node3182;
	wire [4-1:0] node3183;
	wire [4-1:0] node3184;
	wire [4-1:0] node3185;
	wire [4-1:0] node3188;
	wire [4-1:0] node3189;
	wire [4-1:0] node3193;
	wire [4-1:0] node3194;
	wire [4-1:0] node3198;
	wire [4-1:0] node3200;
	wire [4-1:0] node3203;
	wire [4-1:0] node3204;
	wire [4-1:0] node3205;
	wire [4-1:0] node3207;
	wire [4-1:0] node3210;
	wire [4-1:0] node3211;
	wire [4-1:0] node3214;
	wire [4-1:0] node3217;
	wire [4-1:0] node3218;
	wire [4-1:0] node3219;
	wire [4-1:0] node3221;
	wire [4-1:0] node3224;
	wire [4-1:0] node3227;
	wire [4-1:0] node3228;
	wire [4-1:0] node3229;
	wire [4-1:0] node3231;
	wire [4-1:0] node3235;
	wire [4-1:0] node3237;
	wire [4-1:0] node3240;
	wire [4-1:0] node3241;
	wire [4-1:0] node3242;
	wire [4-1:0] node3243;
	wire [4-1:0] node3244;
	wire [4-1:0] node3245;
	wire [4-1:0] node3246;
	wire [4-1:0] node3248;
	wire [4-1:0] node3250;
	wire [4-1:0] node3253;
	wire [4-1:0] node3254;
	wire [4-1:0] node3256;
	wire [4-1:0] node3260;
	wire [4-1:0] node3261;
	wire [4-1:0] node3262;
	wire [4-1:0] node3263;
	wire [4-1:0] node3267;
	wire [4-1:0] node3269;
	wire [4-1:0] node3272;
	wire [4-1:0] node3275;
	wire [4-1:0] node3276;
	wire [4-1:0] node3277;
	wire [4-1:0] node3278;
	wire [4-1:0] node3281;
	wire [4-1:0] node3283;
	wire [4-1:0] node3286;
	wire [4-1:0] node3289;
	wire [4-1:0] node3290;
	wire [4-1:0] node3293;
	wire [4-1:0] node3296;
	wire [4-1:0] node3297;
	wire [4-1:0] node3298;
	wire [4-1:0] node3300;
	wire [4-1:0] node3303;
	wire [4-1:0] node3304;
	wire [4-1:0] node3308;
	wire [4-1:0] node3309;
	wire [4-1:0] node3310;
	wire [4-1:0] node3311;
	wire [4-1:0] node3314;
	wire [4-1:0] node3315;
	wire [4-1:0] node3319;
	wire [4-1:0] node3320;
	wire [4-1:0] node3321;
	wire [4-1:0] node3325;
	wire [4-1:0] node3328;
	wire [4-1:0] node3329;
	wire [4-1:0] node3331;
	wire [4-1:0] node3335;
	wire [4-1:0] node3336;
	wire [4-1:0] node3337;
	wire [4-1:0] node3339;
	wire [4-1:0] node3340;
	wire [4-1:0] node3341;
	wire [4-1:0] node3344;
	wire [4-1:0] node3347;
	wire [4-1:0] node3348;
	wire [4-1:0] node3350;
	wire [4-1:0] node3354;
	wire [4-1:0] node3355;
	wire [4-1:0] node3356;
	wire [4-1:0] node3358;
	wire [4-1:0] node3359;
	wire [4-1:0] node3363;
	wire [4-1:0] node3364;
	wire [4-1:0] node3368;
	wire [4-1:0] node3369;
	wire [4-1:0] node3370;
	wire [4-1:0] node3371;
	wire [4-1:0] node3376;
	wire [4-1:0] node3379;
	wire [4-1:0] node3380;
	wire [4-1:0] node3381;
	wire [4-1:0] node3382;
	wire [4-1:0] node3383;
	wire [4-1:0] node3384;
	wire [4-1:0] node3388;
	wire [4-1:0] node3391;
	wire [4-1:0] node3392;
	wire [4-1:0] node3393;
	wire [4-1:0] node3396;
	wire [4-1:0] node3399;
	wire [4-1:0] node3401;
	wire [4-1:0] node3404;
	wire [4-1:0] node3405;
	wire [4-1:0] node3406;
	wire [4-1:0] node3409;
	wire [4-1:0] node3412;
	wire [4-1:0] node3414;
	wire [4-1:0] node3415;
	wire [4-1:0] node3419;
	wire [4-1:0] node3420;
	wire [4-1:0] node3421;
	wire [4-1:0] node3425;
	wire [4-1:0] node3426;
	wire [4-1:0] node3427;
	wire [4-1:0] node3431;
	wire [4-1:0] node3434;
	wire [4-1:0] node3435;
	wire [4-1:0] node3436;
	wire [4-1:0] node3437;
	wire [4-1:0] node3438;
	wire [4-1:0] node3439;
	wire [4-1:0] node3441;
	wire [4-1:0] node3443;
	wire [4-1:0] node3446;
	wire [4-1:0] node3449;
	wire [4-1:0] node3451;
	wire [4-1:0] node3452;
	wire [4-1:0] node3453;
	wire [4-1:0] node3457;
	wire [4-1:0] node3459;
	wire [4-1:0] node3462;
	wire [4-1:0] node3463;
	wire [4-1:0] node3464;
	wire [4-1:0] node3466;
	wire [4-1:0] node3467;
	wire [4-1:0] node3472;
	wire [4-1:0] node3474;
	wire [4-1:0] node3477;
	wire [4-1:0] node3478;
	wire [4-1:0] node3479;
	wire [4-1:0] node3480;
	wire [4-1:0] node3482;
	wire [4-1:0] node3486;
	wire [4-1:0] node3487;
	wire [4-1:0] node3489;
	wire [4-1:0] node3490;
	wire [4-1:0] node3494;
	wire [4-1:0] node3495;
	wire [4-1:0] node3499;
	wire [4-1:0] node3500;
	wire [4-1:0] node3501;
	wire [4-1:0] node3502;
	wire [4-1:0] node3504;
	wire [4-1:0] node3508;
	wire [4-1:0] node3511;
	wire [4-1:0] node3513;
	wire [4-1:0] node3514;
	wire [4-1:0] node3517;
	wire [4-1:0] node3520;
	wire [4-1:0] node3521;
	wire [4-1:0] node3522;
	wire [4-1:0] node3523;
	wire [4-1:0] node3526;
	wire [4-1:0] node3527;
	wire [4-1:0] node3528;
	wire [4-1:0] node3532;
	wire [4-1:0] node3535;
	wire [4-1:0] node3536;
	wire [4-1:0] node3538;
	wire [4-1:0] node3539;
	wire [4-1:0] node3540;
	wire [4-1:0] node3543;
	wire [4-1:0] node3547;
	wire [4-1:0] node3548;
	wire [4-1:0] node3549;
	wire [4-1:0] node3551;
	wire [4-1:0] node3554;
	wire [4-1:0] node3557;
	wire [4-1:0] node3559;
	wire [4-1:0] node3560;
	wire [4-1:0] node3564;
	wire [4-1:0] node3565;
	wire [4-1:0] node3566;
	wire [4-1:0] node3567;
	wire [4-1:0] node3568;
	wire [4-1:0] node3569;
	wire [4-1:0] node3573;
	wire [4-1:0] node3574;
	wire [4-1:0] node3577;
	wire [4-1:0] node3580;
	wire [4-1:0] node3583;
	wire [4-1:0] node3584;
	wire [4-1:0] node3585;
	wire [4-1:0] node3586;
	wire [4-1:0] node3591;
	wire [4-1:0] node3593;
	wire [4-1:0] node3594;
	wire [4-1:0] node3598;
	wire [4-1:0] node3599;
	wire [4-1:0] node3600;
	wire [4-1:0] node3602;
	wire [4-1:0] node3603;
	wire [4-1:0] node3607;
	wire [4-1:0] node3609;
	wire [4-1:0] node3610;
	wire [4-1:0] node3614;
	wire [4-1:0] node3615;
	wire [4-1:0] node3616;
	wire [4-1:0] node3621;
	wire [4-1:0] node3622;
	wire [4-1:0] node3623;
	wire [4-1:0] node3624;
	wire [4-1:0] node3625;
	wire [4-1:0] node3626;
	wire [4-1:0] node3627;
	wire [4-1:0] node3628;
	wire [4-1:0] node3629;
	wire [4-1:0] node3633;
	wire [4-1:0] node3635;
	wire [4-1:0] node3638;
	wire [4-1:0] node3639;
	wire [4-1:0] node3640;
	wire [4-1:0] node3642;
	wire [4-1:0] node3646;
	wire [4-1:0] node3647;
	wire [4-1:0] node3651;
	wire [4-1:0] node3652;
	wire [4-1:0] node3654;
	wire [4-1:0] node3656;
	wire [4-1:0] node3659;
	wire [4-1:0] node3660;
	wire [4-1:0] node3662;
	wire [4-1:0] node3665;
	wire [4-1:0] node3666;
	wire [4-1:0] node3670;
	wire [4-1:0] node3671;
	wire [4-1:0] node3672;
	wire [4-1:0] node3673;
	wire [4-1:0] node3674;
	wire [4-1:0] node3678;
	wire [4-1:0] node3679;
	wire [4-1:0] node3682;
	wire [4-1:0] node3685;
	wire [4-1:0] node3686;
	wire [4-1:0] node3687;
	wire [4-1:0] node3691;
	wire [4-1:0] node3693;
	wire [4-1:0] node3694;
	wire [4-1:0] node3697;
	wire [4-1:0] node3700;
	wire [4-1:0] node3701;
	wire [4-1:0] node3702;
	wire [4-1:0] node3703;
	wire [4-1:0] node3707;
	wire [4-1:0] node3709;
	wire [4-1:0] node3712;
	wire [4-1:0] node3713;
	wire [4-1:0] node3715;
	wire [4-1:0] node3719;
	wire [4-1:0] node3720;
	wire [4-1:0] node3721;
	wire [4-1:0] node3722;
	wire [4-1:0] node3723;
	wire [4-1:0] node3724;
	wire [4-1:0] node3729;
	wire [4-1:0] node3730;
	wire [4-1:0] node3731;
	wire [4-1:0] node3735;
	wire [4-1:0] node3738;
	wire [4-1:0] node3739;
	wire [4-1:0] node3740;
	wire [4-1:0] node3742;
	wire [4-1:0] node3745;
	wire [4-1:0] node3748;
	wire [4-1:0] node3749;
	wire [4-1:0] node3753;
	wire [4-1:0] node3754;
	wire [4-1:0] node3755;
	wire [4-1:0] node3757;
	wire [4-1:0] node3760;
	wire [4-1:0] node3762;
	wire [4-1:0] node3763;
	wire [4-1:0] node3764;
	wire [4-1:0] node3768;
	wire [4-1:0] node3769;
	wire [4-1:0] node3772;
	wire [4-1:0] node3775;
	wire [4-1:0] node3776;
	wire [4-1:0] node3777;
	wire [4-1:0] node3781;
	wire [4-1:0] node3782;
	wire [4-1:0] node3784;
	wire [4-1:0] node3788;
	wire [4-1:0] node3789;
	wire [4-1:0] node3790;
	wire [4-1:0] node3791;
	wire [4-1:0] node3792;
	wire [4-1:0] node3793;
	wire [4-1:0] node3795;
	wire [4-1:0] node3799;
	wire [4-1:0] node3800;
	wire [4-1:0] node3801;
	wire [4-1:0] node3802;
	wire [4-1:0] node3808;
	wire [4-1:0] node3809;
	wire [4-1:0] node3810;
	wire [4-1:0] node3812;
	wire [4-1:0] node3816;
	wire [4-1:0] node3818;
	wire [4-1:0] node3820;
	wire [4-1:0] node3821;
	wire [4-1:0] node3824;
	wire [4-1:0] node3827;
	wire [4-1:0] node3828;
	wire [4-1:0] node3829;
	wire [4-1:0] node3830;
	wire [4-1:0] node3832;
	wire [4-1:0] node3833;
	wire [4-1:0] node3837;
	wire [4-1:0] node3839;
	wire [4-1:0] node3842;
	wire [4-1:0] node3843;
	wire [4-1:0] node3844;
	wire [4-1:0] node3846;
	wire [4-1:0] node3850;
	wire [4-1:0] node3851;
	wire [4-1:0] node3854;
	wire [4-1:0] node3857;
	wire [4-1:0] node3858;
	wire [4-1:0] node3859;
	wire [4-1:0] node3860;
	wire [4-1:0] node3864;
	wire [4-1:0] node3867;
	wire [4-1:0] node3868;
	wire [4-1:0] node3871;
	wire [4-1:0] node3874;
	wire [4-1:0] node3875;
	wire [4-1:0] node3876;
	wire [4-1:0] node3877;
	wire [4-1:0] node3879;
	wire [4-1:0] node3881;
	wire [4-1:0] node3884;
	wire [4-1:0] node3885;
	wire [4-1:0] node3888;
	wire [4-1:0] node3889;
	wire [4-1:0] node3890;
	wire [4-1:0] node3894;
	wire [4-1:0] node3897;
	wire [4-1:0] node3898;
	wire [4-1:0] node3901;
	wire [4-1:0] node3903;
	wire [4-1:0] node3905;
	wire [4-1:0] node3908;
	wire [4-1:0] node3909;
	wire [4-1:0] node3910;
	wire [4-1:0] node3913;
	wire [4-1:0] node3914;
	wire [4-1:0] node3918;
	wire [4-1:0] node3919;
	wire [4-1:0] node3921;
	wire [4-1:0] node3922;
	wire [4-1:0] node3925;
	wire [4-1:0] node3928;
	wire [4-1:0] node3930;
	wire [4-1:0] node3933;
	wire [4-1:0] node3934;
	wire [4-1:0] node3935;
	wire [4-1:0] node3936;
	wire [4-1:0] node3937;
	wire [4-1:0] node3938;
	wire [4-1:0] node3939;
	wire [4-1:0] node3940;
	wire [4-1:0] node3941;
	wire [4-1:0] node3945;
	wire [4-1:0] node3946;
	wire [4-1:0] node3950;
	wire [4-1:0] node3951;
	wire [4-1:0] node3955;
	wire [4-1:0] node3956;
	wire [4-1:0] node3957;
	wire [4-1:0] node3961;
	wire [4-1:0] node3963;
	wire [4-1:0] node3965;
	wire [4-1:0] node3968;
	wire [4-1:0] node3969;
	wire [4-1:0] node3972;
	wire [4-1:0] node3973;
	wire [4-1:0] node3974;
	wire [4-1:0] node3978;
	wire [4-1:0] node3980;
	wire [4-1:0] node3983;
	wire [4-1:0] node3984;
	wire [4-1:0] node3985;
	wire [4-1:0] node3986;
	wire [4-1:0] node3988;
	wire [4-1:0] node3989;
	wire [4-1:0] node3993;
	wire [4-1:0] node3994;
	wire [4-1:0] node3999;
	wire [4-1:0] node4000;
	wire [4-1:0] node4002;
	wire [4-1:0] node4003;
	wire [4-1:0] node4006;
	wire [4-1:0] node4007;
	wire [4-1:0] node4011;
	wire [4-1:0] node4012;
	wire [4-1:0] node4014;
	wire [4-1:0] node4017;
	wire [4-1:0] node4019;
	wire [4-1:0] node4020;
	wire [4-1:0] node4024;
	wire [4-1:0] node4025;
	wire [4-1:0] node4026;
	wire [4-1:0] node4027;
	wire [4-1:0] node4030;
	wire [4-1:0] node4031;
	wire [4-1:0] node4035;
	wire [4-1:0] node4036;
	wire [4-1:0] node4037;
	wire [4-1:0] node4038;
	wire [4-1:0] node4041;
	wire [4-1:0] node4045;
	wire [4-1:0] node4046;
	wire [4-1:0] node4048;
	wire [4-1:0] node4052;
	wire [4-1:0] node4053;
	wire [4-1:0] node4054;
	wire [4-1:0] node4056;
	wire [4-1:0] node4059;
	wire [4-1:0] node4061;
	wire [4-1:0] node4064;
	wire [4-1:0] node4065;
	wire [4-1:0] node4067;
	wire [4-1:0] node4068;
	wire [4-1:0] node4072;
	wire [4-1:0] node4073;
	wire [4-1:0] node4074;
	wire [4-1:0] node4075;
	wire [4-1:0] node4079;
	wire [4-1:0] node4080;
	wire [4-1:0] node4085;
	wire [4-1:0] node4086;
	wire [4-1:0] node4087;
	wire [4-1:0] node4088;
	wire [4-1:0] node4089;
	wire [4-1:0] node4092;
	wire [4-1:0] node4094;
	wire [4-1:0] node4095;
	wire [4-1:0] node4099;
	wire [4-1:0] node4100;
	wire [4-1:0] node4102;
	wire [4-1:0] node4103;
	wire [4-1:0] node4106;
	wire [4-1:0] node4107;
	wire [4-1:0] node4111;
	wire [4-1:0] node4113;
	wire [4-1:0] node4116;
	wire [4-1:0] node4117;
	wire [4-1:0] node4118;
	wire [4-1:0] node4119;
	wire [4-1:0] node4120;
	wire [4-1:0] node4124;
	wire [4-1:0] node4126;
	wire [4-1:0] node4127;
	wire [4-1:0] node4131;
	wire [4-1:0] node4132;
	wire [4-1:0] node4135;
	wire [4-1:0] node4138;
	wire [4-1:0] node4139;
	wire [4-1:0] node4140;
	wire [4-1:0] node4141;
	wire [4-1:0] node4143;
	wire [4-1:0] node4147;
	wire [4-1:0] node4148;
	wire [4-1:0] node4152;
	wire [4-1:0] node4155;
	wire [4-1:0] node4156;
	wire [4-1:0] node4157;
	wire [4-1:0] node4158;
	wire [4-1:0] node4159;
	wire [4-1:0] node4161;
	wire [4-1:0] node4162;
	wire [4-1:0] node4166;
	wire [4-1:0] node4169;
	wire [4-1:0] node4170;
	wire [4-1:0] node4172;
	wire [4-1:0] node4175;
	wire [4-1:0] node4177;
	wire [4-1:0] node4180;
	wire [4-1:0] node4181;
	wire [4-1:0] node4182;
	wire [4-1:0] node4185;
	wire [4-1:0] node4187;
	wire [4-1:0] node4190;
	wire [4-1:0] node4191;
	wire [4-1:0] node4192;
	wire [4-1:0] node4196;
	wire [4-1:0] node4199;
	wire [4-1:0] node4200;
	wire [4-1:0] node4201;
	wire [4-1:0] node4202;
	wire [4-1:0] node4204;
	wire [4-1:0] node4206;
	wire [4-1:0] node4209;
	wire [4-1:0] node4210;
	wire [4-1:0] node4214;
	wire [4-1:0] node4215;
	wire [4-1:0] node4218;
	wire [4-1:0] node4220;
	wire [4-1:0] node4223;
	wire [4-1:0] node4224;
	wire [4-1:0] node4225;
	wire [4-1:0] node4226;
	wire [4-1:0] node4231;
	wire [4-1:0] node4232;
	wire [4-1:0] node4233;
	wire [4-1:0] node4235;
	wire [4-1:0] node4238;
	wire [4-1:0] node4242;
	wire [4-1:0] node4243;
	wire [4-1:0] node4244;
	wire [4-1:0] node4245;
	wire [4-1:0] node4246;
	wire [4-1:0] node4247;
	wire [4-1:0] node4248;
	wire [4-1:0] node4249;
	wire [4-1:0] node4250;
	wire [4-1:0] node4251;
	wire [4-1:0] node4255;
	wire [4-1:0] node4257;
	wire [4-1:0] node4260;
	wire [4-1:0] node4261;
	wire [4-1:0] node4265;
	wire [4-1:0] node4266;
	wire [4-1:0] node4267;
	wire [4-1:0] node4270;
	wire [4-1:0] node4271;
	wire [4-1:0] node4275;
	wire [4-1:0] node4278;
	wire [4-1:0] node4279;
	wire [4-1:0] node4280;
	wire [4-1:0] node4283;
	wire [4-1:0] node4284;
	wire [4-1:0] node4285;
	wire [4-1:0] node4289;
	wire [4-1:0] node4291;
	wire [4-1:0] node4292;
	wire [4-1:0] node4296;
	wire [4-1:0] node4297;
	wire [4-1:0] node4298;
	wire [4-1:0] node4299;
	wire [4-1:0] node4300;
	wire [4-1:0] node4304;
	wire [4-1:0] node4307;
	wire [4-1:0] node4309;
	wire [4-1:0] node4310;
	wire [4-1:0] node4314;
	wire [4-1:0] node4315;
	wire [4-1:0] node4317;
	wire [4-1:0] node4319;
	wire [4-1:0] node4323;
	wire [4-1:0] node4324;
	wire [4-1:0] node4325;
	wire [4-1:0] node4326;
	wire [4-1:0] node4327;
	wire [4-1:0] node4328;
	wire [4-1:0] node4329;
	wire [4-1:0] node4333;
	wire [4-1:0] node4336;
	wire [4-1:0] node4337;
	wire [4-1:0] node4341;
	wire [4-1:0] node4342;
	wire [4-1:0] node4343;
	wire [4-1:0] node4346;
	wire [4-1:0] node4349;
	wire [4-1:0] node4351;
	wire [4-1:0] node4354;
	wire [4-1:0] node4355;
	wire [4-1:0] node4356;
	wire [4-1:0] node4360;
	wire [4-1:0] node4363;
	wire [4-1:0] node4364;
	wire [4-1:0] node4365;
	wire [4-1:0] node4366;
	wire [4-1:0] node4368;
	wire [4-1:0] node4371;
	wire [4-1:0] node4372;
	wire [4-1:0] node4376;
	wire [4-1:0] node4378;
	wire [4-1:0] node4380;
	wire [4-1:0] node4382;
	wire [4-1:0] node4385;
	wire [4-1:0] node4386;
	wire [4-1:0] node4387;
	wire [4-1:0] node4389;
	wire [4-1:0] node4393;
	wire [4-1:0] node4394;
	wire [4-1:0] node4395;
	wire [4-1:0] node4399;
	wire [4-1:0] node4402;
	wire [4-1:0] node4403;
	wire [4-1:0] node4404;
	wire [4-1:0] node4405;
	wire [4-1:0] node4406;
	wire [4-1:0] node4407;
	wire [4-1:0] node4408;
	wire [4-1:0] node4413;
	wire [4-1:0] node4416;
	wire [4-1:0] node4417;
	wire [4-1:0] node4418;
	wire [4-1:0] node4421;
	wire [4-1:0] node4424;
	wire [4-1:0] node4425;
	wire [4-1:0] node4426;
	wire [4-1:0] node4428;
	wire [4-1:0] node4433;
	wire [4-1:0] node4434;
	wire [4-1:0] node4435;
	wire [4-1:0] node4436;
	wire [4-1:0] node4438;
	wire [4-1:0] node4442;
	wire [4-1:0] node4443;
	wire [4-1:0] node4444;
	wire [4-1:0] node4448;
	wire [4-1:0] node4449;
	wire [4-1:0] node4450;
	wire [4-1:0] node4454;
	wire [4-1:0] node4456;
	wire [4-1:0] node4459;
	wire [4-1:0] node4460;
	wire [4-1:0] node4461;
	wire [4-1:0] node4462;
	wire [4-1:0] node4465;
	wire [4-1:0] node4467;
	wire [4-1:0] node4471;
	wire [4-1:0] node4472;
	wire [4-1:0] node4473;
	wire [4-1:0] node4474;
	wire [4-1:0] node4477;
	wire [4-1:0] node4481;
	wire [4-1:0] node4482;
	wire [4-1:0] node4485;
	wire [4-1:0] node4488;
	wire [4-1:0] node4489;
	wire [4-1:0] node4490;
	wire [4-1:0] node4491;
	wire [4-1:0] node4492;
	wire [4-1:0] node4495;
	wire [4-1:0] node4496;
	wire [4-1:0] node4500;
	wire [4-1:0] node4501;
	wire [4-1:0] node4502;
	wire [4-1:0] node4505;
	wire [4-1:0] node4509;
	wire [4-1:0] node4510;
	wire [4-1:0] node4511;
	wire [4-1:0] node4513;
	wire [4-1:0] node4517;
	wire [4-1:0] node4519;
	wire [4-1:0] node4521;
	wire [4-1:0] node4524;
	wire [4-1:0] node4525;
	wire [4-1:0] node4526;
	wire [4-1:0] node4527;
	wire [4-1:0] node4529;
	wire [4-1:0] node4532;
	wire [4-1:0] node4535;
	wire [4-1:0] node4536;
	wire [4-1:0] node4537;
	wire [4-1:0] node4539;
	wire [4-1:0] node4543;
	wire [4-1:0] node4544;
	wire [4-1:0] node4545;
	wire [4-1:0] node4549;
	wire [4-1:0] node4552;
	wire [4-1:0] node4553;
	wire [4-1:0] node4554;
	wire [4-1:0] node4555;
	wire [4-1:0] node4559;
	wire [4-1:0] node4561;
	wire [4-1:0] node4564;
	wire [4-1:0] node4566;
	wire [4-1:0] node4567;
	wire [4-1:0] node4571;
	wire [4-1:0] node4572;
	wire [4-1:0] node4573;
	wire [4-1:0] node4574;
	wire [4-1:0] node4575;
	wire [4-1:0] node4576;
	wire [4-1:0] node4577;
	wire [4-1:0] node4578;
	wire [4-1:0] node4580;
	wire [4-1:0] node4584;
	wire [4-1:0] node4586;
	wire [4-1:0] node4589;
	wire [4-1:0] node4590;
	wire [4-1:0] node4591;
	wire [4-1:0] node4594;
	wire [4-1:0] node4597;
	wire [4-1:0] node4600;
	wire [4-1:0] node4601;
	wire [4-1:0] node4602;
	wire [4-1:0] node4605;
	wire [4-1:0] node4606;
	wire [4-1:0] node4607;
	wire [4-1:0] node4611;
	wire [4-1:0] node4614;
	wire [4-1:0] node4617;
	wire [4-1:0] node4618;
	wire [4-1:0] node4619;
	wire [4-1:0] node4620;
	wire [4-1:0] node4622;
	wire [4-1:0] node4626;
	wire [4-1:0] node4628;
	wire [4-1:0] node4631;
	wire [4-1:0] node4632;
	wire [4-1:0] node4633;
	wire [4-1:0] node4634;
	wire [4-1:0] node4636;
	wire [4-1:0] node4639;
	wire [4-1:0] node4642;
	wire [4-1:0] node4645;
	wire [4-1:0] node4646;
	wire [4-1:0] node4647;
	wire [4-1:0] node4651;
	wire [4-1:0] node4653;
	wire [4-1:0] node4654;
	wire [4-1:0] node4658;
	wire [4-1:0] node4659;
	wire [4-1:0] node4660;
	wire [4-1:0] node4661;
	wire [4-1:0] node4662;
	wire [4-1:0] node4664;
	wire [4-1:0] node4666;
	wire [4-1:0] node4669;
	wire [4-1:0] node4671;
	wire [4-1:0] node4674;
	wire [4-1:0] node4675;
	wire [4-1:0] node4678;
	wire [4-1:0] node4679;
	wire [4-1:0] node4682;
	wire [4-1:0] node4684;
	wire [4-1:0] node4687;
	wire [4-1:0] node4688;
	wire [4-1:0] node4689;
	wire [4-1:0] node4692;
	wire [4-1:0] node4694;
	wire [4-1:0] node4695;
	wire [4-1:0] node4699;
	wire [4-1:0] node4700;
	wire [4-1:0] node4702;
	wire [4-1:0] node4705;
	wire [4-1:0] node4707;
	wire [4-1:0] node4708;
	wire [4-1:0] node4712;
	wire [4-1:0] node4713;
	wire [4-1:0] node4714;
	wire [4-1:0] node4716;
	wire [4-1:0] node4719;
	wire [4-1:0] node4720;
	wire [4-1:0] node4723;
	wire [4-1:0] node4725;
	wire [4-1:0] node4728;
	wire [4-1:0] node4729;
	wire [4-1:0] node4730;
	wire [4-1:0] node4734;
	wire [4-1:0] node4736;
	wire [4-1:0] node4737;
	wire [4-1:0] node4738;
	wire [4-1:0] node4742;
	wire [4-1:0] node4743;
	wire [4-1:0] node4747;
	wire [4-1:0] node4748;
	wire [4-1:0] node4749;
	wire [4-1:0] node4750;
	wire [4-1:0] node4751;
	wire [4-1:0] node4753;
	wire [4-1:0] node4755;
	wire [4-1:0] node4756;
	wire [4-1:0] node4760;
	wire [4-1:0] node4761;
	wire [4-1:0] node4763;
	wire [4-1:0] node4764;
	wire [4-1:0] node4768;
	wire [4-1:0] node4769;
	wire [4-1:0] node4771;
	wire [4-1:0] node4774;
	wire [4-1:0] node4775;
	wire [4-1:0] node4779;
	wire [4-1:0] node4780;
	wire [4-1:0] node4781;
	wire [4-1:0] node4783;
	wire [4-1:0] node4786;
	wire [4-1:0] node4787;
	wire [4-1:0] node4790;
	wire [4-1:0] node4791;
	wire [4-1:0] node4795;
	wire [4-1:0] node4796;
	wire [4-1:0] node4798;
	wire [4-1:0] node4802;
	wire [4-1:0] node4803;
	wire [4-1:0] node4804;
	wire [4-1:0] node4806;
	wire [4-1:0] node4808;
	wire [4-1:0] node4809;
	wire [4-1:0] node4812;
	wire [4-1:0] node4815;
	wire [4-1:0] node4816;
	wire [4-1:0] node4817;
	wire [4-1:0] node4819;
	wire [4-1:0] node4823;
	wire [4-1:0] node4824;
	wire [4-1:0] node4828;
	wire [4-1:0] node4829;
	wire [4-1:0] node4832;
	wire [4-1:0] node4834;
	wire [4-1:0] node4837;
	wire [4-1:0] node4838;
	wire [4-1:0] node4839;
	wire [4-1:0] node4840;
	wire [4-1:0] node4841;
	wire [4-1:0] node4845;
	wire [4-1:0] node4846;
	wire [4-1:0] node4849;
	wire [4-1:0] node4850;
	wire [4-1:0] node4851;
	wire [4-1:0] node4856;
	wire [4-1:0] node4857;
	wire [4-1:0] node4858;
	wire [4-1:0] node4859;
	wire [4-1:0] node4864;
	wire [4-1:0] node4866;
	wire [4-1:0] node4868;
	wire [4-1:0] node4871;
	wire [4-1:0] node4872;
	wire [4-1:0] node4873;
	wire [4-1:0] node4874;
	wire [4-1:0] node4875;
	wire [4-1:0] node4878;
	wire [4-1:0] node4880;
	wire [4-1:0] node4883;
	wire [4-1:0] node4886;
	wire [4-1:0] node4888;
	wire [4-1:0] node4889;
	wire [4-1:0] node4890;
	wire [4-1:0] node4893;
	wire [4-1:0] node4897;
	wire [4-1:0] node4898;
	wire [4-1:0] node4900;
	wire [4-1:0] node4901;
	wire [4-1:0] node4905;
	wire [4-1:0] node4906;
	wire [4-1:0] node4907;
	wire [4-1:0] node4911;
	wire [4-1:0] node4912;
	wire [4-1:0] node4916;
	wire [4-1:0] node4917;
	wire [4-1:0] node4918;
	wire [4-1:0] node4919;
	wire [4-1:0] node4920;
	wire [4-1:0] node4921;
	wire [4-1:0] node4922;
	wire [4-1:0] node4923;
	wire [4-1:0] node4926;
	wire [4-1:0] node4927;
	wire [4-1:0] node4930;
	wire [4-1:0] node4932;
	wire [4-1:0] node4935;
	wire [4-1:0] node4936;
	wire [4-1:0] node4937;
	wire [4-1:0] node4941;
	wire [4-1:0] node4944;
	wire [4-1:0] node4945;
	wire [4-1:0] node4946;
	wire [4-1:0] node4949;
	wire [4-1:0] node4952;
	wire [4-1:0] node4953;
	wire [4-1:0] node4955;
	wire [4-1:0] node4956;
	wire [4-1:0] node4960;
	wire [4-1:0] node4963;
	wire [4-1:0] node4964;
	wire [4-1:0] node4965;
	wire [4-1:0] node4967;
	wire [4-1:0] node4968;
	wire [4-1:0] node4972;
	wire [4-1:0] node4973;
	wire [4-1:0] node4975;
	wire [4-1:0] node4976;
	wire [4-1:0] node4979;
	wire [4-1:0] node4983;
	wire [4-1:0] node4984;
	wire [4-1:0] node4985;
	wire [4-1:0] node4987;
	wire [4-1:0] node4990;
	wire [4-1:0] node4993;
	wire [4-1:0] node4995;
	wire [4-1:0] node4996;
	wire [4-1:0] node5000;
	wire [4-1:0] node5001;
	wire [4-1:0] node5002;
	wire [4-1:0] node5003;
	wire [4-1:0] node5004;
	wire [4-1:0] node5006;
	wire [4-1:0] node5009;
	wire [4-1:0] node5011;
	wire [4-1:0] node5014;
	wire [4-1:0] node5015;
	wire [4-1:0] node5018;
	wire [4-1:0] node5019;
	wire [4-1:0] node5020;
	wire [4-1:0] node5025;
	wire [4-1:0] node5026;
	wire [4-1:0] node5027;
	wire [4-1:0] node5028;
	wire [4-1:0] node5032;
	wire [4-1:0] node5033;
	wire [4-1:0] node5034;
	wire [4-1:0] node5039;
	wire [4-1:0] node5040;
	wire [4-1:0] node5042;
	wire [4-1:0] node5045;
	wire [4-1:0] node5048;
	wire [4-1:0] node5049;
	wire [4-1:0] node5050;
	wire [4-1:0] node5051;
	wire [4-1:0] node5055;
	wire [4-1:0] node5056;
	wire [4-1:0] node5058;
	wire [4-1:0] node5060;
	wire [4-1:0] node5063;
	wire [4-1:0] node5065;
	wire [4-1:0] node5068;
	wire [4-1:0] node5069;
	wire [4-1:0] node5070;
	wire [4-1:0] node5071;
	wire [4-1:0] node5075;
	wire [4-1:0] node5077;
	wire [4-1:0] node5079;
	wire [4-1:0] node5082;
	wire [4-1:0] node5083;
	wire [4-1:0] node5086;
	wire [4-1:0] node5087;
	wire [4-1:0] node5091;
	wire [4-1:0] node5092;
	wire [4-1:0] node5093;
	wire [4-1:0] node5094;
	wire [4-1:0] node5095;
	wire [4-1:0] node5096;
	wire [4-1:0] node5098;
	wire [4-1:0] node5101;
	wire [4-1:0] node5103;
	wire [4-1:0] node5106;
	wire [4-1:0] node5107;
	wire [4-1:0] node5108;
	wire [4-1:0] node5112;
	wire [4-1:0] node5113;
	wire [4-1:0] node5114;
	wire [4-1:0] node5118;
	wire [4-1:0] node5119;
	wire [4-1:0] node5122;
	wire [4-1:0] node5125;
	wire [4-1:0] node5126;
	wire [4-1:0] node5127;
	wire [4-1:0] node5128;
	wire [4-1:0] node5129;
	wire [4-1:0] node5133;
	wire [4-1:0] node5134;
	wire [4-1:0] node5138;
	wire [4-1:0] node5140;
	wire [4-1:0] node5142;
	wire [4-1:0] node5145;
	wire [4-1:0] node5146;
	wire [4-1:0] node5147;
	wire [4-1:0] node5150;
	wire [4-1:0] node5153;
	wire [4-1:0] node5156;
	wire [4-1:0] node5157;
	wire [4-1:0] node5158;
	wire [4-1:0] node5159;
	wire [4-1:0] node5161;
	wire [4-1:0] node5164;
	wire [4-1:0] node5166;
	wire [4-1:0] node5169;
	wire [4-1:0] node5170;
	wire [4-1:0] node5172;
	wire [4-1:0] node5175;
	wire [4-1:0] node5177;
	wire [4-1:0] node5178;
	wire [4-1:0] node5182;
	wire [4-1:0] node5183;
	wire [4-1:0] node5186;
	wire [4-1:0] node5187;
	wire [4-1:0] node5189;
	wire [4-1:0] node5193;
	wire [4-1:0] node5194;
	wire [4-1:0] node5195;
	wire [4-1:0] node5196;
	wire [4-1:0] node5198;
	wire [4-1:0] node5200;
	wire [4-1:0] node5203;
	wire [4-1:0] node5204;
	wire [4-1:0] node5208;
	wire [4-1:0] node5209;
	wire [4-1:0] node5210;
	wire [4-1:0] node5211;
	wire [4-1:0] node5212;
	wire [4-1:0] node5217;
	wire [4-1:0] node5219;
	wire [4-1:0] node5222;
	wire [4-1:0] node5223;
	wire [4-1:0] node5226;
	wire [4-1:0] node5229;
	wire [4-1:0] node5230;
	wire [4-1:0] node5231;
	wire [4-1:0] node5232;
	wire [4-1:0] node5233;
	wire [4-1:0] node5237;
	wire [4-1:0] node5238;
	wire [4-1:0] node5242;
	wire [4-1:0] node5243;
	wire [4-1:0] node5245;
	wire [4-1:0] node5248;
	wire [4-1:0] node5251;
	wire [4-1:0] node5252;
	wire [4-1:0] node5253;
	wire [4-1:0] node5254;
	wire [4-1:0] node5255;
	wire [4-1:0] node5259;
	wire [4-1:0] node5260;
	wire [4-1:0] node5264;
	wire [4-1:0] node5266;
	wire [4-1:0] node5269;
	wire [4-1:0] node5270;
	wire [4-1:0] node5272;
	wire [4-1:0] node5276;
	wire [4-1:0] node5277;
	wire [4-1:0] node5278;
	wire [4-1:0] node5279;
	wire [4-1:0] node5280;
	wire [4-1:0] node5281;
	wire [4-1:0] node5282;
	wire [4-1:0] node5285;
	wire [4-1:0] node5286;
	wire [4-1:0] node5289;
	wire [4-1:0] node5292;
	wire [4-1:0] node5293;
	wire [4-1:0] node5295;
	wire [4-1:0] node5298;
	wire [4-1:0] node5300;
	wire [4-1:0] node5303;
	wire [4-1:0] node5304;
	wire [4-1:0] node5307;
	wire [4-1:0] node5308;
	wire [4-1:0] node5310;
	wire [4-1:0] node5314;
	wire [4-1:0] node5315;
	wire [4-1:0] node5316;
	wire [4-1:0] node5318;
	wire [4-1:0] node5319;
	wire [4-1:0] node5321;
	wire [4-1:0] node5324;
	wire [4-1:0] node5325;
	wire [4-1:0] node5328;
	wire [4-1:0] node5331;
	wire [4-1:0] node5333;
	wire [4-1:0] node5334;
	wire [4-1:0] node5336;
	wire [4-1:0] node5340;
	wire [4-1:0] node5341;
	wire [4-1:0] node5342;
	wire [4-1:0] node5343;
	wire [4-1:0] node5345;
	wire [4-1:0] node5349;
	wire [4-1:0] node5351;
	wire [4-1:0] node5354;
	wire [4-1:0] node5355;
	wire [4-1:0] node5356;
	wire [4-1:0] node5357;
	wire [4-1:0] node5360;
	wire [4-1:0] node5364;
	wire [4-1:0] node5367;
	wire [4-1:0] node5368;
	wire [4-1:0] node5369;
	wire [4-1:0] node5370;
	wire [4-1:0] node5371;
	wire [4-1:0] node5374;
	wire [4-1:0] node5375;
	wire [4-1:0] node5379;
	wire [4-1:0] node5380;
	wire [4-1:0] node5381;
	wire [4-1:0] node5385;
	wire [4-1:0] node5386;
	wire [4-1:0] node5389;
	wire [4-1:0] node5392;
	wire [4-1:0] node5393;
	wire [4-1:0] node5394;
	wire [4-1:0] node5395;
	wire [4-1:0] node5399;
	wire [4-1:0] node5401;
	wire [4-1:0] node5402;
	wire [4-1:0] node5406;
	wire [4-1:0] node5407;
	wire [4-1:0] node5409;
	wire [4-1:0] node5412;
	wire [4-1:0] node5413;
	wire [4-1:0] node5416;
	wire [4-1:0] node5419;
	wire [4-1:0] node5420;
	wire [4-1:0] node5421;
	wire [4-1:0] node5422;
	wire [4-1:0] node5424;
	wire [4-1:0] node5427;
	wire [4-1:0] node5430;
	wire [4-1:0] node5431;
	wire [4-1:0] node5433;
	wire [4-1:0] node5436;
	wire [4-1:0] node5438;
	wire [4-1:0] node5440;
	wire [4-1:0] node5443;
	wire [4-1:0] node5444;
	wire [4-1:0] node5446;
	wire [4-1:0] node5448;
	wire [4-1:0] node5451;
	wire [4-1:0] node5454;
	wire [4-1:0] node5455;
	wire [4-1:0] node5456;
	wire [4-1:0] node5457;
	wire [4-1:0] node5458;
	wire [4-1:0] node5459;
	wire [4-1:0] node5460;
	wire [4-1:0] node5464;
	wire [4-1:0] node5465;
	wire [4-1:0] node5468;
	wire [4-1:0] node5469;
	wire [4-1:0] node5473;
	wire [4-1:0] node5475;
	wire [4-1:0] node5476;
	wire [4-1:0] node5480;
	wire [4-1:0] node5481;
	wire [4-1:0] node5482;
	wire [4-1:0] node5484;
	wire [4-1:0] node5485;
	wire [4-1:0] node5489;
	wire [4-1:0] node5490;
	wire [4-1:0] node5494;
	wire [4-1:0] node5495;
	wire [4-1:0] node5499;
	wire [4-1:0] node5500;
	wire [4-1:0] node5501;
	wire [4-1:0] node5502;
	wire [4-1:0] node5503;
	wire [4-1:0] node5504;
	wire [4-1:0] node5509;
	wire [4-1:0] node5510;
	wire [4-1:0] node5513;
	wire [4-1:0] node5515;
	wire [4-1:0] node5518;
	wire [4-1:0] node5519;
	wire [4-1:0] node5520;
	wire [4-1:0] node5524;
	wire [4-1:0] node5527;
	wire [4-1:0] node5529;
	wire [4-1:0] node5530;
	wire [4-1:0] node5531;
	wire [4-1:0] node5534;
	wire [4-1:0] node5536;
	wire [4-1:0] node5539;
	wire [4-1:0] node5540;
	wire [4-1:0] node5542;
	wire [4-1:0] node5546;
	wire [4-1:0] node5547;
	wire [4-1:0] node5548;
	wire [4-1:0] node5549;
	wire [4-1:0] node5550;
	wire [4-1:0] node5551;
	wire [4-1:0] node5554;
	wire [4-1:0] node5557;
	wire [4-1:0] node5559;
	wire [4-1:0] node5562;
	wire [4-1:0] node5563;
	wire [4-1:0] node5567;
	wire [4-1:0] node5568;
	wire [4-1:0] node5569;
	wire [4-1:0] node5570;
	wire [4-1:0] node5572;
	wire [4-1:0] node5576;
	wire [4-1:0] node5578;
	wire [4-1:0] node5579;
	wire [4-1:0] node5582;
	wire [4-1:0] node5585;
	wire [4-1:0] node5586;
	wire [4-1:0] node5587;
	wire [4-1:0] node5590;
	wire [4-1:0] node5593;
	wire [4-1:0] node5594;
	wire [4-1:0] node5595;
	wire [4-1:0] node5600;
	wire [4-1:0] node5601;
	wire [4-1:0] node5602;
	wire [4-1:0] node5603;
	wire [4-1:0] node5604;
	wire [4-1:0] node5605;
	wire [4-1:0] node5610;
	wire [4-1:0] node5611;
	wire [4-1:0] node5612;
	wire [4-1:0] node5616;
	wire [4-1:0] node5619;
	wire [4-1:0] node5621;
	wire [4-1:0] node5624;
	wire [4-1:0] node5625;
	wire [4-1:0] node5626;
	wire [4-1:0] node5628;
	wire [4-1:0] node5631;
	wire [4-1:0] node5633;
	wire [4-1:0] node5636;
	wire [4-1:0] node5637;
	wire [4-1:0] node5639;
	wire [4-1:0] node5642;
	wire [4-1:0] node5643;
	wire [4-1:0] node5644;
	wire [4-1:0] node5649;
	wire [4-1:0] node5650;
	wire [4-1:0] node5651;
	wire [4-1:0] node5652;
	wire [4-1:0] node5653;
	wire [4-1:0] node5654;
	wire [4-1:0] node5655;
	wire [4-1:0] node5656;
	wire [4-1:0] node5657;
	wire [4-1:0] node5658;
	wire [4-1:0] node5661;
	wire [4-1:0] node5662;
	wire [4-1:0] node5665;
	wire [4-1:0] node5668;
	wire [4-1:0] node5669;
	wire [4-1:0] node5670;
	wire [4-1:0] node5673;
	wire [4-1:0] node5676;
	wire [4-1:0] node5677;
	wire [4-1:0] node5678;
	wire [4-1:0] node5682;
	wire [4-1:0] node5684;
	wire [4-1:0] node5687;
	wire [4-1:0] node5688;
	wire [4-1:0] node5689;
	wire [4-1:0] node5691;
	wire [4-1:0] node5692;
	wire [4-1:0] node5697;
	wire [4-1:0] node5698;
	wire [4-1:0] node5699;
	wire [4-1:0] node5701;
	wire [4-1:0] node5702;
	wire [4-1:0] node5705;
	wire [4-1:0] node5708;
	wire [4-1:0] node5709;
	wire [4-1:0] node5710;
	wire [4-1:0] node5715;
	wire [4-1:0] node5716;
	wire [4-1:0] node5717;
	wire [4-1:0] node5718;
	wire [4-1:0] node5721;
	wire [4-1:0] node5726;
	wire [4-1:0] node5727;
	wire [4-1:0] node5728;
	wire [4-1:0] node5729;
	wire [4-1:0] node5730;
	wire [4-1:0] node5734;
	wire [4-1:0] node5735;
	wire [4-1:0] node5737;
	wire [4-1:0] node5740;
	wire [4-1:0] node5741;
	wire [4-1:0] node5745;
	wire [4-1:0] node5746;
	wire [4-1:0] node5747;
	wire [4-1:0] node5751;
	wire [4-1:0] node5752;
	wire [4-1:0] node5755;
	wire [4-1:0] node5757;
	wire [4-1:0] node5758;
	wire [4-1:0] node5761;
	wire [4-1:0] node5764;
	wire [4-1:0] node5765;
	wire [4-1:0] node5766;
	wire [4-1:0] node5767;
	wire [4-1:0] node5769;
	wire [4-1:0] node5772;
	wire [4-1:0] node5774;
	wire [4-1:0] node5775;
	wire [4-1:0] node5779;
	wire [4-1:0] node5780;
	wire [4-1:0] node5781;
	wire [4-1:0] node5782;
	wire [4-1:0] node5787;
	wire [4-1:0] node5789;
	wire [4-1:0] node5791;
	wire [4-1:0] node5794;
	wire [4-1:0] node5795;
	wire [4-1:0] node5796;
	wire [4-1:0] node5797;
	wire [4-1:0] node5801;
	wire [4-1:0] node5802;
	wire [4-1:0] node5803;
	wire [4-1:0] node5808;
	wire [4-1:0] node5809;
	wire [4-1:0] node5810;
	wire [4-1:0] node5814;
	wire [4-1:0] node5815;
	wire [4-1:0] node5816;
	wire [4-1:0] node5819;
	wire [4-1:0] node5823;
	wire [4-1:0] node5824;
	wire [4-1:0] node5825;
	wire [4-1:0] node5826;
	wire [4-1:0] node5827;
	wire [4-1:0] node5828;
	wire [4-1:0] node5829;
	wire [4-1:0] node5832;
	wire [4-1:0] node5834;
	wire [4-1:0] node5838;
	wire [4-1:0] node5839;
	wire [4-1:0] node5840;
	wire [4-1:0] node5844;
	wire [4-1:0] node5847;
	wire [4-1:0] node5848;
	wire [4-1:0] node5849;
	wire [4-1:0] node5850;
	wire [4-1:0] node5853;
	wire [4-1:0] node5856;
	wire [4-1:0] node5857;
	wire [4-1:0] node5858;
	wire [4-1:0] node5862;
	wire [4-1:0] node5863;
	wire [4-1:0] node5866;
	wire [4-1:0] node5869;
	wire [4-1:0] node5870;
	wire [4-1:0] node5871;
	wire [4-1:0] node5872;
	wire [4-1:0] node5877;
	wire [4-1:0] node5880;
	wire [4-1:0] node5881;
	wire [4-1:0] node5882;
	wire [4-1:0] node5883;
	wire [4-1:0] node5885;
	wire [4-1:0] node5887;
	wire [4-1:0] node5891;
	wire [4-1:0] node5892;
	wire [4-1:0] node5895;
	wire [4-1:0] node5898;
	wire [4-1:0] node5899;
	wire [4-1:0] node5900;
	wire [4-1:0] node5901;
	wire [4-1:0] node5902;
	wire [4-1:0] node5907;
	wire [4-1:0] node5909;
	wire [4-1:0] node5912;
	wire [4-1:0] node5914;
	wire [4-1:0] node5915;
	wire [4-1:0] node5917;
	wire [4-1:0] node5921;
	wire [4-1:0] node5922;
	wire [4-1:0] node5923;
	wire [4-1:0] node5924;
	wire [4-1:0] node5927;
	wire [4-1:0] node5928;
	wire [4-1:0] node5929;
	wire [4-1:0] node5932;
	wire [4-1:0] node5933;
	wire [4-1:0] node5937;
	wire [4-1:0] node5940;
	wire [4-1:0] node5941;
	wire [4-1:0] node5943;
	wire [4-1:0] node5944;
	wire [4-1:0] node5946;
	wire [4-1:0] node5950;
	wire [4-1:0] node5951;
	wire [4-1:0] node5954;
	wire [4-1:0] node5955;
	wire [4-1:0] node5958;
	wire [4-1:0] node5961;
	wire [4-1:0] node5962;
	wire [4-1:0] node5963;
	wire [4-1:0] node5964;
	wire [4-1:0] node5965;
	wire [4-1:0] node5966;
	wire [4-1:0] node5971;
	wire [4-1:0] node5972;
	wire [4-1:0] node5977;
	wire [4-1:0] node5978;
	wire [4-1:0] node5979;
	wire [4-1:0] node5982;
	wire [4-1:0] node5983;
	wire [4-1:0] node5986;
	wire [4-1:0] node5989;
	wire [4-1:0] node5990;
	wire [4-1:0] node5993;
	wire [4-1:0] node5995;
	wire [4-1:0] node5996;
	wire [4-1:0] node6000;
	wire [4-1:0] node6001;
	wire [4-1:0] node6002;
	wire [4-1:0] node6003;
	wire [4-1:0] node6004;
	wire [4-1:0] node6005;
	wire [4-1:0] node6007;
	wire [4-1:0] node6010;
	wire [4-1:0] node6011;
	wire [4-1:0] node6012;
	wire [4-1:0] node6013;
	wire [4-1:0] node6018;
	wire [4-1:0] node6019;
	wire [4-1:0] node6023;
	wire [4-1:0] node6024;
	wire [4-1:0] node6025;
	wire [4-1:0] node6026;
	wire [4-1:0] node6029;
	wire [4-1:0] node6032;
	wire [4-1:0] node6033;
	wire [4-1:0] node6036;
	wire [4-1:0] node6037;
	wire [4-1:0] node6041;
	wire [4-1:0] node6042;
	wire [4-1:0] node6045;
	wire [4-1:0] node6046;
	wire [4-1:0] node6048;
	wire [4-1:0] node6052;
	wire [4-1:0] node6053;
	wire [4-1:0] node6054;
	wire [4-1:0] node6055;
	wire [4-1:0] node6057;
	wire [4-1:0] node6058;
	wire [4-1:0] node6062;
	wire [4-1:0] node6065;
	wire [4-1:0] node6066;
	wire [4-1:0] node6067;
	wire [4-1:0] node6068;
	wire [4-1:0] node6073;
	wire [4-1:0] node6075;
	wire [4-1:0] node6076;
	wire [4-1:0] node6079;
	wire [4-1:0] node6082;
	wire [4-1:0] node6083;
	wire [4-1:0] node6084;
	wire [4-1:0] node6086;
	wire [4-1:0] node6088;
	wire [4-1:0] node6092;
	wire [4-1:0] node6094;
	wire [4-1:0] node6095;
	wire [4-1:0] node6099;
	wire [4-1:0] node6100;
	wire [4-1:0] node6101;
	wire [4-1:0] node6102;
	wire [4-1:0] node6103;
	wire [4-1:0] node6105;
	wire [4-1:0] node6107;
	wire [4-1:0] node6110;
	wire [4-1:0] node6113;
	wire [4-1:0] node6114;
	wire [4-1:0] node6118;
	wire [4-1:0] node6119;
	wire [4-1:0] node6120;
	wire [4-1:0] node6122;
	wire [4-1:0] node6125;
	wire [4-1:0] node6128;
	wire [4-1:0] node6129;
	wire [4-1:0] node6130;
	wire [4-1:0] node6133;
	wire [4-1:0] node6136;
	wire [4-1:0] node6137;
	wire [4-1:0] node6138;
	wire [4-1:0] node6143;
	wire [4-1:0] node6144;
	wire [4-1:0] node6145;
	wire [4-1:0] node6146;
	wire [4-1:0] node6147;
	wire [4-1:0] node6148;
	wire [4-1:0] node6153;
	wire [4-1:0] node6154;
	wire [4-1:0] node6155;
	wire [4-1:0] node6159;
	wire [4-1:0] node6162;
	wire [4-1:0] node6163;
	wire [4-1:0] node6165;
	wire [4-1:0] node6166;
	wire [4-1:0] node6170;
	wire [4-1:0] node6172;
	wire [4-1:0] node6175;
	wire [4-1:0] node6176;
	wire [4-1:0] node6177;
	wire [4-1:0] node6179;
	wire [4-1:0] node6180;
	wire [4-1:0] node6183;
	wire [4-1:0] node6186;
	wire [4-1:0] node6187;
	wire [4-1:0] node6191;
	wire [4-1:0] node6192;
	wire [4-1:0] node6193;
	wire [4-1:0] node6196;
	wire [4-1:0] node6197;
	wire [4-1:0] node6200;
	wire [4-1:0] node6204;
	wire [4-1:0] node6205;
	wire [4-1:0] node6206;
	wire [4-1:0] node6207;
	wire [4-1:0] node6208;
	wire [4-1:0] node6210;
	wire [4-1:0] node6213;
	wire [4-1:0] node6215;
	wire [4-1:0] node6218;
	wire [4-1:0] node6219;
	wire [4-1:0] node6222;
	wire [4-1:0] node6223;
	wire [4-1:0] node6225;
	wire [4-1:0] node6226;
	wire [4-1:0] node6230;
	wire [4-1:0] node6231;
	wire [4-1:0] node6232;
	wire [4-1:0] node6235;
	wire [4-1:0] node6239;
	wire [4-1:0] node6240;
	wire [4-1:0] node6241;
	wire [4-1:0] node6242;
	wire [4-1:0] node6243;
	wire [4-1:0] node6247;
	wire [4-1:0] node6249;
	wire [4-1:0] node6250;
	wire [4-1:0] node6253;
	wire [4-1:0] node6256;
	wire [4-1:0] node6257;
	wire [4-1:0] node6259;
	wire [4-1:0] node6260;
	wire [4-1:0] node6263;
	wire [4-1:0] node6266;
	wire [4-1:0] node6267;
	wire [4-1:0] node6268;
	wire [4-1:0] node6271;
	wire [4-1:0] node6275;
	wire [4-1:0] node6276;
	wire [4-1:0] node6277;
	wire [4-1:0] node6279;
	wire [4-1:0] node6281;
	wire [4-1:0] node6285;
	wire [4-1:0] node6287;
	wire [4-1:0] node6289;
	wire [4-1:0] node6292;
	wire [4-1:0] node6293;
	wire [4-1:0] node6294;
	wire [4-1:0] node6295;
	wire [4-1:0] node6297;
	wire [4-1:0] node6299;
	wire [4-1:0] node6302;
	wire [4-1:0] node6303;
	wire [4-1:0] node6304;
	wire [4-1:0] node6306;
	wire [4-1:0] node6310;
	wire [4-1:0] node6311;
	wire [4-1:0] node6313;
	wire [4-1:0] node6317;
	wire [4-1:0] node6318;
	wire [4-1:0] node6320;
	wire [4-1:0] node6321;
	wire [4-1:0] node6323;
	wire [4-1:0] node6327;
	wire [4-1:0] node6328;
	wire [4-1:0] node6329;
	wire [4-1:0] node6332;
	wire [4-1:0] node6333;
	wire [4-1:0] node6337;
	wire [4-1:0] node6340;
	wire [4-1:0] node6341;
	wire [4-1:0] node6342;
	wire [4-1:0] node6343;
	wire [4-1:0] node6346;
	wire [4-1:0] node6349;
	wire [4-1:0] node6350;
	wire [4-1:0] node6353;
	wire [4-1:0] node6354;
	wire [4-1:0] node6357;
	wire [4-1:0] node6358;
	wire [4-1:0] node6361;
	wire [4-1:0] node6364;
	wire [4-1:0] node6365;
	wire [4-1:0] node6366;
	wire [4-1:0] node6367;
	wire [4-1:0] node6368;
	wire [4-1:0] node6373;
	wire [4-1:0] node6375;
	wire [4-1:0] node6378;
	wire [4-1:0] node6379;
	wire [4-1:0] node6383;
	wire [4-1:0] node6384;
	wire [4-1:0] node6385;
	wire [4-1:0] node6386;
	wire [4-1:0] node6387;
	wire [4-1:0] node6388;
	wire [4-1:0] node6389;
	wire [4-1:0] node6390;
	wire [4-1:0] node6393;
	wire [4-1:0] node6395;
	wire [4-1:0] node6398;
	wire [4-1:0] node6400;
	wire [4-1:0] node6403;
	wire [4-1:0] node6404;
	wire [4-1:0] node6405;
	wire [4-1:0] node6408;
	wire [4-1:0] node6411;
	wire [4-1:0] node6412;
	wire [4-1:0] node6415;
	wire [4-1:0] node6418;
	wire [4-1:0] node6419;
	wire [4-1:0] node6421;
	wire [4-1:0] node6423;
	wire [4-1:0] node6424;
	wire [4-1:0] node6428;
	wire [4-1:0] node6429;
	wire [4-1:0] node6430;
	wire [4-1:0] node6431;
	wire [4-1:0] node6432;
	wire [4-1:0] node6437;
	wire [4-1:0] node6438;
	wire [4-1:0] node6441;
	wire [4-1:0] node6443;
	wire [4-1:0] node6446;
	wire [4-1:0] node6447;
	wire [4-1:0] node6449;
	wire [4-1:0] node6450;
	wire [4-1:0] node6454;
	wire [4-1:0] node6456;
	wire [4-1:0] node6459;
	wire [4-1:0] node6460;
	wire [4-1:0] node6461;
	wire [4-1:0] node6462;
	wire [4-1:0] node6465;
	wire [4-1:0] node6466;
	wire [4-1:0] node6469;
	wire [4-1:0] node6472;
	wire [4-1:0] node6473;
	wire [4-1:0] node6474;
	wire [4-1:0] node6475;
	wire [4-1:0] node6476;
	wire [4-1:0] node6481;
	wire [4-1:0] node6484;
	wire [4-1:0] node6485;
	wire [4-1:0] node6486;
	wire [4-1:0] node6488;
	wire [4-1:0] node6491;
	wire [4-1:0] node6495;
	wire [4-1:0] node6496;
	wire [4-1:0] node6497;
	wire [4-1:0] node6498;
	wire [4-1:0] node6500;
	wire [4-1:0] node6502;
	wire [4-1:0] node6505;
	wire [4-1:0] node6507;
	wire [4-1:0] node6508;
	wire [4-1:0] node6512;
	wire [4-1:0] node6514;
	wire [4-1:0] node6515;
	wire [4-1:0] node6519;
	wire [4-1:0] node6520;
	wire [4-1:0] node6521;
	wire [4-1:0] node6522;
	wire [4-1:0] node6524;
	wire [4-1:0] node6528;
	wire [4-1:0] node6529;
	wire [4-1:0] node6533;
	wire [4-1:0] node6534;
	wire [4-1:0] node6535;
	wire [4-1:0] node6538;
	wire [4-1:0] node6541;
	wire [4-1:0] node6542;
	wire [4-1:0] node6543;
	wire [4-1:0] node6548;
	wire [4-1:0] node6549;
	wire [4-1:0] node6550;
	wire [4-1:0] node6551;
	wire [4-1:0] node6552;
	wire [4-1:0] node6555;
	wire [4-1:0] node6557;
	wire [4-1:0] node6559;
	wire [4-1:0] node6561;
	wire [4-1:0] node6564;
	wire [4-1:0] node6565;
	wire [4-1:0] node6566;
	wire [4-1:0] node6567;
	wire [4-1:0] node6570;
	wire [4-1:0] node6573;
	wire [4-1:0] node6574;
	wire [4-1:0] node6577;
	wire [4-1:0] node6580;
	wire [4-1:0] node6581;
	wire [4-1:0] node6582;
	wire [4-1:0] node6585;
	wire [4-1:0] node6587;
	wire [4-1:0] node6591;
	wire [4-1:0] node6592;
	wire [4-1:0] node6593;
	wire [4-1:0] node6595;
	wire [4-1:0] node6596;
	wire [4-1:0] node6597;
	wire [4-1:0] node6601;
	wire [4-1:0] node6604;
	wire [4-1:0] node6605;
	wire [4-1:0] node6607;
	wire [4-1:0] node6609;
	wire [4-1:0] node6612;
	wire [4-1:0] node6614;
	wire [4-1:0] node6617;
	wire [4-1:0] node6618;
	wire [4-1:0] node6619;
	wire [4-1:0] node6620;
	wire [4-1:0] node6625;
	wire [4-1:0] node6626;
	wire [4-1:0] node6629;
	wire [4-1:0] node6630;
	wire [4-1:0] node6631;
	wire [4-1:0] node6636;
	wire [4-1:0] node6637;
	wire [4-1:0] node6638;
	wire [4-1:0] node6639;
	wire [4-1:0] node6640;
	wire [4-1:0] node6642;
	wire [4-1:0] node6644;
	wire [4-1:0] node6647;
	wire [4-1:0] node6650;
	wire [4-1:0] node6651;
	wire [4-1:0] node6652;
	wire [4-1:0] node6654;
	wire [4-1:0] node6659;
	wire [4-1:0] node6660;
	wire [4-1:0] node6661;
	wire [4-1:0] node6662;
	wire [4-1:0] node6667;
	wire [4-1:0] node6668;
	wire [4-1:0] node6672;
	wire [4-1:0] node6673;
	wire [4-1:0] node6674;
	wire [4-1:0] node6675;
	wire [4-1:0] node6679;
	wire [4-1:0] node6681;
	wire [4-1:0] node6683;
	wire [4-1:0] node6685;
	wire [4-1:0] node6688;
	wire [4-1:0] node6689;
	wire [4-1:0] node6691;
	wire [4-1:0] node6694;
	wire [4-1:0] node6696;
	wire [4-1:0] node6698;
	wire [4-1:0] node6701;
	wire [4-1:0] node6702;
	wire [4-1:0] node6703;
	wire [4-1:0] node6704;
	wire [4-1:0] node6705;
	wire [4-1:0] node6707;
	wire [4-1:0] node6709;
	wire [4-1:0] node6712;
	wire [4-1:0] node6713;
	wire [4-1:0] node6715;
	wire [4-1:0] node6716;
	wire [4-1:0] node6717;
	wire [4-1:0] node6721;
	wire [4-1:0] node6722;
	wire [4-1:0] node6726;
	wire [4-1:0] node6728;
	wire [4-1:0] node6730;
	wire [4-1:0] node6731;
	wire [4-1:0] node6735;
	wire [4-1:0] node6736;
	wire [4-1:0] node6737;
	wire [4-1:0] node6738;
	wire [4-1:0] node6739;
	wire [4-1:0] node6743;
	wire [4-1:0] node6744;
	wire [4-1:0] node6745;
	wire [4-1:0] node6750;
	wire [4-1:0] node6751;
	wire [4-1:0] node6752;
	wire [4-1:0] node6753;
	wire [4-1:0] node6758;
	wire [4-1:0] node6760;
	wire [4-1:0] node6761;
	wire [4-1:0] node6765;
	wire [4-1:0] node6766;
	wire [4-1:0] node6768;
	wire [4-1:0] node6771;
	wire [4-1:0] node6772;
	wire [4-1:0] node6776;
	wire [4-1:0] node6777;
	wire [4-1:0] node6778;
	wire [4-1:0] node6779;
	wire [4-1:0] node6780;
	wire [4-1:0] node6781;
	wire [4-1:0] node6785;
	wire [4-1:0] node6788;
	wire [4-1:0] node6789;
	wire [4-1:0] node6792;
	wire [4-1:0] node6794;
	wire [4-1:0] node6796;
	wire [4-1:0] node6799;
	wire [4-1:0] node6800;
	wire [4-1:0] node6801;
	wire [4-1:0] node6804;
	wire [4-1:0] node6805;
	wire [4-1:0] node6807;
	wire [4-1:0] node6811;
	wire [4-1:0] node6812;
	wire [4-1:0] node6813;
	wire [4-1:0] node6817;
	wire [4-1:0] node6820;
	wire [4-1:0] node6821;
	wire [4-1:0] node6822;
	wire [4-1:0] node6823;
	wire [4-1:0] node6825;
	wire [4-1:0] node6828;
	wire [4-1:0] node6829;
	wire [4-1:0] node6830;
	wire [4-1:0] node6835;
	wire [4-1:0] node6837;
	wire [4-1:0] node6838;
	wire [4-1:0] node6839;
	wire [4-1:0] node6844;
	wire [4-1:0] node6845;
	wire [4-1:0] node6846;
	wire [4-1:0] node6848;
	wire [4-1:0] node6849;
	wire [4-1:0] node6854;
	wire [4-1:0] node6855;
	wire [4-1:0] node6856;
	wire [4-1:0] node6860;
	wire [4-1:0] node6861;
	wire [4-1:0] node6863;
	wire [4-1:0] node6866;
	wire [4-1:0] node6867;
	wire [4-1:0] node6871;
	wire [4-1:0] node6872;
	wire [4-1:0] node6873;
	wire [4-1:0] node6874;
	wire [4-1:0] node6875;
	wire [4-1:0] node6876;
	wire [4-1:0] node6878;
	wire [4-1:0] node6881;
	wire [4-1:0] node6883;
	wire [4-1:0] node6886;
	wire [4-1:0] node6888;
	wire [4-1:0] node6891;
	wire [4-1:0] node6892;
	wire [4-1:0] node6893;
	wire [4-1:0] node6896;
	wire [4-1:0] node6897;
	wire [4-1:0] node6901;
	wire [4-1:0] node6902;
	wire [4-1:0] node6903;
	wire [4-1:0] node6906;
	wire [4-1:0] node6907;
	wire [4-1:0] node6912;
	wire [4-1:0] node6913;
	wire [4-1:0] node6914;
	wire [4-1:0] node6916;
	wire [4-1:0] node6917;
	wire [4-1:0] node6918;
	wire [4-1:0] node6922;
	wire [4-1:0] node6923;
	wire [4-1:0] node6926;
	wire [4-1:0] node6929;
	wire [4-1:0] node6930;
	wire [4-1:0] node6931;
	wire [4-1:0] node6932;
	wire [4-1:0] node6937;
	wire [4-1:0] node6938;
	wire [4-1:0] node6939;
	wire [4-1:0] node6943;
	wire [4-1:0] node6946;
	wire [4-1:0] node6947;
	wire [4-1:0] node6948;
	wire [4-1:0] node6951;
	wire [4-1:0] node6954;
	wire [4-1:0] node6955;
	wire [4-1:0] node6956;
	wire [4-1:0] node6957;
	wire [4-1:0] node6963;
	wire [4-1:0] node6964;
	wire [4-1:0] node6965;
	wire [4-1:0] node6966;
	wire [4-1:0] node6967;
	wire [4-1:0] node6970;
	wire [4-1:0] node6971;
	wire [4-1:0] node6973;
	wire [4-1:0] node6976;
	wire [4-1:0] node6979;
	wire [4-1:0] node6982;
	wire [4-1:0] node6983;
	wire [4-1:0] node6984;
	wire [4-1:0] node6985;
	wire [4-1:0] node6986;
	wire [4-1:0] node6990;
	wire [4-1:0] node6991;
	wire [4-1:0] node6994;
	wire [4-1:0] node6997;
	wire [4-1:0] node6998;
	wire [4-1:0] node7000;
	wire [4-1:0] node7004;
	wire [4-1:0] node7005;
	wire [4-1:0] node7007;
	wire [4-1:0] node7010;
	wire [4-1:0] node7012;
	wire [4-1:0] node7015;
	wire [4-1:0] node7016;
	wire [4-1:0] node7017;
	wire [4-1:0] node7020;
	wire [4-1:0] node7022;
	wire [4-1:0] node7023;
	wire [4-1:0] node7026;
	wire [4-1:0] node7029;
	wire [4-1:0] node7030;
	wire [4-1:0] node7031;
	wire [4-1:0] node7032;
	wire [4-1:0] node7034;
	wire [4-1:0] node7038;
	wire [4-1:0] node7040;
	wire [4-1:0] node7043;
	wire [4-1:0] node7044;
	wire [4-1:0] node7047;
	wire [4-1:0] node7048;
	wire [4-1:0] node7052;
	wire [4-1:0] node7053;
	wire [4-1:0] node7054;
	wire [4-1:0] node7055;
	wire [4-1:0] node7056;
	wire [4-1:0] node7057;
	wire [4-1:0] node7058;
	wire [4-1:0] node7059;
	wire [4-1:0] node7060;
	wire [4-1:0] node7062;
	wire [4-1:0] node7065;
	wire [4-1:0] node7068;
	wire [4-1:0] node7069;
	wire [4-1:0] node7070;
	wire [4-1:0] node7075;
	wire [4-1:0] node7076;
	wire [4-1:0] node7077;
	wire [4-1:0] node7080;
	wire [4-1:0] node7083;
	wire [4-1:0] node7084;
	wire [4-1:0] node7087;
	wire [4-1:0] node7090;
	wire [4-1:0] node7091;
	wire [4-1:0] node7092;
	wire [4-1:0] node7093;
	wire [4-1:0] node7095;
	wire [4-1:0] node7098;
	wire [4-1:0] node7101;
	wire [4-1:0] node7102;
	wire [4-1:0] node7105;
	wire [4-1:0] node7107;
	wire [4-1:0] node7108;
	wire [4-1:0] node7111;
	wire [4-1:0] node7114;
	wire [4-1:0] node7115;
	wire [4-1:0] node7116;
	wire [4-1:0] node7117;
	wire [4-1:0] node7119;
	wire [4-1:0] node7123;
	wire [4-1:0] node7126;
	wire [4-1:0] node7128;
	wire [4-1:0] node7130;
	wire [4-1:0] node7133;
	wire [4-1:0] node7134;
	wire [4-1:0] node7135;
	wire [4-1:0] node7136;
	wire [4-1:0] node7138;
	wire [4-1:0] node7141;
	wire [4-1:0] node7142;
	wire [4-1:0] node7143;
	wire [4-1:0] node7145;
	wire [4-1:0] node7148;
	wire [4-1:0] node7151;
	wire [4-1:0] node7152;
	wire [4-1:0] node7156;
	wire [4-1:0] node7157;
	wire [4-1:0] node7159;
	wire [4-1:0] node7160;
	wire [4-1:0] node7162;
	wire [4-1:0] node7166;
	wire [4-1:0] node7167;
	wire [4-1:0] node7168;
	wire [4-1:0] node7172;
	wire [4-1:0] node7173;
	wire [4-1:0] node7177;
	wire [4-1:0] node7178;
	wire [4-1:0] node7179;
	wire [4-1:0] node7181;
	wire [4-1:0] node7184;
	wire [4-1:0] node7186;
	wire [4-1:0] node7189;
	wire [4-1:0] node7190;
	wire [4-1:0] node7191;
	wire [4-1:0] node7193;
	wire [4-1:0] node7195;
	wire [4-1:0] node7198;
	wire [4-1:0] node7201;
	wire [4-1:0] node7203;
	wire [4-1:0] node7205;
	wire [4-1:0] node7207;
	wire [4-1:0] node7210;
	wire [4-1:0] node7211;
	wire [4-1:0] node7212;
	wire [4-1:0] node7213;
	wire [4-1:0] node7214;
	wire [4-1:0] node7215;
	wire [4-1:0] node7216;
	wire [4-1:0] node7220;
	wire [4-1:0] node7223;
	wire [4-1:0] node7224;
	wire [4-1:0] node7227;
	wire [4-1:0] node7230;
	wire [4-1:0] node7231;
	wire [4-1:0] node7234;
	wire [4-1:0] node7235;
	wire [4-1:0] node7237;
	wire [4-1:0] node7241;
	wire [4-1:0] node7242;
	wire [4-1:0] node7243;
	wire [4-1:0] node7244;
	wire [4-1:0] node7246;
	wire [4-1:0] node7248;
	wire [4-1:0] node7251;
	wire [4-1:0] node7254;
	wire [4-1:0] node7255;
	wire [4-1:0] node7257;
	wire [4-1:0] node7260;
	wire [4-1:0] node7262;
	wire [4-1:0] node7265;
	wire [4-1:0] node7266;
	wire [4-1:0] node7267;
	wire [4-1:0] node7268;
	wire [4-1:0] node7269;
	wire [4-1:0] node7275;
	wire [4-1:0] node7276;
	wire [4-1:0] node7277;
	wire [4-1:0] node7278;
	wire [4-1:0] node7283;
	wire [4-1:0] node7284;
	wire [4-1:0] node7285;
	wire [4-1:0] node7288;
	wire [4-1:0] node7292;
	wire [4-1:0] node7293;
	wire [4-1:0] node7294;
	wire [4-1:0] node7295;
	wire [4-1:0] node7296;
	wire [4-1:0] node7297;
	wire [4-1:0] node7302;
	wire [4-1:0] node7303;
	wire [4-1:0] node7304;
	wire [4-1:0] node7309;
	wire [4-1:0] node7310;
	wire [4-1:0] node7311;
	wire [4-1:0] node7312;
	wire [4-1:0] node7317;
	wire [4-1:0] node7318;
	wire [4-1:0] node7319;
	wire [4-1:0] node7323;
	wire [4-1:0] node7324;
	wire [4-1:0] node7325;
	wire [4-1:0] node7330;
	wire [4-1:0] node7331;
	wire [4-1:0] node7332;
	wire [4-1:0] node7334;
	wire [4-1:0] node7335;
	wire [4-1:0] node7336;
	wire [4-1:0] node7341;
	wire [4-1:0] node7342;
	wire [4-1:0] node7345;
	wire [4-1:0] node7347;
	wire [4-1:0] node7348;
	wire [4-1:0] node7352;
	wire [4-1:0] node7353;
	wire [4-1:0] node7354;
	wire [4-1:0] node7355;
	wire [4-1:0] node7359;
	wire [4-1:0] node7361;
	wire [4-1:0] node7364;
	wire [4-1:0] node7365;
	wire [4-1:0] node7367;
	wire [4-1:0] node7368;
	wire [4-1:0] node7371;
	wire [4-1:0] node7375;
	wire [4-1:0] node7376;
	wire [4-1:0] node7377;
	wire [4-1:0] node7378;
	wire [4-1:0] node7379;
	wire [4-1:0] node7380;
	wire [4-1:0] node7381;
	wire [4-1:0] node7383;
	wire [4-1:0] node7385;
	wire [4-1:0] node7389;
	wire [4-1:0] node7392;
	wire [4-1:0] node7393;
	wire [4-1:0] node7394;
	wire [4-1:0] node7396;
	wire [4-1:0] node7399;
	wire [4-1:0] node7400;
	wire [4-1:0] node7401;
	wire [4-1:0] node7406;
	wire [4-1:0] node7407;
	wire [4-1:0] node7409;
	wire [4-1:0] node7412;
	wire [4-1:0] node7414;
	wire [4-1:0] node7415;
	wire [4-1:0] node7419;
	wire [4-1:0] node7420;
	wire [4-1:0] node7421;
	wire [4-1:0] node7422;
	wire [4-1:0] node7425;
	wire [4-1:0] node7428;
	wire [4-1:0] node7431;
	wire [4-1:0] node7432;
	wire [4-1:0] node7433;
	wire [4-1:0] node7436;
	wire [4-1:0] node7438;
	wire [4-1:0] node7441;
	wire [4-1:0] node7442;
	wire [4-1:0] node7446;
	wire [4-1:0] node7447;
	wire [4-1:0] node7448;
	wire [4-1:0] node7449;
	wire [4-1:0] node7450;
	wire [4-1:0] node7453;
	wire [4-1:0] node7456;
	wire [4-1:0] node7458;
	wire [4-1:0] node7460;
	wire [4-1:0] node7461;
	wire [4-1:0] node7465;
	wire [4-1:0] node7466;
	wire [4-1:0] node7468;
	wire [4-1:0] node7469;
	wire [4-1:0] node7472;
	wire [4-1:0] node7474;
	wire [4-1:0] node7477;
	wire [4-1:0] node7479;
	wire [4-1:0] node7481;
	wire [4-1:0] node7484;
	wire [4-1:0] node7485;
	wire [4-1:0] node7486;
	wire [4-1:0] node7487;
	wire [4-1:0] node7490;
	wire [4-1:0] node7493;
	wire [4-1:0] node7494;
	wire [4-1:0] node7497;
	wire [4-1:0] node7498;
	wire [4-1:0] node7502;
	wire [4-1:0] node7503;
	wire [4-1:0] node7504;
	wire [4-1:0] node7505;
	wire [4-1:0] node7509;
	wire [4-1:0] node7511;
	wire [4-1:0] node7512;
	wire [4-1:0] node7516;
	wire [4-1:0] node7517;
	wire [4-1:0] node7518;
	wire [4-1:0] node7519;
	wire [4-1:0] node7524;
	wire [4-1:0] node7525;
	wire [4-1:0] node7529;
	wire [4-1:0] node7530;
	wire [4-1:0] node7531;
	wire [4-1:0] node7532;
	wire [4-1:0] node7533;
	wire [4-1:0] node7534;
	wire [4-1:0] node7536;
	wire [4-1:0] node7539;
	wire [4-1:0] node7542;
	wire [4-1:0] node7543;
	wire [4-1:0] node7544;
	wire [4-1:0] node7548;
	wire [4-1:0] node7549;
	wire [4-1:0] node7550;
	wire [4-1:0] node7555;
	wire [4-1:0] node7556;
	wire [4-1:0] node7557;
	wire [4-1:0] node7558;
	wire [4-1:0] node7560;
	wire [4-1:0] node7565;
	wire [4-1:0] node7566;
	wire [4-1:0] node7568;
	wire [4-1:0] node7570;
	wire [4-1:0] node7574;
	wire [4-1:0] node7575;
	wire [4-1:0] node7576;
	wire [4-1:0] node7578;
	wire [4-1:0] node7579;
	wire [4-1:0] node7580;
	wire [4-1:0] node7584;
	wire [4-1:0] node7587;
	wire [4-1:0] node7588;
	wire [4-1:0] node7589;
	wire [4-1:0] node7590;
	wire [4-1:0] node7596;
	wire [4-1:0] node7598;
	wire [4-1:0] node7599;
	wire [4-1:0] node7602;
	wire [4-1:0] node7603;
	wire [4-1:0] node7604;
	wire [4-1:0] node7607;
	wire [4-1:0] node7611;
	wire [4-1:0] node7612;
	wire [4-1:0] node7613;
	wire [4-1:0] node7614;
	wire [4-1:0] node7615;
	wire [4-1:0] node7618;
	wire [4-1:0] node7619;
	wire [4-1:0] node7623;
	wire [4-1:0] node7624;
	wire [4-1:0] node7625;
	wire [4-1:0] node7627;
	wire [4-1:0] node7632;
	wire [4-1:0] node7633;
	wire [4-1:0] node7634;
	wire [4-1:0] node7636;
	wire [4-1:0] node7640;
	wire [4-1:0] node7641;
	wire [4-1:0] node7643;
	wire [4-1:0] node7646;
	wire [4-1:0] node7647;
	wire [4-1:0] node7648;
	wire [4-1:0] node7653;
	wire [4-1:0] node7654;
	wire [4-1:0] node7655;
	wire [4-1:0] node7656;
	wire [4-1:0] node7659;
	wire [4-1:0] node7662;
	wire [4-1:0] node7663;
	wire [4-1:0] node7664;
	wire [4-1:0] node7668;
	wire [4-1:0] node7669;
	wire [4-1:0] node7671;
	wire [4-1:0] node7675;
	wire [4-1:0] node7676;
	wire [4-1:0] node7678;
	wire [4-1:0] node7679;
	wire [4-1:0] node7680;
	wire [4-1:0] node7684;
	wire [4-1:0] node7686;
	wire [4-1:0] node7689;
	wire [4-1:0] node7691;
	wire [4-1:0] node7694;
	wire [4-1:0] node7695;
	wire [4-1:0] node7696;
	wire [4-1:0] node7697;
	wire [4-1:0] node7698;
	wire [4-1:0] node7699;
	wire [4-1:0] node7700;
	wire [4-1:0] node7701;
	wire [4-1:0] node7704;
	wire [4-1:0] node7705;
	wire [4-1:0] node7709;
	wire [4-1:0] node7711;
	wire [4-1:0] node7714;
	wire [4-1:0] node7715;
	wire [4-1:0] node7716;
	wire [4-1:0] node7718;
	wire [4-1:0] node7721;
	wire [4-1:0] node7722;
	wire [4-1:0] node7726;
	wire [4-1:0] node7727;
	wire [4-1:0] node7730;
	wire [4-1:0] node7733;
	wire [4-1:0] node7734;
	wire [4-1:0] node7735;
	wire [4-1:0] node7736;
	wire [4-1:0] node7737;
	wire [4-1:0] node7742;
	wire [4-1:0] node7743;
	wire [4-1:0] node7746;
	wire [4-1:0] node7747;
	wire [4-1:0] node7750;
	wire [4-1:0] node7753;
	wire [4-1:0] node7754;
	wire [4-1:0] node7755;
	wire [4-1:0] node7757;
	wire [4-1:0] node7761;
	wire [4-1:0] node7762;
	wire [4-1:0] node7764;
	wire [4-1:0] node7767;
	wire [4-1:0] node7768;
	wire [4-1:0] node7770;
	wire [4-1:0] node7773;
	wire [4-1:0] node7774;
	wire [4-1:0] node7777;
	wire [4-1:0] node7780;
	wire [4-1:0] node7781;
	wire [4-1:0] node7782;
	wire [4-1:0] node7783;
	wire [4-1:0] node7785;
	wire [4-1:0] node7788;
	wire [4-1:0] node7790;
	wire [4-1:0] node7793;
	wire [4-1:0] node7794;
	wire [4-1:0] node7795;
	wire [4-1:0] node7797;
	wire [4-1:0] node7800;
	wire [4-1:0] node7802;
	wire [4-1:0] node7803;
	wire [4-1:0] node7807;
	wire [4-1:0] node7808;
	wire [4-1:0] node7812;
	wire [4-1:0] node7813;
	wire [4-1:0] node7814;
	wire [4-1:0] node7815;
	wire [4-1:0] node7816;
	wire [4-1:0] node7818;
	wire [4-1:0] node7822;
	wire [4-1:0] node7823;
	wire [4-1:0] node7826;
	wire [4-1:0] node7829;
	wire [4-1:0] node7830;
	wire [4-1:0] node7834;
	wire [4-1:0] node7835;
	wire [4-1:0] node7837;
	wire [4-1:0] node7839;
	wire [4-1:0] node7842;
	wire [4-1:0] node7844;
	wire [4-1:0] node7847;
	wire [4-1:0] node7848;
	wire [4-1:0] node7849;
	wire [4-1:0] node7850;
	wire [4-1:0] node7851;
	wire [4-1:0] node7852;
	wire [4-1:0] node7853;
	wire [4-1:0] node7854;
	wire [4-1:0] node7860;
	wire [4-1:0] node7862;
	wire [4-1:0] node7863;
	wire [4-1:0] node7867;
	wire [4-1:0] node7869;
	wire [4-1:0] node7870;
	wire [4-1:0] node7871;
	wire [4-1:0] node7875;
	wire [4-1:0] node7876;
	wire [4-1:0] node7879;
	wire [4-1:0] node7882;
	wire [4-1:0] node7883;
	wire [4-1:0] node7884;
	wire [4-1:0] node7885;
	wire [4-1:0] node7887;
	wire [4-1:0] node7890;
	wire [4-1:0] node7891;
	wire [4-1:0] node7895;
	wire [4-1:0] node7896;
	wire [4-1:0] node7897;
	wire [4-1:0] node7900;
	wire [4-1:0] node7903;
	wire [4-1:0] node7906;
	wire [4-1:0] node7907;
	wire [4-1:0] node7910;
	wire [4-1:0] node7911;
	wire [4-1:0] node7912;
	wire [4-1:0] node7913;
	wire [4-1:0] node7918;
	wire [4-1:0] node7921;
	wire [4-1:0] node7922;
	wire [4-1:0] node7923;
	wire [4-1:0] node7924;
	wire [4-1:0] node7925;
	wire [4-1:0] node7926;
	wire [4-1:0] node7928;
	wire [4-1:0] node7932;
	wire [4-1:0] node7935;
	wire [4-1:0] node7937;
	wire [4-1:0] node7939;
	wire [4-1:0] node7942;
	wire [4-1:0] node7943;
	wire [4-1:0] node7944;
	wire [4-1:0] node7945;
	wire [4-1:0] node7948;
	wire [4-1:0] node7949;
	wire [4-1:0] node7953;
	wire [4-1:0] node7954;
	wire [4-1:0] node7958;
	wire [4-1:0] node7959;
	wire [4-1:0] node7962;
	wire [4-1:0] node7964;
	wire [4-1:0] node7967;
	wire [4-1:0] node7968;
	wire [4-1:0] node7969;
	wire [4-1:0] node7970;
	wire [4-1:0] node7972;
	wire [4-1:0] node7974;
	wire [4-1:0] node7977;
	wire [4-1:0] node7978;
	wire [4-1:0] node7979;
	wire [4-1:0] node7983;
	wire [4-1:0] node7985;
	wire [4-1:0] node7988;
	wire [4-1:0] node7990;
	wire [4-1:0] node7991;
	wire [4-1:0] node7993;
	wire [4-1:0] node7996;
	wire [4-1:0] node7999;
	wire [4-1:0] node8000;
	wire [4-1:0] node8001;
	wire [4-1:0] node8004;
	wire [4-1:0] node8005;
	wire [4-1:0] node8009;
	wire [4-1:0] node8010;
	wire [4-1:0] node8013;
	wire [4-1:0] node8014;
	wire [4-1:0] node8017;
	wire [4-1:0] node8020;
	wire [4-1:0] node8021;
	wire [4-1:0] node8022;
	wire [4-1:0] node8023;
	wire [4-1:0] node8024;
	wire [4-1:0] node8025;
	wire [4-1:0] node8027;
	wire [4-1:0] node8029;
	wire [4-1:0] node8032;
	wire [4-1:0] node8033;
	wire [4-1:0] node8036;
	wire [4-1:0] node8037;
	wire [4-1:0] node8041;
	wire [4-1:0] node8042;
	wire [4-1:0] node8043;
	wire [4-1:0] node8044;
	wire [4-1:0] node8045;
	wire [4-1:0] node8049;
	wire [4-1:0] node8052;
	wire [4-1:0] node8055;
	wire [4-1:0] node8056;
	wire [4-1:0] node8057;
	wire [4-1:0] node8062;
	wire [4-1:0] node8063;
	wire [4-1:0] node8064;
	wire [4-1:0] node8065;
	wire [4-1:0] node8066;
	wire [4-1:0] node8067;
	wire [4-1:0] node8071;
	wire [4-1:0] node8072;
	wire [4-1:0] node8075;
	wire [4-1:0] node8079;
	wire [4-1:0] node8080;
	wire [4-1:0] node8084;
	wire [4-1:0] node8085;
	wire [4-1:0] node8086;
	wire [4-1:0] node8087;
	wire [4-1:0] node8090;
	wire [4-1:0] node8093;
	wire [4-1:0] node8094;
	wire [4-1:0] node8099;
	wire [4-1:0] node8100;
	wire [4-1:0] node8101;
	wire [4-1:0] node8102;
	wire [4-1:0] node8103;
	wire [4-1:0] node8104;
	wire [4-1:0] node8105;
	wire [4-1:0] node8110;
	wire [4-1:0] node8111;
	wire [4-1:0] node8113;
	wire [4-1:0] node8117;
	wire [4-1:0] node8118;
	wire [4-1:0] node8119;
	wire [4-1:0] node8122;
	wire [4-1:0] node8123;
	wire [4-1:0] node8127;
	wire [4-1:0] node8128;
	wire [4-1:0] node8131;
	wire [4-1:0] node8134;
	wire [4-1:0] node8136;
	wire [4-1:0] node8137;
	wire [4-1:0] node8140;
	wire [4-1:0] node8141;
	wire [4-1:0] node8144;
	wire [4-1:0] node8145;
	wire [4-1:0] node8149;
	wire [4-1:0] node8150;
	wire [4-1:0] node8151;
	wire [4-1:0] node8152;
	wire [4-1:0] node8154;
	wire [4-1:0] node8157;
	wire [4-1:0] node8158;
	wire [4-1:0] node8162;
	wire [4-1:0] node8163;
	wire [4-1:0] node8166;
	wire [4-1:0] node8168;
	wire [4-1:0] node8171;
	wire [4-1:0] node8172;
	wire [4-1:0] node8173;
	wire [4-1:0] node8175;
	wire [4-1:0] node8176;
	wire [4-1:0] node8180;
	wire [4-1:0] node8181;
	wire [4-1:0] node8184;
	wire [4-1:0] node8187;
	wire [4-1:0] node8188;
	wire [4-1:0] node8189;
	wire [4-1:0] node8191;
	wire [4-1:0] node8195;
	wire [4-1:0] node8197;
	wire [4-1:0] node8199;
	wire [4-1:0] node8202;
	wire [4-1:0] node8203;
	wire [4-1:0] node8204;
	wire [4-1:0] node8205;
	wire [4-1:0] node8206;
	wire [4-1:0] node8207;
	wire [4-1:0] node8208;
	wire [4-1:0] node8209;
	wire [4-1:0] node8214;
	wire [4-1:0] node8216;
	wire [4-1:0] node8218;
	wire [4-1:0] node8221;
	wire [4-1:0] node8222;
	wire [4-1:0] node8223;
	wire [4-1:0] node8224;
	wire [4-1:0] node8228;
	wire [4-1:0] node8229;
	wire [4-1:0] node8232;
	wire [4-1:0] node8236;
	wire [4-1:0] node8237;
	wire [4-1:0] node8238;
	wire [4-1:0] node8239;
	wire [4-1:0] node8240;
	wire [4-1:0] node8243;
	wire [4-1:0] node8247;
	wire [4-1:0] node8248;
	wire [4-1:0] node8252;
	wire [4-1:0] node8253;
	wire [4-1:0] node8255;
	wire [4-1:0] node8259;
	wire [4-1:0] node8260;
	wire [4-1:0] node8261;
	wire [4-1:0] node8262;
	wire [4-1:0] node8265;
	wire [4-1:0] node8267;
	wire [4-1:0] node8270;
	wire [4-1:0] node8272;
	wire [4-1:0] node8274;
	wire [4-1:0] node8275;
	wire [4-1:0] node8279;
	wire [4-1:0] node8280;
	wire [4-1:0] node8281;
	wire [4-1:0] node8282;
	wire [4-1:0] node8286;
	wire [4-1:0] node8287;
	wire [4-1:0] node8291;
	wire [4-1:0] node8292;
	wire [4-1:0] node8296;
	wire [4-1:0] node8297;
	wire [4-1:0] node8298;
	wire [4-1:0] node8299;
	wire [4-1:0] node8302;
	wire [4-1:0] node8303;
	wire [4-1:0] node8304;
	wire [4-1:0] node8305;
	wire [4-1:0] node8308;
	wire [4-1:0] node8312;
	wire [4-1:0] node8314;
	wire [4-1:0] node8315;
	wire [4-1:0] node8319;
	wire [4-1:0] node8320;
	wire [4-1:0] node8321;
	wire [4-1:0] node8322;
	wire [4-1:0] node8323;
	wire [4-1:0] node8326;
	wire [4-1:0] node8331;
	wire [4-1:0] node8332;
	wire [4-1:0] node8336;
	wire [4-1:0] node8337;
	wire [4-1:0] node8338;
	wire [4-1:0] node8340;
	wire [4-1:0] node8343;
	wire [4-1:0] node8344;
	wire [4-1:0] node8346;
	wire [4-1:0] node8347;
	wire [4-1:0] node8350;
	wire [4-1:0] node8354;
	wire [4-1:0] node8355;
	wire [4-1:0] node8356;
	wire [4-1:0] node8357;
	wire [4-1:0] node8361;
	wire [4-1:0] node8362;
	wire [4-1:0] node8365;
	wire [4-1:0] node8368;
	wire [4-1:0] node8369;
	wire [4-1:0] node8370;
	wire [4-1:0] node8372;
	wire [4-1:0] node8375;
	wire [4-1:0] node8378;
	wire [4-1:0] node8381;
	wire [4-1:0] node8382;
	wire [4-1:0] node8383;
	wire [4-1:0] node8384;
	wire [4-1:0] node8385;
	wire [4-1:0] node8386;
	wire [4-1:0] node8387;
	wire [4-1:0] node8388;
	wire [4-1:0] node8389;
	wire [4-1:0] node8390;
	wire [4-1:0] node8393;
	wire [4-1:0] node8394;
	wire [4-1:0] node8395;
	wire [4-1:0] node8398;
	wire [4-1:0] node8401;
	wire [4-1:0] node8404;
	wire [4-1:0] node8405;
	wire [4-1:0] node8406;
	wire [4-1:0] node8410;
	wire [4-1:0] node8413;
	wire [4-1:0] node8414;
	wire [4-1:0] node8415;
	wire [4-1:0] node8416;
	wire [4-1:0] node8419;
	wire [4-1:0] node8421;
	wire [4-1:0] node8424;
	wire [4-1:0] node8427;
	wire [4-1:0] node8428;
	wire [4-1:0] node8430;
	wire [4-1:0] node8431;
	wire [4-1:0] node8435;
	wire [4-1:0] node8437;
	wire [4-1:0] node8440;
	wire [4-1:0] node8441;
	wire [4-1:0] node8442;
	wire [4-1:0] node8443;
	wire [4-1:0] node8445;
	wire [4-1:0] node8446;
	wire [4-1:0] node8449;
	wire [4-1:0] node8452;
	wire [4-1:0] node8454;
	wire [4-1:0] node8456;
	wire [4-1:0] node8459;
	wire [4-1:0] node8460;
	wire [4-1:0] node8463;
	wire [4-1:0] node8464;
	wire [4-1:0] node8468;
	wire [4-1:0] node8469;
	wire [4-1:0] node8470;
	wire [4-1:0] node8473;
	wire [4-1:0] node8474;
	wire [4-1:0] node8476;
	wire [4-1:0] node8480;
	wire [4-1:0] node8482;
	wire [4-1:0] node8484;
	wire [4-1:0] node8486;
	wire [4-1:0] node8489;
	wire [4-1:0] node8490;
	wire [4-1:0] node8491;
	wire [4-1:0] node8492;
	wire [4-1:0] node8493;
	wire [4-1:0] node8494;
	wire [4-1:0] node8496;
	wire [4-1:0] node8499;
	wire [4-1:0] node8500;
	wire [4-1:0] node8505;
	wire [4-1:0] node8507;
	wire [4-1:0] node8510;
	wire [4-1:0] node8511;
	wire [4-1:0] node8512;
	wire [4-1:0] node8513;
	wire [4-1:0] node8514;
	wire [4-1:0] node8518;
	wire [4-1:0] node8521;
	wire [4-1:0] node8523;
	wire [4-1:0] node8524;
	wire [4-1:0] node8528;
	wire [4-1:0] node8530;
	wire [4-1:0] node8533;
	wire [4-1:0] node8534;
	wire [4-1:0] node8535;
	wire [4-1:0] node8536;
	wire [4-1:0] node8538;
	wire [4-1:0] node8540;
	wire [4-1:0] node8543;
	wire [4-1:0] node8545;
	wire [4-1:0] node8548;
	wire [4-1:0] node8549;
	wire [4-1:0] node8550;
	wire [4-1:0] node8551;
	wire [4-1:0] node8555;
	wire [4-1:0] node8558;
	wire [4-1:0] node8561;
	wire [4-1:0] node8562;
	wire [4-1:0] node8563;
	wire [4-1:0] node8565;
	wire [4-1:0] node8569;
	wire [4-1:0] node8570;
	wire [4-1:0] node8572;
	wire [4-1:0] node8573;
	wire [4-1:0] node8577;
	wire [4-1:0] node8579;
	wire [4-1:0] node8580;
	wire [4-1:0] node8584;
	wire [4-1:0] node8585;
	wire [4-1:0] node8586;
	wire [4-1:0] node8587;
	wire [4-1:0] node8588;
	wire [4-1:0] node8589;
	wire [4-1:0] node8590;
	wire [4-1:0] node8594;
	wire [4-1:0] node8597;
	wire [4-1:0] node8598;
	wire [4-1:0] node8599;
	wire [4-1:0] node8602;
	wire [4-1:0] node8604;
	wire [4-1:0] node8607;
	wire [4-1:0] node8609;
	wire [4-1:0] node8612;
	wire [4-1:0] node8613;
	wire [4-1:0] node8614;
	wire [4-1:0] node8615;
	wire [4-1:0] node8617;
	wire [4-1:0] node8621;
	wire [4-1:0] node8624;
	wire [4-1:0] node8626;
	wire [4-1:0] node8628;
	wire [4-1:0] node8629;
	wire [4-1:0] node8633;
	wire [4-1:0] node8634;
	wire [4-1:0] node8635;
	wire [4-1:0] node8638;
	wire [4-1:0] node8639;
	wire [4-1:0] node8640;
	wire [4-1:0] node8645;
	wire [4-1:0] node8646;
	wire [4-1:0] node8647;
	wire [4-1:0] node8650;
	wire [4-1:0] node8652;
	wire [4-1:0] node8653;
	wire [4-1:0] node8656;
	wire [4-1:0] node8659;
	wire [4-1:0] node8660;
	wire [4-1:0] node8664;
	wire [4-1:0] node8665;
	wire [4-1:0] node8666;
	wire [4-1:0] node8667;
	wire [4-1:0] node8668;
	wire [4-1:0] node8669;
	wire [4-1:0] node8670;
	wire [4-1:0] node8675;
	wire [4-1:0] node8677;
	wire [4-1:0] node8680;
	wire [4-1:0] node8681;
	wire [4-1:0] node8682;
	wire [4-1:0] node8685;
	wire [4-1:0] node8688;
	wire [4-1:0] node8689;
	wire [4-1:0] node8692;
	wire [4-1:0] node8695;
	wire [4-1:0] node8696;
	wire [4-1:0] node8698;
	wire [4-1:0] node8701;
	wire [4-1:0] node8702;
	wire [4-1:0] node8703;
	wire [4-1:0] node8704;
	wire [4-1:0] node8709;
	wire [4-1:0] node8710;
	wire [4-1:0] node8712;
	wire [4-1:0] node8716;
	wire [4-1:0] node8717;
	wire [4-1:0] node8718;
	wire [4-1:0] node8719;
	wire [4-1:0] node8720;
	wire [4-1:0] node8723;
	wire [4-1:0] node8725;
	wire [4-1:0] node8728;
	wire [4-1:0] node8731;
	wire [4-1:0] node8732;
	wire [4-1:0] node8733;
	wire [4-1:0] node8735;
	wire [4-1:0] node8738;
	wire [4-1:0] node8741;
	wire [4-1:0] node8743;
	wire [4-1:0] node8746;
	wire [4-1:0] node8747;
	wire [4-1:0] node8748;
	wire [4-1:0] node8751;
	wire [4-1:0] node8753;
	wire [4-1:0] node8755;
	wire [4-1:0] node8758;
	wire [4-1:0] node8759;
	wire [4-1:0] node8762;
	wire [4-1:0] node8763;
	wire [4-1:0] node8764;
	wire [4-1:0] node8767;
	wire [4-1:0] node8770;
	wire [4-1:0] node8772;
	wire [4-1:0] node8775;
	wire [4-1:0] node8776;
	wire [4-1:0] node8777;
	wire [4-1:0] node8778;
	wire [4-1:0] node8779;
	wire [4-1:0] node8780;
	wire [4-1:0] node8781;
	wire [4-1:0] node8782;
	wire [4-1:0] node8787;
	wire [4-1:0] node8788;
	wire [4-1:0] node8790;
	wire [4-1:0] node8793;
	wire [4-1:0] node8794;
	wire [4-1:0] node8797;
	wire [4-1:0] node8800;
	wire [4-1:0] node8801;
	wire [4-1:0] node8802;
	wire [4-1:0] node8804;
	wire [4-1:0] node8808;
	wire [4-1:0] node8810;
	wire [4-1:0] node8813;
	wire [4-1:0] node8814;
	wire [4-1:0] node8815;
	wire [4-1:0] node8816;
	wire [4-1:0] node8818;
	wire [4-1:0] node8819;
	wire [4-1:0] node8823;
	wire [4-1:0] node8824;
	wire [4-1:0] node8827;
	wire [4-1:0] node8830;
	wire [4-1:0] node8831;
	wire [4-1:0] node8834;
	wire [4-1:0] node8837;
	wire [4-1:0] node8838;
	wire [4-1:0] node8839;
	wire [4-1:0] node8840;
	wire [4-1:0] node8844;
	wire [4-1:0] node8847;
	wire [4-1:0] node8848;
	wire [4-1:0] node8849;
	wire [4-1:0] node8853;
	wire [4-1:0] node8856;
	wire [4-1:0] node8857;
	wire [4-1:0] node8858;
	wire [4-1:0] node8859;
	wire [4-1:0] node8860;
	wire [4-1:0] node8861;
	wire [4-1:0] node8862;
	wire [4-1:0] node8867;
	wire [4-1:0] node8868;
	wire [4-1:0] node8872;
	wire [4-1:0] node8874;
	wire [4-1:0] node8875;
	wire [4-1:0] node8878;
	wire [4-1:0] node8879;
	wire [4-1:0] node8883;
	wire [4-1:0] node8884;
	wire [4-1:0] node8885;
	wire [4-1:0] node8886;
	wire [4-1:0] node8887;
	wire [4-1:0] node8893;
	wire [4-1:0] node8894;
	wire [4-1:0] node8895;
	wire [4-1:0] node8898;
	wire [4-1:0] node8901;
	wire [4-1:0] node8902;
	wire [4-1:0] node8903;
	wire [4-1:0] node8908;
	wire [4-1:0] node8909;
	wire [4-1:0] node8910;
	wire [4-1:0] node8911;
	wire [4-1:0] node8913;
	wire [4-1:0] node8916;
	wire [4-1:0] node8918;
	wire [4-1:0] node8921;
	wire [4-1:0] node8923;
	wire [4-1:0] node8926;
	wire [4-1:0] node8927;
	wire [4-1:0] node8928;
	wire [4-1:0] node8929;
	wire [4-1:0] node8930;
	wire [4-1:0] node8934;
	wire [4-1:0] node8935;
	wire [4-1:0] node8939;
	wire [4-1:0] node8940;
	wire [4-1:0] node8941;
	wire [4-1:0] node8944;
	wire [4-1:0] node8948;
	wire [4-1:0] node8950;
	wire [4-1:0] node8952;
	wire [4-1:0] node8953;
	wire [4-1:0] node8957;
	wire [4-1:0] node8958;
	wire [4-1:0] node8959;
	wire [4-1:0] node8960;
	wire [4-1:0] node8961;
	wire [4-1:0] node8962;
	wire [4-1:0] node8963;
	wire [4-1:0] node8964;
	wire [4-1:0] node8970;
	wire [4-1:0] node8971;
	wire [4-1:0] node8973;
	wire [4-1:0] node8976;
	wire [4-1:0] node8979;
	wire [4-1:0] node8980;
	wire [4-1:0] node8981;
	wire [4-1:0] node8984;
	wire [4-1:0] node8987;
	wire [4-1:0] node8989;
	wire [4-1:0] node8991;
	wire [4-1:0] node8992;
	wire [4-1:0] node8996;
	wire [4-1:0] node8997;
	wire [4-1:0] node8998;
	wire [4-1:0] node8999;
	wire [4-1:0] node9001;
	wire [4-1:0] node9004;
	wire [4-1:0] node9007;
	wire [4-1:0] node9008;
	wire [4-1:0] node9010;
	wire [4-1:0] node9011;
	wire [4-1:0] node9015;
	wire [4-1:0] node9017;
	wire [4-1:0] node9018;
	wire [4-1:0] node9022;
	wire [4-1:0] node9023;
	wire [4-1:0] node9024;
	wire [4-1:0] node9025;
	wire [4-1:0] node9028;
	wire [4-1:0] node9031;
	wire [4-1:0] node9032;
	wire [4-1:0] node9036;
	wire [4-1:0] node9039;
	wire [4-1:0] node9040;
	wire [4-1:0] node9041;
	wire [4-1:0] node9042;
	wire [4-1:0] node9043;
	wire [4-1:0] node9044;
	wire [4-1:0] node9045;
	wire [4-1:0] node9048;
	wire [4-1:0] node9051;
	wire [4-1:0] node9054;
	wire [4-1:0] node9055;
	wire [4-1:0] node9059;
	wire [4-1:0] node9060;
	wire [4-1:0] node9062;
	wire [4-1:0] node9064;
	wire [4-1:0] node9067;
	wire [4-1:0] node9069;
	wire [4-1:0] node9071;
	wire [4-1:0] node9074;
	wire [4-1:0] node9075;
	wire [4-1:0] node9077;
	wire [4-1:0] node9079;
	wire [4-1:0] node9081;
	wire [4-1:0] node9084;
	wire [4-1:0] node9086;
	wire [4-1:0] node9088;
	wire [4-1:0] node9090;
	wire [4-1:0] node9093;
	wire [4-1:0] node9094;
	wire [4-1:0] node9095;
	wire [4-1:0] node9096;
	wire [4-1:0] node9098;
	wire [4-1:0] node9102;
	wire [4-1:0] node9103;
	wire [4-1:0] node9105;
	wire [4-1:0] node9106;
	wire [4-1:0] node9110;
	wire [4-1:0] node9111;
	wire [4-1:0] node9113;
	wire [4-1:0] node9116;
	wire [4-1:0] node9117;
	wire [4-1:0] node9121;
	wire [4-1:0] node9122;
	wire [4-1:0] node9124;
	wire [4-1:0] node9126;
	wire [4-1:0] node9129;
	wire [4-1:0] node9130;
	wire [4-1:0] node9132;
	wire [4-1:0] node9133;
	wire [4-1:0] node9138;
	wire [4-1:0] node9139;
	wire [4-1:0] node9140;
	wire [4-1:0] node9141;
	wire [4-1:0] node9142;
	wire [4-1:0] node9143;
	wire [4-1:0] node9144;
	wire [4-1:0] node9145;
	wire [4-1:0] node9147;
	wire [4-1:0] node9151;
	wire [4-1:0] node9153;
	wire [4-1:0] node9154;
	wire [4-1:0] node9157;
	wire [4-1:0] node9160;
	wire [4-1:0] node9161;
	wire [4-1:0] node9164;
	wire [4-1:0] node9165;
	wire [4-1:0] node9167;
	wire [4-1:0] node9171;
	wire [4-1:0] node9172;
	wire [4-1:0] node9173;
	wire [4-1:0] node9174;
	wire [4-1:0] node9177;
	wire [4-1:0] node9180;
	wire [4-1:0] node9181;
	wire [4-1:0] node9182;
	wire [4-1:0] node9183;
	wire [4-1:0] node9186;
	wire [4-1:0] node9189;
	wire [4-1:0] node9190;
	wire [4-1:0] node9194;
	wire [4-1:0] node9196;
	wire [4-1:0] node9198;
	wire [4-1:0] node9201;
	wire [4-1:0] node9202;
	wire [4-1:0] node9203;
	wire [4-1:0] node9205;
	wire [4-1:0] node9206;
	wire [4-1:0] node9211;
	wire [4-1:0] node9213;
	wire [4-1:0] node9216;
	wire [4-1:0] node9217;
	wire [4-1:0] node9218;
	wire [4-1:0] node9219;
	wire [4-1:0] node9220;
	wire [4-1:0] node9223;
	wire [4-1:0] node9224;
	wire [4-1:0] node9228;
	wire [4-1:0] node9229;
	wire [4-1:0] node9230;
	wire [4-1:0] node9234;
	wire [4-1:0] node9235;
	wire [4-1:0] node9239;
	wire [4-1:0] node9240;
	wire [4-1:0] node9241;
	wire [4-1:0] node9243;
	wire [4-1:0] node9245;
	wire [4-1:0] node9248;
	wire [4-1:0] node9251;
	wire [4-1:0] node9252;
	wire [4-1:0] node9253;
	wire [4-1:0] node9257;
	wire [4-1:0] node9258;
	wire [4-1:0] node9261;
	wire [4-1:0] node9262;
	wire [4-1:0] node9266;
	wire [4-1:0] node9267;
	wire [4-1:0] node9268;
	wire [4-1:0] node9270;
	wire [4-1:0] node9273;
	wire [4-1:0] node9275;
	wire [4-1:0] node9276;
	wire [4-1:0] node9277;
	wire [4-1:0] node9282;
	wire [4-1:0] node9283;
	wire [4-1:0] node9284;
	wire [4-1:0] node9285;
	wire [4-1:0] node9289;
	wire [4-1:0] node9291;
	wire [4-1:0] node9293;
	wire [4-1:0] node9296;
	wire [4-1:0] node9297;
	wire [4-1:0] node9298;
	wire [4-1:0] node9299;
	wire [4-1:0] node9302;
	wire [4-1:0] node9307;
	wire [4-1:0] node9308;
	wire [4-1:0] node9309;
	wire [4-1:0] node9310;
	wire [4-1:0] node9311;
	wire [4-1:0] node9312;
	wire [4-1:0] node9314;
	wire [4-1:0] node9316;
	wire [4-1:0] node9319;
	wire [4-1:0] node9322;
	wire [4-1:0] node9324;
	wire [4-1:0] node9327;
	wire [4-1:0] node9328;
	wire [4-1:0] node9330;
	wire [4-1:0] node9331;
	wire [4-1:0] node9332;
	wire [4-1:0] node9335;
	wire [4-1:0] node9339;
	wire [4-1:0] node9341;
	wire [4-1:0] node9343;
	wire [4-1:0] node9346;
	wire [4-1:0] node9347;
	wire [4-1:0] node9348;
	wire [4-1:0] node9349;
	wire [4-1:0] node9350;
	wire [4-1:0] node9351;
	wire [4-1:0] node9357;
	wire [4-1:0] node9359;
	wire [4-1:0] node9360;
	wire [4-1:0] node9364;
	wire [4-1:0] node9365;
	wire [4-1:0] node9366;
	wire [4-1:0] node9367;
	wire [4-1:0] node9368;
	wire [4-1:0] node9372;
	wire [4-1:0] node9373;
	wire [4-1:0] node9377;
	wire [4-1:0] node9380;
	wire [4-1:0] node9381;
	wire [4-1:0] node9382;
	wire [4-1:0] node9387;
	wire [4-1:0] node9388;
	wire [4-1:0] node9389;
	wire [4-1:0] node9390;
	wire [4-1:0] node9391;
	wire [4-1:0] node9392;
	wire [4-1:0] node9393;
	wire [4-1:0] node9398;
	wire [4-1:0] node9401;
	wire [4-1:0] node9402;
	wire [4-1:0] node9403;
	wire [4-1:0] node9405;
	wire [4-1:0] node9408;
	wire [4-1:0] node9411;
	wire [4-1:0] node9413;
	wire [4-1:0] node9416;
	wire [4-1:0] node9417;
	wire [4-1:0] node9418;
	wire [4-1:0] node9422;
	wire [4-1:0] node9423;
	wire [4-1:0] node9424;
	wire [4-1:0] node9426;
	wire [4-1:0] node9431;
	wire [4-1:0] node9432;
	wire [4-1:0] node9433;
	wire [4-1:0] node9434;
	wire [4-1:0] node9437;
	wire [4-1:0] node9438;
	wire [4-1:0] node9440;
	wire [4-1:0] node9444;
	wire [4-1:0] node9445;
	wire [4-1:0] node9446;
	wire [4-1:0] node9450;
	wire [4-1:0] node9451;
	wire [4-1:0] node9452;
	wire [4-1:0] node9455;
	wire [4-1:0] node9459;
	wire [4-1:0] node9460;
	wire [4-1:0] node9461;
	wire [4-1:0] node9462;
	wire [4-1:0] node9463;
	wire [4-1:0] node9467;
	wire [4-1:0] node9468;
	wire [4-1:0] node9472;
	wire [4-1:0] node9475;
	wire [4-1:0] node9476;
	wire [4-1:0] node9480;
	wire [4-1:0] node9481;
	wire [4-1:0] node9482;
	wire [4-1:0] node9483;
	wire [4-1:0] node9484;
	wire [4-1:0] node9485;
	wire [4-1:0] node9486;
	wire [4-1:0] node9487;
	wire [4-1:0] node9491;
	wire [4-1:0] node9494;
	wire [4-1:0] node9495;
	wire [4-1:0] node9497;
	wire [4-1:0] node9501;
	wire [4-1:0] node9502;
	wire [4-1:0] node9503;
	wire [4-1:0] node9504;
	wire [4-1:0] node9507;
	wire [4-1:0] node9508;
	wire [4-1:0] node9513;
	wire [4-1:0] node9514;
	wire [4-1:0] node9515;
	wire [4-1:0] node9518;
	wire [4-1:0] node9521;
	wire [4-1:0] node9522;
	wire [4-1:0] node9525;
	wire [4-1:0] node9528;
	wire [4-1:0] node9529;
	wire [4-1:0] node9530;
	wire [4-1:0] node9531;
	wire [4-1:0] node9534;
	wire [4-1:0] node9536;
	wire [4-1:0] node9539;
	wire [4-1:0] node9540;
	wire [4-1:0] node9542;
	wire [4-1:0] node9544;
	wire [4-1:0] node9548;
	wire [4-1:0] node9549;
	wire [4-1:0] node9550;
	wire [4-1:0] node9552;
	wire [4-1:0] node9555;
	wire [4-1:0] node9557;
	wire [4-1:0] node9559;
	wire [4-1:0] node9562;
	wire [4-1:0] node9563;
	wire [4-1:0] node9564;
	wire [4-1:0] node9565;
	wire [4-1:0] node9570;
	wire [4-1:0] node9571;
	wire [4-1:0] node9575;
	wire [4-1:0] node9576;
	wire [4-1:0] node9577;
	wire [4-1:0] node9578;
	wire [4-1:0] node9579;
	wire [4-1:0] node9581;
	wire [4-1:0] node9582;
	wire [4-1:0] node9586;
	wire [4-1:0] node9587;
	wire [4-1:0] node9590;
	wire [4-1:0] node9593;
	wire [4-1:0] node9594;
	wire [4-1:0] node9596;
	wire [4-1:0] node9598;
	wire [4-1:0] node9601;
	wire [4-1:0] node9602;
	wire [4-1:0] node9605;
	wire [4-1:0] node9608;
	wire [4-1:0] node9609;
	wire [4-1:0] node9610;
	wire [4-1:0] node9613;
	wire [4-1:0] node9616;
	wire [4-1:0] node9618;
	wire [4-1:0] node9619;
	wire [4-1:0] node9620;
	wire [4-1:0] node9625;
	wire [4-1:0] node9626;
	wire [4-1:0] node9627;
	wire [4-1:0] node9628;
	wire [4-1:0] node9631;
	wire [4-1:0] node9634;
	wire [4-1:0] node9635;
	wire [4-1:0] node9637;
	wire [4-1:0] node9640;
	wire [4-1:0] node9642;
	wire [4-1:0] node9645;
	wire [4-1:0] node9646;
	wire [4-1:0] node9647;
	wire [4-1:0] node9649;
	wire [4-1:0] node9652;
	wire [4-1:0] node9655;
	wire [4-1:0] node9656;
	wire [4-1:0] node9658;
	wire [4-1:0] node9661;
	wire [4-1:0] node9662;
	wire [4-1:0] node9663;
	wire [4-1:0] node9668;
	wire [4-1:0] node9669;
	wire [4-1:0] node9670;
	wire [4-1:0] node9671;
	wire [4-1:0] node9672;
	wire [4-1:0] node9673;
	wire [4-1:0] node9674;
	wire [4-1:0] node9675;
	wire [4-1:0] node9679;
	wire [4-1:0] node9680;
	wire [4-1:0] node9684;
	wire [4-1:0] node9686;
	wire [4-1:0] node9689;
	wire [4-1:0] node9691;
	wire [4-1:0] node9692;
	wire [4-1:0] node9693;
	wire [4-1:0] node9698;
	wire [4-1:0] node9699;
	wire [4-1:0] node9700;
	wire [4-1:0] node9701;
	wire [4-1:0] node9703;
	wire [4-1:0] node9707;
	wire [4-1:0] node9709;
	wire [4-1:0] node9712;
	wire [4-1:0] node9713;
	wire [4-1:0] node9714;
	wire [4-1:0] node9715;
	wire [4-1:0] node9719;
	wire [4-1:0] node9721;
	wire [4-1:0] node9725;
	wire [4-1:0] node9726;
	wire [4-1:0] node9727;
	wire [4-1:0] node9729;
	wire [4-1:0] node9732;
	wire [4-1:0] node9735;
	wire [4-1:0] node9736;
	wire [4-1:0] node9737;
	wire [4-1:0] node9741;
	wire [4-1:0] node9742;
	wire [4-1:0] node9746;
	wire [4-1:0] node9747;
	wire [4-1:0] node9748;
	wire [4-1:0] node9749;
	wire [4-1:0] node9750;
	wire [4-1:0] node9751;
	wire [4-1:0] node9753;
	wire [4-1:0] node9757;
	wire [4-1:0] node9760;
	wire [4-1:0] node9762;
	wire [4-1:0] node9763;
	wire [4-1:0] node9767;
	wire [4-1:0] node9768;
	wire [4-1:0] node9769;
	wire [4-1:0] node9773;
	wire [4-1:0] node9774;
	wire [4-1:0] node9777;
	wire [4-1:0] node9779;
	wire [4-1:0] node9782;
	wire [4-1:0] node9783;
	wire [4-1:0] node9784;
	wire [4-1:0] node9786;
	wire [4-1:0] node9787;
	wire [4-1:0] node9788;
	wire [4-1:0] node9793;
	wire [4-1:0] node9794;
	wire [4-1:0] node9796;
	wire [4-1:0] node9797;
	wire [4-1:0] node9801;
	wire [4-1:0] node9803;
	wire [4-1:0] node9806;
	wire [4-1:0] node9807;
	wire [4-1:0] node9808;
	wire [4-1:0] node9809;
	wire [4-1:0] node9810;
	wire [4-1:0] node9813;
	wire [4-1:0] node9817;
	wire [4-1:0] node9819;
	wire [4-1:0] node9822;
	wire [4-1:0] node9823;
	wire [4-1:0] node9825;
	wire [4-1:0] node9827;
	wire [4-1:0] node9830;
	wire [4-1:0] node9831;
	wire [4-1:0] node9832;
	wire [4-1:0] node9837;
	wire [4-1:0] node9838;
	wire [4-1:0] node9839;
	wire [4-1:0] node9840;
	wire [4-1:0] node9841;
	wire [4-1:0] node9842;
	wire [4-1:0] node9843;
	wire [4-1:0] node9844;
	wire [4-1:0] node9845;
	wire [4-1:0] node9849;
	wire [4-1:0] node9850;
	wire [4-1:0] node9851;
	wire [4-1:0] node9854;
	wire [4-1:0] node9855;
	wire [4-1:0] node9860;
	wire [4-1:0] node9861;
	wire [4-1:0] node9862;
	wire [4-1:0] node9863;
	wire [4-1:0] node9866;
	wire [4-1:0] node9869;
	wire [4-1:0] node9870;
	wire [4-1:0] node9871;
	wire [4-1:0] node9875;
	wire [4-1:0] node9878;
	wire [4-1:0] node9879;
	wire [4-1:0] node9880;
	wire [4-1:0] node9884;
	wire [4-1:0] node9885;
	wire [4-1:0] node9888;
	wire [4-1:0] node9891;
	wire [4-1:0] node9892;
	wire [4-1:0] node9893;
	wire [4-1:0] node9894;
	wire [4-1:0] node9895;
	wire [4-1:0] node9898;
	wire [4-1:0] node9899;
	wire [4-1:0] node9903;
	wire [4-1:0] node9904;
	wire [4-1:0] node9908;
	wire [4-1:0] node9910;
	wire [4-1:0] node9911;
	wire [4-1:0] node9915;
	wire [4-1:0] node9916;
	wire [4-1:0] node9917;
	wire [4-1:0] node9920;
	wire [4-1:0] node9921;
	wire [4-1:0] node9925;
	wire [4-1:0] node9927;
	wire [4-1:0] node9929;
	wire [4-1:0] node9932;
	wire [4-1:0] node9933;
	wire [4-1:0] node9934;
	wire [4-1:0] node9935;
	wire [4-1:0] node9936;
	wire [4-1:0] node9937;
	wire [4-1:0] node9938;
	wire [4-1:0] node9944;
	wire [4-1:0] node9946;
	wire [4-1:0] node9947;
	wire [4-1:0] node9950;
	wire [4-1:0] node9953;
	wire [4-1:0] node9954;
	wire [4-1:0] node9955;
	wire [4-1:0] node9959;
	wire [4-1:0] node9960;
	wire [4-1:0] node9961;
	wire [4-1:0] node9966;
	wire [4-1:0] node9967;
	wire [4-1:0] node9968;
	wire [4-1:0] node9969;
	wire [4-1:0] node9970;
	wire [4-1:0] node9974;
	wire [4-1:0] node9976;
	wire [4-1:0] node9979;
	wire [4-1:0] node9980;
	wire [4-1:0] node9982;
	wire [4-1:0] node9986;
	wire [4-1:0] node9987;
	wire [4-1:0] node9988;
	wire [4-1:0] node9989;
	wire [4-1:0] node9993;
	wire [4-1:0] node9995;
	wire [4-1:0] node9998;
	wire [4-1:0] node9999;
	wire [4-1:0] node10003;
	wire [4-1:0] node10004;
	wire [4-1:0] node10005;
	wire [4-1:0] node10006;
	wire [4-1:0] node10007;
	wire [4-1:0] node10008;
	wire [4-1:0] node10009;
	wire [4-1:0] node10015;
	wire [4-1:0] node10016;
	wire [4-1:0] node10017;
	wire [4-1:0] node10019;
	wire [4-1:0] node10022;
	wire [4-1:0] node10023;
	wire [4-1:0] node10027;
	wire [4-1:0] node10029;
	wire [4-1:0] node10030;
	wire [4-1:0] node10031;
	wire [4-1:0] node10036;
	wire [4-1:0] node10037;
	wire [4-1:0] node10038;
	wire [4-1:0] node10039;
	wire [4-1:0] node10041;
	wire [4-1:0] node10043;
	wire [4-1:0] node10047;
	wire [4-1:0] node10048;
	wire [4-1:0] node10052;
	wire [4-1:0] node10053;
	wire [4-1:0] node10054;
	wire [4-1:0] node10057;
	wire [4-1:0] node10060;
	wire [4-1:0] node10061;
	wire [4-1:0] node10062;
	wire [4-1:0] node10066;
	wire [4-1:0] node10067;
	wire [4-1:0] node10071;
	wire [4-1:0] node10072;
	wire [4-1:0] node10073;
	wire [4-1:0] node10074;
	wire [4-1:0] node10075;
	wire [4-1:0] node10076;
	wire [4-1:0] node10080;
	wire [4-1:0] node10082;
	wire [4-1:0] node10083;
	wire [4-1:0] node10087;
	wire [4-1:0] node10089;
	wire [4-1:0] node10091;
	wire [4-1:0] node10092;
	wire [4-1:0] node10096;
	wire [4-1:0] node10097;
	wire [4-1:0] node10098;
	wire [4-1:0] node10101;
	wire [4-1:0] node10104;
	wire [4-1:0] node10105;
	wire [4-1:0] node10106;
	wire [4-1:0] node10108;
	wire [4-1:0] node10112;
	wire [4-1:0] node10114;
	wire [4-1:0] node10117;
	wire [4-1:0] node10118;
	wire [4-1:0] node10119;
	wire [4-1:0] node10120;
	wire [4-1:0] node10123;
	wire [4-1:0] node10126;
	wire [4-1:0] node10127;
	wire [4-1:0] node10130;
	wire [4-1:0] node10133;
	wire [4-1:0] node10134;
	wire [4-1:0] node10136;
	wire [4-1:0] node10139;
	wire [4-1:0] node10140;
	wire [4-1:0] node10141;
	wire [4-1:0] node10143;
	wire [4-1:0] node10147;
	wire [4-1:0] node10149;
	wire [4-1:0] node10150;
	wire [4-1:0] node10154;
	wire [4-1:0] node10155;
	wire [4-1:0] node10156;
	wire [4-1:0] node10157;
	wire [4-1:0] node10158;
	wire [4-1:0] node10159;
	wire [4-1:0] node10160;
	wire [4-1:0] node10163;
	wire [4-1:0] node10166;
	wire [4-1:0] node10167;
	wire [4-1:0] node10168;
	wire [4-1:0] node10173;
	wire [4-1:0] node10174;
	wire [4-1:0] node10175;
	wire [4-1:0] node10178;
	wire [4-1:0] node10180;
	wire [4-1:0] node10183;
	wire [4-1:0] node10184;
	wire [4-1:0] node10187;
	wire [4-1:0] node10188;
	wire [4-1:0] node10192;
	wire [4-1:0] node10193;
	wire [4-1:0] node10194;
	wire [4-1:0] node10195;
	wire [4-1:0] node10196;
	wire [4-1:0] node10201;
	wire [4-1:0] node10203;
	wire [4-1:0] node10205;
	wire [4-1:0] node10207;
	wire [4-1:0] node10210;
	wire [4-1:0] node10211;
	wire [4-1:0] node10213;
	wire [4-1:0] node10214;
	wire [4-1:0] node10215;
	wire [4-1:0] node10220;
	wire [4-1:0] node10221;
	wire [4-1:0] node10224;
	wire [4-1:0] node10225;
	wire [4-1:0] node10226;
	wire [4-1:0] node10231;
	wire [4-1:0] node10232;
	wire [4-1:0] node10233;
	wire [4-1:0] node10234;
	wire [4-1:0] node10235;
	wire [4-1:0] node10237;
	wire [4-1:0] node10238;
	wire [4-1:0] node10242;
	wire [4-1:0] node10244;
	wire [4-1:0] node10247;
	wire [4-1:0] node10248;
	wire [4-1:0] node10249;
	wire [4-1:0] node10251;
	wire [4-1:0] node10254;
	wire [4-1:0] node10256;
	wire [4-1:0] node10259;
	wire [4-1:0] node10262;
	wire [4-1:0] node10263;
	wire [4-1:0] node10265;
	wire [4-1:0] node10266;
	wire [4-1:0] node10270;
	wire [4-1:0] node10271;
	wire [4-1:0] node10272;
	wire [4-1:0] node10276;
	wire [4-1:0] node10277;
	wire [4-1:0] node10281;
	wire [4-1:0] node10282;
	wire [4-1:0] node10283;
	wire [4-1:0] node10286;
	wire [4-1:0] node10287;
	wire [4-1:0] node10288;
	wire [4-1:0] node10291;
	wire [4-1:0] node10294;
	wire [4-1:0] node10295;
	wire [4-1:0] node10299;
	wire [4-1:0] node10300;
	wire [4-1:0] node10302;
	wire [4-1:0] node10303;
	wire [4-1:0] node10306;
	wire [4-1:0] node10309;
	wire [4-1:0] node10310;
	wire [4-1:0] node10311;
	wire [4-1:0] node10316;
	wire [4-1:0] node10317;
	wire [4-1:0] node10318;
	wire [4-1:0] node10319;
	wire [4-1:0] node10320;
	wire [4-1:0] node10322;
	wire [4-1:0] node10325;
	wire [4-1:0] node10326;
	wire [4-1:0] node10327;
	wire [4-1:0] node10328;
	wire [4-1:0] node10331;
	wire [4-1:0] node10335;
	wire [4-1:0] node10337;
	wire [4-1:0] node10340;
	wire [4-1:0] node10341;
	wire [4-1:0] node10342;
	wire [4-1:0] node10344;
	wire [4-1:0] node10348;
	wire [4-1:0] node10349;
	wire [4-1:0] node10351;
	wire [4-1:0] node10354;
	wire [4-1:0] node10356;
	wire [4-1:0] node10359;
	wire [4-1:0] node10360;
	wire [4-1:0] node10361;
	wire [4-1:0] node10362;
	wire [4-1:0] node10364;
	wire [4-1:0] node10368;
	wire [4-1:0] node10369;
	wire [4-1:0] node10371;
	wire [4-1:0] node10373;
	wire [4-1:0] node10376;
	wire [4-1:0] node10377;
	wire [4-1:0] node10378;
	wire [4-1:0] node10383;
	wire [4-1:0] node10384;
	wire [4-1:0] node10385;
	wire [4-1:0] node10388;
	wire [4-1:0] node10391;
	wire [4-1:0] node10393;
	wire [4-1:0] node10396;
	wire [4-1:0] node10397;
	wire [4-1:0] node10398;
	wire [4-1:0] node10399;
	wire [4-1:0] node10400;
	wire [4-1:0] node10402;
	wire [4-1:0] node10405;
	wire [4-1:0] node10407;
	wire [4-1:0] node10408;
	wire [4-1:0] node10412;
	wire [4-1:0] node10413;
	wire [4-1:0] node10415;
	wire [4-1:0] node10417;
	wire [4-1:0] node10420;
	wire [4-1:0] node10421;
	wire [4-1:0] node10425;
	wire [4-1:0] node10426;
	wire [4-1:0] node10427;
	wire [4-1:0] node10428;
	wire [4-1:0] node10429;
	wire [4-1:0] node10432;
	wire [4-1:0] node10436;
	wire [4-1:0] node10438;
	wire [4-1:0] node10441;
	wire [4-1:0] node10442;
	wire [4-1:0] node10443;
	wire [4-1:0] node10444;
	wire [4-1:0] node10450;
	wire [4-1:0] node10451;
	wire [4-1:0] node10452;
	wire [4-1:0] node10453;
	wire [4-1:0] node10454;
	wire [4-1:0] node10455;
	wire [4-1:0] node10461;
	wire [4-1:0] node10463;
	wire [4-1:0] node10464;
	wire [4-1:0] node10466;
	wire [4-1:0] node10469;
	wire [4-1:0] node10472;
	wire [4-1:0] node10473;
	wire [4-1:0] node10474;
	wire [4-1:0] node10475;
	wire [4-1:0] node10476;
	wire [4-1:0] node10481;
	wire [4-1:0] node10484;
	wire [4-1:0] node10486;
	wire [4-1:0] node10488;
	wire [4-1:0] node10490;
	wire [4-1:0] node10493;
	wire [4-1:0] node10494;
	wire [4-1:0] node10495;
	wire [4-1:0] node10496;
	wire [4-1:0] node10497;
	wire [4-1:0] node10498;
	wire [4-1:0] node10499;
	wire [4-1:0] node10500;
	wire [4-1:0] node10501;
	wire [4-1:0] node10503;
	wire [4-1:0] node10507;
	wire [4-1:0] node10509;
	wire [4-1:0] node10512;
	wire [4-1:0] node10513;
	wire [4-1:0] node10516;
	wire [4-1:0] node10519;
	wire [4-1:0] node10520;
	wire [4-1:0] node10522;
	wire [4-1:0] node10523;
	wire [4-1:0] node10526;
	wire [4-1:0] node10528;
	wire [4-1:0] node10531;
	wire [4-1:0] node10532;
	wire [4-1:0] node10536;
	wire [4-1:0] node10537;
	wire [4-1:0] node10538;
	wire [4-1:0] node10539;
	wire [4-1:0] node10542;
	wire [4-1:0] node10543;
	wire [4-1:0] node10546;
	wire [4-1:0] node10549;
	wire [4-1:0] node10550;
	wire [4-1:0] node10551;
	wire [4-1:0] node10553;
	wire [4-1:0] node10557;
	wire [4-1:0] node10559;
	wire [4-1:0] node10560;
	wire [4-1:0] node10564;
	wire [4-1:0] node10565;
	wire [4-1:0] node10566;
	wire [4-1:0] node10567;
	wire [4-1:0] node10568;
	wire [4-1:0] node10571;
	wire [4-1:0] node10574;
	wire [4-1:0] node10577;
	wire [4-1:0] node10580;
	wire [4-1:0] node10581;
	wire [4-1:0] node10584;
	wire [4-1:0] node10585;
	wire [4-1:0] node10587;
	wire [4-1:0] node10591;
	wire [4-1:0] node10592;
	wire [4-1:0] node10593;
	wire [4-1:0] node10594;
	wire [4-1:0] node10595;
	wire [4-1:0] node10596;
	wire [4-1:0] node10600;
	wire [4-1:0] node10603;
	wire [4-1:0] node10605;
	wire [4-1:0] node10607;
	wire [4-1:0] node10609;
	wire [4-1:0] node10612;
	wire [4-1:0] node10613;
	wire [4-1:0] node10615;
	wire [4-1:0] node10616;
	wire [4-1:0] node10617;
	wire [4-1:0] node10621;
	wire [4-1:0] node10623;
	wire [4-1:0] node10626;
	wire [4-1:0] node10628;
	wire [4-1:0] node10631;
	wire [4-1:0] node10632;
	wire [4-1:0] node10633;
	wire [4-1:0] node10634;
	wire [4-1:0] node10636;
	wire [4-1:0] node10637;
	wire [4-1:0] node10642;
	wire [4-1:0] node10644;
	wire [4-1:0] node10646;
	wire [4-1:0] node10648;
	wire [4-1:0] node10651;
	wire [4-1:0] node10652;
	wire [4-1:0] node10653;
	wire [4-1:0] node10656;
	wire [4-1:0] node10657;
	wire [4-1:0] node10660;
	wire [4-1:0] node10661;
	wire [4-1:0] node10664;
	wire [4-1:0] node10667;
	wire [4-1:0] node10668;
	wire [4-1:0] node10671;
	wire [4-1:0] node10673;
	wire [4-1:0] node10675;
	wire [4-1:0] node10678;
	wire [4-1:0] node10679;
	wire [4-1:0] node10680;
	wire [4-1:0] node10681;
	wire [4-1:0] node10682;
	wire [4-1:0] node10683;
	wire [4-1:0] node10687;
	wire [4-1:0] node10689;
	wire [4-1:0] node10691;
	wire [4-1:0] node10692;
	wire [4-1:0] node10696;
	wire [4-1:0] node10697;
	wire [4-1:0] node10698;
	wire [4-1:0] node10699;
	wire [4-1:0] node10701;
	wire [4-1:0] node10705;
	wire [4-1:0] node10706;
	wire [4-1:0] node10710;
	wire [4-1:0] node10711;
	wire [4-1:0] node10712;
	wire [4-1:0] node10716;
	wire [4-1:0] node10718;
	wire [4-1:0] node10719;
	wire [4-1:0] node10723;
	wire [4-1:0] node10724;
	wire [4-1:0] node10725;
	wire [4-1:0] node10726;
	wire [4-1:0] node10727;
	wire [4-1:0] node10728;
	wire [4-1:0] node10732;
	wire [4-1:0] node10736;
	wire [4-1:0] node10737;
	wire [4-1:0] node10738;
	wire [4-1:0] node10742;
	wire [4-1:0] node10743;
	wire [4-1:0] node10747;
	wire [4-1:0] node10748;
	wire [4-1:0] node10749;
	wire [4-1:0] node10752;
	wire [4-1:0] node10754;
	wire [4-1:0] node10755;
	wire [4-1:0] node10759;
	wire [4-1:0] node10761;
	wire [4-1:0] node10762;
	wire [4-1:0] node10766;
	wire [4-1:0] node10767;
	wire [4-1:0] node10768;
	wire [4-1:0] node10769;
	wire [4-1:0] node10770;
	wire [4-1:0] node10772;
	wire [4-1:0] node10773;
	wire [4-1:0] node10777;
	wire [4-1:0] node10780;
	wire [4-1:0] node10781;
	wire [4-1:0] node10783;
	wire [4-1:0] node10787;
	wire [4-1:0] node10788;
	wire [4-1:0] node10789;
	wire [4-1:0] node10791;
	wire [4-1:0] node10794;
	wire [4-1:0] node10797;
	wire [4-1:0] node10798;
	wire [4-1:0] node10799;
	wire [4-1:0] node10800;
	wire [4-1:0] node10803;
	wire [4-1:0] node10807;
	wire [4-1:0] node10808;
	wire [4-1:0] node10811;
	wire [4-1:0] node10814;
	wire [4-1:0] node10815;
	wire [4-1:0] node10816;
	wire [4-1:0] node10817;
	wire [4-1:0] node10819;
	wire [4-1:0] node10820;
	wire [4-1:0] node10825;
	wire [4-1:0] node10826;
	wire [4-1:0] node10829;
	wire [4-1:0] node10832;
	wire [4-1:0] node10833;
	wire [4-1:0] node10834;
	wire [4-1:0] node10836;
	wire [4-1:0] node10839;
	wire [4-1:0] node10840;
	wire [4-1:0] node10844;
	wire [4-1:0] node10845;
	wire [4-1:0] node10846;
	wire [4-1:0] node10847;
	wire [4-1:0] node10852;
	wire [4-1:0] node10853;
	wire [4-1:0] node10855;
	wire [4-1:0] node10859;
	wire [4-1:0] node10860;
	wire [4-1:0] node10861;
	wire [4-1:0] node10862;
	wire [4-1:0] node10863;
	wire [4-1:0] node10864;
	wire [4-1:0] node10865;
	wire [4-1:0] node10867;
	wire [4-1:0] node10870;
	wire [4-1:0] node10871;
	wire [4-1:0] node10873;
	wire [4-1:0] node10876;
	wire [4-1:0] node10879;
	wire [4-1:0] node10880;
	wire [4-1:0] node10883;
	wire [4-1:0] node10886;
	wire [4-1:0] node10887;
	wire [4-1:0] node10889;
	wire [4-1:0] node10892;
	wire [4-1:0] node10893;
	wire [4-1:0] node10896;
	wire [4-1:0] node10898;
	wire [4-1:0] node10901;
	wire [4-1:0] node10902;
	wire [4-1:0] node10903;
	wire [4-1:0] node10904;
	wire [4-1:0] node10905;
	wire [4-1:0] node10910;
	wire [4-1:0] node10913;
	wire [4-1:0] node10914;
	wire [4-1:0] node10916;
	wire [4-1:0] node10917;
	wire [4-1:0] node10920;
	wire [4-1:0] node10921;
	wire [4-1:0] node10925;
	wire [4-1:0] node10926;
	wire [4-1:0] node10929;
	wire [4-1:0] node10930;
	wire [4-1:0] node10931;
	wire [4-1:0] node10935;
	wire [4-1:0] node10937;
	wire [4-1:0] node10940;
	wire [4-1:0] node10941;
	wire [4-1:0] node10942;
	wire [4-1:0] node10943;
	wire [4-1:0] node10944;
	wire [4-1:0] node10945;
	wire [4-1:0] node10947;
	wire [4-1:0] node10950;
	wire [4-1:0] node10952;
	wire [4-1:0] node10955;
	wire [4-1:0] node10958;
	wire [4-1:0] node10959;
	wire [4-1:0] node10963;
	wire [4-1:0] node10964;
	wire [4-1:0] node10965;
	wire [4-1:0] node10967;
	wire [4-1:0] node10968;
	wire [4-1:0] node10972;
	wire [4-1:0] node10973;
	wire [4-1:0] node10975;
	wire [4-1:0] node10979;
	wire [4-1:0] node10980;
	wire [4-1:0] node10981;
	wire [4-1:0] node10984;
	wire [4-1:0] node10987;
	wire [4-1:0] node10988;
	wire [4-1:0] node10992;
	wire [4-1:0] node10993;
	wire [4-1:0] node10994;
	wire [4-1:0] node10995;
	wire [4-1:0] node10996;
	wire [4-1:0] node11000;
	wire [4-1:0] node11002;
	wire [4-1:0] node11005;
	wire [4-1:0] node11006;
	wire [4-1:0] node11008;
	wire [4-1:0] node11009;
	wire [4-1:0] node11013;
	wire [4-1:0] node11015;
	wire [4-1:0] node11018;
	wire [4-1:0] node11019;
	wire [4-1:0] node11020;
	wire [4-1:0] node11021;
	wire [4-1:0] node11025;
	wire [4-1:0] node11028;
	wire [4-1:0] node11029;
	wire [4-1:0] node11030;
	wire [4-1:0] node11034;
	wire [4-1:0] node11037;
	wire [4-1:0] node11038;
	wire [4-1:0] node11039;
	wire [4-1:0] node11040;
	wire [4-1:0] node11041;
	wire [4-1:0] node11042;
	wire [4-1:0] node11043;
	wire [4-1:0] node11045;
	wire [4-1:0] node11049;
	wire [4-1:0] node11051;
	wire [4-1:0] node11054;
	wire [4-1:0] node11055;
	wire [4-1:0] node11056;
	wire [4-1:0] node11060;
	wire [4-1:0] node11061;
	wire [4-1:0] node11064;
	wire [4-1:0] node11066;
	wire [4-1:0] node11069;
	wire [4-1:0] node11070;
	wire [4-1:0] node11071;
	wire [4-1:0] node11072;
	wire [4-1:0] node11075;
	wire [4-1:0] node11078;
	wire [4-1:0] node11079;
	wire [4-1:0] node11081;
	wire [4-1:0] node11085;
	wire [4-1:0] node11086;
	wire [4-1:0] node11089;
	wire [4-1:0] node11090;
	wire [4-1:0] node11091;
	wire [4-1:0] node11096;
	wire [4-1:0] node11097;
	wire [4-1:0] node11098;
	wire [4-1:0] node11099;
	wire [4-1:0] node11100;
	wire [4-1:0] node11101;
	wire [4-1:0] node11106;
	wire [4-1:0] node11109;
	wire [4-1:0] node11110;
	wire [4-1:0] node11111;
	wire [4-1:0] node11114;
	wire [4-1:0] node11117;
	wire [4-1:0] node11118;
	wire [4-1:0] node11120;
	wire [4-1:0] node11123;
	wire [4-1:0] node11125;
	wire [4-1:0] node11128;
	wire [4-1:0] node11129;
	wire [4-1:0] node11130;
	wire [4-1:0] node11131;
	wire [4-1:0] node11132;
	wire [4-1:0] node11138;
	wire [4-1:0] node11139;
	wire [4-1:0] node11143;
	wire [4-1:0] node11144;
	wire [4-1:0] node11145;
	wire [4-1:0] node11146;
	wire [4-1:0] node11147;
	wire [4-1:0] node11148;
	wire [4-1:0] node11151;
	wire [4-1:0] node11152;
	wire [4-1:0] node11155;
	wire [4-1:0] node11158;
	wire [4-1:0] node11160;
	wire [4-1:0] node11163;
	wire [4-1:0] node11165;
	wire [4-1:0] node11166;
	wire [4-1:0] node11169;
	wire [4-1:0] node11172;
	wire [4-1:0] node11173;
	wire [4-1:0] node11174;
	wire [4-1:0] node11175;
	wire [4-1:0] node11177;
	wire [4-1:0] node11180;
	wire [4-1:0] node11182;
	wire [4-1:0] node11185;
	wire [4-1:0] node11187;
	wire [4-1:0] node11190;
	wire [4-1:0] node11191;
	wire [4-1:0] node11192;
	wire [4-1:0] node11196;
	wire [4-1:0] node11199;
	wire [4-1:0] node11200;
	wire [4-1:0] node11201;
	wire [4-1:0] node11202;
	wire [4-1:0] node11204;
	wire [4-1:0] node11205;
	wire [4-1:0] node11209;
	wire [4-1:0] node11210;
	wire [4-1:0] node11213;
	wire [4-1:0] node11214;
	wire [4-1:0] node11218;
	wire [4-1:0] node11219;
	wire [4-1:0] node11220;
	wire [4-1:0] node11221;
	wire [4-1:0] node11224;
	wire [4-1:0] node11228;
	wire [4-1:0] node11229;
	wire [4-1:0] node11233;
	wire [4-1:0] node11234;
	wire [4-1:0] node11235;
	wire [4-1:0] node11238;
	wire [4-1:0] node11240;
	wire [4-1:0] node11243;
	wire [4-1:0] node11244;
	wire [4-1:0] node11245;
	wire [4-1:0] node11247;
	wire [4-1:0] node11250;
	wire [4-1:0] node11254;
	wire [4-1:0] node11255;
	wire [4-1:0] node11256;
	wire [4-1:0] node11257;
	wire [4-1:0] node11258;
	wire [4-1:0] node11259;
	wire [4-1:0] node11260;
	wire [4-1:0] node11261;
	wire [4-1:0] node11262;
	wire [4-1:0] node11263;
	wire [4-1:0] node11264;
	wire [4-1:0] node11265;
	wire [4-1:0] node11267;
	wire [4-1:0] node11270;
	wire [4-1:0] node11271;
	wire [4-1:0] node11275;
	wire [4-1:0] node11276;
	wire [4-1:0] node11277;
	wire [4-1:0] node11278;
	wire [4-1:0] node11282;
	wire [4-1:0] node11285;
	wire [4-1:0] node11286;
	wire [4-1:0] node11287;
	wire [4-1:0] node11290;
	wire [4-1:0] node11293;
	wire [4-1:0] node11296;
	wire [4-1:0] node11297;
	wire [4-1:0] node11298;
	wire [4-1:0] node11301;
	wire [4-1:0] node11304;
	wire [4-1:0] node11306;
	wire [4-1:0] node11307;
	wire [4-1:0] node11310;
	wire [4-1:0] node11311;
	wire [4-1:0] node11315;
	wire [4-1:0] node11316;
	wire [4-1:0] node11317;
	wire [4-1:0] node11319;
	wire [4-1:0] node11320;
	wire [4-1:0] node11324;
	wire [4-1:0] node11325;
	wire [4-1:0] node11326;
	wire [4-1:0] node11331;
	wire [4-1:0] node11332;
	wire [4-1:0] node11333;
	wire [4-1:0] node11335;
	wire [4-1:0] node11339;
	wire [4-1:0] node11340;
	wire [4-1:0] node11341;
	wire [4-1:0] node11344;
	wire [4-1:0] node11347;
	wire [4-1:0] node11350;
	wire [4-1:0] node11351;
	wire [4-1:0] node11352;
	wire [4-1:0] node11353;
	wire [4-1:0] node11355;
	wire [4-1:0] node11356;
	wire [4-1:0] node11359;
	wire [4-1:0] node11362;
	wire [4-1:0] node11363;
	wire [4-1:0] node11364;
	wire [4-1:0] node11368;
	wire [4-1:0] node11369;
	wire [4-1:0] node11372;
	wire [4-1:0] node11374;
	wire [4-1:0] node11377;
	wire [4-1:0] node11378;
	wire [4-1:0] node11379;
	wire [4-1:0] node11381;
	wire [4-1:0] node11384;
	wire [4-1:0] node11387;
	wire [4-1:0] node11388;
	wire [4-1:0] node11389;
	wire [4-1:0] node11393;
	wire [4-1:0] node11396;
	wire [4-1:0] node11397;
	wire [4-1:0] node11398;
	wire [4-1:0] node11399;
	wire [4-1:0] node11401;
	wire [4-1:0] node11405;
	wire [4-1:0] node11406;
	wire [4-1:0] node11407;
	wire [4-1:0] node11411;
	wire [4-1:0] node11414;
	wire [4-1:0] node11415;
	wire [4-1:0] node11416;
	wire [4-1:0] node11417;
	wire [4-1:0] node11420;
	wire [4-1:0] node11423;
	wire [4-1:0] node11426;
	wire [4-1:0] node11428;
	wire [4-1:0] node11429;
	wire [4-1:0] node11433;
	wire [4-1:0] node11434;
	wire [4-1:0] node11435;
	wire [4-1:0] node11436;
	wire [4-1:0] node11437;
	wire [4-1:0] node11438;
	wire [4-1:0] node11440;
	wire [4-1:0] node11443;
	wire [4-1:0] node11446;
	wire [4-1:0] node11448;
	wire [4-1:0] node11449;
	wire [4-1:0] node11453;
	wire [4-1:0] node11454;
	wire [4-1:0] node11456;
	wire [4-1:0] node11459;
	wire [4-1:0] node11460;
	wire [4-1:0] node11462;
	wire [4-1:0] node11465;
	wire [4-1:0] node11466;
	wire [4-1:0] node11467;
	wire [4-1:0] node11471;
	wire [4-1:0] node11472;
	wire [4-1:0] node11476;
	wire [4-1:0] node11477;
	wire [4-1:0] node11478;
	wire [4-1:0] node11479;
	wire [4-1:0] node11482;
	wire [4-1:0] node11483;
	wire [4-1:0] node11484;
	wire [4-1:0] node11487;
	wire [4-1:0] node11490;
	wire [4-1:0] node11491;
	wire [4-1:0] node11495;
	wire [4-1:0] node11497;
	wire [4-1:0] node11499;
	wire [4-1:0] node11501;
	wire [4-1:0] node11504;
	wire [4-1:0] node11505;
	wire [4-1:0] node11506;
	wire [4-1:0] node11509;
	wire [4-1:0] node11512;
	wire [4-1:0] node11513;
	wire [4-1:0] node11515;
	wire [4-1:0] node11519;
	wire [4-1:0] node11520;
	wire [4-1:0] node11521;
	wire [4-1:0] node11522;
	wire [4-1:0] node11524;
	wire [4-1:0] node11527;
	wire [4-1:0] node11528;
	wire [4-1:0] node11531;
	wire [4-1:0] node11534;
	wire [4-1:0] node11535;
	wire [4-1:0] node11536;
	wire [4-1:0] node11537;
	wire [4-1:0] node11541;
	wire [4-1:0] node11542;
	wire [4-1:0] node11544;
	wire [4-1:0] node11548;
	wire [4-1:0] node11550;
	wire [4-1:0] node11553;
	wire [4-1:0] node11554;
	wire [4-1:0] node11556;
	wire [4-1:0] node11557;
	wire [4-1:0] node11558;
	wire [4-1:0] node11563;
	wire [4-1:0] node11564;
	wire [4-1:0] node11566;
	wire [4-1:0] node11568;
	wire [4-1:0] node11571;
	wire [4-1:0] node11572;
	wire [4-1:0] node11575;
	wire [4-1:0] node11578;
	wire [4-1:0] node11579;
	wire [4-1:0] node11580;
	wire [4-1:0] node11581;
	wire [4-1:0] node11582;
	wire [4-1:0] node11583;
	wire [4-1:0] node11584;
	wire [4-1:0] node11588;
	wire [4-1:0] node11589;
	wire [4-1:0] node11592;
	wire [4-1:0] node11593;
	wire [4-1:0] node11596;
	wire [4-1:0] node11597;
	wire [4-1:0] node11601;
	wire [4-1:0] node11602;
	wire [4-1:0] node11603;
	wire [4-1:0] node11604;
	wire [4-1:0] node11605;
	wire [4-1:0] node11609;
	wire [4-1:0] node11612;
	wire [4-1:0] node11613;
	wire [4-1:0] node11616;
	wire [4-1:0] node11617;
	wire [4-1:0] node11621;
	wire [4-1:0] node11622;
	wire [4-1:0] node11623;
	wire [4-1:0] node11627;
	wire [4-1:0] node11628;
	wire [4-1:0] node11629;
	wire [4-1:0] node11633;
	wire [4-1:0] node11636;
	wire [4-1:0] node11637;
	wire [4-1:0] node11638;
	wire [4-1:0] node11640;
	wire [4-1:0] node11641;
	wire [4-1:0] node11642;
	wire [4-1:0] node11648;
	wire [4-1:0] node11649;
	wire [4-1:0] node11650;
	wire [4-1:0] node11651;
	wire [4-1:0] node11654;
	wire [4-1:0] node11655;
	wire [4-1:0] node11659;
	wire [4-1:0] node11660;
	wire [4-1:0] node11664;
	wire [4-1:0] node11666;
	wire [4-1:0] node11669;
	wire [4-1:0] node11670;
	wire [4-1:0] node11671;
	wire [4-1:0] node11672;
	wire [4-1:0] node11673;
	wire [4-1:0] node11676;
	wire [4-1:0] node11677;
	wire [4-1:0] node11681;
	wire [4-1:0] node11684;
	wire [4-1:0] node11685;
	wire [4-1:0] node11686;
	wire [4-1:0] node11690;
	wire [4-1:0] node11691;
	wire [4-1:0] node11693;
	wire [4-1:0] node11696;
	wire [4-1:0] node11697;
	wire [4-1:0] node11698;
	wire [4-1:0] node11702;
	wire [4-1:0] node11703;
	wire [4-1:0] node11706;
	wire [4-1:0] node11709;
	wire [4-1:0] node11710;
	wire [4-1:0] node11711;
	wire [4-1:0] node11714;
	wire [4-1:0] node11716;
	wire [4-1:0] node11717;
	wire [4-1:0] node11719;
	wire [4-1:0] node11723;
	wire [4-1:0] node11724;
	wire [4-1:0] node11725;
	wire [4-1:0] node11727;
	wire [4-1:0] node11731;
	wire [4-1:0] node11732;
	wire [4-1:0] node11736;
	wire [4-1:0] node11737;
	wire [4-1:0] node11738;
	wire [4-1:0] node11739;
	wire [4-1:0] node11740;
	wire [4-1:0] node11741;
	wire [4-1:0] node11742;
	wire [4-1:0] node11744;
	wire [4-1:0] node11748;
	wire [4-1:0] node11749;
	wire [4-1:0] node11754;
	wire [4-1:0] node11755;
	wire [4-1:0] node11756;
	wire [4-1:0] node11758;
	wire [4-1:0] node11759;
	wire [4-1:0] node11762;
	wire [4-1:0] node11765;
	wire [4-1:0] node11768;
	wire [4-1:0] node11769;
	wire [4-1:0] node11773;
	wire [4-1:0] node11774;
	wire [4-1:0] node11775;
	wire [4-1:0] node11776;
	wire [4-1:0] node11777;
	wire [4-1:0] node11778;
	wire [4-1:0] node11782;
	wire [4-1:0] node11784;
	wire [4-1:0] node11788;
	wire [4-1:0] node11789;
	wire [4-1:0] node11791;
	wire [4-1:0] node11795;
	wire [4-1:0] node11796;
	wire [4-1:0] node11798;
	wire [4-1:0] node11799;
	wire [4-1:0] node11800;
	wire [4-1:0] node11803;
	wire [4-1:0] node11807;
	wire [4-1:0] node11809;
	wire [4-1:0] node11810;
	wire [4-1:0] node11814;
	wire [4-1:0] node11815;
	wire [4-1:0] node11816;
	wire [4-1:0] node11817;
	wire [4-1:0] node11818;
	wire [4-1:0] node11821;
	wire [4-1:0] node11824;
	wire [4-1:0] node11825;
	wire [4-1:0] node11826;
	wire [4-1:0] node11830;
	wire [4-1:0] node11833;
	wire [4-1:0] node11834;
	wire [4-1:0] node11835;
	wire [4-1:0] node11838;
	wire [4-1:0] node11841;
	wire [4-1:0] node11842;
	wire [4-1:0] node11844;
	wire [4-1:0] node11847;
	wire [4-1:0] node11849;
	wire [4-1:0] node11850;
	wire [4-1:0] node11853;
	wire [4-1:0] node11856;
	wire [4-1:0] node11857;
	wire [4-1:0] node11858;
	wire [4-1:0] node11859;
	wire [4-1:0] node11861;
	wire [4-1:0] node11865;
	wire [4-1:0] node11868;
	wire [4-1:0] node11869;
	wire [4-1:0] node11870;
	wire [4-1:0] node11872;
	wire [4-1:0] node11875;
	wire [4-1:0] node11876;
	wire [4-1:0] node11880;
	wire [4-1:0] node11882;
	wire [4-1:0] node11885;
	wire [4-1:0] node11886;
	wire [4-1:0] node11887;
	wire [4-1:0] node11888;
	wire [4-1:0] node11889;
	wire [4-1:0] node11890;
	wire [4-1:0] node11891;
	wire [4-1:0] node11892;
	wire [4-1:0] node11893;
	wire [4-1:0] node11896;
	wire [4-1:0] node11899;
	wire [4-1:0] node11902;
	wire [4-1:0] node11903;
	wire [4-1:0] node11907;
	wire [4-1:0] node11908;
	wire [4-1:0] node11909;
	wire [4-1:0] node11910;
	wire [4-1:0] node11911;
	wire [4-1:0] node11914;
	wire [4-1:0] node11918;
	wire [4-1:0] node11921;
	wire [4-1:0] node11922;
	wire [4-1:0] node11924;
	wire [4-1:0] node11926;
	wire [4-1:0] node11929;
	wire [4-1:0] node11932;
	wire [4-1:0] node11933;
	wire [4-1:0] node11934;
	wire [4-1:0] node11935;
	wire [4-1:0] node11937;
	wire [4-1:0] node11940;
	wire [4-1:0] node11943;
	wire [4-1:0] node11944;
	wire [4-1:0] node11946;
	wire [4-1:0] node11948;
	wire [4-1:0] node11952;
	wire [4-1:0] node11953;
	wire [4-1:0] node11954;
	wire [4-1:0] node11955;
	wire [4-1:0] node11956;
	wire [4-1:0] node11962;
	wire [4-1:0] node11964;
	wire [4-1:0] node11967;
	wire [4-1:0] node11968;
	wire [4-1:0] node11969;
	wire [4-1:0] node11970;
	wire [4-1:0] node11971;
	wire [4-1:0] node11972;
	wire [4-1:0] node11975;
	wire [4-1:0] node11977;
	wire [4-1:0] node11980;
	wire [4-1:0] node11982;
	wire [4-1:0] node11983;
	wire [4-1:0] node11987;
	wire [4-1:0] node11988;
	wire [4-1:0] node11991;
	wire [4-1:0] node11992;
	wire [4-1:0] node11996;
	wire [4-1:0] node11997;
	wire [4-1:0] node11998;
	wire [4-1:0] node12000;
	wire [4-1:0] node12003;
	wire [4-1:0] node12005;
	wire [4-1:0] node12008;
	wire [4-1:0] node12009;
	wire [4-1:0] node12012;
	wire [4-1:0] node12015;
	wire [4-1:0] node12016;
	wire [4-1:0] node12017;
	wire [4-1:0] node12019;
	wire [4-1:0] node12020;
	wire [4-1:0] node12021;
	wire [4-1:0] node12025;
	wire [4-1:0] node12026;
	wire [4-1:0] node12030;
	wire [4-1:0] node12032;
	wire [4-1:0] node12033;
	wire [4-1:0] node12036;
	wire [4-1:0] node12039;
	wire [4-1:0] node12040;
	wire [4-1:0] node12041;
	wire [4-1:0] node12042;
	wire [4-1:0] node12045;
	wire [4-1:0] node12049;
	wire [4-1:0] node12051;
	wire [4-1:0] node12053;
	wire [4-1:0] node12056;
	wire [4-1:0] node12057;
	wire [4-1:0] node12058;
	wire [4-1:0] node12059;
	wire [4-1:0] node12060;
	wire [4-1:0] node12061;
	wire [4-1:0] node12062;
	wire [4-1:0] node12063;
	wire [4-1:0] node12067;
	wire [4-1:0] node12071;
	wire [4-1:0] node12072;
	wire [4-1:0] node12074;
	wire [4-1:0] node12077;
	wire [4-1:0] node12078;
	wire [4-1:0] node12082;
	wire [4-1:0] node12083;
	wire [4-1:0] node12084;
	wire [4-1:0] node12085;
	wire [4-1:0] node12086;
	wire [4-1:0] node12092;
	wire [4-1:0] node12094;
	wire [4-1:0] node12096;
	wire [4-1:0] node12099;
	wire [4-1:0] node12100;
	wire [4-1:0] node12101;
	wire [4-1:0] node12103;
	wire [4-1:0] node12104;
	wire [4-1:0] node12108;
	wire [4-1:0] node12110;
	wire [4-1:0] node12112;
	wire [4-1:0] node12114;
	wire [4-1:0] node12117;
	wire [4-1:0] node12118;
	wire [4-1:0] node12119;
	wire [4-1:0] node12121;
	wire [4-1:0] node12125;
	wire [4-1:0] node12126;
	wire [4-1:0] node12127;
	wire [4-1:0] node12129;
	wire [4-1:0] node12132;
	wire [4-1:0] node12136;
	wire [4-1:0] node12137;
	wire [4-1:0] node12138;
	wire [4-1:0] node12139;
	wire [4-1:0] node12140;
	wire [4-1:0] node12141;
	wire [4-1:0] node12144;
	wire [4-1:0] node12145;
	wire [4-1:0] node12149;
	wire [4-1:0] node12151;
	wire [4-1:0] node12154;
	wire [4-1:0] node12155;
	wire [4-1:0] node12158;
	wire [4-1:0] node12159;
	wire [4-1:0] node12162;
	wire [4-1:0] node12165;
	wire [4-1:0] node12166;
	wire [4-1:0] node12167;
	wire [4-1:0] node12168;
	wire [4-1:0] node12171;
	wire [4-1:0] node12172;
	wire [4-1:0] node12176;
	wire [4-1:0] node12177;
	wire [4-1:0] node12180;
	wire [4-1:0] node12181;
	wire [4-1:0] node12185;
	wire [4-1:0] node12186;
	wire [4-1:0] node12188;
	wire [4-1:0] node12189;
	wire [4-1:0] node12193;
	wire [4-1:0] node12196;
	wire [4-1:0] node12197;
	wire [4-1:0] node12198;
	wire [4-1:0] node12200;
	wire [4-1:0] node12201;
	wire [4-1:0] node12203;
	wire [4-1:0] node12206;
	wire [4-1:0] node12209;
	wire [4-1:0] node12210;
	wire [4-1:0] node12212;
	wire [4-1:0] node12216;
	wire [4-1:0] node12217;
	wire [4-1:0] node12219;
	wire [4-1:0] node12220;
	wire [4-1:0] node12224;
	wire [4-1:0] node12225;
	wire [4-1:0] node12228;
	wire [4-1:0] node12229;
	wire [4-1:0] node12233;
	wire [4-1:0] node12234;
	wire [4-1:0] node12235;
	wire [4-1:0] node12236;
	wire [4-1:0] node12237;
	wire [4-1:0] node12238;
	wire [4-1:0] node12239;
	wire [4-1:0] node12240;
	wire [4-1:0] node12244;
	wire [4-1:0] node12245;
	wire [4-1:0] node12247;
	wire [4-1:0] node12251;
	wire [4-1:0] node12253;
	wire [4-1:0] node12254;
	wire [4-1:0] node12257;
	wire [4-1:0] node12259;
	wire [4-1:0] node12262;
	wire [4-1:0] node12263;
	wire [4-1:0] node12264;
	wire [4-1:0] node12265;
	wire [4-1:0] node12270;
	wire [4-1:0] node12271;
	wire [4-1:0] node12273;
	wire [4-1:0] node12274;
	wire [4-1:0] node12278;
	wire [4-1:0] node12281;
	wire [4-1:0] node12282;
	wire [4-1:0] node12283;
	wire [4-1:0] node12284;
	wire [4-1:0] node12286;
	wire [4-1:0] node12290;
	wire [4-1:0] node12291;
	wire [4-1:0] node12292;
	wire [4-1:0] node12296;
	wire [4-1:0] node12299;
	wire [4-1:0] node12300;
	wire [4-1:0] node12302;
	wire [4-1:0] node12304;
	wire [4-1:0] node12305;
	wire [4-1:0] node12308;
	wire [4-1:0] node12311;
	wire [4-1:0] node12312;
	wire [4-1:0] node12313;
	wire [4-1:0] node12316;
	wire [4-1:0] node12320;
	wire [4-1:0] node12321;
	wire [4-1:0] node12322;
	wire [4-1:0] node12323;
	wire [4-1:0] node12326;
	wire [4-1:0] node12327;
	wire [4-1:0] node12330;
	wire [4-1:0] node12331;
	wire [4-1:0] node12335;
	wire [4-1:0] node12336;
	wire [4-1:0] node12337;
	wire [4-1:0] node12341;
	wire [4-1:0] node12342;
	wire [4-1:0] node12344;
	wire [4-1:0] node12347;
	wire [4-1:0] node12350;
	wire [4-1:0] node12351;
	wire [4-1:0] node12352;
	wire [4-1:0] node12353;
	wire [4-1:0] node12355;
	wire [4-1:0] node12358;
	wire [4-1:0] node12359;
	wire [4-1:0] node12362;
	wire [4-1:0] node12364;
	wire [4-1:0] node12367;
	wire [4-1:0] node12368;
	wire [4-1:0] node12369;
	wire [4-1:0] node12370;
	wire [4-1:0] node12374;
	wire [4-1:0] node12378;
	wire [4-1:0] node12379;
	wire [4-1:0] node12380;
	wire [4-1:0] node12382;
	wire [4-1:0] node12384;
	wire [4-1:0] node12387;
	wire [4-1:0] node12388;
	wire [4-1:0] node12392;
	wire [4-1:0] node12393;
	wire [4-1:0] node12395;
	wire [4-1:0] node12398;
	wire [4-1:0] node12400;
	wire [4-1:0] node12403;
	wire [4-1:0] node12404;
	wire [4-1:0] node12405;
	wire [4-1:0] node12406;
	wire [4-1:0] node12407;
	wire [4-1:0] node12409;
	wire [4-1:0] node12410;
	wire [4-1:0] node12414;
	wire [4-1:0] node12415;
	wire [4-1:0] node12418;
	wire [4-1:0] node12420;
	wire [4-1:0] node12422;
	wire [4-1:0] node12425;
	wire [4-1:0] node12426;
	wire [4-1:0] node12427;
	wire [4-1:0] node12428;
	wire [4-1:0] node12430;
	wire [4-1:0] node12433;
	wire [4-1:0] node12435;
	wire [4-1:0] node12439;
	wire [4-1:0] node12441;
	wire [4-1:0] node12442;
	wire [4-1:0] node12443;
	wire [4-1:0] node12448;
	wire [4-1:0] node12449;
	wire [4-1:0] node12450;
	wire [4-1:0] node12451;
	wire [4-1:0] node12452;
	wire [4-1:0] node12454;
	wire [4-1:0] node12458;
	wire [4-1:0] node12460;
	wire [4-1:0] node12463;
	wire [4-1:0] node12464;
	wire [4-1:0] node12466;
	wire [4-1:0] node12469;
	wire [4-1:0] node12471;
	wire [4-1:0] node12474;
	wire [4-1:0] node12475;
	wire [4-1:0] node12477;
	wire [4-1:0] node12478;
	wire [4-1:0] node12480;
	wire [4-1:0] node12484;
	wire [4-1:0] node12486;
	wire [4-1:0] node12489;
	wire [4-1:0] node12490;
	wire [4-1:0] node12491;
	wire [4-1:0] node12492;
	wire [4-1:0] node12494;
	wire [4-1:0] node12496;
	wire [4-1:0] node12499;
	wire [4-1:0] node12500;
	wire [4-1:0] node12501;
	wire [4-1:0] node12502;
	wire [4-1:0] node12506;
	wire [4-1:0] node12507;
	wire [4-1:0] node12511;
	wire [4-1:0] node12513;
	wire [4-1:0] node12516;
	wire [4-1:0] node12517;
	wire [4-1:0] node12518;
	wire [4-1:0] node12519;
	wire [4-1:0] node12522;
	wire [4-1:0] node12523;
	wire [4-1:0] node12527;
	wire [4-1:0] node12528;
	wire [4-1:0] node12529;
	wire [4-1:0] node12532;
	wire [4-1:0] node12537;
	wire [4-1:0] node12538;
	wire [4-1:0] node12539;
	wire [4-1:0] node12540;
	wire [4-1:0] node12544;
	wire [4-1:0] node12546;
	wire [4-1:0] node12549;
	wire [4-1:0] node12550;
	wire [4-1:0] node12551;
	wire [4-1:0] node12552;
	wire [4-1:0] node12557;
	wire [4-1:0] node12559;
	wire [4-1:0] node12562;
	wire [4-1:0] node12563;
	wire [4-1:0] node12564;
	wire [4-1:0] node12565;
	wire [4-1:0] node12566;
	wire [4-1:0] node12567;
	wire [4-1:0] node12568;
	wire [4-1:0] node12569;
	wire [4-1:0] node12571;
	wire [4-1:0] node12572;
	wire [4-1:0] node12573;
	wire [4-1:0] node12578;
	wire [4-1:0] node12579;
	wire [4-1:0] node12582;
	wire [4-1:0] node12583;
	wire [4-1:0] node12585;
	wire [4-1:0] node12588;
	wire [4-1:0] node12591;
	wire [4-1:0] node12592;
	wire [4-1:0] node12593;
	wire [4-1:0] node12595;
	wire [4-1:0] node12598;
	wire [4-1:0] node12599;
	wire [4-1:0] node12601;
	wire [4-1:0] node12604;
	wire [4-1:0] node12605;
	wire [4-1:0] node12609;
	wire [4-1:0] node12610;
	wire [4-1:0] node12611;
	wire [4-1:0] node12616;
	wire [4-1:0] node12617;
	wire [4-1:0] node12618;
	wire [4-1:0] node12619;
	wire [4-1:0] node12620;
	wire [4-1:0] node12624;
	wire [4-1:0] node12627;
	wire [4-1:0] node12628;
	wire [4-1:0] node12629;
	wire [4-1:0] node12631;
	wire [4-1:0] node12634;
	wire [4-1:0] node12637;
	wire [4-1:0] node12638;
	wire [4-1:0] node12642;
	wire [4-1:0] node12643;
	wire [4-1:0] node12644;
	wire [4-1:0] node12645;
	wire [4-1:0] node12648;
	wire [4-1:0] node12650;
	wire [4-1:0] node12653;
	wire [4-1:0] node12655;
	wire [4-1:0] node12658;
	wire [4-1:0] node12659;
	wire [4-1:0] node12661;
	wire [4-1:0] node12662;
	wire [4-1:0] node12666;
	wire [4-1:0] node12667;
	wire [4-1:0] node12670;
	wire [4-1:0] node12673;
	wire [4-1:0] node12674;
	wire [4-1:0] node12675;
	wire [4-1:0] node12676;
	wire [4-1:0] node12677;
	wire [4-1:0] node12679;
	wire [4-1:0] node12682;
	wire [4-1:0] node12683;
	wire [4-1:0] node12687;
	wire [4-1:0] node12688;
	wire [4-1:0] node12691;
	wire [4-1:0] node12693;
	wire [4-1:0] node12695;
	wire [4-1:0] node12698;
	wire [4-1:0] node12699;
	wire [4-1:0] node12700;
	wire [4-1:0] node12702;
	wire [4-1:0] node12705;
	wire [4-1:0] node12708;
	wire [4-1:0] node12709;
	wire [4-1:0] node12710;
	wire [4-1:0] node12712;
	wire [4-1:0] node12715;
	wire [4-1:0] node12717;
	wire [4-1:0] node12720;
	wire [4-1:0] node12721;
	wire [4-1:0] node12725;
	wire [4-1:0] node12726;
	wire [4-1:0] node12727;
	wire [4-1:0] node12728;
	wire [4-1:0] node12731;
	wire [4-1:0] node12734;
	wire [4-1:0] node12735;
	wire [4-1:0] node12736;
	wire [4-1:0] node12738;
	wire [4-1:0] node12742;
	wire [4-1:0] node12743;
	wire [4-1:0] node12746;
	wire [4-1:0] node12749;
	wire [4-1:0] node12750;
	wire [4-1:0] node12751;
	wire [4-1:0] node12752;
	wire [4-1:0] node12753;
	wire [4-1:0] node12758;
	wire [4-1:0] node12760;
	wire [4-1:0] node12761;
	wire [4-1:0] node12765;
	wire [4-1:0] node12767;
	wire [4-1:0] node12769;
	wire [4-1:0] node12772;
	wire [4-1:0] node12773;
	wire [4-1:0] node12774;
	wire [4-1:0] node12775;
	wire [4-1:0] node12776;
	wire [4-1:0] node12777;
	wire [4-1:0] node12778;
	wire [4-1:0] node12779;
	wire [4-1:0] node12784;
	wire [4-1:0] node12786;
	wire [4-1:0] node12789;
	wire [4-1:0] node12790;
	wire [4-1:0] node12792;
	wire [4-1:0] node12793;
	wire [4-1:0] node12797;
	wire [4-1:0] node12798;
	wire [4-1:0] node12801;
	wire [4-1:0] node12803;
	wire [4-1:0] node12806;
	wire [4-1:0] node12807;
	wire [4-1:0] node12808;
	wire [4-1:0] node12809;
	wire [4-1:0] node12812;
	wire [4-1:0] node12815;
	wire [4-1:0] node12816;
	wire [4-1:0] node12818;
	wire [4-1:0] node12822;
	wire [4-1:0] node12823;
	wire [4-1:0] node12824;
	wire [4-1:0] node12825;
	wire [4-1:0] node12829;
	wire [4-1:0] node12831;
	wire [4-1:0] node12834;
	wire [4-1:0] node12836;
	wire [4-1:0] node12837;
	wire [4-1:0] node12841;
	wire [4-1:0] node12842;
	wire [4-1:0] node12843;
	wire [4-1:0] node12844;
	wire [4-1:0] node12845;
	wire [4-1:0] node12846;
	wire [4-1:0] node12850;
	wire [4-1:0] node12853;
	wire [4-1:0] node12855;
	wire [4-1:0] node12857;
	wire [4-1:0] node12860;
	wire [4-1:0] node12861;
	wire [4-1:0] node12862;
	wire [4-1:0] node12863;
	wire [4-1:0] node12866;
	wire [4-1:0] node12869;
	wire [4-1:0] node12872;
	wire [4-1:0] node12873;
	wire [4-1:0] node12876;
	wire [4-1:0] node12879;
	wire [4-1:0] node12880;
	wire [4-1:0] node12881;
	wire [4-1:0] node12883;
	wire [4-1:0] node12885;
	wire [4-1:0] node12889;
	wire [4-1:0] node12890;
	wire [4-1:0] node12891;
	wire [4-1:0] node12893;
	wire [4-1:0] node12897;
	wire [4-1:0] node12898;
	wire [4-1:0] node12900;
	wire [4-1:0] node12903;
	wire [4-1:0] node12906;
	wire [4-1:0] node12907;
	wire [4-1:0] node12908;
	wire [4-1:0] node12909;
	wire [4-1:0] node12911;
	wire [4-1:0] node12912;
	wire [4-1:0] node12916;
	wire [4-1:0] node12917;
	wire [4-1:0] node12918;
	wire [4-1:0] node12920;
	wire [4-1:0] node12924;
	wire [4-1:0] node12925;
	wire [4-1:0] node12928;
	wire [4-1:0] node12930;
	wire [4-1:0] node12933;
	wire [4-1:0] node12934;
	wire [4-1:0] node12936;
	wire [4-1:0] node12939;
	wire [4-1:0] node12940;
	wire [4-1:0] node12941;
	wire [4-1:0] node12943;
	wire [4-1:0] node12947;
	wire [4-1:0] node12950;
	wire [4-1:0] node12951;
	wire [4-1:0] node12953;
	wire [4-1:0] node12954;
	wire [4-1:0] node12955;
	wire [4-1:0] node12959;
	wire [4-1:0] node12960;
	wire [4-1:0] node12964;
	wire [4-1:0] node12965;
	wire [4-1:0] node12967;
	wire [4-1:0] node12968;
	wire [4-1:0] node12971;
	wire [4-1:0] node12972;
	wire [4-1:0] node12975;
	wire [4-1:0] node12978;
	wire [4-1:0] node12979;
	wire [4-1:0] node12982;
	wire [4-1:0] node12983;
	wire [4-1:0] node12987;
	wire [4-1:0] node12988;
	wire [4-1:0] node12989;
	wire [4-1:0] node12990;
	wire [4-1:0] node12991;
	wire [4-1:0] node12992;
	wire [4-1:0] node12993;
	wire [4-1:0] node12997;
	wire [4-1:0] node13000;
	wire [4-1:0] node13001;
	wire [4-1:0] node13002;
	wire [4-1:0] node13003;
	wire [4-1:0] node13008;
	wire [4-1:0] node13011;
	wire [4-1:0] node13012;
	wire [4-1:0] node13013;
	wire [4-1:0] node13014;
	wire [4-1:0] node13015;
	wire [4-1:0] node13016;
	wire [4-1:0] node13021;
	wire [4-1:0] node13023;
	wire [4-1:0] node13026;
	wire [4-1:0] node13027;
	wire [4-1:0] node13028;
	wire [4-1:0] node13031;
	wire [4-1:0] node13034;
	wire [4-1:0] node13036;
	wire [4-1:0] node13039;
	wire [4-1:0] node13040;
	wire [4-1:0] node13041;
	wire [4-1:0] node13043;
	wire [4-1:0] node13046;
	wire [4-1:0] node13047;
	wire [4-1:0] node13051;
	wire [4-1:0] node13052;
	wire [4-1:0] node13054;
	wire [4-1:0] node13057;
	wire [4-1:0] node13060;
	wire [4-1:0] node13061;
	wire [4-1:0] node13062;
	wire [4-1:0] node13064;
	wire [4-1:0] node13065;
	wire [4-1:0] node13069;
	wire [4-1:0] node13070;
	wire [4-1:0] node13071;
	wire [4-1:0] node13074;
	wire [4-1:0] node13076;
	wire [4-1:0] node13079;
	wire [4-1:0] node13080;
	wire [4-1:0] node13082;
	wire [4-1:0] node13083;
	wire [4-1:0] node13087;
	wire [4-1:0] node13088;
	wire [4-1:0] node13092;
	wire [4-1:0] node13093;
	wire [4-1:0] node13094;
	wire [4-1:0] node13095;
	wire [4-1:0] node13098;
	wire [4-1:0] node13101;
	wire [4-1:0] node13102;
	wire [4-1:0] node13103;
	wire [4-1:0] node13104;
	wire [4-1:0] node13108;
	wire [4-1:0] node13110;
	wire [4-1:0] node13114;
	wire [4-1:0] node13116;
	wire [4-1:0] node13118;
	wire [4-1:0] node13121;
	wire [4-1:0] node13122;
	wire [4-1:0] node13123;
	wire [4-1:0] node13124;
	wire [4-1:0] node13125;
	wire [4-1:0] node13127;
	wire [4-1:0] node13129;
	wire [4-1:0] node13132;
	wire [4-1:0] node13134;
	wire [4-1:0] node13135;
	wire [4-1:0] node13139;
	wire [4-1:0] node13140;
	wire [4-1:0] node13141;
	wire [4-1:0] node13143;
	wire [4-1:0] node13148;
	wire [4-1:0] node13149;
	wire [4-1:0] node13150;
	wire [4-1:0] node13152;
	wire [4-1:0] node13153;
	wire [4-1:0] node13154;
	wire [4-1:0] node13158;
	wire [4-1:0] node13160;
	wire [4-1:0] node13163;
	wire [4-1:0] node13165;
	wire [4-1:0] node13166;
	wire [4-1:0] node13170;
	wire [4-1:0] node13171;
	wire [4-1:0] node13172;
	wire [4-1:0] node13176;
	wire [4-1:0] node13177;
	wire [4-1:0] node13179;
	wire [4-1:0] node13183;
	wire [4-1:0] node13184;
	wire [4-1:0] node13185;
	wire [4-1:0] node13186;
	wire [4-1:0] node13187;
	wire [4-1:0] node13189;
	wire [4-1:0] node13190;
	wire [4-1:0] node13195;
	wire [4-1:0] node13197;
	wire [4-1:0] node13200;
	wire [4-1:0] node13202;
	wire [4-1:0] node13203;
	wire [4-1:0] node13207;
	wire [4-1:0] node13208;
	wire [4-1:0] node13209;
	wire [4-1:0] node13210;
	wire [4-1:0] node13211;
	wire [4-1:0] node13215;
	wire [4-1:0] node13217;
	wire [4-1:0] node13218;
	wire [4-1:0] node13222;
	wire [4-1:0] node13224;
	wire [4-1:0] node13227;
	wire [4-1:0] node13228;
	wire [4-1:0] node13230;
	wire [4-1:0] node13232;
	wire [4-1:0] node13235;
	wire [4-1:0] node13237;
	wire [4-1:0] node13240;
	wire [4-1:0] node13241;
	wire [4-1:0] node13242;
	wire [4-1:0] node13243;
	wire [4-1:0] node13244;
	wire [4-1:0] node13245;
	wire [4-1:0] node13246;
	wire [4-1:0] node13247;
	wire [4-1:0] node13250;
	wire [4-1:0] node13251;
	wire [4-1:0] node13255;
	wire [4-1:0] node13256;
	wire [4-1:0] node13258;
	wire [4-1:0] node13261;
	wire [4-1:0] node13262;
	wire [4-1:0] node13264;
	wire [4-1:0] node13267;
	wire [4-1:0] node13270;
	wire [4-1:0] node13271;
	wire [4-1:0] node13272;
	wire [4-1:0] node13276;
	wire [4-1:0] node13277;
	wire [4-1:0] node13278;
	wire [4-1:0] node13282;
	wire [4-1:0] node13285;
	wire [4-1:0] node13286;
	wire [4-1:0] node13287;
	wire [4-1:0] node13288;
	wire [4-1:0] node13289;
	wire [4-1:0] node13293;
	wire [4-1:0] node13294;
	wire [4-1:0] node13298;
	wire [4-1:0] node13299;
	wire [4-1:0] node13301;
	wire [4-1:0] node13304;
	wire [4-1:0] node13305;
	wire [4-1:0] node13309;
	wire [4-1:0] node13310;
	wire [4-1:0] node13311;
	wire [4-1:0] node13314;
	wire [4-1:0] node13317;
	wire [4-1:0] node13318;
	wire [4-1:0] node13319;
	wire [4-1:0] node13320;
	wire [4-1:0] node13324;
	wire [4-1:0] node13325;
	wire [4-1:0] node13329;
	wire [4-1:0] node13331;
	wire [4-1:0] node13334;
	wire [4-1:0] node13335;
	wire [4-1:0] node13336;
	wire [4-1:0] node13337;
	wire [4-1:0] node13338;
	wire [4-1:0] node13342;
	wire [4-1:0] node13345;
	wire [4-1:0] node13346;
	wire [4-1:0] node13348;
	wire [4-1:0] node13349;
	wire [4-1:0] node13354;
	wire [4-1:0] node13355;
	wire [4-1:0] node13356;
	wire [4-1:0] node13357;
	wire [4-1:0] node13360;
	wire [4-1:0] node13361;
	wire [4-1:0] node13362;
	wire [4-1:0] node13367;
	wire [4-1:0] node13368;
	wire [4-1:0] node13371;
	wire [4-1:0] node13372;
	wire [4-1:0] node13374;
	wire [4-1:0] node13378;
	wire [4-1:0] node13379;
	wire [4-1:0] node13380;
	wire [4-1:0] node13381;
	wire [4-1:0] node13382;
	wire [4-1:0] node13387;
	wire [4-1:0] node13389;
	wire [4-1:0] node13390;
	wire [4-1:0] node13393;
	wire [4-1:0] node13396;
	wire [4-1:0] node13398;
	wire [4-1:0] node13400;
	wire [4-1:0] node13403;
	wire [4-1:0] node13404;
	wire [4-1:0] node13405;
	wire [4-1:0] node13406;
	wire [4-1:0] node13407;
	wire [4-1:0] node13410;
	wire [4-1:0] node13411;
	wire [4-1:0] node13412;
	wire [4-1:0] node13414;
	wire [4-1:0] node13417;
	wire [4-1:0] node13419;
	wire [4-1:0] node13423;
	wire [4-1:0] node13424;
	wire [4-1:0] node13425;
	wire [4-1:0] node13428;
	wire [4-1:0] node13429;
	wire [4-1:0] node13432;
	wire [4-1:0] node13434;
	wire [4-1:0] node13437;
	wire [4-1:0] node13439;
	wire [4-1:0] node13440;
	wire [4-1:0] node13441;
	wire [4-1:0] node13446;
	wire [4-1:0] node13447;
	wire [4-1:0] node13448;
	wire [4-1:0] node13449;
	wire [4-1:0] node13451;
	wire [4-1:0] node13454;
	wire [4-1:0] node13455;
	wire [4-1:0] node13456;
	wire [4-1:0] node13460;
	wire [4-1:0] node13461;
	wire [4-1:0] node13465;
	wire [4-1:0] node13466;
	wire [4-1:0] node13468;
	wire [4-1:0] node13471;
	wire [4-1:0] node13473;
	wire [4-1:0] node13474;
	wire [4-1:0] node13478;
	wire [4-1:0] node13479;
	wire [4-1:0] node13480;
	wire [4-1:0] node13481;
	wire [4-1:0] node13484;
	wire [4-1:0] node13487;
	wire [4-1:0] node13488;
	wire [4-1:0] node13489;
	wire [4-1:0] node13494;
	wire [4-1:0] node13496;
	wire [4-1:0] node13499;
	wire [4-1:0] node13500;
	wire [4-1:0] node13501;
	wire [4-1:0] node13502;
	wire [4-1:0] node13503;
	wire [4-1:0] node13504;
	wire [4-1:0] node13507;
	wire [4-1:0] node13509;
	wire [4-1:0] node13513;
	wire [4-1:0] node13514;
	wire [4-1:0] node13515;
	wire [4-1:0] node13517;
	wire [4-1:0] node13522;
	wire [4-1:0] node13523;
	wire [4-1:0] node13525;
	wire [4-1:0] node13526;
	wire [4-1:0] node13528;
	wire [4-1:0] node13532;
	wire [4-1:0] node13533;
	wire [4-1:0] node13534;
	wire [4-1:0] node13539;
	wire [4-1:0] node13540;
	wire [4-1:0] node13541;
	wire [4-1:0] node13544;
	wire [4-1:0] node13545;
	wire [4-1:0] node13548;
	wire [4-1:0] node13549;
	wire [4-1:0] node13550;
	wire [4-1:0] node13554;
	wire [4-1:0] node13556;
	wire [4-1:0] node13559;
	wire [4-1:0] node13560;
	wire [4-1:0] node13561;
	wire [4-1:0] node13562;
	wire [4-1:0] node13563;
	wire [4-1:0] node13569;
	wire [4-1:0] node13572;
	wire [4-1:0] node13573;
	wire [4-1:0] node13574;
	wire [4-1:0] node13575;
	wire [4-1:0] node13576;
	wire [4-1:0] node13577;
	wire [4-1:0] node13578;
	wire [4-1:0] node13579;
	wire [4-1:0] node13584;
	wire [4-1:0] node13585;
	wire [4-1:0] node13586;
	wire [4-1:0] node13589;
	wire [4-1:0] node13592;
	wire [4-1:0] node13593;
	wire [4-1:0] node13597;
	wire [4-1:0] node13598;
	wire [4-1:0] node13599;
	wire [4-1:0] node13601;
	wire [4-1:0] node13603;
	wire [4-1:0] node13607;
	wire [4-1:0] node13608;
	wire [4-1:0] node13609;
	wire [4-1:0] node13614;
	wire [4-1:0] node13615;
	wire [4-1:0] node13616;
	wire [4-1:0] node13617;
	wire [4-1:0] node13619;
	wire [4-1:0] node13621;
	wire [4-1:0] node13624;
	wire [4-1:0] node13627;
	wire [4-1:0] node13629;
	wire [4-1:0] node13630;
	wire [4-1:0] node13631;
	wire [4-1:0] node13636;
	wire [4-1:0] node13637;
	wire [4-1:0] node13638;
	wire [4-1:0] node13639;
	wire [4-1:0] node13642;
	wire [4-1:0] node13645;
	wire [4-1:0] node13646;
	wire [4-1:0] node13650;
	wire [4-1:0] node13651;
	wire [4-1:0] node13652;
	wire [4-1:0] node13655;
	wire [4-1:0] node13656;
	wire [4-1:0] node13661;
	wire [4-1:0] node13662;
	wire [4-1:0] node13663;
	wire [4-1:0] node13664;
	wire [4-1:0] node13665;
	wire [4-1:0] node13667;
	wire [4-1:0] node13668;
	wire [4-1:0] node13673;
	wire [4-1:0] node13674;
	wire [4-1:0] node13676;
	wire [4-1:0] node13679;
	wire [4-1:0] node13681;
	wire [4-1:0] node13684;
	wire [4-1:0] node13685;
	wire [4-1:0] node13686;
	wire [4-1:0] node13689;
	wire [4-1:0] node13690;
	wire [4-1:0] node13694;
	wire [4-1:0] node13697;
	wire [4-1:0] node13698;
	wire [4-1:0] node13699;
	wire [4-1:0] node13700;
	wire [4-1:0] node13702;
	wire [4-1:0] node13703;
	wire [4-1:0] node13707;
	wire [4-1:0] node13710;
	wire [4-1:0] node13711;
	wire [4-1:0] node13712;
	wire [4-1:0] node13717;
	wire [4-1:0] node13718;
	wire [4-1:0] node13719;
	wire [4-1:0] node13720;
	wire [4-1:0] node13721;
	wire [4-1:0] node13727;
	wire [4-1:0] node13729;
	wire [4-1:0] node13732;
	wire [4-1:0] node13733;
	wire [4-1:0] node13734;
	wire [4-1:0] node13735;
	wire [4-1:0] node13736;
	wire [4-1:0] node13738;
	wire [4-1:0] node13739;
	wire [4-1:0] node13743;
	wire [4-1:0] node13744;
	wire [4-1:0] node13745;
	wire [4-1:0] node13749;
	wire [4-1:0] node13752;
	wire [4-1:0] node13753;
	wire [4-1:0] node13754;
	wire [4-1:0] node13755;
	wire [4-1:0] node13756;
	wire [4-1:0] node13761;
	wire [4-1:0] node13764;
	wire [4-1:0] node13765;
	wire [4-1:0] node13768;
	wire [4-1:0] node13770;
	wire [4-1:0] node13771;
	wire [4-1:0] node13775;
	wire [4-1:0] node13776;
	wire [4-1:0] node13777;
	wire [4-1:0] node13778;
	wire [4-1:0] node13780;
	wire [4-1:0] node13784;
	wire [4-1:0] node13785;
	wire [4-1:0] node13787;
	wire [4-1:0] node13788;
	wire [4-1:0] node13791;
	wire [4-1:0] node13794;
	wire [4-1:0] node13795;
	wire [4-1:0] node13799;
	wire [4-1:0] node13800;
	wire [4-1:0] node13801;
	wire [4-1:0] node13804;
	wire [4-1:0] node13806;
	wire [4-1:0] node13809;
	wire [4-1:0] node13810;
	wire [4-1:0] node13811;
	wire [4-1:0] node13815;
	wire [4-1:0] node13818;
	wire [4-1:0] node13819;
	wire [4-1:0] node13820;
	wire [4-1:0] node13821;
	wire [4-1:0] node13822;
	wire [4-1:0] node13823;
	wire [4-1:0] node13824;
	wire [4-1:0] node13830;
	wire [4-1:0] node13831;
	wire [4-1:0] node13835;
	wire [4-1:0] node13836;
	wire [4-1:0] node13837;
	wire [4-1:0] node13840;
	wire [4-1:0] node13841;
	wire [4-1:0] node13844;
	wire [4-1:0] node13847;
	wire [4-1:0] node13850;
	wire [4-1:0] node13851;
	wire [4-1:0] node13852;
	wire [4-1:0] node13853;
	wire [4-1:0] node13854;
	wire [4-1:0] node13857;
	wire [4-1:0] node13858;
	wire [4-1:0] node13862;
	wire [4-1:0] node13864;
	wire [4-1:0] node13867;
	wire [4-1:0] node13869;
	wire [4-1:0] node13871;
	wire [4-1:0] node13872;
	wire [4-1:0] node13876;
	wire [4-1:0] node13877;
	wire [4-1:0] node13879;
	wire [4-1:0] node13880;
	wire [4-1:0] node13881;
	wire [4-1:0] node13886;
	wire [4-1:0] node13887;
	wire [4-1:0] node13890;
	wire [4-1:0] node13893;
	wire [4-1:0] node13894;
	wire [4-1:0] node13895;
	wire [4-1:0] node13896;
	wire [4-1:0] node13897;
	wire [4-1:0] node13898;
	wire [4-1:0] node13899;
	wire [4-1:0] node13900;
	wire [4-1:0] node13901;
	wire [4-1:0] node13902;
	wire [4-1:0] node13903;
	wire [4-1:0] node13907;
	wire [4-1:0] node13909;
	wire [4-1:0] node13912;
	wire [4-1:0] node13913;
	wire [4-1:0] node13914;
	wire [4-1:0] node13917;
	wire [4-1:0] node13918;
	wire [4-1:0] node13922;
	wire [4-1:0] node13923;
	wire [4-1:0] node13926;
	wire [4-1:0] node13927;
	wire [4-1:0] node13931;
	wire [4-1:0] node13932;
	wire [4-1:0] node13933;
	wire [4-1:0] node13934;
	wire [4-1:0] node13938;
	wire [4-1:0] node13939;
	wire [4-1:0] node13942;
	wire [4-1:0] node13944;
	wire [4-1:0] node13947;
	wire [4-1:0] node13949;
	wire [4-1:0] node13952;
	wire [4-1:0] node13953;
	wire [4-1:0] node13954;
	wire [4-1:0] node13955;
	wire [4-1:0] node13958;
	wire [4-1:0] node13961;
	wire [4-1:0] node13963;
	wire [4-1:0] node13964;
	wire [4-1:0] node13966;
	wire [4-1:0] node13970;
	wire [4-1:0] node13972;
	wire [4-1:0] node13973;
	wire [4-1:0] node13977;
	wire [4-1:0] node13978;
	wire [4-1:0] node13979;
	wire [4-1:0] node13980;
	wire [4-1:0] node13982;
	wire [4-1:0] node13983;
	wire [4-1:0] node13984;
	wire [4-1:0] node13987;
	wire [4-1:0] node13991;
	wire [4-1:0] node13993;
	wire [4-1:0] node13996;
	wire [4-1:0] node13997;
	wire [4-1:0] node13998;
	wire [4-1:0] node14001;
	wire [4-1:0] node14003;
	wire [4-1:0] node14006;
	wire [4-1:0] node14007;
	wire [4-1:0] node14008;
	wire [4-1:0] node14011;
	wire [4-1:0] node14012;
	wire [4-1:0] node14015;
	wire [4-1:0] node14019;
	wire [4-1:0] node14020;
	wire [4-1:0] node14021;
	wire [4-1:0] node14023;
	wire [4-1:0] node14025;
	wire [4-1:0] node14028;
	wire [4-1:0] node14029;
	wire [4-1:0] node14030;
	wire [4-1:0] node14034;
	wire [4-1:0] node14036;
	wire [4-1:0] node14039;
	wire [4-1:0] node14040;
	wire [4-1:0] node14041;
	wire [4-1:0] node14042;
	wire [4-1:0] node14043;
	wire [4-1:0] node14048;
	wire [4-1:0] node14050;
	wire [4-1:0] node14053;
	wire [4-1:0] node14054;
	wire [4-1:0] node14055;
	wire [4-1:0] node14056;
	wire [4-1:0] node14061;
	wire [4-1:0] node14063;
	wire [4-1:0] node14064;
	wire [4-1:0] node14068;
	wire [4-1:0] node14069;
	wire [4-1:0] node14070;
	wire [4-1:0] node14071;
	wire [4-1:0] node14072;
	wire [4-1:0] node14073;
	wire [4-1:0] node14074;
	wire [4-1:0] node14078;
	wire [4-1:0] node14079;
	wire [4-1:0] node14083;
	wire [4-1:0] node14086;
	wire [4-1:0] node14087;
	wire [4-1:0] node14088;
	wire [4-1:0] node14089;
	wire [4-1:0] node14093;
	wire [4-1:0] node14094;
	wire [4-1:0] node14095;
	wire [4-1:0] node14098;
	wire [4-1:0] node14101;
	wire [4-1:0] node14104;
	wire [4-1:0] node14106;
	wire [4-1:0] node14109;
	wire [4-1:0] node14110;
	wire [4-1:0] node14111;
	wire [4-1:0] node14113;
	wire [4-1:0] node14116;
	wire [4-1:0] node14117;
	wire [4-1:0] node14121;
	wire [4-1:0] node14122;
	wire [4-1:0] node14123;
	wire [4-1:0] node14124;
	wire [4-1:0] node14128;
	wire [4-1:0] node14130;
	wire [4-1:0] node14133;
	wire [4-1:0] node14134;
	wire [4-1:0] node14135;
	wire [4-1:0] node14138;
	wire [4-1:0] node14139;
	wire [4-1:0] node14143;
	wire [4-1:0] node14146;
	wire [4-1:0] node14147;
	wire [4-1:0] node14148;
	wire [4-1:0] node14149;
	wire [4-1:0] node14150;
	wire [4-1:0] node14152;
	wire [4-1:0] node14153;
	wire [4-1:0] node14156;
	wire [4-1:0] node14159;
	wire [4-1:0] node14160;
	wire [4-1:0] node14164;
	wire [4-1:0] node14165;
	wire [4-1:0] node14167;
	wire [4-1:0] node14170;
	wire [4-1:0] node14173;
	wire [4-1:0] node14174;
	wire [4-1:0] node14175;
	wire [4-1:0] node14177;
	wire [4-1:0] node14180;
	wire [4-1:0] node14181;
	wire [4-1:0] node14185;
	wire [4-1:0] node14186;
	wire [4-1:0] node14189;
	wire [4-1:0] node14190;
	wire [4-1:0] node14194;
	wire [4-1:0] node14195;
	wire [4-1:0] node14196;
	wire [4-1:0] node14197;
	wire [4-1:0] node14199;
	wire [4-1:0] node14202;
	wire [4-1:0] node14203;
	wire [4-1:0] node14207;
	wire [4-1:0] node14208;
	wire [4-1:0] node14210;
	wire [4-1:0] node14213;
	wire [4-1:0] node14214;
	wire [4-1:0] node14217;
	wire [4-1:0] node14220;
	wire [4-1:0] node14221;
	wire [4-1:0] node14222;
	wire [4-1:0] node14224;
	wire [4-1:0] node14227;
	wire [4-1:0] node14228;
	wire [4-1:0] node14231;
	wire [4-1:0] node14234;
	wire [4-1:0] node14236;
	wire [4-1:0] node14238;
	wire [4-1:0] node14239;
	wire [4-1:0] node14243;
	wire [4-1:0] node14244;
	wire [4-1:0] node14245;
	wire [4-1:0] node14246;
	wire [4-1:0] node14247;
	wire [4-1:0] node14248;
	wire [4-1:0] node14249;
	wire [4-1:0] node14250;
	wire [4-1:0] node14252;
	wire [4-1:0] node14256;
	wire [4-1:0] node14257;
	wire [4-1:0] node14258;
	wire [4-1:0] node14261;
	wire [4-1:0] node14265;
	wire [4-1:0] node14266;
	wire [4-1:0] node14268;
	wire [4-1:0] node14271;
	wire [4-1:0] node14274;
	wire [4-1:0] node14275;
	wire [4-1:0] node14276;
	wire [4-1:0] node14278;
	wire [4-1:0] node14282;
	wire [4-1:0] node14283;
	wire [4-1:0] node14286;
	wire [4-1:0] node14289;
	wire [4-1:0] node14290;
	wire [4-1:0] node14291;
	wire [4-1:0] node14292;
	wire [4-1:0] node14295;
	wire [4-1:0] node14298;
	wire [4-1:0] node14300;
	wire [4-1:0] node14302;
	wire [4-1:0] node14305;
	wire [4-1:0] node14306;
	wire [4-1:0] node14309;
	wire [4-1:0] node14310;
	wire [4-1:0] node14312;
	wire [4-1:0] node14314;
	wire [4-1:0] node14318;
	wire [4-1:0] node14319;
	wire [4-1:0] node14320;
	wire [4-1:0] node14321;
	wire [4-1:0] node14322;
	wire [4-1:0] node14324;
	wire [4-1:0] node14325;
	wire [4-1:0] node14328;
	wire [4-1:0] node14331;
	wire [4-1:0] node14334;
	wire [4-1:0] node14335;
	wire [4-1:0] node14337;
	wire [4-1:0] node14341;
	wire [4-1:0] node14342;
	wire [4-1:0] node14344;
	wire [4-1:0] node14345;
	wire [4-1:0] node14346;
	wire [4-1:0] node14351;
	wire [4-1:0] node14354;
	wire [4-1:0] node14355;
	wire [4-1:0] node14356;
	wire [4-1:0] node14358;
	wire [4-1:0] node14361;
	wire [4-1:0] node14363;
	wire [4-1:0] node14365;
	wire [4-1:0] node14366;
	wire [4-1:0] node14370;
	wire [4-1:0] node14371;
	wire [4-1:0] node14372;
	wire [4-1:0] node14373;
	wire [4-1:0] node14374;
	wire [4-1:0] node14377;
	wire [4-1:0] node14380;
	wire [4-1:0] node14381;
	wire [4-1:0] node14385;
	wire [4-1:0] node14388;
	wire [4-1:0] node14390;
	wire [4-1:0] node14393;
	wire [4-1:0] node14394;
	wire [4-1:0] node14395;
	wire [4-1:0] node14396;
	wire [4-1:0] node14397;
	wire [4-1:0] node14398;
	wire [4-1:0] node14400;
	wire [4-1:0] node14403;
	wire [4-1:0] node14405;
	wire [4-1:0] node14408;
	wire [4-1:0] node14410;
	wire [4-1:0] node14412;
	wire [4-1:0] node14415;
	wire [4-1:0] node14416;
	wire [4-1:0] node14417;
	wire [4-1:0] node14421;
	wire [4-1:0] node14423;
	wire [4-1:0] node14424;
	wire [4-1:0] node14425;
	wire [4-1:0] node14428;
	wire [4-1:0] node14432;
	wire [4-1:0] node14433;
	wire [4-1:0] node14434;
	wire [4-1:0] node14435;
	wire [4-1:0] node14438;
	wire [4-1:0] node14441;
	wire [4-1:0] node14442;
	wire [4-1:0] node14444;
	wire [4-1:0] node14447;
	wire [4-1:0] node14448;
	wire [4-1:0] node14452;
	wire [4-1:0] node14453;
	wire [4-1:0] node14455;
	wire [4-1:0] node14456;
	wire [4-1:0] node14459;
	wire [4-1:0] node14461;
	wire [4-1:0] node14464;
	wire [4-1:0] node14465;
	wire [4-1:0] node14466;
	wire [4-1:0] node14467;
	wire [4-1:0] node14473;
	wire [4-1:0] node14474;
	wire [4-1:0] node14475;
	wire [4-1:0] node14476;
	wire [4-1:0] node14477;
	wire [4-1:0] node14479;
	wire [4-1:0] node14480;
	wire [4-1:0] node14483;
	wire [4-1:0] node14487;
	wire [4-1:0] node14488;
	wire [4-1:0] node14489;
	wire [4-1:0] node14492;
	wire [4-1:0] node14495;
	wire [4-1:0] node14496;
	wire [4-1:0] node14499;
	wire [4-1:0] node14502;
	wire [4-1:0] node14503;
	wire [4-1:0] node14504;
	wire [4-1:0] node14506;
	wire [4-1:0] node14509;
	wire [4-1:0] node14510;
	wire [4-1:0] node14512;
	wire [4-1:0] node14515;
	wire [4-1:0] node14517;
	wire [4-1:0] node14520;
	wire [4-1:0] node14521;
	wire [4-1:0] node14523;
	wire [4-1:0] node14526;
	wire [4-1:0] node14528;
	wire [4-1:0] node14529;
	wire [4-1:0] node14533;
	wire [4-1:0] node14534;
	wire [4-1:0] node14535;
	wire [4-1:0] node14536;
	wire [4-1:0] node14538;
	wire [4-1:0] node14540;
	wire [4-1:0] node14543;
	wire [4-1:0] node14544;
	wire [4-1:0] node14545;
	wire [4-1:0] node14549;
	wire [4-1:0] node14552;
	wire [4-1:0] node14553;
	wire [4-1:0] node14555;
	wire [4-1:0] node14559;
	wire [4-1:0] node14560;
	wire [4-1:0] node14561;
	wire [4-1:0] node14562;
	wire [4-1:0] node14566;
	wire [4-1:0] node14567;
	wire [4-1:0] node14568;
	wire [4-1:0] node14573;
	wire [4-1:0] node14575;
	wire [4-1:0] node14576;
	wire [4-1:0] node14579;
	wire [4-1:0] node14581;
	wire [4-1:0] node14584;
	wire [4-1:0] node14585;
	wire [4-1:0] node14586;
	wire [4-1:0] node14587;
	wire [4-1:0] node14588;
	wire [4-1:0] node14589;
	wire [4-1:0] node14590;
	wire [4-1:0] node14591;
	wire [4-1:0] node14594;
	wire [4-1:0] node14596;
	wire [4-1:0] node14599;
	wire [4-1:0] node14600;
	wire [4-1:0] node14601;
	wire [4-1:0] node14604;
	wire [4-1:0] node14608;
	wire [4-1:0] node14609;
	wire [4-1:0] node14610;
	wire [4-1:0] node14611;
	wire [4-1:0] node14613;
	wire [4-1:0] node14618;
	wire [4-1:0] node14619;
	wire [4-1:0] node14620;
	wire [4-1:0] node14624;
	wire [4-1:0] node14625;
	wire [4-1:0] node14626;
	wire [4-1:0] node14629;
	wire [4-1:0] node14633;
	wire [4-1:0] node14634;
	wire [4-1:0] node14635;
	wire [4-1:0] node14636;
	wire [4-1:0] node14638;
	wire [4-1:0] node14639;
	wire [4-1:0] node14643;
	wire [4-1:0] node14645;
	wire [4-1:0] node14648;
	wire [4-1:0] node14649;
	wire [4-1:0] node14650;
	wire [4-1:0] node14652;
	wire [4-1:0] node14656;
	wire [4-1:0] node14658;
	wire [4-1:0] node14661;
	wire [4-1:0] node14662;
	wire [4-1:0] node14663;
	wire [4-1:0] node14664;
	wire [4-1:0] node14667;
	wire [4-1:0] node14671;
	wire [4-1:0] node14672;
	wire [4-1:0] node14673;
	wire [4-1:0] node14674;
	wire [4-1:0] node14680;
	wire [4-1:0] node14681;
	wire [4-1:0] node14682;
	wire [4-1:0] node14683;
	wire [4-1:0] node14685;
	wire [4-1:0] node14687;
	wire [4-1:0] node14688;
	wire [4-1:0] node14692;
	wire [4-1:0] node14693;
	wire [4-1:0] node14695;
	wire [4-1:0] node14696;
	wire [4-1:0] node14699;
	wire [4-1:0] node14702;
	wire [4-1:0] node14705;
	wire [4-1:0] node14706;
	wire [4-1:0] node14708;
	wire [4-1:0] node14709;
	wire [4-1:0] node14713;
	wire [4-1:0] node14714;
	wire [4-1:0] node14716;
	wire [4-1:0] node14717;
	wire [4-1:0] node14722;
	wire [4-1:0] node14723;
	wire [4-1:0] node14724;
	wire [4-1:0] node14725;
	wire [4-1:0] node14727;
	wire [4-1:0] node14728;
	wire [4-1:0] node14732;
	wire [4-1:0] node14733;
	wire [4-1:0] node14734;
	wire [4-1:0] node14739;
	wire [4-1:0] node14740;
	wire [4-1:0] node14741;
	wire [4-1:0] node14742;
	wire [4-1:0] node14746;
	wire [4-1:0] node14750;
	wire [4-1:0] node14751;
	wire [4-1:0] node14752;
	wire [4-1:0] node14753;
	wire [4-1:0] node14758;
	wire [4-1:0] node14759;
	wire [4-1:0] node14762;
	wire [4-1:0] node14765;
	wire [4-1:0] node14766;
	wire [4-1:0] node14767;
	wire [4-1:0] node14768;
	wire [4-1:0] node14769;
	wire [4-1:0] node14770;
	wire [4-1:0] node14771;
	wire [4-1:0] node14773;
	wire [4-1:0] node14778;
	wire [4-1:0] node14779;
	wire [4-1:0] node14781;
	wire [4-1:0] node14785;
	wire [4-1:0] node14786;
	wire [4-1:0] node14787;
	wire [4-1:0] node14788;
	wire [4-1:0] node14790;
	wire [4-1:0] node14795;
	wire [4-1:0] node14796;
	wire [4-1:0] node14797;
	wire [4-1:0] node14802;
	wire [4-1:0] node14803;
	wire [4-1:0] node14804;
	wire [4-1:0] node14805;
	wire [4-1:0] node14806;
	wire [4-1:0] node14810;
	wire [4-1:0] node14812;
	wire [4-1:0] node14814;
	wire [4-1:0] node14817;
	wire [4-1:0] node14818;
	wire [4-1:0] node14819;
	wire [4-1:0] node14820;
	wire [4-1:0] node14824;
	wire [4-1:0] node14826;
	wire [4-1:0] node14830;
	wire [4-1:0] node14831;
	wire [4-1:0] node14832;
	wire [4-1:0] node14835;
	wire [4-1:0] node14837;
	wire [4-1:0] node14838;
	wire [4-1:0] node14842;
	wire [4-1:0] node14843;
	wire [4-1:0] node14844;
	wire [4-1:0] node14848;
	wire [4-1:0] node14849;
	wire [4-1:0] node14852;
	wire [4-1:0] node14854;
	wire [4-1:0] node14857;
	wire [4-1:0] node14858;
	wire [4-1:0] node14859;
	wire [4-1:0] node14860;
	wire [4-1:0] node14861;
	wire [4-1:0] node14864;
	wire [4-1:0] node14865;
	wire [4-1:0] node14869;
	wire [4-1:0] node14870;
	wire [4-1:0] node14871;
	wire [4-1:0] node14872;
	wire [4-1:0] node14876;
	wire [4-1:0] node14880;
	wire [4-1:0] node14881;
	wire [4-1:0] node14882;
	wire [4-1:0] node14883;
	wire [4-1:0] node14886;
	wire [4-1:0] node14889;
	wire [4-1:0] node14891;
	wire [4-1:0] node14892;
	wire [4-1:0] node14896;
	wire [4-1:0] node14898;
	wire [4-1:0] node14900;
	wire [4-1:0] node14903;
	wire [4-1:0] node14904;
	wire [4-1:0] node14905;
	wire [4-1:0] node14906;
	wire [4-1:0] node14907;
	wire [4-1:0] node14908;
	wire [4-1:0] node14913;
	wire [4-1:0] node14914;
	wire [4-1:0] node14918;
	wire [4-1:0] node14919;
	wire [4-1:0] node14920;
	wire [4-1:0] node14921;
	wire [4-1:0] node14927;
	wire [4-1:0] node14928;
	wire [4-1:0] node14929;
	wire [4-1:0] node14932;
	wire [4-1:0] node14935;
	wire [4-1:0] node14936;
	wire [4-1:0] node14938;
	wire [4-1:0] node14941;
	wire [4-1:0] node14943;
	wire [4-1:0] node14946;
	wire [4-1:0] node14947;
	wire [4-1:0] node14948;
	wire [4-1:0] node14949;
	wire [4-1:0] node14950;
	wire [4-1:0] node14951;
	wire [4-1:0] node14952;
	wire [4-1:0] node14953;
	wire [4-1:0] node14957;
	wire [4-1:0] node14958;
	wire [4-1:0] node14962;
	wire [4-1:0] node14964;
	wire [4-1:0] node14967;
	wire [4-1:0] node14968;
	wire [4-1:0] node14969;
	wire [4-1:0] node14970;
	wire [4-1:0] node14972;
	wire [4-1:0] node14976;
	wire [4-1:0] node14979;
	wire [4-1:0] node14980;
	wire [4-1:0] node14981;
	wire [4-1:0] node14983;
	wire [4-1:0] node14986;
	wire [4-1:0] node14988;
	wire [4-1:0] node14991;
	wire [4-1:0] node14992;
	wire [4-1:0] node14996;
	wire [4-1:0] node14997;
	wire [4-1:0] node14999;
	wire [4-1:0] node15000;
	wire [4-1:0] node15002;
	wire [4-1:0] node15005;
	wire [4-1:0] node15006;
	wire [4-1:0] node15010;
	wire [4-1:0] node15011;
	wire [4-1:0] node15012;
	wire [4-1:0] node15013;
	wire [4-1:0] node15014;
	wire [4-1:0] node15017;
	wire [4-1:0] node15022;
	wire [4-1:0] node15023;
	wire [4-1:0] node15024;
	wire [4-1:0] node15029;
	wire [4-1:0] node15030;
	wire [4-1:0] node15031;
	wire [4-1:0] node15032;
	wire [4-1:0] node15034;
	wire [4-1:0] node15036;
	wire [4-1:0] node15037;
	wire [4-1:0] node15040;
	wire [4-1:0] node15043;
	wire [4-1:0] node15045;
	wire [4-1:0] node15047;
	wire [4-1:0] node15050;
	wire [4-1:0] node15051;
	wire [4-1:0] node15052;
	wire [4-1:0] node15054;
	wire [4-1:0] node15056;
	wire [4-1:0] node15060;
	wire [4-1:0] node15061;
	wire [4-1:0] node15063;
	wire [4-1:0] node15065;
	wire [4-1:0] node15068;
	wire [4-1:0] node15069;
	wire [4-1:0] node15070;
	wire [4-1:0] node15074;
	wire [4-1:0] node15076;
	wire [4-1:0] node15079;
	wire [4-1:0] node15080;
	wire [4-1:0] node15081;
	wire [4-1:0] node15082;
	wire [4-1:0] node15084;
	wire [4-1:0] node15085;
	wire [4-1:0] node15088;
	wire [4-1:0] node15091;
	wire [4-1:0] node15094;
	wire [4-1:0] node15095;
	wire [4-1:0] node15096;
	wire [4-1:0] node15098;
	wire [4-1:0] node15101;
	wire [4-1:0] node15102;
	wire [4-1:0] node15106;
	wire [4-1:0] node15109;
	wire [4-1:0] node15110;
	wire [4-1:0] node15111;
	wire [4-1:0] node15112;
	wire [4-1:0] node15114;
	wire [4-1:0] node15118;
	wire [4-1:0] node15120;
	wire [4-1:0] node15123;
	wire [4-1:0] node15124;
	wire [4-1:0] node15126;
	wire [4-1:0] node15129;
	wire [4-1:0] node15130;
	wire [4-1:0] node15133;
	wire [4-1:0] node15136;
	wire [4-1:0] node15137;
	wire [4-1:0] node15138;
	wire [4-1:0] node15139;
	wire [4-1:0] node15140;
	wire [4-1:0] node15141;
	wire [4-1:0] node15142;
	wire [4-1:0] node15143;
	wire [4-1:0] node15148;
	wire [4-1:0] node15150;
	wire [4-1:0] node15153;
	wire [4-1:0] node15155;
	wire [4-1:0] node15157;
	wire [4-1:0] node15160;
	wire [4-1:0] node15161;
	wire [4-1:0] node15163;
	wire [4-1:0] node15166;
	wire [4-1:0] node15168;
	wire [4-1:0] node15169;
	wire [4-1:0] node15173;
	wire [4-1:0] node15174;
	wire [4-1:0] node15175;
	wire [4-1:0] node15176;
	wire [4-1:0] node15180;
	wire [4-1:0] node15182;
	wire [4-1:0] node15183;
	wire [4-1:0] node15184;
	wire [4-1:0] node15189;
	wire [4-1:0] node15190;
	wire [4-1:0] node15191;
	wire [4-1:0] node15193;
	wire [4-1:0] node15195;
	wire [4-1:0] node15198;
	wire [4-1:0] node15201;
	wire [4-1:0] node15202;
	wire [4-1:0] node15204;
	wire [4-1:0] node15207;
	wire [4-1:0] node15208;
	wire [4-1:0] node15209;
	wire [4-1:0] node15214;
	wire [4-1:0] node15215;
	wire [4-1:0] node15216;
	wire [4-1:0] node15217;
	wire [4-1:0] node15219;
	wire [4-1:0] node15221;
	wire [4-1:0] node15224;
	wire [4-1:0] node15225;
	wire [4-1:0] node15227;
	wire [4-1:0] node15230;
	wire [4-1:0] node15233;
	wire [4-1:0] node15234;
	wire [4-1:0] node15235;
	wire [4-1:0] node15237;
	wire [4-1:0] node15241;
	wire [4-1:0] node15243;
	wire [4-1:0] node15245;
	wire [4-1:0] node15248;
	wire [4-1:0] node15249;
	wire [4-1:0] node15250;
	wire [4-1:0] node15251;
	wire [4-1:0] node15252;
	wire [4-1:0] node15253;
	wire [4-1:0] node15257;
	wire [4-1:0] node15258;
	wire [4-1:0] node15262;
	wire [4-1:0] node15265;
	wire [4-1:0] node15266;
	wire [4-1:0] node15269;
	wire [4-1:0] node15271;
	wire [4-1:0] node15274;
	wire [4-1:0] node15275;
	wire [4-1:0] node15276;
	wire [4-1:0] node15280;
	wire [4-1:0] node15282;
	wire [4-1:0] node15284;
	wire [4-1:0] node15287;
	wire [4-1:0] node15288;
	wire [4-1:0] node15289;
	wire [4-1:0] node15290;
	wire [4-1:0] node15291;
	wire [4-1:0] node15292;
	wire [4-1:0] node15293;
	wire [4-1:0] node15294;
	wire [4-1:0] node15295;
	wire [4-1:0] node15297;
	wire [4-1:0] node15299;
	wire [4-1:0] node15302;
	wire [4-1:0] node15304;
	wire [4-1:0] node15305;
	wire [4-1:0] node15308;
	wire [4-1:0] node15311;
	wire [4-1:0] node15312;
	wire [4-1:0] node15313;
	wire [4-1:0] node15316;
	wire [4-1:0] node15319;
	wire [4-1:0] node15321;
	wire [4-1:0] node15324;
	wire [4-1:0] node15325;
	wire [4-1:0] node15326;
	wire [4-1:0] node15327;
	wire [4-1:0] node15328;
	wire [4-1:0] node15332;
	wire [4-1:0] node15333;
	wire [4-1:0] node15338;
	wire [4-1:0] node15339;
	wire [4-1:0] node15341;
	wire [4-1:0] node15342;
	wire [4-1:0] node15346;
	wire [4-1:0] node15349;
	wire [4-1:0] node15350;
	wire [4-1:0] node15351;
	wire [4-1:0] node15352;
	wire [4-1:0] node15353;
	wire [4-1:0] node15357;
	wire [4-1:0] node15358;
	wire [4-1:0] node15359;
	wire [4-1:0] node15363;
	wire [4-1:0] node15366;
	wire [4-1:0] node15367;
	wire [4-1:0] node15369;
	wire [4-1:0] node15372;
	wire [4-1:0] node15373;
	wire [4-1:0] node15377;
	wire [4-1:0] node15378;
	wire [4-1:0] node15379;
	wire [4-1:0] node15380;
	wire [4-1:0] node15382;
	wire [4-1:0] node15385;
	wire [4-1:0] node15387;
	wire [4-1:0] node15390;
	wire [4-1:0] node15393;
	wire [4-1:0] node15394;
	wire [4-1:0] node15396;
	wire [4-1:0] node15400;
	wire [4-1:0] node15401;
	wire [4-1:0] node15402;
	wire [4-1:0] node15403;
	wire [4-1:0] node15404;
	wire [4-1:0] node15406;
	wire [4-1:0] node15409;
	wire [4-1:0] node15410;
	wire [4-1:0] node15413;
	wire [4-1:0] node15415;
	wire [4-1:0] node15418;
	wire [4-1:0] node15421;
	wire [4-1:0] node15422;
	wire [4-1:0] node15424;
	wire [4-1:0] node15425;
	wire [4-1:0] node15429;
	wire [4-1:0] node15430;
	wire [4-1:0] node15433;
	wire [4-1:0] node15435;
	wire [4-1:0] node15437;
	wire [4-1:0] node15440;
	wire [4-1:0] node15441;
	wire [4-1:0] node15442;
	wire [4-1:0] node15443;
	wire [4-1:0] node15444;
	wire [4-1:0] node15448;
	wire [4-1:0] node15450;
	wire [4-1:0] node15453;
	wire [4-1:0] node15454;
	wire [4-1:0] node15455;
	wire [4-1:0] node15458;
	wire [4-1:0] node15461;
	wire [4-1:0] node15463;
	wire [4-1:0] node15466;
	wire [4-1:0] node15467;
	wire [4-1:0] node15469;
	wire [4-1:0] node15470;
	wire [4-1:0] node15474;
	wire [4-1:0] node15476;
	wire [4-1:0] node15477;
	wire [4-1:0] node15478;
	wire [4-1:0] node15481;
	wire [4-1:0] node15485;
	wire [4-1:0] node15486;
	wire [4-1:0] node15487;
	wire [4-1:0] node15488;
	wire [4-1:0] node15489;
	wire [4-1:0] node15490;
	wire [4-1:0] node15491;
	wire [4-1:0] node15493;
	wire [4-1:0] node15497;
	wire [4-1:0] node15498;
	wire [4-1:0] node15502;
	wire [4-1:0] node15503;
	wire [4-1:0] node15506;
	wire [4-1:0] node15509;
	wire [4-1:0] node15510;
	wire [4-1:0] node15512;
	wire [4-1:0] node15514;
	wire [4-1:0] node15515;
	wire [4-1:0] node15519;
	wire [4-1:0] node15522;
	wire [4-1:0] node15523;
	wire [4-1:0] node15524;
	wire [4-1:0] node15525;
	wire [4-1:0] node15527;
	wire [4-1:0] node15530;
	wire [4-1:0] node15531;
	wire [4-1:0] node15534;
	wire [4-1:0] node15535;
	wire [4-1:0] node15539;
	wire [4-1:0] node15541;
	wire [4-1:0] node15544;
	wire [4-1:0] node15545;
	wire [4-1:0] node15546;
	wire [4-1:0] node15550;
	wire [4-1:0] node15553;
	wire [4-1:0] node15554;
	wire [4-1:0] node15555;
	wire [4-1:0] node15556;
	wire [4-1:0] node15557;
	wire [4-1:0] node15561;
	wire [4-1:0] node15562;
	wire [4-1:0] node15563;
	wire [4-1:0] node15567;
	wire [4-1:0] node15569;
	wire [4-1:0] node15570;
	wire [4-1:0] node15574;
	wire [4-1:0] node15575;
	wire [4-1:0] node15576;
	wire [4-1:0] node15578;
	wire [4-1:0] node15582;
	wire [4-1:0] node15583;
	wire [4-1:0] node15584;
	wire [4-1:0] node15587;
	wire [4-1:0] node15589;
	wire [4-1:0] node15592;
	wire [4-1:0] node15594;
	wire [4-1:0] node15596;
	wire [4-1:0] node15599;
	wire [4-1:0] node15600;
	wire [4-1:0] node15601;
	wire [4-1:0] node15602;
	wire [4-1:0] node15604;
	wire [4-1:0] node15605;
	wire [4-1:0] node15608;
	wire [4-1:0] node15612;
	wire [4-1:0] node15613;
	wire [4-1:0] node15614;
	wire [4-1:0] node15619;
	wire [4-1:0] node15620;
	wire [4-1:0] node15622;
	wire [4-1:0] node15624;
	wire [4-1:0] node15625;
	wire [4-1:0] node15629;
	wire [4-1:0] node15630;
	wire [4-1:0] node15633;
	wire [4-1:0] node15634;
	wire [4-1:0] node15635;
	wire [4-1:0] node15640;
	wire [4-1:0] node15641;
	wire [4-1:0] node15642;
	wire [4-1:0] node15643;
	wire [4-1:0] node15644;
	wire [4-1:0] node15645;
	wire [4-1:0] node15646;
	wire [4-1:0] node15648;
	wire [4-1:0] node15649;
	wire [4-1:0] node15653;
	wire [4-1:0] node15655;
	wire [4-1:0] node15656;
	wire [4-1:0] node15660;
	wire [4-1:0] node15661;
	wire [4-1:0] node15663;
	wire [4-1:0] node15667;
	wire [4-1:0] node15668;
	wire [4-1:0] node15669;
	wire [4-1:0] node15670;
	wire [4-1:0] node15673;
	wire [4-1:0] node15676;
	wire [4-1:0] node15677;
	wire [4-1:0] node15678;
	wire [4-1:0] node15682;
	wire [4-1:0] node15685;
	wire [4-1:0] node15686;
	wire [4-1:0] node15687;
	wire [4-1:0] node15690;
	wire [4-1:0] node15693;
	wire [4-1:0] node15694;
	wire [4-1:0] node15698;
	wire [4-1:0] node15699;
	wire [4-1:0] node15700;
	wire [4-1:0] node15702;
	wire [4-1:0] node15705;
	wire [4-1:0] node15707;
	wire [4-1:0] node15709;
	wire [4-1:0] node15712;
	wire [4-1:0] node15713;
	wire [4-1:0] node15715;
	wire [4-1:0] node15717;
	wire [4-1:0] node15720;
	wire [4-1:0] node15721;
	wire [4-1:0] node15725;
	wire [4-1:0] node15726;
	wire [4-1:0] node15727;
	wire [4-1:0] node15730;
	wire [4-1:0] node15731;
	wire [4-1:0] node15733;
	wire [4-1:0] node15734;
	wire [4-1:0] node15738;
	wire [4-1:0] node15740;
	wire [4-1:0] node15741;
	wire [4-1:0] node15744;
	wire [4-1:0] node15747;
	wire [4-1:0] node15748;
	wire [4-1:0] node15749;
	wire [4-1:0] node15750;
	wire [4-1:0] node15752;
	wire [4-1:0] node15753;
	wire [4-1:0] node15757;
	wire [4-1:0] node15760;
	wire [4-1:0] node15761;
	wire [4-1:0] node15762;
	wire [4-1:0] node15763;
	wire [4-1:0] node15766;
	wire [4-1:0] node15770;
	wire [4-1:0] node15771;
	wire [4-1:0] node15772;
	wire [4-1:0] node15776;
	wire [4-1:0] node15777;
	wire [4-1:0] node15781;
	wire [4-1:0] node15782;
	wire [4-1:0] node15783;
	wire [4-1:0] node15784;
	wire [4-1:0] node15786;
	wire [4-1:0] node15790;
	wire [4-1:0] node15793;
	wire [4-1:0] node15794;
	wire [4-1:0] node15795;
	wire [4-1:0] node15796;
	wire [4-1:0] node15801;
	wire [4-1:0] node15803;
	wire [4-1:0] node15806;
	wire [4-1:0] node15807;
	wire [4-1:0] node15808;
	wire [4-1:0] node15809;
	wire [4-1:0] node15810;
	wire [4-1:0] node15811;
	wire [4-1:0] node15812;
	wire [4-1:0] node15813;
	wire [4-1:0] node15816;
	wire [4-1:0] node15820;
	wire [4-1:0] node15821;
	wire [4-1:0] node15824;
	wire [4-1:0] node15827;
	wire [4-1:0] node15829;
	wire [4-1:0] node15831;
	wire [4-1:0] node15834;
	wire [4-1:0] node15835;
	wire [4-1:0] node15836;
	wire [4-1:0] node15838;
	wire [4-1:0] node15841;
	wire [4-1:0] node15844;
	wire [4-1:0] node15845;
	wire [4-1:0] node15847;
	wire [4-1:0] node15848;
	wire [4-1:0] node15851;
	wire [4-1:0] node15855;
	wire [4-1:0] node15856;
	wire [4-1:0] node15857;
	wire [4-1:0] node15858;
	wire [4-1:0] node15861;
	wire [4-1:0] node15864;
	wire [4-1:0] node15865;
	wire [4-1:0] node15868;
	wire [4-1:0] node15871;
	wire [4-1:0] node15872;
	wire [4-1:0] node15873;
	wire [4-1:0] node15876;
	wire [4-1:0] node15879;
	wire [4-1:0] node15881;
	wire [4-1:0] node15884;
	wire [4-1:0] node15885;
	wire [4-1:0] node15886;
	wire [4-1:0] node15887;
	wire [4-1:0] node15888;
	wire [4-1:0] node15890;
	wire [4-1:0] node15892;
	wire [4-1:0] node15895;
	wire [4-1:0] node15898;
	wire [4-1:0] node15900;
	wire [4-1:0] node15903;
	wire [4-1:0] node15905;
	wire [4-1:0] node15906;
	wire [4-1:0] node15908;
	wire [4-1:0] node15911;
	wire [4-1:0] node15912;
	wire [4-1:0] node15915;
	wire [4-1:0] node15917;
	wire [4-1:0] node15920;
	wire [4-1:0] node15921;
	wire [4-1:0] node15922;
	wire [4-1:0] node15923;
	wire [4-1:0] node15927;
	wire [4-1:0] node15928;
	wire [4-1:0] node15932;
	wire [4-1:0] node15933;
	wire [4-1:0] node15934;
	wire [4-1:0] node15937;
	wire [4-1:0] node15940;
	wire [4-1:0] node15942;
	wire [4-1:0] node15945;
	wire [4-1:0] node15946;
	wire [4-1:0] node15947;
	wire [4-1:0] node15948;
	wire [4-1:0] node15949;
	wire [4-1:0] node15950;
	wire [4-1:0] node15951;
	wire [4-1:0] node15952;
	wire [4-1:0] node15954;
	wire [4-1:0] node15957;
	wire [4-1:0] node15959;
	wire [4-1:0] node15960;
	wire [4-1:0] node15964;
	wire [4-1:0] node15965;
	wire [4-1:0] node15966;
	wire [4-1:0] node15969;
	wire [4-1:0] node15973;
	wire [4-1:0] node15974;
	wire [4-1:0] node15976;
	wire [4-1:0] node15978;
	wire [4-1:0] node15981;
	wire [4-1:0] node15982;
	wire [4-1:0] node15986;
	wire [4-1:0] node15987;
	wire [4-1:0] node15988;
	wire [4-1:0] node15989;
	wire [4-1:0] node15991;
	wire [4-1:0] node15992;
	wire [4-1:0] node15996;
	wire [4-1:0] node15999;
	wire [4-1:0] node16000;
	wire [4-1:0] node16001;
	wire [4-1:0] node16005;
	wire [4-1:0] node16007;
	wire [4-1:0] node16010;
	wire [4-1:0] node16011;
	wire [4-1:0] node16013;
	wire [4-1:0] node16015;
	wire [4-1:0] node16017;
	wire [4-1:0] node16020;
	wire [4-1:0] node16021;
	wire [4-1:0] node16024;
	wire [4-1:0] node16025;
	wire [4-1:0] node16027;
	wire [4-1:0] node16031;
	wire [4-1:0] node16032;
	wire [4-1:0] node16033;
	wire [4-1:0] node16034;
	wire [4-1:0] node16035;
	wire [4-1:0] node16036;
	wire [4-1:0] node16039;
	wire [4-1:0] node16040;
	wire [4-1:0] node16043;
	wire [4-1:0] node16046;
	wire [4-1:0] node16047;
	wire [4-1:0] node16048;
	wire [4-1:0] node16053;
	wire [4-1:0] node16054;
	wire [4-1:0] node16055;
	wire [4-1:0] node16057;
	wire [4-1:0] node16060;
	wire [4-1:0] node16063;
	wire [4-1:0] node16064;
	wire [4-1:0] node16066;
	wire [4-1:0] node16069;
	wire [4-1:0] node16072;
	wire [4-1:0] node16073;
	wire [4-1:0] node16074;
	wire [4-1:0] node16075;
	wire [4-1:0] node16078;
	wire [4-1:0] node16081;
	wire [4-1:0] node16084;
	wire [4-1:0] node16085;
	wire [4-1:0] node16086;
	wire [4-1:0] node16091;
	wire [4-1:0] node16092;
	wire [4-1:0] node16093;
	wire [4-1:0] node16094;
	wire [4-1:0] node16096;
	wire [4-1:0] node16098;
	wire [4-1:0] node16101;
	wire [4-1:0] node16103;
	wire [4-1:0] node16105;
	wire [4-1:0] node16108;
	wire [4-1:0] node16109;
	wire [4-1:0] node16110;
	wire [4-1:0] node16114;
	wire [4-1:0] node16116;
	wire [4-1:0] node16119;
	wire [4-1:0] node16120;
	wire [4-1:0] node16121;
	wire [4-1:0] node16123;
	wire [4-1:0] node16125;
	wire [4-1:0] node16128;
	wire [4-1:0] node16131;
	wire [4-1:0] node16132;
	wire [4-1:0] node16135;
	wire [4-1:0] node16137;
	wire [4-1:0] node16139;
	wire [4-1:0] node16142;
	wire [4-1:0] node16143;
	wire [4-1:0] node16144;
	wire [4-1:0] node16145;
	wire [4-1:0] node16146;
	wire [4-1:0] node16147;
	wire [4-1:0] node16148;
	wire [4-1:0] node16149;
	wire [4-1:0] node16155;
	wire [4-1:0] node16156;
	wire [4-1:0] node16157;
	wire [4-1:0] node16158;
	wire [4-1:0] node16161;
	wire [4-1:0] node16165;
	wire [4-1:0] node16167;
	wire [4-1:0] node16170;
	wire [4-1:0] node16171;
	wire [4-1:0] node16172;
	wire [4-1:0] node16173;
	wire [4-1:0] node16174;
	wire [4-1:0] node16178;
	wire [4-1:0] node16179;
	wire [4-1:0] node16183;
	wire [4-1:0] node16186;
	wire [4-1:0] node16187;
	wire [4-1:0] node16188;
	wire [4-1:0] node16193;
	wire [4-1:0] node16194;
	wire [4-1:0] node16195;
	wire [4-1:0] node16196;
	wire [4-1:0] node16198;
	wire [4-1:0] node16199;
	wire [4-1:0] node16203;
	wire [4-1:0] node16206;
	wire [4-1:0] node16207;
	wire [4-1:0] node16211;
	wire [4-1:0] node16212;
	wire [4-1:0] node16213;
	wire [4-1:0] node16216;
	wire [4-1:0] node16217;
	wire [4-1:0] node16219;
	wire [4-1:0] node16223;
	wire [4-1:0] node16224;
	wire [4-1:0] node16225;
	wire [4-1:0] node16229;
	wire [4-1:0] node16232;
	wire [4-1:0] node16233;
	wire [4-1:0] node16234;
	wire [4-1:0] node16235;
	wire [4-1:0] node16236;
	wire [4-1:0] node16239;
	wire [4-1:0] node16240;
	wire [4-1:0] node16241;
	wire [4-1:0] node16246;
	wire [4-1:0] node16247;
	wire [4-1:0] node16248;
	wire [4-1:0] node16251;
	wire [4-1:0] node16255;
	wire [4-1:0] node16256;
	wire [4-1:0] node16257;
	wire [4-1:0] node16258;
	wire [4-1:0] node16260;
	wire [4-1:0] node16263;
	wire [4-1:0] node16264;
	wire [4-1:0] node16267;
	wire [4-1:0] node16270;
	wire [4-1:0] node16272;
	wire [4-1:0] node16275;
	wire [4-1:0] node16278;
	wire [4-1:0] node16279;
	wire [4-1:0] node16280;
	wire [4-1:0] node16282;
	wire [4-1:0] node16284;
	wire [4-1:0] node16285;
	wire [4-1:0] node16289;
	wire [4-1:0] node16290;
	wire [4-1:0] node16291;
	wire [4-1:0] node16295;
	wire [4-1:0] node16296;
	wire [4-1:0] node16298;
	wire [4-1:0] node16301;
	wire [4-1:0] node16304;
	wire [4-1:0] node16305;
	wire [4-1:0] node16306;
	wire [4-1:0] node16307;
	wire [4-1:0] node16309;
	wire [4-1:0] node16313;
	wire [4-1:0] node16316;
	wire [4-1:0] node16317;
	wire [4-1:0] node16318;
	wire [4-1:0] node16319;
	wire [4-1:0] node16325;
	wire [4-1:0] node16326;
	wire [4-1:0] node16327;
	wire [4-1:0] node16328;
	wire [4-1:0] node16329;
	wire [4-1:0] node16330;
	wire [4-1:0] node16331;
	wire [4-1:0] node16332;
	wire [4-1:0] node16336;
	wire [4-1:0] node16339;
	wire [4-1:0] node16341;
	wire [4-1:0] node16344;
	wire [4-1:0] node16345;
	wire [4-1:0] node16346;
	wire [4-1:0] node16350;
	wire [4-1:0] node16351;
	wire [4-1:0] node16352;
	wire [4-1:0] node16354;
	wire [4-1:0] node16359;
	wire [4-1:0] node16360;
	wire [4-1:0] node16361;
	wire [4-1:0] node16362;
	wire [4-1:0] node16363;
	wire [4-1:0] node16364;
	wire [4-1:0] node16367;
	wire [4-1:0] node16371;
	wire [4-1:0] node16373;
	wire [4-1:0] node16374;
	wire [4-1:0] node16378;
	wire [4-1:0] node16379;
	wire [4-1:0] node16380;
	wire [4-1:0] node16384;
	wire [4-1:0] node16385;
	wire [4-1:0] node16389;
	wire [4-1:0] node16390;
	wire [4-1:0] node16391;
	wire [4-1:0] node16392;
	wire [4-1:0] node16393;
	wire [4-1:0] node16397;
	wire [4-1:0] node16400;
	wire [4-1:0] node16401;
	wire [4-1:0] node16405;
	wire [4-1:0] node16406;
	wire [4-1:0] node16408;
	wire [4-1:0] node16410;
	wire [4-1:0] node16413;
	wire [4-1:0] node16414;
	wire [4-1:0] node16417;
	wire [4-1:0] node16420;
	wire [4-1:0] node16421;
	wire [4-1:0] node16422;
	wire [4-1:0] node16423;
	wire [4-1:0] node16424;
	wire [4-1:0] node16426;
	wire [4-1:0] node16427;
	wire [4-1:0] node16432;
	wire [4-1:0] node16433;
	wire [4-1:0] node16436;
	wire [4-1:0] node16437;
	wire [4-1:0] node16440;
	wire [4-1:0] node16443;
	wire [4-1:0] node16444;
	wire [4-1:0] node16445;
	wire [4-1:0] node16446;
	wire [4-1:0] node16447;
	wire [4-1:0] node16452;
	wire [4-1:0] node16453;
	wire [4-1:0] node16457;
	wire [4-1:0] node16458;
	wire [4-1:0] node16459;
	wire [4-1:0] node16462;
	wire [4-1:0] node16464;
	wire [4-1:0] node16467;
	wire [4-1:0] node16468;
	wire [4-1:0] node16471;
	wire [4-1:0] node16473;
	wire [4-1:0] node16476;
	wire [4-1:0] node16477;
	wire [4-1:0] node16478;
	wire [4-1:0] node16480;
	wire [4-1:0] node16482;
	wire [4-1:0] node16483;
	wire [4-1:0] node16487;
	wire [4-1:0] node16489;
	wire [4-1:0] node16491;
	wire [4-1:0] node16493;
	wire [4-1:0] node16496;
	wire [4-1:0] node16497;
	wire [4-1:0] node16498;
	wire [4-1:0] node16499;
	wire [4-1:0] node16503;
	wire [4-1:0] node16506;
	wire [4-1:0] node16507;
	wire [4-1:0] node16510;
	wire [4-1:0] node16513;
	wire [4-1:0] node16514;
	wire [4-1:0] node16515;
	wire [4-1:0] node16516;
	wire [4-1:0] node16517;
	wire [4-1:0] node16518;
	wire [4-1:0] node16521;
	wire [4-1:0] node16522;
	wire [4-1:0] node16526;
	wire [4-1:0] node16527;
	wire [4-1:0] node16531;
	wire [4-1:0] node16532;
	wire [4-1:0] node16533;
	wire [4-1:0] node16535;
	wire [4-1:0] node16539;
	wire [4-1:0] node16540;
	wire [4-1:0] node16541;
	wire [4-1:0] node16543;
	wire [4-1:0] node16548;
	wire [4-1:0] node16549;
	wire [4-1:0] node16550;
	wire [4-1:0] node16551;
	wire [4-1:0] node16553;
	wire [4-1:0] node16554;
	wire [4-1:0] node16558;
	wire [4-1:0] node16559;
	wire [4-1:0] node16563;
	wire [4-1:0] node16565;
	wire [4-1:0] node16566;
	wire [4-1:0] node16567;
	wire [4-1:0] node16572;
	wire [4-1:0] node16573;
	wire [4-1:0] node16574;
	wire [4-1:0] node16575;
	wire [4-1:0] node16578;
	wire [4-1:0] node16579;
	wire [4-1:0] node16584;
	wire [4-1:0] node16586;
	wire [4-1:0] node16587;
	wire [4-1:0] node16588;
	wire [4-1:0] node16593;
	wire [4-1:0] node16594;
	wire [4-1:0] node16595;
	wire [4-1:0] node16596;
	wire [4-1:0] node16597;
	wire [4-1:0] node16598;
	wire [4-1:0] node16600;
	wire [4-1:0] node16604;
	wire [4-1:0] node16607;
	wire [4-1:0] node16608;
	wire [4-1:0] node16610;
	wire [4-1:0] node16613;
	wire [4-1:0] node16615;
	wire [4-1:0] node16618;
	wire [4-1:0] node16619;
	wire [4-1:0] node16620;
	wire [4-1:0] node16621;
	wire [4-1:0] node16625;
	wire [4-1:0] node16627;
	wire [4-1:0] node16629;
	wire [4-1:0] node16632;
	wire [4-1:0] node16633;
	wire [4-1:0] node16634;
	wire [4-1:0] node16636;
	wire [4-1:0] node16640;
	wire [4-1:0] node16641;
	wire [4-1:0] node16643;
	wire [4-1:0] node16647;
	wire [4-1:0] node16648;
	wire [4-1:0] node16649;
	wire [4-1:0] node16650;
	wire [4-1:0] node16653;
	wire [4-1:0] node16655;
	wire [4-1:0] node16658;
	wire [4-1:0] node16659;
	wire [4-1:0] node16661;
	wire [4-1:0] node16664;
	wire [4-1:0] node16665;
	wire [4-1:0] node16666;
	wire [4-1:0] node16671;
	wire [4-1:0] node16672;
	wire [4-1:0] node16675;
	wire [4-1:0] node16676;
	wire [4-1:0] node16679;
	wire [4-1:0] node16680;
	wire [4-1:0] node16684;
	wire [4-1:0] node16685;
	wire [4-1:0] node16686;
	wire [4-1:0] node16687;
	wire [4-1:0] node16688;
	wire [4-1:0] node16689;
	wire [4-1:0] node16690;
	wire [4-1:0] node16691;
	wire [4-1:0] node16692;
	wire [4-1:0] node16693;
	wire [4-1:0] node16695;
	wire [4-1:0] node16697;
	wire [4-1:0] node16700;
	wire [4-1:0] node16701;
	wire [4-1:0] node16702;
	wire [4-1:0] node16704;
	wire [4-1:0] node16707;
	wire [4-1:0] node16710;
	wire [4-1:0] node16713;
	wire [4-1:0] node16714;
	wire [4-1:0] node16715;
	wire [4-1:0] node16718;
	wire [4-1:0] node16721;
	wire [4-1:0] node16722;
	wire [4-1:0] node16723;
	wire [4-1:0] node16724;
	wire [4-1:0] node16727;
	wire [4-1:0] node16732;
	wire [4-1:0] node16733;
	wire [4-1:0] node16734;
	wire [4-1:0] node16735;
	wire [4-1:0] node16736;
	wire [4-1:0] node16739;
	wire [4-1:0] node16742;
	wire [4-1:0] node16743;
	wire [4-1:0] node16745;
	wire [4-1:0] node16749;
	wire [4-1:0] node16750;
	wire [4-1:0] node16751;
	wire [4-1:0] node16752;
	wire [4-1:0] node16757;
	wire [4-1:0] node16758;
	wire [4-1:0] node16762;
	wire [4-1:0] node16763;
	wire [4-1:0] node16764;
	wire [4-1:0] node16766;
	wire [4-1:0] node16768;
	wire [4-1:0] node16771;
	wire [4-1:0] node16773;
	wire [4-1:0] node16775;
	wire [4-1:0] node16778;
	wire [4-1:0] node16780;
	wire [4-1:0] node16781;
	wire [4-1:0] node16785;
	wire [4-1:0] node16786;
	wire [4-1:0] node16787;
	wire [4-1:0] node16788;
	wire [4-1:0] node16789;
	wire [4-1:0] node16790;
	wire [4-1:0] node16794;
	wire [4-1:0] node16796;
	wire [4-1:0] node16797;
	wire [4-1:0] node16802;
	wire [4-1:0] node16804;
	wire [4-1:0] node16805;
	wire [4-1:0] node16807;
	wire [4-1:0] node16811;
	wire [4-1:0] node16812;
	wire [4-1:0] node16813;
	wire [4-1:0] node16815;
	wire [4-1:0] node16818;
	wire [4-1:0] node16819;
	wire [4-1:0] node16820;
	wire [4-1:0] node16821;
	wire [4-1:0] node16824;
	wire [4-1:0] node16829;
	wire [4-1:0] node16830;
	wire [4-1:0] node16831;
	wire [4-1:0] node16833;
	wire [4-1:0] node16834;
	wire [4-1:0] node16838;
	wire [4-1:0] node16840;
	wire [4-1:0] node16843;
	wire [4-1:0] node16845;
	wire [4-1:0] node16847;
	wire [4-1:0] node16849;
	wire [4-1:0] node16852;
	wire [4-1:0] node16853;
	wire [4-1:0] node16854;
	wire [4-1:0] node16855;
	wire [4-1:0] node16856;
	wire [4-1:0] node16857;
	wire [4-1:0] node16859;
	wire [4-1:0] node16861;
	wire [4-1:0] node16864;
	wire [4-1:0] node16865;
	wire [4-1:0] node16869;
	wire [4-1:0] node16871;
	wire [4-1:0] node16872;
	wire [4-1:0] node16873;
	wire [4-1:0] node16878;
	wire [4-1:0] node16879;
	wire [4-1:0] node16881;
	wire [4-1:0] node16883;
	wire [4-1:0] node16884;
	wire [4-1:0] node16887;
	wire [4-1:0] node16890;
	wire [4-1:0] node16891;
	wire [4-1:0] node16892;
	wire [4-1:0] node16897;
	wire [4-1:0] node16898;
	wire [4-1:0] node16899;
	wire [4-1:0] node16900;
	wire [4-1:0] node16901;
	wire [4-1:0] node16902;
	wire [4-1:0] node16907;
	wire [4-1:0] node16910;
	wire [4-1:0] node16911;
	wire [4-1:0] node16912;
	wire [4-1:0] node16913;
	wire [4-1:0] node16917;
	wire [4-1:0] node16920;
	wire [4-1:0] node16922;
	wire [4-1:0] node16925;
	wire [4-1:0] node16926;
	wire [4-1:0] node16927;
	wire [4-1:0] node16929;
	wire [4-1:0] node16931;
	wire [4-1:0] node16935;
	wire [4-1:0] node16936;
	wire [4-1:0] node16937;
	wire [4-1:0] node16940;
	wire [4-1:0] node16943;
	wire [4-1:0] node16945;
	wire [4-1:0] node16948;
	wire [4-1:0] node16949;
	wire [4-1:0] node16950;
	wire [4-1:0] node16951;
	wire [4-1:0] node16952;
	wire [4-1:0] node16955;
	wire [4-1:0] node16956;
	wire [4-1:0] node16960;
	wire [4-1:0] node16962;
	wire [4-1:0] node16965;
	wire [4-1:0] node16966;
	wire [4-1:0] node16967;
	wire [4-1:0] node16969;
	wire [4-1:0] node16970;
	wire [4-1:0] node16975;
	wire [4-1:0] node16976;
	wire [4-1:0] node16977;
	wire [4-1:0] node16981;
	wire [4-1:0] node16982;
	wire [4-1:0] node16986;
	wire [4-1:0] node16987;
	wire [4-1:0] node16988;
	wire [4-1:0] node16989;
	wire [4-1:0] node16990;
	wire [4-1:0] node16993;
	wire [4-1:0] node16994;
	wire [4-1:0] node16998;
	wire [4-1:0] node16999;
	wire [4-1:0] node17003;
	wire [4-1:0] node17004;
	wire [4-1:0] node17005;
	wire [4-1:0] node17008;
	wire [4-1:0] node17012;
	wire [4-1:0] node17013;
	wire [4-1:0] node17014;
	wire [4-1:0] node17016;
	wire [4-1:0] node17017;
	wire [4-1:0] node17020;
	wire [4-1:0] node17023;
	wire [4-1:0] node17026;
	wire [4-1:0] node17027;
	wire [4-1:0] node17030;
	wire [4-1:0] node17033;
	wire [4-1:0] node17034;
	wire [4-1:0] node17035;
	wire [4-1:0] node17036;
	wire [4-1:0] node17037;
	wire [4-1:0] node17038;
	wire [4-1:0] node17039;
	wire [4-1:0] node17040;
	wire [4-1:0] node17044;
	wire [4-1:0] node17045;
	wire [4-1:0] node17048;
	wire [4-1:0] node17051;
	wire [4-1:0] node17054;
	wire [4-1:0] node17055;
	wire [4-1:0] node17056;
	wire [4-1:0] node17057;
	wire [4-1:0] node17058;
	wire [4-1:0] node17062;
	wire [4-1:0] node17064;
	wire [4-1:0] node17068;
	wire [4-1:0] node17069;
	wire [4-1:0] node17070;
	wire [4-1:0] node17073;
	wire [4-1:0] node17076;
	wire [4-1:0] node17077;
	wire [4-1:0] node17079;
	wire [4-1:0] node17083;
	wire [4-1:0] node17084;
	wire [4-1:0] node17085;
	wire [4-1:0] node17086;
	wire [4-1:0] node17089;
	wire [4-1:0] node17090;
	wire [4-1:0] node17091;
	wire [4-1:0] node17096;
	wire [4-1:0] node17097;
	wire [4-1:0] node17099;
	wire [4-1:0] node17100;
	wire [4-1:0] node17104;
	wire [4-1:0] node17105;
	wire [4-1:0] node17109;
	wire [4-1:0] node17110;
	wire [4-1:0] node17111;
	wire [4-1:0] node17115;
	wire [4-1:0] node17116;
	wire [4-1:0] node17117;
	wire [4-1:0] node17119;
	wire [4-1:0] node17123;
	wire [4-1:0] node17124;
	wire [4-1:0] node17128;
	wire [4-1:0] node17129;
	wire [4-1:0] node17130;
	wire [4-1:0] node17131;
	wire [4-1:0] node17132;
	wire [4-1:0] node17133;
	wire [4-1:0] node17134;
	wire [4-1:0] node17140;
	wire [4-1:0] node17141;
	wire [4-1:0] node17142;
	wire [4-1:0] node17146;
	wire [4-1:0] node17148;
	wire [4-1:0] node17151;
	wire [4-1:0] node17152;
	wire [4-1:0] node17153;
	wire [4-1:0] node17155;
	wire [4-1:0] node17159;
	wire [4-1:0] node17160;
	wire [4-1:0] node17162;
	wire [4-1:0] node17164;
	wire [4-1:0] node17168;
	wire [4-1:0] node17169;
	wire [4-1:0] node17170;
	wire [4-1:0] node17171;
	wire [4-1:0] node17173;
	wire [4-1:0] node17175;
	wire [4-1:0] node17179;
	wire [4-1:0] node17180;
	wire [4-1:0] node17181;
	wire [4-1:0] node17185;
	wire [4-1:0] node17187;
	wire [4-1:0] node17189;
	wire [4-1:0] node17192;
	wire [4-1:0] node17193;
	wire [4-1:0] node17194;
	wire [4-1:0] node17195;
	wire [4-1:0] node17200;
	wire [4-1:0] node17201;
	wire [4-1:0] node17205;
	wire [4-1:0] node17206;
	wire [4-1:0] node17207;
	wire [4-1:0] node17208;
	wire [4-1:0] node17209;
	wire [4-1:0] node17210;
	wire [4-1:0] node17211;
	wire [4-1:0] node17215;
	wire [4-1:0] node17218;
	wire [4-1:0] node17219;
	wire [4-1:0] node17220;
	wire [4-1:0] node17221;
	wire [4-1:0] node17227;
	wire [4-1:0] node17228;
	wire [4-1:0] node17229;
	wire [4-1:0] node17231;
	wire [4-1:0] node17234;
	wire [4-1:0] node17235;
	wire [4-1:0] node17237;
	wire [4-1:0] node17241;
	wire [4-1:0] node17243;
	wire [4-1:0] node17246;
	wire [4-1:0] node17247;
	wire [4-1:0] node17248;
	wire [4-1:0] node17250;
	wire [4-1:0] node17253;
	wire [4-1:0] node17254;
	wire [4-1:0] node17255;
	wire [4-1:0] node17258;
	wire [4-1:0] node17261;
	wire [4-1:0] node17263;
	wire [4-1:0] node17266;
	wire [4-1:0] node17267;
	wire [4-1:0] node17269;
	wire [4-1:0] node17272;
	wire [4-1:0] node17273;
	wire [4-1:0] node17276;
	wire [4-1:0] node17279;
	wire [4-1:0] node17280;
	wire [4-1:0] node17281;
	wire [4-1:0] node17282;
	wire [4-1:0] node17283;
	wire [4-1:0] node17284;
	wire [4-1:0] node17286;
	wire [4-1:0] node17290;
	wire [4-1:0] node17291;
	wire [4-1:0] node17295;
	wire [4-1:0] node17297;
	wire [4-1:0] node17299;
	wire [4-1:0] node17302;
	wire [4-1:0] node17303;
	wire [4-1:0] node17304;
	wire [4-1:0] node17305;
	wire [4-1:0] node17309;
	wire [4-1:0] node17312;
	wire [4-1:0] node17314;
	wire [4-1:0] node17315;
	wire [4-1:0] node17319;
	wire [4-1:0] node17320;
	wire [4-1:0] node17321;
	wire [4-1:0] node17322;
	wire [4-1:0] node17323;
	wire [4-1:0] node17326;
	wire [4-1:0] node17328;
	wire [4-1:0] node17331;
	wire [4-1:0] node17334;
	wire [4-1:0] node17335;
	wire [4-1:0] node17336;
	wire [4-1:0] node17340;
	wire [4-1:0] node17342;
	wire [4-1:0] node17345;
	wire [4-1:0] node17346;
	wire [4-1:0] node17348;
	wire [4-1:0] node17349;
	wire [4-1:0] node17352;
	wire [4-1:0] node17355;
	wire [4-1:0] node17356;
	wire [4-1:0] node17360;
	wire [4-1:0] node17361;
	wire [4-1:0] node17362;
	wire [4-1:0] node17363;
	wire [4-1:0] node17364;
	wire [4-1:0] node17365;
	wire [4-1:0] node17366;
	wire [4-1:0] node17367;
	wire [4-1:0] node17369;
	wire [4-1:0] node17371;
	wire [4-1:0] node17374;
	wire [4-1:0] node17376;
	wire [4-1:0] node17377;
	wire [4-1:0] node17381;
	wire [4-1:0] node17383;
	wire [4-1:0] node17386;
	wire [4-1:0] node17387;
	wire [4-1:0] node17388;
	wire [4-1:0] node17389;
	wire [4-1:0] node17391;
	wire [4-1:0] node17394;
	wire [4-1:0] node17395;
	wire [4-1:0] node17399;
	wire [4-1:0] node17401;
	wire [4-1:0] node17404;
	wire [4-1:0] node17405;
	wire [4-1:0] node17406;
	wire [4-1:0] node17410;
	wire [4-1:0] node17413;
	wire [4-1:0] node17414;
	wire [4-1:0] node17415;
	wire [4-1:0] node17416;
	wire [4-1:0] node17419;
	wire [4-1:0] node17420;
	wire [4-1:0] node17423;
	wire [4-1:0] node17426;
	wire [4-1:0] node17427;
	wire [4-1:0] node17429;
	wire [4-1:0] node17430;
	wire [4-1:0] node17434;
	wire [4-1:0] node17437;
	wire [4-1:0] node17438;
	wire [4-1:0] node17439;
	wire [4-1:0] node17440;
	wire [4-1:0] node17444;
	wire [4-1:0] node17445;
	wire [4-1:0] node17448;
	wire [4-1:0] node17450;
	wire [4-1:0] node17453;
	wire [4-1:0] node17455;
	wire [4-1:0] node17456;
	wire [4-1:0] node17460;
	wire [4-1:0] node17461;
	wire [4-1:0] node17462;
	wire [4-1:0] node17463;
	wire [4-1:0] node17464;
	wire [4-1:0] node17467;
	wire [4-1:0] node17470;
	wire [4-1:0] node17471;
	wire [4-1:0] node17472;
	wire [4-1:0] node17473;
	wire [4-1:0] node17477;
	wire [4-1:0] node17480;
	wire [4-1:0] node17483;
	wire [4-1:0] node17484;
	wire [4-1:0] node17485;
	wire [4-1:0] node17488;
	wire [4-1:0] node17490;
	wire [4-1:0] node17493;
	wire [4-1:0] node17494;
	wire [4-1:0] node17498;
	wire [4-1:0] node17499;
	wire [4-1:0] node17500;
	wire [4-1:0] node17501;
	wire [4-1:0] node17502;
	wire [4-1:0] node17506;
	wire [4-1:0] node17509;
	wire [4-1:0] node17510;
	wire [4-1:0] node17512;
	wire [4-1:0] node17514;
	wire [4-1:0] node17517;
	wire [4-1:0] node17518;
	wire [4-1:0] node17520;
	wire [4-1:0] node17523;
	wire [4-1:0] node17525;
	wire [4-1:0] node17528;
	wire [4-1:0] node17529;
	wire [4-1:0] node17532;
	wire [4-1:0] node17533;
	wire [4-1:0] node17534;
	wire [4-1:0] node17537;
	wire [4-1:0] node17539;
	wire [4-1:0] node17543;
	wire [4-1:0] node17544;
	wire [4-1:0] node17545;
	wire [4-1:0] node17546;
	wire [4-1:0] node17547;
	wire [4-1:0] node17550;
	wire [4-1:0] node17553;
	wire [4-1:0] node17554;
	wire [4-1:0] node17555;
	wire [4-1:0] node17558;
	wire [4-1:0] node17559;
	wire [4-1:0] node17560;
	wire [4-1:0] node17565;
	wire [4-1:0] node17566;
	wire [4-1:0] node17567;
	wire [4-1:0] node17569;
	wire [4-1:0] node17573;
	wire [4-1:0] node17574;
	wire [4-1:0] node17575;
	wire [4-1:0] node17579;
	wire [4-1:0] node17582;
	wire [4-1:0] node17583;
	wire [4-1:0] node17584;
	wire [4-1:0] node17585;
	wire [4-1:0] node17587;
	wire [4-1:0] node17588;
	wire [4-1:0] node17592;
	wire [4-1:0] node17594;
	wire [4-1:0] node17597;
	wire [4-1:0] node17598;
	wire [4-1:0] node17601;
	wire [4-1:0] node17602;
	wire [4-1:0] node17606;
	wire [4-1:0] node17607;
	wire [4-1:0] node17608;
	wire [4-1:0] node17609;
	wire [4-1:0] node17610;
	wire [4-1:0] node17614;
	wire [4-1:0] node17616;
	wire [4-1:0] node17619;
	wire [4-1:0] node17622;
	wire [4-1:0] node17623;
	wire [4-1:0] node17624;
	wire [4-1:0] node17627;
	wire [4-1:0] node17629;
	wire [4-1:0] node17632;
	wire [4-1:0] node17634;
	wire [4-1:0] node17637;
	wire [4-1:0] node17638;
	wire [4-1:0] node17639;
	wire [4-1:0] node17640;
	wire [4-1:0] node17642;
	wire [4-1:0] node17644;
	wire [4-1:0] node17645;
	wire [4-1:0] node17649;
	wire [4-1:0] node17650;
	wire [4-1:0] node17653;
	wire [4-1:0] node17656;
	wire [4-1:0] node17657;
	wire [4-1:0] node17658;
	wire [4-1:0] node17661;
	wire [4-1:0] node17662;
	wire [4-1:0] node17666;
	wire [4-1:0] node17667;
	wire [4-1:0] node17668;
	wire [4-1:0] node17671;
	wire [4-1:0] node17675;
	wire [4-1:0] node17676;
	wire [4-1:0] node17677;
	wire [4-1:0] node17679;
	wire [4-1:0] node17682;
	wire [4-1:0] node17683;
	wire [4-1:0] node17685;
	wire [4-1:0] node17688;
	wire [4-1:0] node17691;
	wire [4-1:0] node17692;
	wire [4-1:0] node17693;
	wire [4-1:0] node17694;
	wire [4-1:0] node17695;
	wire [4-1:0] node17701;
	wire [4-1:0] node17702;
	wire [4-1:0] node17703;
	wire [4-1:0] node17705;
	wire [4-1:0] node17710;
	wire [4-1:0] node17711;
	wire [4-1:0] node17712;
	wire [4-1:0] node17713;
	wire [4-1:0] node17714;
	wire [4-1:0] node17715;
	wire [4-1:0] node17717;
	wire [4-1:0] node17718;
	wire [4-1:0] node17720;
	wire [4-1:0] node17723;
	wire [4-1:0] node17724;
	wire [4-1:0] node17727;
	wire [4-1:0] node17730;
	wire [4-1:0] node17732;
	wire [4-1:0] node17733;
	wire [4-1:0] node17737;
	wire [4-1:0] node17738;
	wire [4-1:0] node17739;
	wire [4-1:0] node17740;
	wire [4-1:0] node17743;
	wire [4-1:0] node17744;
	wire [4-1:0] node17749;
	wire [4-1:0] node17750;
	wire [4-1:0] node17753;
	wire [4-1:0] node17755;
	wire [4-1:0] node17756;
	wire [4-1:0] node17760;
	wire [4-1:0] node17761;
	wire [4-1:0] node17762;
	wire [4-1:0] node17763;
	wire [4-1:0] node17765;
	wire [4-1:0] node17766;
	wire [4-1:0] node17770;
	wire [4-1:0] node17771;
	wire [4-1:0] node17775;
	wire [4-1:0] node17776;
	wire [4-1:0] node17778;
	wire [4-1:0] node17781;
	wire [4-1:0] node17783;
	wire [4-1:0] node17786;
	wire [4-1:0] node17787;
	wire [4-1:0] node17788;
	wire [4-1:0] node17790;
	wire [4-1:0] node17793;
	wire [4-1:0] node17794;
	wire [4-1:0] node17797;
	wire [4-1:0] node17800;
	wire [4-1:0] node17801;
	wire [4-1:0] node17802;
	wire [4-1:0] node17804;
	wire [4-1:0] node17809;
	wire [4-1:0] node17810;
	wire [4-1:0] node17811;
	wire [4-1:0] node17812;
	wire [4-1:0] node17813;
	wire [4-1:0] node17814;
	wire [4-1:0] node17818;
	wire [4-1:0] node17819;
	wire [4-1:0] node17823;
	wire [4-1:0] node17824;
	wire [4-1:0] node17827;
	wire [4-1:0] node17829;
	wire [4-1:0] node17830;
	wire [4-1:0] node17833;
	wire [4-1:0] node17836;
	wire [4-1:0] node17837;
	wire [4-1:0] node17838;
	wire [4-1:0] node17839;
	wire [4-1:0] node17840;
	wire [4-1:0] node17845;
	wire [4-1:0] node17846;
	wire [4-1:0] node17848;
	wire [4-1:0] node17852;
	wire [4-1:0] node17853;
	wire [4-1:0] node17854;
	wire [4-1:0] node17858;
	wire [4-1:0] node17859;
	wire [4-1:0] node17860;
	wire [4-1:0] node17865;
	wire [4-1:0] node17866;
	wire [4-1:0] node17867;
	wire [4-1:0] node17868;
	wire [4-1:0] node17870;
	wire [4-1:0] node17874;
	wire [4-1:0] node17875;
	wire [4-1:0] node17877;
	wire [4-1:0] node17881;
	wire [4-1:0] node17882;
	wire [4-1:0] node17883;
	wire [4-1:0] node17884;
	wire [4-1:0] node17887;
	wire [4-1:0] node17890;
	wire [4-1:0] node17892;
	wire [4-1:0] node17895;
	wire [4-1:0] node17896;
	wire [4-1:0] node17897;
	wire [4-1:0] node17900;
	wire [4-1:0] node17901;
	wire [4-1:0] node17904;
	wire [4-1:0] node17907;
	wire [4-1:0] node17908;
	wire [4-1:0] node17910;
	wire [4-1:0] node17914;
	wire [4-1:0] node17915;
	wire [4-1:0] node17916;
	wire [4-1:0] node17917;
	wire [4-1:0] node17918;
	wire [4-1:0] node17919;
	wire [4-1:0] node17920;
	wire [4-1:0] node17921;
	wire [4-1:0] node17925;
	wire [4-1:0] node17926;
	wire [4-1:0] node17929;
	wire [4-1:0] node17932;
	wire [4-1:0] node17933;
	wire [4-1:0] node17934;
	wire [4-1:0] node17937;
	wire [4-1:0] node17940;
	wire [4-1:0] node17941;
	wire [4-1:0] node17944;
	wire [4-1:0] node17947;
	wire [4-1:0] node17950;
	wire [4-1:0] node17951;
	wire [4-1:0] node17954;
	wire [4-1:0] node17955;
	wire [4-1:0] node17956;
	wire [4-1:0] node17960;
	wire [4-1:0] node17962;
	wire [4-1:0] node17963;
	wire [4-1:0] node17966;
	wire [4-1:0] node17969;
	wire [4-1:0] node17970;
	wire [4-1:0] node17971;
	wire [4-1:0] node17972;
	wire [4-1:0] node17973;
	wire [4-1:0] node17974;
	wire [4-1:0] node17978;
	wire [4-1:0] node17979;
	wire [4-1:0] node17982;
	wire [4-1:0] node17985;
	wire [4-1:0] node17986;
	wire [4-1:0] node17989;
	wire [4-1:0] node17991;
	wire [4-1:0] node17994;
	wire [4-1:0] node17995;
	wire [4-1:0] node17997;
	wire [4-1:0] node17999;
	wire [4-1:0] node18002;
	wire [4-1:0] node18005;
	wire [4-1:0] node18006;
	wire [4-1:0] node18007;
	wire [4-1:0] node18011;
	wire [4-1:0] node18012;
	wire [4-1:0] node18013;
	wire [4-1:0] node18014;
	wire [4-1:0] node18018;
	wire [4-1:0] node18019;
	wire [4-1:0] node18023;
	wire [4-1:0] node18024;
	wire [4-1:0] node18026;
	wire [4-1:0] node18029;
	wire [4-1:0] node18030;
	wire [4-1:0] node18033;
	wire [4-1:0] node18036;
	wire [4-1:0] node18037;
	wire [4-1:0] node18038;
	wire [4-1:0] node18039;
	wire [4-1:0] node18040;
	wire [4-1:0] node18041;
	wire [4-1:0] node18042;
	wire [4-1:0] node18046;
	wire [4-1:0] node18048;
	wire [4-1:0] node18051;
	wire [4-1:0] node18054;
	wire [4-1:0] node18055;
	wire [4-1:0] node18056;
	wire [4-1:0] node18060;
	wire [4-1:0] node18062;
	wire [4-1:0] node18063;
	wire [4-1:0] node18067;
	wire [4-1:0] node18068;
	wire [4-1:0] node18069;
	wire [4-1:0] node18071;
	wire [4-1:0] node18074;
	wire [4-1:0] node18075;
	wire [4-1:0] node18078;
	wire [4-1:0] node18080;
	wire [4-1:0] node18083;
	wire [4-1:0] node18084;
	wire [4-1:0] node18087;
	wire [4-1:0] node18088;
	wire [4-1:0] node18089;
	wire [4-1:0] node18094;
	wire [4-1:0] node18095;
	wire [4-1:0] node18096;
	wire [4-1:0] node18097;
	wire [4-1:0] node18099;
	wire [4-1:0] node18102;
	wire [4-1:0] node18104;
	wire [4-1:0] node18105;
	wire [4-1:0] node18109;
	wire [4-1:0] node18111;
	wire [4-1:0] node18112;
	wire [4-1:0] node18115;
	wire [4-1:0] node18118;
	wire [4-1:0] node18119;
	wire [4-1:0] node18120;
	wire [4-1:0] node18121;
	wire [4-1:0] node18125;
	wire [4-1:0] node18126;
	wire [4-1:0] node18127;
	wire [4-1:0] node18132;
	wire [4-1:0] node18133;
	wire [4-1:0] node18135;
	wire [4-1:0] node18137;
	wire [4-1:0] node18140;
	wire [4-1:0] node18141;
	wire [4-1:0] node18144;
	wire [4-1:0] node18146;
	wire [4-1:0] node18149;
	wire [4-1:0] node18150;
	wire [4-1:0] node18151;
	wire [4-1:0] node18152;
	wire [4-1:0] node18153;
	wire [4-1:0] node18154;
	wire [4-1:0] node18155;
	wire [4-1:0] node18156;
	wire [4-1:0] node18158;
	wire [4-1:0] node18160;
	wire [4-1:0] node18163;
	wire [4-1:0] node18164;
	wire [4-1:0] node18166;
	wire [4-1:0] node18167;
	wire [4-1:0] node18171;
	wire [4-1:0] node18172;
	wire [4-1:0] node18176;
	wire [4-1:0] node18177;
	wire [4-1:0] node18178;
	wire [4-1:0] node18179;
	wire [4-1:0] node18183;
	wire [4-1:0] node18184;
	wire [4-1:0] node18186;
	wire [4-1:0] node18190;
	wire [4-1:0] node18191;
	wire [4-1:0] node18194;
	wire [4-1:0] node18197;
	wire [4-1:0] node18198;
	wire [4-1:0] node18199;
	wire [4-1:0] node18200;
	wire [4-1:0] node18201;
	wire [4-1:0] node18206;
	wire [4-1:0] node18208;
	wire [4-1:0] node18211;
	wire [4-1:0] node18212;
	wire [4-1:0] node18214;
	wire [4-1:0] node18216;
	wire [4-1:0] node18219;
	wire [4-1:0] node18220;
	wire [4-1:0] node18222;
	wire [4-1:0] node18225;
	wire [4-1:0] node18226;
	wire [4-1:0] node18229;
	wire [4-1:0] node18232;
	wire [4-1:0] node18233;
	wire [4-1:0] node18234;
	wire [4-1:0] node18235;
	wire [4-1:0] node18236;
	wire [4-1:0] node18237;
	wire [4-1:0] node18238;
	wire [4-1:0] node18242;
	wire [4-1:0] node18245;
	wire [4-1:0] node18248;
	wire [4-1:0] node18249;
	wire [4-1:0] node18252;
	wire [4-1:0] node18253;
	wire [4-1:0] node18254;
	wire [4-1:0] node18258;
	wire [4-1:0] node18261;
	wire [4-1:0] node18262;
	wire [4-1:0] node18263;
	wire [4-1:0] node18265;
	wire [4-1:0] node18266;
	wire [4-1:0] node18269;
	wire [4-1:0] node18272;
	wire [4-1:0] node18274;
	wire [4-1:0] node18277;
	wire [4-1:0] node18278;
	wire [4-1:0] node18280;
	wire [4-1:0] node18281;
	wire [4-1:0] node18284;
	wire [4-1:0] node18288;
	wire [4-1:0] node18289;
	wire [4-1:0] node18290;
	wire [4-1:0] node18291;
	wire [4-1:0] node18292;
	wire [4-1:0] node18294;
	wire [4-1:0] node18298;
	wire [4-1:0] node18299;
	wire [4-1:0] node18302;
	wire [4-1:0] node18303;
	wire [4-1:0] node18307;
	wire [4-1:0] node18309;
	wire [4-1:0] node18310;
	wire [4-1:0] node18313;
	wire [4-1:0] node18316;
	wire [4-1:0] node18317;
	wire [4-1:0] node18318;
	wire [4-1:0] node18319;
	wire [4-1:0] node18320;
	wire [4-1:0] node18324;
	wire [4-1:0] node18326;
	wire [4-1:0] node18329;
	wire [4-1:0] node18331;
	wire [4-1:0] node18334;
	wire [4-1:0] node18335;
	wire [4-1:0] node18338;
	wire [4-1:0] node18341;
	wire [4-1:0] node18342;
	wire [4-1:0] node18343;
	wire [4-1:0] node18344;
	wire [4-1:0] node18345;
	wire [4-1:0] node18346;
	wire [4-1:0] node18347;
	wire [4-1:0] node18348;
	wire [4-1:0] node18352;
	wire [4-1:0] node18355;
	wire [4-1:0] node18358;
	wire [4-1:0] node18359;
	wire [4-1:0] node18360;
	wire [4-1:0] node18363;
	wire [4-1:0] node18364;
	wire [4-1:0] node18369;
	wire [4-1:0] node18370;
	wire [4-1:0] node18371;
	wire [4-1:0] node18374;
	wire [4-1:0] node18377;
	wire [4-1:0] node18380;
	wire [4-1:0] node18381;
	wire [4-1:0] node18382;
	wire [4-1:0] node18383;
	wire [4-1:0] node18384;
	wire [4-1:0] node18385;
	wire [4-1:0] node18389;
	wire [4-1:0] node18391;
	wire [4-1:0] node18394;
	wire [4-1:0] node18396;
	wire [4-1:0] node18397;
	wire [4-1:0] node18401;
	wire [4-1:0] node18402;
	wire [4-1:0] node18404;
	wire [4-1:0] node18405;
	wire [4-1:0] node18410;
	wire [4-1:0] node18411;
	wire [4-1:0] node18412;
	wire [4-1:0] node18414;
	wire [4-1:0] node18417;
	wire [4-1:0] node18419;
	wire [4-1:0] node18422;
	wire [4-1:0] node18423;
	wire [4-1:0] node18425;
	wire [4-1:0] node18428;
	wire [4-1:0] node18429;
	wire [4-1:0] node18431;
	wire [4-1:0] node18435;
	wire [4-1:0] node18436;
	wire [4-1:0] node18437;
	wire [4-1:0] node18438;
	wire [4-1:0] node18439;
	wire [4-1:0] node18442;
	wire [4-1:0] node18444;
	wire [4-1:0] node18445;
	wire [4-1:0] node18449;
	wire [4-1:0] node18450;
	wire [4-1:0] node18453;
	wire [4-1:0] node18454;
	wire [4-1:0] node18455;
	wire [4-1:0] node18458;
	wire [4-1:0] node18462;
	wire [4-1:0] node18463;
	wire [4-1:0] node18464;
	wire [4-1:0] node18468;
	wire [4-1:0] node18469;
	wire [4-1:0] node18472;
	wire [4-1:0] node18474;
	wire [4-1:0] node18477;
	wire [4-1:0] node18478;
	wire [4-1:0] node18479;
	wire [4-1:0] node18480;
	wire [4-1:0] node18481;
	wire [4-1:0] node18482;
	wire [4-1:0] node18485;
	wire [4-1:0] node18489;
	wire [4-1:0] node18491;
	wire [4-1:0] node18493;
	wire [4-1:0] node18496;
	wire [4-1:0] node18497;
	wire [4-1:0] node18499;
	wire [4-1:0] node18500;
	wire [4-1:0] node18504;
	wire [4-1:0] node18505;
	wire [4-1:0] node18506;
	wire [4-1:0] node18511;
	wire [4-1:0] node18512;
	wire [4-1:0] node18515;
	wire [4-1:0] node18516;
	wire [4-1:0] node18517;
	wire [4-1:0] node18518;
	wire [4-1:0] node18524;
	wire [4-1:0] node18525;
	wire [4-1:0] node18526;
	wire [4-1:0] node18527;
	wire [4-1:0] node18528;
	wire [4-1:0] node18529;
	wire [4-1:0] node18530;
	wire [4-1:0] node18532;
	wire [4-1:0] node18535;
	wire [4-1:0] node18537;
	wire [4-1:0] node18540;
	wire [4-1:0] node18541;
	wire [4-1:0] node18542;
	wire [4-1:0] node18543;
	wire [4-1:0] node18548;
	wire [4-1:0] node18551;
	wire [4-1:0] node18552;
	wire [4-1:0] node18554;
	wire [4-1:0] node18556;
	wire [4-1:0] node18558;
	wire [4-1:0] node18561;
	wire [4-1:0] node18562;
	wire [4-1:0] node18563;
	wire [4-1:0] node18567;
	wire [4-1:0] node18570;
	wire [4-1:0] node18571;
	wire [4-1:0] node18572;
	wire [4-1:0] node18573;
	wire [4-1:0] node18574;
	wire [4-1:0] node18575;
	wire [4-1:0] node18579;
	wire [4-1:0] node18582;
	wire [4-1:0] node18583;
	wire [4-1:0] node18587;
	wire [4-1:0] node18588;
	wire [4-1:0] node18589;
	wire [4-1:0] node18593;
	wire [4-1:0] node18596;
	wire [4-1:0] node18598;
	wire [4-1:0] node18599;
	wire [4-1:0] node18600;
	wire [4-1:0] node18602;
	wire [4-1:0] node18606;
	wire [4-1:0] node18609;
	wire [4-1:0] node18610;
	wire [4-1:0] node18611;
	wire [4-1:0] node18612;
	wire [4-1:0] node18613;
	wire [4-1:0] node18614;
	wire [4-1:0] node18619;
	wire [4-1:0] node18620;
	wire [4-1:0] node18623;
	wire [4-1:0] node18624;
	wire [4-1:0] node18627;
	wire [4-1:0] node18630;
	wire [4-1:0] node18631;
	wire [4-1:0] node18634;
	wire [4-1:0] node18636;
	wire [4-1:0] node18638;
	wire [4-1:0] node18639;
	wire [4-1:0] node18642;
	wire [4-1:0] node18645;
	wire [4-1:0] node18646;
	wire [4-1:0] node18647;
	wire [4-1:0] node18648;
	wire [4-1:0] node18653;
	wire [4-1:0] node18654;
	wire [4-1:0] node18655;
	wire [4-1:0] node18656;
	wire [4-1:0] node18658;
	wire [4-1:0] node18663;
	wire [4-1:0] node18664;
	wire [4-1:0] node18665;
	wire [4-1:0] node18669;
	wire [4-1:0] node18670;
	wire [4-1:0] node18674;
	wire [4-1:0] node18675;
	wire [4-1:0] node18676;
	wire [4-1:0] node18677;
	wire [4-1:0] node18678;
	wire [4-1:0] node18679;
	wire [4-1:0] node18680;
	wire [4-1:0] node18681;
	wire [4-1:0] node18686;
	wire [4-1:0] node18688;
	wire [4-1:0] node18691;
	wire [4-1:0] node18692;
	wire [4-1:0] node18693;
	wire [4-1:0] node18697;
	wire [4-1:0] node18698;
	wire [4-1:0] node18700;
	wire [4-1:0] node18704;
	wire [4-1:0] node18705;
	wire [4-1:0] node18708;
	wire [4-1:0] node18709;
	wire [4-1:0] node18712;
	wire [4-1:0] node18714;
	wire [4-1:0] node18717;
	wire [4-1:0] node18718;
	wire [4-1:0] node18719;
	wire [4-1:0] node18721;
	wire [4-1:0] node18722;
	wire [4-1:0] node18725;
	wire [4-1:0] node18726;
	wire [4-1:0] node18730;
	wire [4-1:0] node18732;
	wire [4-1:0] node18733;
	wire [4-1:0] node18735;
	wire [4-1:0] node18738;
	wire [4-1:0] node18741;
	wire [4-1:0] node18742;
	wire [4-1:0] node18743;
	wire [4-1:0] node18745;
	wire [4-1:0] node18746;
	wire [4-1:0] node18749;
	wire [4-1:0] node18752;
	wire [4-1:0] node18755;
	wire [4-1:0] node18758;
	wire [4-1:0] node18759;
	wire [4-1:0] node18760;
	wire [4-1:0] node18761;
	wire [4-1:0] node18762;
	wire [4-1:0] node18763;
	wire [4-1:0] node18767;
	wire [4-1:0] node18770;
	wire [4-1:0] node18771;
	wire [4-1:0] node18772;
	wire [4-1:0] node18776;
	wire [4-1:0] node18777;
	wire [4-1:0] node18779;
	wire [4-1:0] node18782;
	wire [4-1:0] node18785;
	wire [4-1:0] node18786;
	wire [4-1:0] node18787;
	wire [4-1:0] node18788;
	wire [4-1:0] node18789;
	wire [4-1:0] node18794;
	wire [4-1:0] node18796;
	wire [4-1:0] node18799;
	wire [4-1:0] node18800;
	wire [4-1:0] node18801;
	wire [4-1:0] node18803;
	wire [4-1:0] node18807;
	wire [4-1:0] node18810;
	wire [4-1:0] node18811;
	wire [4-1:0] node18812;
	wire [4-1:0] node18815;
	wire [4-1:0] node18816;
	wire [4-1:0] node18817;
	wire [4-1:0] node18821;
	wire [4-1:0] node18822;
	wire [4-1:0] node18823;
	wire [4-1:0] node18827;
	wire [4-1:0] node18830;
	wire [4-1:0] node18831;
	wire [4-1:0] node18832;
	wire [4-1:0] node18834;
	wire [4-1:0] node18836;
	wire [4-1:0] node18839;
	wire [4-1:0] node18840;
	wire [4-1:0] node18841;
	wire [4-1:0] node18845;
	wire [4-1:0] node18846;
	wire [4-1:0] node18850;
	wire [4-1:0] node18851;
	wire [4-1:0] node18852;
	wire [4-1:0] node18853;
	wire [4-1:0] node18858;
	wire [4-1:0] node18860;
	wire [4-1:0] node18862;
	wire [4-1:0] node18865;
	wire [4-1:0] node18866;
	wire [4-1:0] node18867;
	wire [4-1:0] node18868;
	wire [4-1:0] node18869;
	wire [4-1:0] node18870;
	wire [4-1:0] node18871;
	wire [4-1:0] node18872;
	wire [4-1:0] node18874;
	wire [4-1:0] node18877;
	wire [4-1:0] node18880;
	wire [4-1:0] node18881;
	wire [4-1:0] node18882;
	wire [4-1:0] node18884;
	wire [4-1:0] node18888;
	wire [4-1:0] node18891;
	wire [4-1:0] node18892;
	wire [4-1:0] node18893;
	wire [4-1:0] node18896;
	wire [4-1:0] node18899;
	wire [4-1:0] node18901;
	wire [4-1:0] node18904;
	wire [4-1:0] node18905;
	wire [4-1:0] node18906;
	wire [4-1:0] node18907;
	wire [4-1:0] node18909;
	wire [4-1:0] node18910;
	wire [4-1:0] node18915;
	wire [4-1:0] node18917;
	wire [4-1:0] node18919;
	wire [4-1:0] node18922;
	wire [4-1:0] node18923;
	wire [4-1:0] node18924;
	wire [4-1:0] node18926;
	wire [4-1:0] node18927;
	wire [4-1:0] node18931;
	wire [4-1:0] node18934;
	wire [4-1:0] node18936;
	wire [4-1:0] node18937;
	wire [4-1:0] node18940;
	wire [4-1:0] node18941;
	wire [4-1:0] node18945;
	wire [4-1:0] node18946;
	wire [4-1:0] node18947;
	wire [4-1:0] node18948;
	wire [4-1:0] node18949;
	wire [4-1:0] node18951;
	wire [4-1:0] node18953;
	wire [4-1:0] node18956;
	wire [4-1:0] node18958;
	wire [4-1:0] node18961;
	wire [4-1:0] node18962;
	wire [4-1:0] node18963;
	wire [4-1:0] node18967;
	wire [4-1:0] node18968;
	wire [4-1:0] node18969;
	wire [4-1:0] node18974;
	wire [4-1:0] node18975;
	wire [4-1:0] node18976;
	wire [4-1:0] node18979;
	wire [4-1:0] node18981;
	wire [4-1:0] node18983;
	wire [4-1:0] node18986;
	wire [4-1:0] node18988;
	wire [4-1:0] node18989;
	wire [4-1:0] node18990;
	wire [4-1:0] node18993;
	wire [4-1:0] node18997;
	wire [4-1:0] node18998;
	wire [4-1:0] node18999;
	wire [4-1:0] node19000;
	wire [4-1:0] node19002;
	wire [4-1:0] node19005;
	wire [4-1:0] node19007;
	wire [4-1:0] node19010;
	wire [4-1:0] node19011;
	wire [4-1:0] node19014;
	wire [4-1:0] node19016;
	wire [4-1:0] node19017;
	wire [4-1:0] node19021;
	wire [4-1:0] node19022;
	wire [4-1:0] node19023;
	wire [4-1:0] node19024;
	wire [4-1:0] node19029;
	wire [4-1:0] node19030;
	wire [4-1:0] node19031;
	wire [4-1:0] node19032;
	wire [4-1:0] node19035;
	wire [4-1:0] node19038;
	wire [4-1:0] node19040;
	wire [4-1:0] node19043;
	wire [4-1:0] node19044;
	wire [4-1:0] node19048;
	wire [4-1:0] node19049;
	wire [4-1:0] node19050;
	wire [4-1:0] node19051;
	wire [4-1:0] node19052;
	wire [4-1:0] node19053;
	wire [4-1:0] node19054;
	wire [4-1:0] node19058;
	wire [4-1:0] node19060;
	wire [4-1:0] node19063;
	wire [4-1:0] node19064;
	wire [4-1:0] node19067;
	wire [4-1:0] node19068;
	wire [4-1:0] node19072;
	wire [4-1:0] node19073;
	wire [4-1:0] node19074;
	wire [4-1:0] node19078;
	wire [4-1:0] node19079;
	wire [4-1:0] node19083;
	wire [4-1:0] node19084;
	wire [4-1:0] node19085;
	wire [4-1:0] node19086;
	wire [4-1:0] node19088;
	wire [4-1:0] node19089;
	wire [4-1:0] node19092;
	wire [4-1:0] node19095;
	wire [4-1:0] node19097;
	wire [4-1:0] node19098;
	wire [4-1:0] node19101;
	wire [4-1:0] node19104;
	wire [4-1:0] node19105;
	wire [4-1:0] node19106;
	wire [4-1:0] node19109;
	wire [4-1:0] node19112;
	wire [4-1:0] node19114;
	wire [4-1:0] node19117;
	wire [4-1:0] node19118;
	wire [4-1:0] node19119;
	wire [4-1:0] node19120;
	wire [4-1:0] node19123;
	wire [4-1:0] node19126;
	wire [4-1:0] node19128;
	wire [4-1:0] node19129;
	wire [4-1:0] node19133;
	wire [4-1:0] node19135;
	wire [4-1:0] node19136;
	wire [4-1:0] node19139;
	wire [4-1:0] node19142;
	wire [4-1:0] node19143;
	wire [4-1:0] node19144;
	wire [4-1:0] node19145;
	wire [4-1:0] node19146;
	wire [4-1:0] node19147;
	wire [4-1:0] node19151;
	wire [4-1:0] node19152;
	wire [4-1:0] node19156;
	wire [4-1:0] node19157;
	wire [4-1:0] node19160;
	wire [4-1:0] node19163;
	wire [4-1:0] node19164;
	wire [4-1:0] node19165;
	wire [4-1:0] node19167;
	wire [4-1:0] node19171;
	wire [4-1:0] node19172;
	wire [4-1:0] node19173;
	wire [4-1:0] node19178;
	wire [4-1:0] node19179;
	wire [4-1:0] node19180;
	wire [4-1:0] node19182;
	wire [4-1:0] node19184;
	wire [4-1:0] node19187;
	wire [4-1:0] node19188;
	wire [4-1:0] node19190;
	wire [4-1:0] node19194;
	wire [4-1:0] node19195;
	wire [4-1:0] node19196;
	wire [4-1:0] node19197;
	wire [4-1:0] node19198;
	wire [4-1:0] node19203;
	wire [4-1:0] node19206;
	wire [4-1:0] node19207;
	wire [4-1:0] node19208;
	wire [4-1:0] node19213;
	wire [4-1:0] node19214;
	wire [4-1:0] node19215;
	wire [4-1:0] node19216;
	wire [4-1:0] node19217;
	wire [4-1:0] node19218;
	wire [4-1:0] node19219;
	wire [4-1:0] node19220;
	wire [4-1:0] node19222;
	wire [4-1:0] node19225;
	wire [4-1:0] node19226;
	wire [4-1:0] node19230;
	wire [4-1:0] node19233;
	wire [4-1:0] node19234;
	wire [4-1:0] node19237;
	wire [4-1:0] node19240;
	wire [4-1:0] node19241;
	wire [4-1:0] node19242;
	wire [4-1:0] node19243;
	wire [4-1:0] node19244;
	wire [4-1:0] node19247;
	wire [4-1:0] node19250;
	wire [4-1:0] node19253;
	wire [4-1:0] node19254;
	wire [4-1:0] node19256;
	wire [4-1:0] node19260;
	wire [4-1:0] node19261;
	wire [4-1:0] node19263;
	wire [4-1:0] node19266;
	wire [4-1:0] node19267;
	wire [4-1:0] node19270;
	wire [4-1:0] node19273;
	wire [4-1:0] node19274;
	wire [4-1:0] node19275;
	wire [4-1:0] node19276;
	wire [4-1:0] node19277;
	wire [4-1:0] node19280;
	wire [4-1:0] node19283;
	wire [4-1:0] node19286;
	wire [4-1:0] node19287;
	wire [4-1:0] node19290;
	wire [4-1:0] node19291;
	wire [4-1:0] node19294;
	wire [4-1:0] node19297;
	wire [4-1:0] node19298;
	wire [4-1:0] node19300;
	wire [4-1:0] node19303;
	wire [4-1:0] node19305;
	wire [4-1:0] node19306;
	wire [4-1:0] node19310;
	wire [4-1:0] node19311;
	wire [4-1:0] node19312;
	wire [4-1:0] node19313;
	wire [4-1:0] node19314;
	wire [4-1:0] node19315;
	wire [4-1:0] node19318;
	wire [4-1:0] node19320;
	wire [4-1:0] node19323;
	wire [4-1:0] node19324;
	wire [4-1:0] node19325;
	wire [4-1:0] node19329;
	wire [4-1:0] node19332;
	wire [4-1:0] node19333;
	wire [4-1:0] node19334;
	wire [4-1:0] node19337;
	wire [4-1:0] node19340;
	wire [4-1:0] node19341;
	wire [4-1:0] node19342;
	wire [4-1:0] node19346;
	wire [4-1:0] node19349;
	wire [4-1:0] node19350;
	wire [4-1:0] node19351;
	wire [4-1:0] node19352;
	wire [4-1:0] node19356;
	wire [4-1:0] node19358;
	wire [4-1:0] node19359;
	wire [4-1:0] node19363;
	wire [4-1:0] node19364;
	wire [4-1:0] node19366;
	wire [4-1:0] node19369;
	wire [4-1:0] node19371;
	wire [4-1:0] node19374;
	wire [4-1:0] node19375;
	wire [4-1:0] node19376;
	wire [4-1:0] node19377;
	wire [4-1:0] node19378;
	wire [4-1:0] node19383;
	wire [4-1:0] node19384;
	wire [4-1:0] node19386;
	wire [4-1:0] node19388;
	wire [4-1:0] node19391;
	wire [4-1:0] node19394;
	wire [4-1:0] node19395;
	wire [4-1:0] node19396;
	wire [4-1:0] node19399;
	wire [4-1:0] node19400;
	wire [4-1:0] node19401;
	wire [4-1:0] node19404;
	wire [4-1:0] node19408;
	wire [4-1:0] node19409;
	wire [4-1:0] node19410;
	wire [4-1:0] node19412;
	wire [4-1:0] node19415;
	wire [4-1:0] node19418;
	wire [4-1:0] node19419;
	wire [4-1:0] node19420;
	wire [4-1:0] node19424;
	wire [4-1:0] node19426;
	wire [4-1:0] node19429;
	wire [4-1:0] node19430;
	wire [4-1:0] node19431;
	wire [4-1:0] node19432;
	wire [4-1:0] node19433;
	wire [4-1:0] node19434;
	wire [4-1:0] node19436;
	wire [4-1:0] node19438;
	wire [4-1:0] node19441;
	wire [4-1:0] node19442;
	wire [4-1:0] node19445;
	wire [4-1:0] node19448;
	wire [4-1:0] node19449;
	wire [4-1:0] node19451;
	wire [4-1:0] node19454;
	wire [4-1:0] node19456;
	wire [4-1:0] node19457;
	wire [4-1:0] node19461;
	wire [4-1:0] node19462;
	wire [4-1:0] node19463;
	wire [4-1:0] node19464;
	wire [4-1:0] node19467;
	wire [4-1:0] node19471;
	wire [4-1:0] node19472;
	wire [4-1:0] node19476;
	wire [4-1:0] node19477;
	wire [4-1:0] node19478;
	wire [4-1:0] node19479;
	wire [4-1:0] node19480;
	wire [4-1:0] node19483;
	wire [4-1:0] node19487;
	wire [4-1:0] node19489;
	wire [4-1:0] node19491;
	wire [4-1:0] node19494;
	wire [4-1:0] node19495;
	wire [4-1:0] node19496;
	wire [4-1:0] node19499;
	wire [4-1:0] node19502;
	wire [4-1:0] node19503;
	wire [4-1:0] node19505;
	wire [4-1:0] node19508;
	wire [4-1:0] node19509;
	wire [4-1:0] node19512;
	wire [4-1:0] node19515;
	wire [4-1:0] node19516;
	wire [4-1:0] node19517;
	wire [4-1:0] node19518;
	wire [4-1:0] node19519;
	wire [4-1:0] node19522;
	wire [4-1:0] node19523;
	wire [4-1:0] node19525;
	wire [4-1:0] node19528;
	wire [4-1:0] node19530;
	wire [4-1:0] node19533;
	wire [4-1:0] node19534;
	wire [4-1:0] node19535;
	wire [4-1:0] node19536;
	wire [4-1:0] node19541;
	wire [4-1:0] node19543;
	wire [4-1:0] node19544;
	wire [4-1:0] node19548;
	wire [4-1:0] node19549;
	wire [4-1:0] node19550;
	wire [4-1:0] node19552;
	wire [4-1:0] node19554;
	wire [4-1:0] node19557;
	wire [4-1:0] node19558;
	wire [4-1:0] node19562;
	wire [4-1:0] node19565;
	wire [4-1:0] node19566;
	wire [4-1:0] node19567;
	wire [4-1:0] node19568;
	wire [4-1:0] node19570;
	wire [4-1:0] node19574;
	wire [4-1:0] node19575;
	wire [4-1:0] node19577;
	wire [4-1:0] node19580;
	wire [4-1:0] node19581;
	wire [4-1:0] node19585;
	wire [4-1:0] node19586;
	wire [4-1:0] node19588;
	wire [4-1:0] node19589;
	wire [4-1:0] node19590;
	wire [4-1:0] node19594;
	wire [4-1:0] node19596;
	wire [4-1:0] node19599;
	wire [4-1:0] node19600;
	wire [4-1:0] node19603;
	wire [4-1:0] node19604;
	wire [4-1:0] node19608;
	wire [4-1:0] node19609;
	wire [4-1:0] node19610;
	wire [4-1:0] node19611;
	wire [4-1:0] node19612;
	wire [4-1:0] node19613;
	wire [4-1:0] node19614;
	wire [4-1:0] node19615;
	wire [4-1:0] node19616;
	wire [4-1:0] node19617;
	wire [4-1:0] node19618;
	wire [4-1:0] node19620;
	wire [4-1:0] node19624;
	wire [4-1:0] node19625;
	wire [4-1:0] node19629;
	wire [4-1:0] node19631;
	wire [4-1:0] node19634;
	wire [4-1:0] node19635;
	wire [4-1:0] node19636;
	wire [4-1:0] node19637;
	wire [4-1:0] node19640;
	wire [4-1:0] node19643;
	wire [4-1:0] node19644;
	wire [4-1:0] node19649;
	wire [4-1:0] node19650;
	wire [4-1:0] node19651;
	wire [4-1:0] node19652;
	wire [4-1:0] node19653;
	wire [4-1:0] node19654;
	wire [4-1:0] node19659;
	wire [4-1:0] node19662;
	wire [4-1:0] node19664;
	wire [4-1:0] node19667;
	wire [4-1:0] node19668;
	wire [4-1:0] node19669;
	wire [4-1:0] node19671;
	wire [4-1:0] node19673;
	wire [4-1:0] node19677;
	wire [4-1:0] node19678;
	wire [4-1:0] node19680;
	wire [4-1:0] node19681;
	wire [4-1:0] node19686;
	wire [4-1:0] node19687;
	wire [4-1:0] node19688;
	wire [4-1:0] node19689;
	wire [4-1:0] node19690;
	wire [4-1:0] node19694;
	wire [4-1:0] node19695;
	wire [4-1:0] node19696;
	wire [4-1:0] node19700;
	wire [4-1:0] node19701;
	wire [4-1:0] node19705;
	wire [4-1:0] node19706;
	wire [4-1:0] node19708;
	wire [4-1:0] node19710;
	wire [4-1:0] node19713;
	wire [4-1:0] node19714;
	wire [4-1:0] node19717;
	wire [4-1:0] node19720;
	wire [4-1:0] node19721;
	wire [4-1:0] node19722;
	wire [4-1:0] node19723;
	wire [4-1:0] node19725;
	wire [4-1:0] node19727;
	wire [4-1:0] node19730;
	wire [4-1:0] node19731;
	wire [4-1:0] node19735;
	wire [4-1:0] node19736;
	wire [4-1:0] node19739;
	wire [4-1:0] node19742;
	wire [4-1:0] node19743;
	wire [4-1:0] node19745;
	wire [4-1:0] node19747;
	wire [4-1:0] node19748;
	wire [4-1:0] node19752;
	wire [4-1:0] node19753;
	wire [4-1:0] node19755;
	wire [4-1:0] node19758;
	wire [4-1:0] node19760;
	wire [4-1:0] node19761;
	wire [4-1:0] node19765;
	wire [4-1:0] node19766;
	wire [4-1:0] node19767;
	wire [4-1:0] node19768;
	wire [4-1:0] node19769;
	wire [4-1:0] node19770;
	wire [4-1:0] node19771;
	wire [4-1:0] node19776;
	wire [4-1:0] node19777;
	wire [4-1:0] node19778;
	wire [4-1:0] node19782;
	wire [4-1:0] node19785;
	wire [4-1:0] node19786;
	wire [4-1:0] node19787;
	wire [4-1:0] node19791;
	wire [4-1:0] node19792;
	wire [4-1:0] node19796;
	wire [4-1:0] node19797;
	wire [4-1:0] node19798;
	wire [4-1:0] node19800;
	wire [4-1:0] node19802;
	wire [4-1:0] node19803;
	wire [4-1:0] node19807;
	wire [4-1:0] node19808;
	wire [4-1:0] node19812;
	wire [4-1:0] node19813;
	wire [4-1:0] node19814;
	wire [4-1:0] node19818;
	wire [4-1:0] node19819;
	wire [4-1:0] node19821;
	wire [4-1:0] node19824;
	wire [4-1:0] node19825;
	wire [4-1:0] node19829;
	wire [4-1:0] node19830;
	wire [4-1:0] node19831;
	wire [4-1:0] node19832;
	wire [4-1:0] node19833;
	wire [4-1:0] node19834;
	wire [4-1:0] node19838;
	wire [4-1:0] node19840;
	wire [4-1:0] node19843;
	wire [4-1:0] node19844;
	wire [4-1:0] node19845;
	wire [4-1:0] node19849;
	wire [4-1:0] node19851;
	wire [4-1:0] node19853;
	wire [4-1:0] node19856;
	wire [4-1:0] node19857;
	wire [4-1:0] node19858;
	wire [4-1:0] node19859;
	wire [4-1:0] node19863;
	wire [4-1:0] node19864;
	wire [4-1:0] node19867;
	wire [4-1:0] node19870;
	wire [4-1:0] node19873;
	wire [4-1:0] node19874;
	wire [4-1:0] node19875;
	wire [4-1:0] node19877;
	wire [4-1:0] node19878;
	wire [4-1:0] node19879;
	wire [4-1:0] node19884;
	wire [4-1:0] node19886;
	wire [4-1:0] node19887;
	wire [4-1:0] node19888;
	wire [4-1:0] node19891;
	wire [4-1:0] node19895;
	wire [4-1:0] node19896;
	wire [4-1:0] node19897;
	wire [4-1:0] node19898;
	wire [4-1:0] node19899;
	wire [4-1:0] node19902;
	wire [4-1:0] node19907;
	wire [4-1:0] node19909;
	wire [4-1:0] node19912;
	wire [4-1:0] node19913;
	wire [4-1:0] node19914;
	wire [4-1:0] node19915;
	wire [4-1:0] node19916;
	wire [4-1:0] node19917;
	wire [4-1:0] node19919;
	wire [4-1:0] node19922;
	wire [4-1:0] node19923;
	wire [4-1:0] node19924;
	wire [4-1:0] node19928;
	wire [4-1:0] node19931;
	wire [4-1:0] node19932;
	wire [4-1:0] node19935;
	wire [4-1:0] node19936;
	wire [4-1:0] node19938;
	wire [4-1:0] node19941;
	wire [4-1:0] node19944;
	wire [4-1:0] node19945;
	wire [4-1:0] node19946;
	wire [4-1:0] node19947;
	wire [4-1:0] node19948;
	wire [4-1:0] node19951;
	wire [4-1:0] node19952;
	wire [4-1:0] node19956;
	wire [4-1:0] node19958;
	wire [4-1:0] node19961;
	wire [4-1:0] node19962;
	wire [4-1:0] node19965;
	wire [4-1:0] node19968;
	wire [4-1:0] node19969;
	wire [4-1:0] node19970;
	wire [4-1:0] node19973;
	wire [4-1:0] node19974;
	wire [4-1:0] node19975;
	wire [4-1:0] node19980;
	wire [4-1:0] node19981;
	wire [4-1:0] node19984;
	wire [4-1:0] node19985;
	wire [4-1:0] node19987;
	wire [4-1:0] node19990;
	wire [4-1:0] node19991;
	wire [4-1:0] node19994;
	wire [4-1:0] node19997;
	wire [4-1:0] node19998;
	wire [4-1:0] node19999;
	wire [4-1:0] node20000;
	wire [4-1:0] node20001;
	wire [4-1:0] node20003;
	wire [4-1:0] node20004;
	wire [4-1:0] node20008;
	wire [4-1:0] node20010;
	wire [4-1:0] node20011;
	wire [4-1:0] node20014;
	wire [4-1:0] node20017;
	wire [4-1:0] node20019;
	wire [4-1:0] node20020;
	wire [4-1:0] node20021;
	wire [4-1:0] node20025;
	wire [4-1:0] node20028;
	wire [4-1:0] node20029;
	wire [4-1:0] node20030;
	wire [4-1:0] node20032;
	wire [4-1:0] node20034;
	wire [4-1:0] node20037;
	wire [4-1:0] node20039;
	wire [4-1:0] node20040;
	wire [4-1:0] node20045;
	wire [4-1:0] node20046;
	wire [4-1:0] node20047;
	wire [4-1:0] node20048;
	wire [4-1:0] node20050;
	wire [4-1:0] node20054;
	wire [4-1:0] node20055;
	wire [4-1:0] node20056;
	wire [4-1:0] node20059;
	wire [4-1:0] node20060;
	wire [4-1:0] node20065;
	wire [4-1:0] node20066;
	wire [4-1:0] node20068;
	wire [4-1:0] node20071;
	wire [4-1:0] node20072;
	wire [4-1:0] node20075;
	wire [4-1:0] node20078;
	wire [4-1:0] node20079;
	wire [4-1:0] node20080;
	wire [4-1:0] node20081;
	wire [4-1:0] node20082;
	wire [4-1:0] node20083;
	wire [4-1:0] node20084;
	wire [4-1:0] node20088;
	wire [4-1:0] node20091;
	wire [4-1:0] node20092;
	wire [4-1:0] node20095;
	wire [4-1:0] node20096;
	wire [4-1:0] node20097;
	wire [4-1:0] node20100;
	wire [4-1:0] node20104;
	wire [4-1:0] node20105;
	wire [4-1:0] node20108;
	wire [4-1:0] node20109;
	wire [4-1:0] node20111;
	wire [4-1:0] node20114;
	wire [4-1:0] node20115;
	wire [4-1:0] node20118;
	wire [4-1:0] node20119;
	wire [4-1:0] node20123;
	wire [4-1:0] node20124;
	wire [4-1:0] node20125;
	wire [4-1:0] node20126;
	wire [4-1:0] node20127;
	wire [4-1:0] node20128;
	wire [4-1:0] node20132;
	wire [4-1:0] node20136;
	wire [4-1:0] node20137;
	wire [4-1:0] node20138;
	wire [4-1:0] node20141;
	wire [4-1:0] node20142;
	wire [4-1:0] node20146;
	wire [4-1:0] node20147;
	wire [4-1:0] node20151;
	wire [4-1:0] node20152;
	wire [4-1:0] node20153;
	wire [4-1:0] node20154;
	wire [4-1:0] node20155;
	wire [4-1:0] node20160;
	wire [4-1:0] node20161;
	wire [4-1:0] node20163;
	wire [4-1:0] node20167;
	wire [4-1:0] node20168;
	wire [4-1:0] node20171;
	wire [4-1:0] node20172;
	wire [4-1:0] node20173;
	wire [4-1:0] node20176;
	wire [4-1:0] node20180;
	wire [4-1:0] node20181;
	wire [4-1:0] node20182;
	wire [4-1:0] node20183;
	wire [4-1:0] node20184;
	wire [4-1:0] node20185;
	wire [4-1:0] node20189;
	wire [4-1:0] node20191;
	wire [4-1:0] node20194;
	wire [4-1:0] node20195;
	wire [4-1:0] node20196;
	wire [4-1:0] node20198;
	wire [4-1:0] node20201;
	wire [4-1:0] node20204;
	wire [4-1:0] node20206;
	wire [4-1:0] node20209;
	wire [4-1:0] node20210;
	wire [4-1:0] node20211;
	wire [4-1:0] node20214;
	wire [4-1:0] node20215;
	wire [4-1:0] node20217;
	wire [4-1:0] node20221;
	wire [4-1:0] node20222;
	wire [4-1:0] node20223;
	wire [4-1:0] node20227;
	wire [4-1:0] node20229;
	wire [4-1:0] node20232;
	wire [4-1:0] node20233;
	wire [4-1:0] node20234;
	wire [4-1:0] node20235;
	wire [4-1:0] node20237;
	wire [4-1:0] node20240;
	wire [4-1:0] node20243;
	wire [4-1:0] node20244;
	wire [4-1:0] node20246;
	wire [4-1:0] node20250;
	wire [4-1:0] node20251;
	wire [4-1:0] node20252;
	wire [4-1:0] node20253;
	wire [4-1:0] node20256;
	wire [4-1:0] node20259;
	wire [4-1:0] node20261;
	wire [4-1:0] node20262;
	wire [4-1:0] node20266;
	wire [4-1:0] node20267;
	wire [4-1:0] node20268;
	wire [4-1:0] node20270;
	wire [4-1:0] node20273;
	wire [4-1:0] node20274;
	wire [4-1:0] node20278;
	wire [4-1:0] node20280;
	wire [4-1:0] node20283;
	wire [4-1:0] node20284;
	wire [4-1:0] node20285;
	wire [4-1:0] node20286;
	wire [4-1:0] node20287;
	wire [4-1:0] node20288;
	wire [4-1:0] node20289;
	wire [4-1:0] node20290;
	wire [4-1:0] node20293;
	wire [4-1:0] node20296;
	wire [4-1:0] node20297;
	wire [4-1:0] node20300;
	wire [4-1:0] node20303;
	wire [4-1:0] node20304;
	wire [4-1:0] node20305;
	wire [4-1:0] node20306;
	wire [4-1:0] node20308;
	wire [4-1:0] node20311;
	wire [4-1:0] node20313;
	wire [4-1:0] node20317;
	wire [4-1:0] node20318;
	wire [4-1:0] node20321;
	wire [4-1:0] node20322;
	wire [4-1:0] node20326;
	wire [4-1:0] node20327;
	wire [4-1:0] node20328;
	wire [4-1:0] node20329;
	wire [4-1:0] node20331;
	wire [4-1:0] node20334;
	wire [4-1:0] node20335;
	wire [4-1:0] node20337;
	wire [4-1:0] node20340;
	wire [4-1:0] node20343;
	wire [4-1:0] node20344;
	wire [4-1:0] node20345;
	wire [4-1:0] node20348;
	wire [4-1:0] node20351;
	wire [4-1:0] node20352;
	wire [4-1:0] node20356;
	wire [4-1:0] node20357;
	wire [4-1:0] node20358;
	wire [4-1:0] node20360;
	wire [4-1:0] node20362;
	wire [4-1:0] node20365;
	wire [4-1:0] node20366;
	wire [4-1:0] node20370;
	wire [4-1:0] node20372;
	wire [4-1:0] node20374;
	wire [4-1:0] node20377;
	wire [4-1:0] node20378;
	wire [4-1:0] node20379;
	wire [4-1:0] node20380;
	wire [4-1:0] node20381;
	wire [4-1:0] node20384;
	wire [4-1:0] node20386;
	wire [4-1:0] node20389;
	wire [4-1:0] node20390;
	wire [4-1:0] node20393;
	wire [4-1:0] node20396;
	wire [4-1:0] node20397;
	wire [4-1:0] node20398;
	wire [4-1:0] node20400;
	wire [4-1:0] node20403;
	wire [4-1:0] node20405;
	wire [4-1:0] node20406;
	wire [4-1:0] node20410;
	wire [4-1:0] node20411;
	wire [4-1:0] node20414;
	wire [4-1:0] node20416;
	wire [4-1:0] node20417;
	wire [4-1:0] node20421;
	wire [4-1:0] node20422;
	wire [4-1:0] node20423;
	wire [4-1:0] node20424;
	wire [4-1:0] node20426;
	wire [4-1:0] node20429;
	wire [4-1:0] node20430;
	wire [4-1:0] node20432;
	wire [4-1:0] node20436;
	wire [4-1:0] node20437;
	wire [4-1:0] node20438;
	wire [4-1:0] node20442;
	wire [4-1:0] node20445;
	wire [4-1:0] node20446;
	wire [4-1:0] node20447;
	wire [4-1:0] node20450;
	wire [4-1:0] node20451;
	wire [4-1:0] node20454;
	wire [4-1:0] node20455;
	wire [4-1:0] node20458;
	wire [4-1:0] node20461;
	wire [4-1:0] node20463;
	wire [4-1:0] node20465;
	wire [4-1:0] node20468;
	wire [4-1:0] node20469;
	wire [4-1:0] node20470;
	wire [4-1:0] node20471;
	wire [4-1:0] node20472;
	wire [4-1:0] node20473;
	wire [4-1:0] node20475;
	wire [4-1:0] node20478;
	wire [4-1:0] node20479;
	wire [4-1:0] node20480;
	wire [4-1:0] node20484;
	wire [4-1:0] node20486;
	wire [4-1:0] node20489;
	wire [4-1:0] node20490;
	wire [4-1:0] node20493;
	wire [4-1:0] node20495;
	wire [4-1:0] node20498;
	wire [4-1:0] node20499;
	wire [4-1:0] node20500;
	wire [4-1:0] node20503;
	wire [4-1:0] node20504;
	wire [4-1:0] node20507;
	wire [4-1:0] node20510;
	wire [4-1:0] node20513;
	wire [4-1:0] node20514;
	wire [4-1:0] node20515;
	wire [4-1:0] node20516;
	wire [4-1:0] node20517;
	wire [4-1:0] node20520;
	wire [4-1:0] node20523;
	wire [4-1:0] node20526;
	wire [4-1:0] node20527;
	wire [4-1:0] node20528;
	wire [4-1:0] node20530;
	wire [4-1:0] node20533;
	wire [4-1:0] node20535;
	wire [4-1:0] node20538;
	wire [4-1:0] node20539;
	wire [4-1:0] node20540;
	wire [4-1:0] node20543;
	wire [4-1:0] node20547;
	wire [4-1:0] node20548;
	wire [4-1:0] node20549;
	wire [4-1:0] node20552;
	wire [4-1:0] node20553;
	wire [4-1:0] node20554;
	wire [4-1:0] node20559;
	wire [4-1:0] node20560;
	wire [4-1:0] node20561;
	wire [4-1:0] node20564;
	wire [4-1:0] node20568;
	wire [4-1:0] node20569;
	wire [4-1:0] node20570;
	wire [4-1:0] node20571;
	wire [4-1:0] node20572;
	wire [4-1:0] node20573;
	wire [4-1:0] node20575;
	wire [4-1:0] node20579;
	wire [4-1:0] node20580;
	wire [4-1:0] node20581;
	wire [4-1:0] node20584;
	wire [4-1:0] node20588;
	wire [4-1:0] node20589;
	wire [4-1:0] node20592;
	wire [4-1:0] node20595;
	wire [4-1:0] node20596;
	wire [4-1:0] node20598;
	wire [4-1:0] node20599;
	wire [4-1:0] node20603;
	wire [4-1:0] node20604;
	wire [4-1:0] node20607;
	wire [4-1:0] node20610;
	wire [4-1:0] node20611;
	wire [4-1:0] node20612;
	wire [4-1:0] node20613;
	wire [4-1:0] node20615;
	wire [4-1:0] node20618;
	wire [4-1:0] node20620;
	wire [4-1:0] node20621;
	wire [4-1:0] node20626;
	wire [4-1:0] node20627;
	wire [4-1:0] node20628;
	wire [4-1:0] node20631;
	wire [4-1:0] node20632;
	wire [4-1:0] node20634;
	wire [4-1:0] node20637;
	wire [4-1:0] node20638;
	wire [4-1:0] node20642;
	wire [4-1:0] node20644;
	wire [4-1:0] node20647;
	wire [4-1:0] node20648;
	wire [4-1:0] node20649;
	wire [4-1:0] node20650;
	wire [4-1:0] node20651;
	wire [4-1:0] node20652;
	wire [4-1:0] node20653;
	wire [4-1:0] node20654;
	wire [4-1:0] node20655;
	wire [4-1:0] node20660;
	wire [4-1:0] node20663;
	wire [4-1:0] node20664;
	wire [4-1:0] node20668;
	wire [4-1:0] node20669;
	wire [4-1:0] node20672;
	wire [4-1:0] node20673;
	wire [4-1:0] node20676;
	wire [4-1:0] node20677;
	wire [4-1:0] node20681;
	wire [4-1:0] node20682;
	wire [4-1:0] node20683;
	wire [4-1:0] node20684;
	wire [4-1:0] node20685;
	wire [4-1:0] node20690;
	wire [4-1:0] node20691;
	wire [4-1:0] node20692;
	wire [4-1:0] node20695;
	wire [4-1:0] node20698;
	wire [4-1:0] node20701;
	wire [4-1:0] node20702;
	wire [4-1:0] node20703;
	wire [4-1:0] node20704;
	wire [4-1:0] node20705;
	wire [4-1:0] node20709;
	wire [4-1:0] node20710;
	wire [4-1:0] node20714;
	wire [4-1:0] node20715;
	wire [4-1:0] node20718;
	wire [4-1:0] node20719;
	wire [4-1:0] node20723;
	wire [4-1:0] node20725;
	wire [4-1:0] node20728;
	wire [4-1:0] node20729;
	wire [4-1:0] node20730;
	wire [4-1:0] node20731;
	wire [4-1:0] node20732;
	wire [4-1:0] node20733;
	wire [4-1:0] node20737;
	wire [4-1:0] node20738;
	wire [4-1:0] node20742;
	wire [4-1:0] node20743;
	wire [4-1:0] node20745;
	wire [4-1:0] node20748;
	wire [4-1:0] node20749;
	wire [4-1:0] node20753;
	wire [4-1:0] node20754;
	wire [4-1:0] node20755;
	wire [4-1:0] node20758;
	wire [4-1:0] node20759;
	wire [4-1:0] node20760;
	wire [4-1:0] node20764;
	wire [4-1:0] node20766;
	wire [4-1:0] node20769;
	wire [4-1:0] node20770;
	wire [4-1:0] node20773;
	wire [4-1:0] node20774;
	wire [4-1:0] node20777;
	wire [4-1:0] node20779;
	wire [4-1:0] node20782;
	wire [4-1:0] node20783;
	wire [4-1:0] node20784;
	wire [4-1:0] node20785;
	wire [4-1:0] node20786;
	wire [4-1:0] node20789;
	wire [4-1:0] node20790;
	wire [4-1:0] node20793;
	wire [4-1:0] node20796;
	wire [4-1:0] node20797;
	wire [4-1:0] node20798;
	wire [4-1:0] node20803;
	wire [4-1:0] node20804;
	wire [4-1:0] node20805;
	wire [4-1:0] node20810;
	wire [4-1:0] node20811;
	wire [4-1:0] node20812;
	wire [4-1:0] node20813;
	wire [4-1:0] node20814;
	wire [4-1:0] node20818;
	wire [4-1:0] node20819;
	wire [4-1:0] node20823;
	wire [4-1:0] node20824;
	wire [4-1:0] node20827;
	wire [4-1:0] node20830;
	wire [4-1:0] node20831;
	wire [4-1:0] node20833;
	wire [4-1:0] node20836;
	wire [4-1:0] node20837;
	wire [4-1:0] node20841;
	wire [4-1:0] node20842;
	wire [4-1:0] node20843;
	wire [4-1:0] node20844;
	wire [4-1:0] node20845;
	wire [4-1:0] node20846;
	wire [4-1:0] node20850;
	wire [4-1:0] node20851;
	wire [4-1:0] node20853;
	wire [4-1:0] node20856;
	wire [4-1:0] node20857;
	wire [4-1:0] node20859;
	wire [4-1:0] node20862;
	wire [4-1:0] node20864;
	wire [4-1:0] node20867;
	wire [4-1:0] node20868;
	wire [4-1:0] node20869;
	wire [4-1:0] node20870;
	wire [4-1:0] node20874;
	wire [4-1:0] node20875;
	wire [4-1:0] node20876;
	wire [4-1:0] node20881;
	wire [4-1:0] node20882;
	wire [4-1:0] node20883;
	wire [4-1:0] node20885;
	wire [4-1:0] node20889;
	wire [4-1:0] node20890;
	wire [4-1:0] node20891;
	wire [4-1:0] node20896;
	wire [4-1:0] node20897;
	wire [4-1:0] node20898;
	wire [4-1:0] node20899;
	wire [4-1:0] node20900;
	wire [4-1:0] node20904;
	wire [4-1:0] node20905;
	wire [4-1:0] node20906;
	wire [4-1:0] node20910;
	wire [4-1:0] node20912;
	wire [4-1:0] node20915;
	wire [4-1:0] node20916;
	wire [4-1:0] node20919;
	wire [4-1:0] node20921;
	wire [4-1:0] node20924;
	wire [4-1:0] node20925;
	wire [4-1:0] node20926;
	wire [4-1:0] node20929;
	wire [4-1:0] node20932;
	wire [4-1:0] node20934;
	wire [4-1:0] node20935;
	wire [4-1:0] node20939;
	wire [4-1:0] node20940;
	wire [4-1:0] node20941;
	wire [4-1:0] node20942;
	wire [4-1:0] node20944;
	wire [4-1:0] node20946;
	wire [4-1:0] node20949;
	wire [4-1:0] node20950;
	wire [4-1:0] node20952;
	wire [4-1:0] node20954;
	wire [4-1:0] node20957;
	wire [4-1:0] node20959;
	wire [4-1:0] node20960;
	wire [4-1:0] node20964;
	wire [4-1:0] node20965;
	wire [4-1:0] node20966;
	wire [4-1:0] node20968;
	wire [4-1:0] node20971;
	wire [4-1:0] node20973;
	wire [4-1:0] node20976;
	wire [4-1:0] node20978;
	wire [4-1:0] node20979;
	wire [4-1:0] node20983;
	wire [4-1:0] node20984;
	wire [4-1:0] node20985;
	wire [4-1:0] node20986;
	wire [4-1:0] node20989;
	wire [4-1:0] node20991;
	wire [4-1:0] node20992;
	wire [4-1:0] node20995;
	wire [4-1:0] node20998;
	wire [4-1:0] node20999;
	wire [4-1:0] node21000;
	wire [4-1:0] node21004;
	wire [4-1:0] node21007;
	wire [4-1:0] node21008;
	wire [4-1:0] node21009;
	wire [4-1:0] node21011;
	wire [4-1:0] node21015;
	wire [4-1:0] node21016;
	wire [4-1:0] node21018;
	wire [4-1:0] node21021;
	wire [4-1:0] node21023;
	wire [4-1:0] node21024;
	wire [4-1:0] node21027;
	wire [4-1:0] node21030;
	wire [4-1:0] node21031;
	wire [4-1:0] node21032;
	wire [4-1:0] node21033;
	wire [4-1:0] node21034;
	wire [4-1:0] node21035;
	wire [4-1:0] node21036;
	wire [4-1:0] node21037;
	wire [4-1:0] node21038;
	wire [4-1:0] node21039;
	wire [4-1:0] node21042;
	wire [4-1:0] node21044;
	wire [4-1:0] node21047;
	wire [4-1:0] node21050;
	wire [4-1:0] node21052;
	wire [4-1:0] node21055;
	wire [4-1:0] node21056;
	wire [4-1:0] node21057;
	wire [4-1:0] node21058;
	wire [4-1:0] node21061;
	wire [4-1:0] node21064;
	wire [4-1:0] node21065;
	wire [4-1:0] node21066;
	wire [4-1:0] node21071;
	wire [4-1:0] node21072;
	wire [4-1:0] node21075;
	wire [4-1:0] node21076;
	wire [4-1:0] node21078;
	wire [4-1:0] node21081;
	wire [4-1:0] node21082;
	wire [4-1:0] node21086;
	wire [4-1:0] node21087;
	wire [4-1:0] node21088;
	wire [4-1:0] node21089;
	wire [4-1:0] node21090;
	wire [4-1:0] node21091;
	wire [4-1:0] node21096;
	wire [4-1:0] node21099;
	wire [4-1:0] node21100;
	wire [4-1:0] node21102;
	wire [4-1:0] node21105;
	wire [4-1:0] node21106;
	wire [4-1:0] node21108;
	wire [4-1:0] node21111;
	wire [4-1:0] node21114;
	wire [4-1:0] node21115;
	wire [4-1:0] node21116;
	wire [4-1:0] node21117;
	wire [4-1:0] node21120;
	wire [4-1:0] node21123;
	wire [4-1:0] node21126;
	wire [4-1:0] node21128;
	wire [4-1:0] node21131;
	wire [4-1:0] node21132;
	wire [4-1:0] node21133;
	wire [4-1:0] node21134;
	wire [4-1:0] node21136;
	wire [4-1:0] node21139;
	wire [4-1:0] node21141;
	wire [4-1:0] node21142;
	wire [4-1:0] node21146;
	wire [4-1:0] node21147;
	wire [4-1:0] node21148;
	wire [4-1:0] node21149;
	wire [4-1:0] node21150;
	wire [4-1:0] node21155;
	wire [4-1:0] node21156;
	wire [4-1:0] node21159;
	wire [4-1:0] node21160;
	wire [4-1:0] node21164;
	wire [4-1:0] node21165;
	wire [4-1:0] node21166;
	wire [4-1:0] node21167;
	wire [4-1:0] node21172;
	wire [4-1:0] node21174;
	wire [4-1:0] node21177;
	wire [4-1:0] node21178;
	wire [4-1:0] node21179;
	wire [4-1:0] node21180;
	wire [4-1:0] node21182;
	wire [4-1:0] node21184;
	wire [4-1:0] node21187;
	wire [4-1:0] node21188;
	wire [4-1:0] node21190;
	wire [4-1:0] node21194;
	wire [4-1:0] node21195;
	wire [4-1:0] node21196;
	wire [4-1:0] node21201;
	wire [4-1:0] node21202;
	wire [4-1:0] node21203;
	wire [4-1:0] node21208;
	wire [4-1:0] node21209;
	wire [4-1:0] node21210;
	wire [4-1:0] node21211;
	wire [4-1:0] node21212;
	wire [4-1:0] node21213;
	wire [4-1:0] node21215;
	wire [4-1:0] node21216;
	wire [4-1:0] node21220;
	wire [4-1:0] node21221;
	wire [4-1:0] node21225;
	wire [4-1:0] node21226;
	wire [4-1:0] node21229;
	wire [4-1:0] node21232;
	wire [4-1:0] node21233;
	wire [4-1:0] node21234;
	wire [4-1:0] node21236;
	wire [4-1:0] node21239;
	wire [4-1:0] node21240;
	wire [4-1:0] node21241;
	wire [4-1:0] node21246;
	wire [4-1:0] node21247;
	wire [4-1:0] node21248;
	wire [4-1:0] node21252;
	wire [4-1:0] node21253;
	wire [4-1:0] node21255;
	wire [4-1:0] node21259;
	wire [4-1:0] node21260;
	wire [4-1:0] node21261;
	wire [4-1:0] node21262;
	wire [4-1:0] node21263;
	wire [4-1:0] node21264;
	wire [4-1:0] node21269;
	wire [4-1:0] node21271;
	wire [4-1:0] node21274;
	wire [4-1:0] node21275;
	wire [4-1:0] node21276;
	wire [4-1:0] node21279;
	wire [4-1:0] node21280;
	wire [4-1:0] node21284;
	wire [4-1:0] node21285;
	wire [4-1:0] node21288;
	wire [4-1:0] node21291;
	wire [4-1:0] node21292;
	wire [4-1:0] node21293;
	wire [4-1:0] node21294;
	wire [4-1:0] node21295;
	wire [4-1:0] node21298;
	wire [4-1:0] node21303;
	wire [4-1:0] node21304;
	wire [4-1:0] node21307;
	wire [4-1:0] node21308;
	wire [4-1:0] node21312;
	wire [4-1:0] node21313;
	wire [4-1:0] node21314;
	wire [4-1:0] node21315;
	wire [4-1:0] node21316;
	wire [4-1:0] node21319;
	wire [4-1:0] node21320;
	wire [4-1:0] node21322;
	wire [4-1:0] node21326;
	wire [4-1:0] node21327;
	wire [4-1:0] node21328;
	wire [4-1:0] node21331;
	wire [4-1:0] node21334;
	wire [4-1:0] node21336;
	wire [4-1:0] node21339;
	wire [4-1:0] node21340;
	wire [4-1:0] node21341;
	wire [4-1:0] node21342;
	wire [4-1:0] node21343;
	wire [4-1:0] node21348;
	wire [4-1:0] node21349;
	wire [4-1:0] node21351;
	wire [4-1:0] node21354;
	wire [4-1:0] node21355;
	wire [4-1:0] node21358;
	wire [4-1:0] node21361;
	wire [4-1:0] node21362;
	wire [4-1:0] node21364;
	wire [4-1:0] node21365;
	wire [4-1:0] node21369;
	wire [4-1:0] node21372;
	wire [4-1:0] node21373;
	wire [4-1:0] node21374;
	wire [4-1:0] node21376;
	wire [4-1:0] node21377;
	wire [4-1:0] node21379;
	wire [4-1:0] node21382;
	wire [4-1:0] node21384;
	wire [4-1:0] node21387;
	wire [4-1:0] node21388;
	wire [4-1:0] node21391;
	wire [4-1:0] node21394;
	wire [4-1:0] node21395;
	wire [4-1:0] node21396;
	wire [4-1:0] node21399;
	wire [4-1:0] node21400;
	wire [4-1:0] node21404;
	wire [4-1:0] node21406;
	wire [4-1:0] node21408;
	wire [4-1:0] node21411;
	wire [4-1:0] node21412;
	wire [4-1:0] node21413;
	wire [4-1:0] node21414;
	wire [4-1:0] node21415;
	wire [4-1:0] node21416;
	wire [4-1:0] node21417;
	wire [4-1:0] node21418;
	wire [4-1:0] node21423;
	wire [4-1:0] node21424;
	wire [4-1:0] node21425;
	wire [4-1:0] node21426;
	wire [4-1:0] node21430;
	wire [4-1:0] node21433;
	wire [4-1:0] node21435;
	wire [4-1:0] node21438;
	wire [4-1:0] node21439;
	wire [4-1:0] node21440;
	wire [4-1:0] node21441;
	wire [4-1:0] node21446;
	wire [4-1:0] node21447;
	wire [4-1:0] node21448;
	wire [4-1:0] node21450;
	wire [4-1:0] node21453;
	wire [4-1:0] node21457;
	wire [4-1:0] node21458;
	wire [4-1:0] node21459;
	wire [4-1:0] node21460;
	wire [4-1:0] node21462;
	wire [4-1:0] node21464;
	wire [4-1:0] node21467;
	wire [4-1:0] node21469;
	wire [4-1:0] node21471;
	wire [4-1:0] node21474;
	wire [4-1:0] node21475;
	wire [4-1:0] node21478;
	wire [4-1:0] node21481;
	wire [4-1:0] node21482;
	wire [4-1:0] node21484;
	wire [4-1:0] node21485;
	wire [4-1:0] node21486;
	wire [4-1:0] node21489;
	wire [4-1:0] node21493;
	wire [4-1:0] node21495;
	wire [4-1:0] node21496;
	wire [4-1:0] node21500;
	wire [4-1:0] node21501;
	wire [4-1:0] node21502;
	wire [4-1:0] node21503;
	wire [4-1:0] node21504;
	wire [4-1:0] node21506;
	wire [4-1:0] node21510;
	wire [4-1:0] node21511;
	wire [4-1:0] node21512;
	wire [4-1:0] node21513;
	wire [4-1:0] node21518;
	wire [4-1:0] node21520;
	wire [4-1:0] node21523;
	wire [4-1:0] node21524;
	wire [4-1:0] node21526;
	wire [4-1:0] node21527;
	wire [4-1:0] node21530;
	wire [4-1:0] node21533;
	wire [4-1:0] node21534;
	wire [4-1:0] node21536;
	wire [4-1:0] node21537;
	wire [4-1:0] node21540;
	wire [4-1:0] node21543;
	wire [4-1:0] node21544;
	wire [4-1:0] node21548;
	wire [4-1:0] node21549;
	wire [4-1:0] node21550;
	wire [4-1:0] node21551;
	wire [4-1:0] node21554;
	wire [4-1:0] node21557;
	wire [4-1:0] node21558;
	wire [4-1:0] node21560;
	wire [4-1:0] node21561;
	wire [4-1:0] node21566;
	wire [4-1:0] node21567;
	wire [4-1:0] node21569;
	wire [4-1:0] node21572;
	wire [4-1:0] node21573;
	wire [4-1:0] node21576;
	wire [4-1:0] node21577;
	wire [4-1:0] node21578;
	wire [4-1:0] node21583;
	wire [4-1:0] node21584;
	wire [4-1:0] node21585;
	wire [4-1:0] node21586;
	wire [4-1:0] node21587;
	wire [4-1:0] node21588;
	wire [4-1:0] node21591;
	wire [4-1:0] node21593;
	wire [4-1:0] node21596;
	wire [4-1:0] node21597;
	wire [4-1:0] node21598;
	wire [4-1:0] node21602;
	wire [4-1:0] node21603;
	wire [4-1:0] node21607;
	wire [4-1:0] node21608;
	wire [4-1:0] node21609;
	wire [4-1:0] node21612;
	wire [4-1:0] node21613;
	wire [4-1:0] node21614;
	wire [4-1:0] node21618;
	wire [4-1:0] node21619;
	wire [4-1:0] node21622;
	wire [4-1:0] node21625;
	wire [4-1:0] node21627;
	wire [4-1:0] node21629;
	wire [4-1:0] node21631;
	wire [4-1:0] node21634;
	wire [4-1:0] node21635;
	wire [4-1:0] node21636;
	wire [4-1:0] node21637;
	wire [4-1:0] node21638;
	wire [4-1:0] node21641;
	wire [4-1:0] node21644;
	wire [4-1:0] node21647;
	wire [4-1:0] node21648;
	wire [4-1:0] node21649;
	wire [4-1:0] node21651;
	wire [4-1:0] node21655;
	wire [4-1:0] node21656;
	wire [4-1:0] node21659;
	wire [4-1:0] node21661;
	wire [4-1:0] node21664;
	wire [4-1:0] node21665;
	wire [4-1:0] node21666;
	wire [4-1:0] node21667;
	wire [4-1:0] node21670;
	wire [4-1:0] node21672;
	wire [4-1:0] node21676;
	wire [4-1:0] node21677;
	wire [4-1:0] node21679;
	wire [4-1:0] node21680;
	wire [4-1:0] node21684;
	wire [4-1:0] node21686;
	wire [4-1:0] node21688;
	wire [4-1:0] node21691;
	wire [4-1:0] node21692;
	wire [4-1:0] node21693;
	wire [4-1:0] node21694;
	wire [4-1:0] node21696;
	wire [4-1:0] node21697;
	wire [4-1:0] node21701;
	wire [4-1:0] node21702;
	wire [4-1:0] node21703;
	wire [4-1:0] node21704;
	wire [4-1:0] node21709;
	wire [4-1:0] node21712;
	wire [4-1:0] node21713;
	wire [4-1:0] node21714;
	wire [4-1:0] node21717;
	wire [4-1:0] node21718;
	wire [4-1:0] node21722;
	wire [4-1:0] node21723;
	wire [4-1:0] node21724;
	wire [4-1:0] node21728;
	wire [4-1:0] node21730;
	wire [4-1:0] node21733;
	wire [4-1:0] node21734;
	wire [4-1:0] node21735;
	wire [4-1:0] node21736;
	wire [4-1:0] node21739;
	wire [4-1:0] node21741;
	wire [4-1:0] node21744;
	wire [4-1:0] node21745;
	wire [4-1:0] node21747;
	wire [4-1:0] node21749;
	wire [4-1:0] node21753;
	wire [4-1:0] node21754;
	wire [4-1:0] node21755;
	wire [4-1:0] node21757;
	wire [4-1:0] node21760;
	wire [4-1:0] node21762;
	wire [4-1:0] node21765;
	wire [4-1:0] node21766;
	wire [4-1:0] node21767;
	wire [4-1:0] node21771;
	wire [4-1:0] node21774;
	wire [4-1:0] node21775;
	wire [4-1:0] node21776;
	wire [4-1:0] node21777;
	wire [4-1:0] node21778;
	wire [4-1:0] node21779;
	wire [4-1:0] node21780;
	wire [4-1:0] node21781;
	wire [4-1:0] node21783;
	wire [4-1:0] node21786;
	wire [4-1:0] node21788;
	wire [4-1:0] node21789;
	wire [4-1:0] node21792;
	wire [4-1:0] node21795;
	wire [4-1:0] node21796;
	wire [4-1:0] node21799;
	wire [4-1:0] node21802;
	wire [4-1:0] node21803;
	wire [4-1:0] node21804;
	wire [4-1:0] node21808;
	wire [4-1:0] node21809;
	wire [4-1:0] node21811;
	wire [4-1:0] node21815;
	wire [4-1:0] node21816;
	wire [4-1:0] node21817;
	wire [4-1:0] node21818;
	wire [4-1:0] node21820;
	wire [4-1:0] node21821;
	wire [4-1:0] node21826;
	wire [4-1:0] node21828;
	wire [4-1:0] node21831;
	wire [4-1:0] node21832;
	wire [4-1:0] node21833;
	wire [4-1:0] node21834;
	wire [4-1:0] node21838;
	wire [4-1:0] node21839;
	wire [4-1:0] node21840;
	wire [4-1:0] node21843;
	wire [4-1:0] node21847;
	wire [4-1:0] node21849;
	wire [4-1:0] node21850;
	wire [4-1:0] node21851;
	wire [4-1:0] node21854;
	wire [4-1:0] node21858;
	wire [4-1:0] node21859;
	wire [4-1:0] node21860;
	wire [4-1:0] node21861;
	wire [4-1:0] node21862;
	wire [4-1:0] node21865;
	wire [4-1:0] node21867;
	wire [4-1:0] node21868;
	wire [4-1:0] node21872;
	wire [4-1:0] node21873;
	wire [4-1:0] node21876;
	wire [4-1:0] node21879;
	wire [4-1:0] node21880;
	wire [4-1:0] node21881;
	wire [4-1:0] node21884;
	wire [4-1:0] node21885;
	wire [4-1:0] node21887;
	wire [4-1:0] node21891;
	wire [4-1:0] node21893;
	wire [4-1:0] node21894;
	wire [4-1:0] node21898;
	wire [4-1:0] node21899;
	wire [4-1:0] node21900;
	wire [4-1:0] node21901;
	wire [4-1:0] node21902;
	wire [4-1:0] node21903;
	wire [4-1:0] node21908;
	wire [4-1:0] node21909;
	wire [4-1:0] node21912;
	wire [4-1:0] node21913;
	wire [4-1:0] node21917;
	wire [4-1:0] node21918;
	wire [4-1:0] node21919;
	wire [4-1:0] node21922;
	wire [4-1:0] node21926;
	wire [4-1:0] node21927;
	wire [4-1:0] node21928;
	wire [4-1:0] node21931;
	wire [4-1:0] node21934;
	wire [4-1:0] node21935;
	wire [4-1:0] node21938;
	wire [4-1:0] node21940;
	wire [4-1:0] node21943;
	wire [4-1:0] node21944;
	wire [4-1:0] node21945;
	wire [4-1:0] node21946;
	wire [4-1:0] node21947;
	wire [4-1:0] node21949;
	wire [4-1:0] node21950;
	wire [4-1:0] node21951;
	wire [4-1:0] node21956;
	wire [4-1:0] node21957;
	wire [4-1:0] node21958;
	wire [4-1:0] node21959;
	wire [4-1:0] node21964;
	wire [4-1:0] node21966;
	wire [4-1:0] node21969;
	wire [4-1:0] node21970;
	wire [4-1:0] node21971;
	wire [4-1:0] node21975;
	wire [4-1:0] node21976;
	wire [4-1:0] node21977;
	wire [4-1:0] node21978;
	wire [4-1:0] node21983;
	wire [4-1:0] node21986;
	wire [4-1:0] node21987;
	wire [4-1:0] node21988;
	wire [4-1:0] node21989;
	wire [4-1:0] node21990;
	wire [4-1:0] node21992;
	wire [4-1:0] node21996;
	wire [4-1:0] node21998;
	wire [4-1:0] node21999;
	wire [4-1:0] node22003;
	wire [4-1:0] node22004;
	wire [4-1:0] node22006;
	wire [4-1:0] node22008;
	wire [4-1:0] node22011;
	wire [4-1:0] node22012;
	wire [4-1:0] node22016;
	wire [4-1:0] node22017;
	wire [4-1:0] node22018;
	wire [4-1:0] node22019;
	wire [4-1:0] node22020;
	wire [4-1:0] node22024;
	wire [4-1:0] node22025;
	wire [4-1:0] node22029;
	wire [4-1:0] node22030;
	wire [4-1:0] node22033;
	wire [4-1:0] node22034;
	wire [4-1:0] node22038;
	wire [4-1:0] node22040;
	wire [4-1:0] node22042;
	wire [4-1:0] node22043;
	wire [4-1:0] node22047;
	wire [4-1:0] node22048;
	wire [4-1:0] node22049;
	wire [4-1:0] node22050;
	wire [4-1:0] node22051;
	wire [4-1:0] node22053;
	wire [4-1:0] node22057;
	wire [4-1:0] node22058;
	wire [4-1:0] node22060;
	wire [4-1:0] node22063;
	wire [4-1:0] node22064;
	wire [4-1:0] node22068;
	wire [4-1:0] node22069;
	wire [4-1:0] node22070;
	wire [4-1:0] node22072;
	wire [4-1:0] node22073;
	wire [4-1:0] node22077;
	wire [4-1:0] node22078;
	wire [4-1:0] node22080;
	wire [4-1:0] node22084;
	wire [4-1:0] node22086;
	wire [4-1:0] node22087;
	wire [4-1:0] node22090;
	wire [4-1:0] node22093;
	wire [4-1:0] node22094;
	wire [4-1:0] node22095;
	wire [4-1:0] node22096;
	wire [4-1:0] node22097;
	wire [4-1:0] node22100;
	wire [4-1:0] node22104;
	wire [4-1:0] node22105;
	wire [4-1:0] node22107;
	wire [4-1:0] node22111;
	wire [4-1:0] node22112;
	wire [4-1:0] node22113;
	wire [4-1:0] node22115;
	wire [4-1:0] node22119;
	wire [4-1:0] node22120;
	wire [4-1:0] node22121;
	wire [4-1:0] node22126;
	wire [4-1:0] node22127;
	wire [4-1:0] node22128;
	wire [4-1:0] node22129;
	wire [4-1:0] node22130;
	wire [4-1:0] node22131;
	wire [4-1:0] node22132;
	wire [4-1:0] node22134;
	wire [4-1:0] node22137;
	wire [4-1:0] node22139;
	wire [4-1:0] node22142;
	wire [4-1:0] node22143;
	wire [4-1:0] node22144;
	wire [4-1:0] node22146;
	wire [4-1:0] node22151;
	wire [4-1:0] node22152;
	wire [4-1:0] node22153;
	wire [4-1:0] node22156;
	wire [4-1:0] node22158;
	wire [4-1:0] node22159;
	wire [4-1:0] node22163;
	wire [4-1:0] node22165;
	wire [4-1:0] node22168;
	wire [4-1:0] node22169;
	wire [4-1:0] node22170;
	wire [4-1:0] node22171;
	wire [4-1:0] node22175;
	wire [4-1:0] node22176;
	wire [4-1:0] node22177;
	wire [4-1:0] node22179;
	wire [4-1:0] node22183;
	wire [4-1:0] node22186;
	wire [4-1:0] node22187;
	wire [4-1:0] node22188;
	wire [4-1:0] node22189;
	wire [4-1:0] node22190;
	wire [4-1:0] node22195;
	wire [4-1:0] node22198;
	wire [4-1:0] node22199;
	wire [4-1:0] node22201;
	wire [4-1:0] node22202;
	wire [4-1:0] node22206;
	wire [4-1:0] node22208;
	wire [4-1:0] node22210;
	wire [4-1:0] node22213;
	wire [4-1:0] node22214;
	wire [4-1:0] node22215;
	wire [4-1:0] node22216;
	wire [4-1:0] node22217;
	wire [4-1:0] node22218;
	wire [4-1:0] node22219;
	wire [4-1:0] node22224;
	wire [4-1:0] node22227;
	wire [4-1:0] node22228;
	wire [4-1:0] node22231;
	wire [4-1:0] node22233;
	wire [4-1:0] node22235;
	wire [4-1:0] node22238;
	wire [4-1:0] node22239;
	wire [4-1:0] node22240;
	wire [4-1:0] node22243;
	wire [4-1:0] node22244;
	wire [4-1:0] node22248;
	wire [4-1:0] node22249;
	wire [4-1:0] node22251;
	wire [4-1:0] node22255;
	wire [4-1:0] node22256;
	wire [4-1:0] node22257;
	wire [4-1:0] node22258;
	wire [4-1:0] node22261;
	wire [4-1:0] node22264;
	wire [4-1:0] node22266;
	wire [4-1:0] node22269;
	wire [4-1:0] node22270;
	wire [4-1:0] node22271;
	wire [4-1:0] node22275;
	wire [4-1:0] node22276;
	wire [4-1:0] node22280;
	wire [4-1:0] node22281;
	wire [4-1:0] node22282;
	wire [4-1:0] node22283;
	wire [4-1:0] node22284;
	wire [4-1:0] node22285;
	wire [4-1:0] node22287;
	wire [4-1:0] node22288;
	wire [4-1:0] node22293;
	wire [4-1:0] node22294;
	wire [4-1:0] node22295;
	wire [4-1:0] node22297;
	wire [4-1:0] node22301;
	wire [4-1:0] node22302;
	wire [4-1:0] node22303;
	wire [4-1:0] node22308;
	wire [4-1:0] node22309;
	wire [4-1:0] node22310;
	wire [4-1:0] node22314;
	wire [4-1:0] node22315;
	wire [4-1:0] node22316;
	wire [4-1:0] node22318;
	wire [4-1:0] node22322;
	wire [4-1:0] node22323;
	wire [4-1:0] node22327;
	wire [4-1:0] node22328;
	wire [4-1:0] node22329;
	wire [4-1:0] node22330;
	wire [4-1:0] node22332;
	wire [4-1:0] node22333;
	wire [4-1:0] node22336;
	wire [4-1:0] node22340;
	wire [4-1:0] node22341;
	wire [4-1:0] node22344;
	wire [4-1:0] node22347;
	wire [4-1:0] node22348;
	wire [4-1:0] node22351;
	wire [4-1:0] node22352;
	wire [4-1:0] node22353;
	wire [4-1:0] node22355;
	wire [4-1:0] node22359;
	wire [4-1:0] node22360;
	wire [4-1:0] node22364;
	wire [4-1:0] node22365;
	wire [4-1:0] node22366;
	wire [4-1:0] node22367;
	wire [4-1:0] node22368;
	wire [4-1:0] node22369;
	wire [4-1:0] node22370;
	wire [4-1:0] node22373;
	wire [4-1:0] node22376;
	wire [4-1:0] node22378;
	wire [4-1:0] node22381;
	wire [4-1:0] node22382;
	wire [4-1:0] node22383;
	wire [4-1:0] node22386;
	wire [4-1:0] node22389;
	wire [4-1:0] node22392;
	wire [4-1:0] node22393;
	wire [4-1:0] node22397;
	wire [4-1:0] node22398;
	wire [4-1:0] node22400;
	wire [4-1:0] node22402;
	wire [4-1:0] node22403;
	wire [4-1:0] node22407;
	wire [4-1:0] node22408;
	wire [4-1:0] node22412;
	wire [4-1:0] node22413;
	wire [4-1:0] node22414;
	wire [4-1:0] node22415;
	wire [4-1:0] node22417;
	wire [4-1:0] node22421;
	wire [4-1:0] node22422;
	wire [4-1:0] node22424;
	wire [4-1:0] node22427;
	wire [4-1:0] node22428;
	wire [4-1:0] node22432;
	wire [4-1:0] node22433;
	wire [4-1:0] node22435;
	wire [4-1:0] node22438;
	wire [4-1:0] node22439;
	wire [4-1:0] node22442;

	assign outp = (inp[13]) ? node11254 : node1;
		assign node1 = (inp[9]) ? node5649 : node2;
			assign node2 = (inp[4]) ? node2920 : node3;
				assign node3 = (inp[12]) ? node1461 : node4;
					assign node4 = (inp[10]) ? node798 : node5;
						assign node5 = (inp[14]) ? node405 : node6;
							assign node6 = (inp[8]) ? node222 : node7;
								assign node7 = (inp[0]) ? node123 : node8;
									assign node8 = (inp[15]) ? node74 : node9;
										assign node9 = (inp[3]) ? node41 : node10;
											assign node10 = (inp[1]) ? node24 : node11;
												assign node11 = (inp[5]) ? node19 : node12;
													assign node12 = (inp[2]) ? 4'b1111 : node13;
														assign node13 = (inp[11]) ? 4'b0111 : node14;
															assign node14 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node19 = (inp[11]) ? 4'b0110 : node20;
														assign node20 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node24 = (inp[5]) ? node30 : node25;
													assign node25 = (inp[7]) ? node27 : 4'b1110;
														assign node27 = (inp[6]) ? 4'b1111 : 4'b0111;
													assign node30 = (inp[11]) ? node34 : node31;
														assign node31 = (inp[7]) ? 4'b1110 : 4'b0110;
														assign node34 = (inp[6]) ? node38 : node35;
															assign node35 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node38 = (inp[2]) ? 4'b0110 : 4'b1110;
											assign node41 = (inp[5]) ? node55 : node42;
												assign node42 = (inp[1]) ? node46 : node43;
													assign node43 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node46 = (inp[7]) ? node52 : node47;
														assign node47 = (inp[2]) ? node49 : 4'b0111;
															assign node49 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node52 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node55 = (inp[11]) ? node67 : node56;
													assign node56 = (inp[2]) ? node62 : node57;
														assign node57 = (inp[6]) ? node59 : 4'b1101;
															assign node59 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node62 = (inp[6]) ? node64 : 4'b0101;
															assign node64 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node67 = (inp[6]) ? node71 : node68;
														assign node68 = (inp[2]) ? 4'b1101 : 4'b0101;
														assign node71 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node74 = (inp[5]) ? node96 : node75;
											assign node75 = (inp[3]) ? node83 : node76;
												assign node76 = (inp[7]) ? node80 : node77;
													assign node77 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node80 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node83 = (inp[7]) ? node93 : node84;
													assign node84 = (inp[2]) ? node90 : node85;
														assign node85 = (inp[1]) ? 4'b1101 : node86;
															assign node86 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node90 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node93 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node96 = (inp[3]) ? node108 : node97;
												assign node97 = (inp[11]) ? node103 : node98;
													assign node98 = (inp[7]) ? 4'b1101 : node99;
														assign node99 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node103 = (inp[1]) ? node105 : 4'b1100;
														assign node105 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node108 = (inp[11]) ? node114 : node109;
													assign node109 = (inp[1]) ? node111 : 4'b1110;
														assign node111 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node114 = (inp[6]) ? 4'b1111 : node115;
														assign node115 = (inp[2]) ? node119 : node116;
															assign node116 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node119 = (inp[1]) ? 4'b1111 : 4'b0110;
									assign node123 = (inp[15]) ? node177 : node124;
										assign node124 = (inp[3]) ? node150 : node125;
											assign node125 = (inp[6]) ? node137 : node126;
												assign node126 = (inp[11]) ? node134 : node127;
													assign node127 = (inp[7]) ? node131 : node128;
														assign node128 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node131 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node134 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node137 = (inp[11]) ? node145 : node138;
													assign node138 = (inp[7]) ? node142 : node139;
														assign node139 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node142 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node145 = (inp[7]) ? node147 : 4'b1101;
														assign node147 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node150 = (inp[5]) ? node166 : node151;
												assign node151 = (inp[6]) ? node159 : node152;
													assign node152 = (inp[11]) ? node154 : 4'b1101;
														assign node154 = (inp[2]) ? node156 : 4'b0101;
															assign node156 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node159 = (inp[1]) ? node161 : 4'b0100;
														assign node161 = (inp[7]) ? 4'b1101 : node162;
															assign node162 = (inp[11]) ? 4'b1100 : 4'b0100;
												assign node166 = (inp[7]) ? node168 : 4'b1110;
													assign node168 = (inp[2]) ? 4'b0111 : node169;
														assign node169 = (inp[11]) ? node173 : node170;
															assign node170 = (inp[6]) ? 4'b0110 : 4'b1110;
															assign node173 = (inp[6]) ? 4'b1110 : 4'b0110;
										assign node177 = (inp[5]) ? node201 : node178;
											assign node178 = (inp[6]) ? node190 : node179;
												assign node179 = (inp[11]) ? node183 : node180;
													assign node180 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node183 = (inp[1]) ? node185 : 4'b0111;
														assign node185 = (inp[2]) ? 4'b0110 : node186;
															assign node186 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node190 = (inp[11]) ? node196 : node191;
													assign node191 = (inp[2]) ? node193 : 4'b0110;
														assign node193 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node196 = (inp[7]) ? node198 : 4'b1110;
														assign node198 = (inp[2]) ? 4'b0111 : 4'b1110;
											assign node201 = (inp[3]) ? node211 : node202;
												assign node202 = (inp[2]) ? node206 : node203;
													assign node203 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node206 = (inp[7]) ? node208 : 4'b1110;
														assign node208 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node211 = (inp[7]) ? node217 : node212;
													assign node212 = (inp[2]) ? 4'b0100 : node213;
														assign node213 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node217 = (inp[1]) ? node219 : 4'b1101;
														assign node219 = (inp[6]) ? 4'b0101 : 4'b1101;
								assign node222 = (inp[3]) ? node306 : node223;
									assign node223 = (inp[2]) ? node257 : node224;
										assign node224 = (inp[7]) ? node244 : node225;
											assign node225 = (inp[0]) ? node237 : node226;
												assign node226 = (inp[15]) ? node232 : node227;
													assign node227 = (inp[11]) ? node229 : 4'b1110;
														assign node229 = (inp[6]) ? 4'b1110 : 4'b0110;
													assign node232 = (inp[1]) ? 4'b0100 : node233;
														assign node233 = (inp[5]) ? 4'b1100 : 4'b0100;
												assign node237 = (inp[15]) ? 4'b1110 : node238;
													assign node238 = (inp[5]) ? 4'b1100 : node239;
														assign node239 = (inp[11]) ? 4'b0100 : 4'b1100;
											assign node244 = (inp[15]) ? node252 : node245;
												assign node245 = (inp[0]) ? 4'b1101 : node246;
													assign node246 = (inp[1]) ? node248 : 4'b1111;
														assign node248 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node252 = (inp[0]) ? 4'b0111 : node253;
													assign node253 = (inp[1]) ? 4'b1101 : 4'b0101;
										assign node257 = (inp[7]) ? node277 : node258;
											assign node258 = (inp[1]) ? node264 : node259;
												assign node259 = (inp[11]) ? 4'b0111 : node260;
													assign node260 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node264 = (inp[0]) ? node268 : node265;
													assign node265 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node268 = (inp[15]) ? node274 : node269;
														assign node269 = (inp[11]) ? node271 : 4'b0101;
															assign node271 = (inp[6]) ? 4'b0101 : 4'b1101;
														assign node274 = (inp[6]) ? 4'b1111 : 4'b0111;
											assign node277 = (inp[11]) ? node289 : node278;
												assign node278 = (inp[1]) ? node282 : node279;
													assign node279 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node282 = (inp[6]) ? 4'b1110 : node283;
														assign node283 = (inp[0]) ? 4'b0110 : node284;
															assign node284 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node289 = (inp[1]) ? node297 : node290;
													assign node290 = (inp[6]) ? 4'b1110 : node291;
														assign node291 = (inp[15]) ? node293 : 4'b0100;
															assign node293 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node297 = (inp[6]) ? 4'b0100 : node298;
														assign node298 = (inp[0]) ? node302 : node299;
															assign node299 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node302 = (inp[15]) ? 4'b1110 : 4'b1100;
									assign node306 = (inp[6]) ? node360 : node307;
										assign node307 = (inp[1]) ? node337 : node308;
											assign node308 = (inp[11]) ? node318 : node309;
												assign node309 = (inp[15]) ? node315 : node310;
													assign node310 = (inp[5]) ? node312 : 4'b1100;
														assign node312 = (inp[0]) ? 4'b1111 : 4'b1100;
													assign node315 = (inp[7]) ? 4'b1111 : 4'b1101;
												assign node318 = (inp[5]) ? node330 : node319;
													assign node319 = (inp[7]) ? node327 : node320;
														assign node320 = (inp[2]) ? node324 : node321;
															assign node321 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node324 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node327 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node330 = (inp[15]) ? node334 : node331;
														assign node331 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node334 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node337 = (inp[11]) ? node347 : node338;
												assign node338 = (inp[7]) ? node340 : 4'b1110;
													assign node340 = (inp[2]) ? 4'b0100 : node341;
														assign node341 = (inp[0]) ? node343 : 4'b0101;
															assign node343 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node347 = (inp[0]) ? node357 : node348;
													assign node348 = (inp[5]) ? node354 : node349;
														assign node349 = (inp[7]) ? node351 : 4'b1101;
															assign node351 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node354 = (inp[2]) ? 4'b1101 : 4'b0100;
													assign node357 = (inp[15]) ? 4'b1111 : 4'b1101;
										assign node360 = (inp[11]) ? node374 : node361;
											assign node361 = (inp[5]) ? node371 : node362;
												assign node362 = (inp[0]) ? node366 : node363;
													assign node363 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node366 = (inp[15]) ? node368 : 4'b1100;
														assign node368 = (inp[1]) ? 4'b1111 : 4'b0111;
												assign node371 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node374 = (inp[1]) ? node394 : node375;
												assign node375 = (inp[15]) ? node383 : node376;
													assign node376 = (inp[0]) ? node378 : 4'b1111;
														assign node378 = (inp[7]) ? node380 : 4'b1110;
															assign node380 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node383 = (inp[2]) ? node387 : node384;
														assign node384 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node387 = (inp[5]) ? node391 : node388;
															assign node388 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node391 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node394 = (inp[15]) ? node398 : node395;
													assign node395 = (inp[7]) ? 4'b0101 : 4'b0111;
													assign node398 = (inp[7]) ? node402 : node399;
														assign node399 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node402 = (inp[0]) ? 4'b0110 : 4'b0100;
							assign node405 = (inp[2]) ? node595 : node406;
								assign node406 = (inp[7]) ? node490 : node407;
									assign node407 = (inp[8]) ? node445 : node408;
										assign node408 = (inp[5]) ? node426 : node409;
											assign node409 = (inp[11]) ? node417 : node410;
												assign node410 = (inp[6]) ? 4'b0110 : node411;
													assign node411 = (inp[15]) ? 4'b1110 : node412;
														assign node412 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node417 = (inp[6]) ? 4'b1110 : node418;
													assign node418 = (inp[0]) ? node422 : node419;
														assign node419 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node422 = (inp[15]) ? 4'b0110 : 4'b0100;
											assign node426 = (inp[11]) ? node442 : node427;
												assign node427 = (inp[6]) ? node435 : node428;
													assign node428 = (inp[15]) ? node430 : 4'b1110;
														assign node430 = (inp[1]) ? node432 : 4'b1100;
															assign node432 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node435 = (inp[1]) ? 4'b0110 : node436;
														assign node436 = (inp[3]) ? node438 : 4'b0100;
															assign node438 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node442 = (inp[6]) ? 4'b1100 : 4'b0100;
										assign node445 = (inp[5]) ? node469 : node446;
											assign node446 = (inp[11]) ? node462 : node447;
												assign node447 = (inp[15]) ? node451 : node448;
													assign node448 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node451 = (inp[0]) ? node457 : node452;
														assign node452 = (inp[1]) ? 4'b0101 : node453;
															assign node453 = (inp[6]) ? 4'b0101 : 4'b1101;
														assign node457 = (inp[3]) ? node459 : 4'b1111;
															assign node459 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node462 = (inp[0]) ? node466 : node463;
													assign node463 = (inp[15]) ? 4'b1101 : 4'b0111;
													assign node466 = (inp[15]) ? 4'b0111 : 4'b1101;
											assign node469 = (inp[0]) ? node481 : node470;
												assign node470 = (inp[11]) ? node476 : node471;
													assign node471 = (inp[15]) ? node473 : 4'b1111;
														assign node473 = (inp[1]) ? 4'b1111 : 4'b0111;
													assign node476 = (inp[1]) ? 4'b0111 : node477;
														assign node477 = (inp[6]) ? 4'b1111 : 4'b0111;
												assign node481 = (inp[1]) ? 4'b0101 : node482;
													assign node482 = (inp[6]) ? node484 : 4'b1111;
														assign node484 = (inp[11]) ? 4'b1111 : node485;
															assign node485 = (inp[3]) ? 4'b0101 : 4'b0111;
									assign node490 = (inp[8]) ? node544 : node491;
										assign node491 = (inp[0]) ? node519 : node492;
											assign node492 = (inp[6]) ? node512 : node493;
												assign node493 = (inp[15]) ? node503 : node494;
													assign node494 = (inp[5]) ? node498 : node495;
														assign node495 = (inp[3]) ? 4'b1111 : 4'b0111;
														assign node498 = (inp[3]) ? node500 : 4'b1111;
															assign node500 = (inp[1]) ? 4'b0101 : 4'b0101;
													assign node503 = (inp[3]) ? node509 : node504;
														assign node504 = (inp[5]) ? 4'b0101 : node505;
															assign node505 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node509 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node512 = (inp[5]) ? node514 : 4'b1101;
													assign node514 = (inp[11]) ? node516 : 4'b1111;
														assign node516 = (inp[1]) ? 4'b0111 : 4'b1111;
											assign node519 = (inp[15]) ? node529 : node520;
												assign node520 = (inp[5]) ? node526 : node521;
													assign node521 = (inp[3]) ? node523 : 4'b1101;
														assign node523 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node526 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node529 = (inp[3]) ? node537 : node530;
													assign node530 = (inp[11]) ? 4'b0111 : node531;
														assign node531 = (inp[6]) ? 4'b1111 : node532;
															assign node532 = (inp[1]) ? 4'b0111 : 4'b1111;
													assign node537 = (inp[5]) ? node539 : 4'b1111;
														assign node539 = (inp[6]) ? node541 : 4'b1101;
															assign node541 = (inp[1]) ? 4'b1101 : 4'b0101;
										assign node544 = (inp[1]) ? node572 : node545;
											assign node545 = (inp[6]) ? node557 : node546;
												assign node546 = (inp[11]) ? node552 : node547;
													assign node547 = (inp[15]) ? node549 : 4'b1110;
														assign node549 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node552 = (inp[0]) ? 4'b0100 : node553;
														assign node553 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node557 = (inp[0]) ? node567 : node558;
													assign node558 = (inp[15]) ? node564 : node559;
														assign node559 = (inp[3]) ? node561 : 4'b1110;
															assign node561 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node564 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node567 = (inp[3]) ? 4'b1100 : node568;
														assign node568 = (inp[5]) ? 4'b1110 : 4'b1100;
											assign node572 = (inp[0]) ? node586 : node573;
												assign node573 = (inp[15]) ? node579 : node574;
													assign node574 = (inp[3]) ? 4'b0100 : node575;
														assign node575 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node579 = (inp[3]) ? node581 : 4'b1100;
														assign node581 = (inp[5]) ? node583 : 4'b1100;
															assign node583 = (inp[6]) ? 4'b1110 : 4'b0110;
												assign node586 = (inp[15]) ? 4'b0110 : node587;
													assign node587 = (inp[3]) ? 4'b1100 : node588;
														assign node588 = (inp[11]) ? node590 : 4'b0100;
															assign node590 = (inp[6]) ? 4'b0100 : 4'b1100;
								assign node595 = (inp[5]) ? node691 : node596;
									assign node596 = (inp[15]) ? node644 : node597;
										assign node597 = (inp[0]) ? node625 : node598;
											assign node598 = (inp[6]) ? node612 : node599;
												assign node599 = (inp[11]) ? node607 : node600;
													assign node600 = (inp[7]) ? node602 : 4'b1110;
														assign node602 = (inp[1]) ? node604 : 4'b1110;
															assign node604 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node607 = (inp[8]) ? 4'b0110 : node608;
														assign node608 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node612 = (inp[7]) ? node620 : node613;
													assign node613 = (inp[8]) ? node615 : 4'b1110;
														assign node615 = (inp[1]) ? 4'b0111 : node616;
															assign node616 = (inp[11]) ? 4'b1111 : 4'b0111;
													assign node620 = (inp[8]) ? 4'b1110 : node621;
														assign node621 = (inp[3]) ? 4'b0111 : 4'b1111;
											assign node625 = (inp[7]) ? node637 : node626;
												assign node626 = (inp[8]) ? node628 : 4'b1100;
													assign node628 = (inp[1]) ? node630 : 4'b1101;
														assign node630 = (inp[6]) ? node634 : node631;
															assign node631 = (inp[3]) ? 4'b0101 : 4'b1101;
															assign node634 = (inp[3]) ? 4'b1101 : 4'b0101;
												assign node637 = (inp[8]) ? node639 : 4'b0101;
													assign node639 = (inp[1]) ? 4'b1100 : node640;
														assign node640 = (inp[11]) ? 4'b1100 : 4'b0100;
										assign node644 = (inp[0]) ? node668 : node645;
											assign node645 = (inp[11]) ? node655 : node646;
												assign node646 = (inp[6]) ? node652 : node647;
													assign node647 = (inp[1]) ? node649 : 4'b1101;
														assign node649 = (inp[7]) ? 4'b0101 : 4'b1100;
													assign node652 = (inp[1]) ? 4'b1101 : 4'b0101;
												assign node655 = (inp[6]) ? node665 : node656;
													assign node656 = (inp[1]) ? 4'b1101 : node657;
														assign node657 = (inp[7]) ? node661 : node658;
															assign node658 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node661 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node665 = (inp[3]) ? 4'b0101 : 4'b1101;
											assign node668 = (inp[1]) ? node680 : node669;
												assign node669 = (inp[11]) ? node675 : node670;
													assign node670 = (inp[8]) ? node672 : 4'b1111;
														assign node672 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node675 = (inp[8]) ? node677 : 4'b1110;
														assign node677 = (inp[6]) ? 4'b1111 : 4'b0111;
												assign node680 = (inp[3]) ? node686 : node681;
													assign node681 = (inp[6]) ? node683 : 4'b0111;
														assign node683 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node686 = (inp[7]) ? 4'b1110 : node687;
														assign node687 = (inp[8]) ? 4'b0111 : 4'b0110;
									assign node691 = (inp[6]) ? node743 : node692;
										assign node692 = (inp[11]) ? node716 : node693;
											assign node693 = (inp[1]) ? node701 : node694;
												assign node694 = (inp[8]) ? 4'b1111 : node695;
													assign node695 = (inp[0]) ? node697 : 4'b1101;
														assign node697 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node701 = (inp[8]) ? node709 : node702;
													assign node702 = (inp[15]) ? node704 : 4'b0101;
														assign node704 = (inp[3]) ? node706 : 4'b0111;
															assign node706 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node709 = (inp[15]) ? node711 : 4'b0101;
														assign node711 = (inp[0]) ? node713 : 4'b0110;
															assign node713 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node716 = (inp[1]) ? node730 : node717;
												assign node717 = (inp[15]) ? node723 : node718;
													assign node718 = (inp[7]) ? node720 : 4'b0111;
														assign node720 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node723 = (inp[0]) ? node725 : 4'b0110;
														assign node725 = (inp[3]) ? node727 : 4'b0110;
															assign node727 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node730 = (inp[8]) ? node736 : node731;
													assign node731 = (inp[7]) ? 4'b1111 : node732;
														assign node732 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node736 = (inp[7]) ? 4'b1110 : node737;
														assign node737 = (inp[0]) ? node739 : 4'b1111;
															assign node739 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node743 = (inp[0]) ? node775 : node744;
											assign node744 = (inp[15]) ? node760 : node745;
												assign node745 = (inp[3]) ? node753 : node746;
													assign node746 = (inp[1]) ? node748 : 4'b1111;
														assign node748 = (inp[7]) ? node750 : 4'b1110;
															assign node750 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node753 = (inp[8]) ? 4'b1100 : node754;
														assign node754 = (inp[7]) ? 4'b0101 : node755;
															assign node755 = (inp[11]) ? 4'b1100 : 4'b0100;
												assign node760 = (inp[3]) ? node768 : node761;
													assign node761 = (inp[8]) ? 4'b1101 : node762;
														assign node762 = (inp[7]) ? node764 : 4'b0100;
															assign node764 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node768 = (inp[8]) ? 4'b0111 : node769;
														assign node769 = (inp[11]) ? 4'b1111 : node770;
															assign node770 = (inp[1]) ? 4'b1111 : 4'b0111;
											assign node775 = (inp[11]) ? node787 : node776;
												assign node776 = (inp[1]) ? node780 : node777;
													assign node777 = (inp[3]) ? 4'b0111 : 4'b0110;
													assign node780 = (inp[7]) ? node784 : node781;
														assign node781 = (inp[8]) ? 4'b1111 : 4'b0110;
														assign node784 = (inp[15]) ? 4'b1110 : 4'b1111;
												assign node787 = (inp[1]) ? 4'b0110 : node788;
													assign node788 = (inp[8]) ? 4'b1111 : node789;
														assign node789 = (inp[3]) ? node793 : node790;
															assign node790 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node793 = (inp[15]) ? 4'b1100 : 4'b1110;
						assign node798 = (inp[6]) ? node1132 : node799;
							assign node799 = (inp[11]) ? node963 : node800;
								assign node800 = (inp[1]) ? node886 : node801;
									assign node801 = (inp[3]) ? node845 : node802;
										assign node802 = (inp[14]) ? node830 : node803;
											assign node803 = (inp[8]) ? node819 : node804;
												assign node804 = (inp[2]) ? node812 : node805;
													assign node805 = (inp[7]) ? node807 : 4'b1111;
														assign node807 = (inp[15]) ? node809 : 4'b1100;
															assign node809 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node812 = (inp[5]) ? 4'b1110 : node813;
														assign node813 = (inp[0]) ? 4'b1100 : node814;
															assign node814 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node819 = (inp[0]) ? node823 : node820;
													assign node820 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node823 = (inp[15]) ? 4'b1111 : node824;
														assign node824 = (inp[7]) ? 4'b1100 : node825;
															assign node825 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node830 = (inp[2]) ? node836 : node831;
												assign node831 = (inp[8]) ? node833 : 4'b1101;
													assign node833 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node836 = (inp[7]) ? node840 : node837;
													assign node837 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node840 = (inp[0]) ? node842 : 4'b1111;
														assign node842 = (inp[15]) ? 4'b1110 : 4'b1100;
										assign node845 = (inp[14]) ? node861 : node846;
											assign node846 = (inp[2]) ? node852 : node847;
												assign node847 = (inp[5]) ? 4'b1111 : node848;
													assign node848 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node852 = (inp[5]) ? node854 : 4'b1111;
													assign node854 = (inp[0]) ? node856 : 4'b1100;
														assign node856 = (inp[15]) ? node858 : 4'b1111;
															assign node858 = (inp[7]) ? 4'b1101 : 4'b1100;
											assign node861 = (inp[7]) ? node873 : node862;
												assign node862 = (inp[8]) ? node868 : node863;
													assign node863 = (inp[0]) ? 4'b1100 : node864;
														assign node864 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node868 = (inp[15]) ? node870 : 4'b1101;
														assign node870 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node873 = (inp[8]) ? node877 : node874;
													assign node874 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node877 = (inp[0]) ? 4'b1110 : node878;
														assign node878 = (inp[5]) ? node882 : node879;
															assign node879 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node882 = (inp[15]) ? 4'b1110 : 4'b1100;
									assign node886 = (inp[7]) ? node922 : node887;
										assign node887 = (inp[8]) ? node903 : node888;
											assign node888 = (inp[2]) ? node894 : node889;
												assign node889 = (inp[5]) ? node891 : 4'b1110;
													assign node891 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node894 = (inp[0]) ? node898 : node895;
													assign node895 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node898 = (inp[15]) ? node900 : 4'b1100;
														assign node900 = (inp[3]) ? 4'b1100 : 4'b1110;
											assign node903 = (inp[2]) ? node913 : node904;
												assign node904 = (inp[14]) ? node908 : node905;
													assign node905 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node908 = (inp[5]) ? 4'b0111 : node909;
														assign node909 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node913 = (inp[14]) ? 4'b0111 : node914;
													assign node914 = (inp[15]) ? node916 : 4'b0111;
														assign node916 = (inp[3]) ? node918 : 4'b0101;
															assign node918 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node922 = (inp[8]) ? node946 : node923;
											assign node923 = (inp[14]) ? node933 : node924;
												assign node924 = (inp[2]) ? node928 : node925;
													assign node925 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node928 = (inp[3]) ? node930 : 4'b0111;
														assign node930 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node933 = (inp[5]) ? node941 : node934;
													assign node934 = (inp[0]) ? node938 : node935;
														assign node935 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node938 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node941 = (inp[3]) ? node943 : 4'b0101;
														assign node943 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node946 = (inp[15]) ? node954 : node947;
												assign node947 = (inp[0]) ? node951 : node948;
													assign node948 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node951 = (inp[3]) ? 4'b0101 : 4'b0100;
												assign node954 = (inp[5]) ? node956 : 4'b0110;
													assign node956 = (inp[14]) ? node958 : 4'b0110;
														assign node958 = (inp[3]) ? node960 : 4'b0100;
															assign node960 = (inp[0]) ? 4'b0100 : 4'b0110;
								assign node963 = (inp[1]) ? node1053 : node964;
									assign node964 = (inp[15]) ? node1010 : node965;
										assign node965 = (inp[0]) ? node985 : node966;
											assign node966 = (inp[3]) ? node974 : node967;
												assign node967 = (inp[8]) ? 4'b0111 : node968;
													assign node968 = (inp[14]) ? 4'b0110 : node969;
														assign node969 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node974 = (inp[5]) ? node978 : node975;
													assign node975 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node978 = (inp[2]) ? node980 : 4'b0101;
														assign node980 = (inp[14]) ? node982 : 4'b0100;
															assign node982 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node985 = (inp[8]) ? node993 : node986;
												assign node986 = (inp[7]) ? 4'b0101 : node987;
													assign node987 = (inp[3]) ? node989 : 4'b0100;
														assign node989 = (inp[14]) ? 4'b0110 : 4'b0100;
												assign node993 = (inp[2]) ? node1005 : node994;
													assign node994 = (inp[5]) ? node1000 : node995;
														assign node995 = (inp[14]) ? 4'b0100 : node996;
															assign node996 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node1000 = (inp[14]) ? 4'b0101 : node1001;
															assign node1001 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node1005 = (inp[5]) ? 4'b0111 : node1006;
														assign node1006 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node1010 = (inp[0]) ? node1028 : node1011;
											assign node1011 = (inp[3]) ? node1021 : node1012;
												assign node1012 = (inp[5]) ? node1014 : 4'b0101;
													assign node1014 = (inp[2]) ? 4'b0100 : node1015;
														assign node1015 = (inp[14]) ? 4'b0101 : node1016;
															assign node1016 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node1021 = (inp[5]) ? 4'b0111 : node1022;
													assign node1022 = (inp[7]) ? node1024 : 4'b0100;
														assign node1024 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node1028 = (inp[14]) ? node1046 : node1029;
												assign node1029 = (inp[5]) ? node1039 : node1030;
													assign node1030 = (inp[3]) ? node1032 : 4'b0111;
														assign node1032 = (inp[8]) ? node1036 : node1033;
															assign node1033 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node1036 = (inp[2]) ? 4'b0110 : 4'b0110;
													assign node1039 = (inp[3]) ? 4'b0101 : node1040;
														assign node1040 = (inp[7]) ? 4'b0110 : node1041;
															assign node1041 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node1046 = (inp[8]) ? node1050 : node1047;
													assign node1047 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node1050 = (inp[7]) ? 4'b0110 : 4'b0111;
									assign node1053 = (inp[8]) ? node1085 : node1054;
										assign node1054 = (inp[7]) ? node1068 : node1055;
											assign node1055 = (inp[3]) ? node1061 : node1056;
												assign node1056 = (inp[15]) ? 4'b0100 : node1057;
													assign node1057 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node1061 = (inp[15]) ? node1063 : 4'b0110;
													assign node1063 = (inp[0]) ? node1065 : 4'b0101;
														assign node1065 = (inp[14]) ? 4'b0110 : 4'b0111;
											assign node1068 = (inp[14]) ? node1078 : node1069;
												assign node1069 = (inp[2]) ? node1075 : node1070;
													assign node1070 = (inp[3]) ? 4'b0110 : node1071;
														assign node1071 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node1075 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node1078 = (inp[3]) ? node1080 : 4'b1001;
													assign node1080 = (inp[2]) ? 4'b1001 : node1081;
														assign node1081 = (inp[5]) ? 4'b1001 : 4'b1011;
										assign node1085 = (inp[7]) ? node1103 : node1086;
											assign node1086 = (inp[2]) ? node1096 : node1087;
												assign node1087 = (inp[14]) ? node1093 : node1088;
													assign node1088 = (inp[15]) ? 4'b0100 : node1089;
														assign node1089 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node1093 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node1096 = (inp[15]) ? node1100 : node1097;
													assign node1097 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node1100 = (inp[0]) ? 4'b1011 : 4'b1001;
											assign node1103 = (inp[2]) ? node1119 : node1104;
												assign node1104 = (inp[14]) ? node1114 : node1105;
													assign node1105 = (inp[15]) ? node1111 : node1106;
														assign node1106 = (inp[3]) ? 4'b1001 : node1107;
															assign node1107 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node1111 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node1114 = (inp[3]) ? node1116 : 4'b1000;
														assign node1116 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node1119 = (inp[0]) ? node1125 : node1120;
													assign node1120 = (inp[14]) ? 4'b1010 : node1121;
														assign node1121 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node1125 = (inp[15]) ? node1129 : node1126;
														assign node1126 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node1129 = (inp[3]) ? 4'b1000 : 4'b1010;
							assign node1132 = (inp[11]) ? node1280 : node1133;
								assign node1133 = (inp[1]) ? node1199 : node1134;
									assign node1134 = (inp[15]) ? node1170 : node1135;
										assign node1135 = (inp[0]) ? node1159 : node1136;
											assign node1136 = (inp[5]) ? node1148 : node1137;
												assign node1137 = (inp[7]) ? node1141 : node1138;
													assign node1138 = (inp[3]) ? 4'b0110 : 4'b0111;
													assign node1141 = (inp[2]) ? 4'b0111 : node1142;
														assign node1142 = (inp[14]) ? 4'b0110 : node1143;
															assign node1143 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node1148 = (inp[3]) ? node1152 : node1149;
													assign node1149 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node1152 = (inp[14]) ? 4'b0101 : node1153;
														assign node1153 = (inp[7]) ? node1155 : 4'b0100;
															assign node1155 = (inp[8]) ? 4'b0101 : 4'b0100;
											assign node1159 = (inp[3]) ? 4'b0111 : node1160;
												assign node1160 = (inp[8]) ? 4'b0100 : node1161;
													assign node1161 = (inp[2]) ? 4'b0101 : node1162;
														assign node1162 = (inp[5]) ? node1164 : 4'b0100;
															assign node1164 = (inp[7]) ? 4'b0101 : 4'b0100;
										assign node1170 = (inp[0]) ? node1186 : node1171;
											assign node1171 = (inp[7]) ? node1175 : node1172;
												assign node1172 = (inp[8]) ? 4'b0101 : 4'b0110;
												assign node1175 = (inp[8]) ? node1181 : node1176;
													assign node1176 = (inp[2]) ? 4'b0101 : node1177;
														assign node1177 = (inp[3]) ? 4'b0101 : 4'b0100;
													assign node1181 = (inp[14]) ? 4'b0100 : node1182;
														assign node1182 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node1186 = (inp[3]) ? node1196 : node1187;
												assign node1187 = (inp[8]) ? node1189 : 4'b0111;
													assign node1189 = (inp[2]) ? 4'b0111 : node1190;
														assign node1190 = (inp[7]) ? node1192 : 4'b0110;
															assign node1192 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node1196 = (inp[2]) ? 4'b0110 : 4'b0101;
									assign node1199 = (inp[7]) ? node1247 : node1200;
										assign node1200 = (inp[8]) ? node1220 : node1201;
											assign node1201 = (inp[2]) ? node1215 : node1202;
												assign node1202 = (inp[14]) ? node1212 : node1203;
													assign node1203 = (inp[5]) ? 4'b0101 : node1204;
														assign node1204 = (inp[15]) ? node1208 : node1205;
															assign node1205 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node1208 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node1212 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node1215 = (inp[0]) ? node1217 : 4'b0100;
													assign node1217 = (inp[15]) ? 4'b0110 : 4'b0100;
											assign node1220 = (inp[2]) ? node1234 : node1221;
												assign node1221 = (inp[14]) ? node1229 : node1222;
													assign node1222 = (inp[15]) ? node1224 : 4'b0110;
														assign node1224 = (inp[5]) ? node1226 : 4'b0100;
															assign node1226 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node1229 = (inp[5]) ? 4'b1001 : node1230;
														assign node1230 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node1234 = (inp[14]) ? 4'b1001 : node1235;
													assign node1235 = (inp[0]) ? node1239 : node1236;
														assign node1236 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node1239 = (inp[5]) ? node1243 : node1240;
															assign node1240 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node1243 = (inp[3]) ? 4'b1001 : 4'b1001;
										assign node1247 = (inp[8]) ? node1263 : node1248;
											assign node1248 = (inp[14]) ? node1256 : node1249;
												assign node1249 = (inp[2]) ? node1253 : node1250;
													assign node1250 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node1253 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node1256 = (inp[0]) ? 4'b1011 : node1257;
													assign node1257 = (inp[3]) ? node1259 : 4'b1011;
														assign node1259 = (inp[2]) ? 4'b1001 : 4'b1011;
											assign node1263 = (inp[2]) ? node1273 : node1264;
												assign node1264 = (inp[14]) ? node1270 : node1265;
													assign node1265 = (inp[3]) ? 4'b1001 : node1266;
														assign node1266 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node1270 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node1273 = (inp[0]) ? 4'b1000 : node1274;
													assign node1274 = (inp[15]) ? node1276 : 4'b1010;
														assign node1276 = (inp[5]) ? 4'b1010 : 4'b1000;
								assign node1280 = (inp[1]) ? node1372 : node1281;
									assign node1281 = (inp[5]) ? node1321 : node1282;
										assign node1282 = (inp[7]) ? node1304 : node1283;
											assign node1283 = (inp[14]) ? node1293 : node1284;
												assign node1284 = (inp[0]) ? node1290 : node1285;
													assign node1285 = (inp[2]) ? 4'b1011 : node1286;
														assign node1286 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node1290 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node1293 = (inp[8]) ? node1297 : node1294;
													assign node1294 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node1297 = (inp[3]) ? node1299 : 4'b1001;
														assign node1299 = (inp[15]) ? node1301 : 4'b1011;
															assign node1301 = (inp[0]) ? 4'b1011 : 4'b1001;
											assign node1304 = (inp[14]) ? node1316 : node1305;
												assign node1305 = (inp[8]) ? node1311 : node1306;
													assign node1306 = (inp[0]) ? 4'b1011 : node1307;
														assign node1307 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node1311 = (inp[3]) ? node1313 : 4'b1001;
														assign node1313 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node1316 = (inp[8]) ? 4'b1010 : node1317;
													assign node1317 = (inp[15]) ? 4'b1011 : 4'b1001;
										assign node1321 = (inp[3]) ? node1355 : node1322;
											assign node1322 = (inp[2]) ? node1340 : node1323;
												assign node1323 = (inp[7]) ? node1329 : node1324;
													assign node1324 = (inp[0]) ? 4'b1000 : node1325;
														assign node1325 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node1329 = (inp[14]) ? node1333 : node1330;
														assign node1330 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node1333 = (inp[15]) ? node1337 : node1334;
															assign node1334 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node1337 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node1340 = (inp[7]) ? node1348 : node1341;
													assign node1341 = (inp[8]) ? node1343 : 4'b1010;
														assign node1343 = (inp[0]) ? 4'b1011 : node1344;
															assign node1344 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node1348 = (inp[15]) ? node1352 : node1349;
														assign node1349 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node1352 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node1355 = (inp[7]) ? node1359 : node1356;
												assign node1356 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node1359 = (inp[15]) ? node1369 : node1360;
													assign node1360 = (inp[0]) ? node1362 : 4'b1001;
														assign node1362 = (inp[8]) ? node1366 : node1363;
															assign node1363 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node1366 = (inp[2]) ? 4'b1010 : 4'b1010;
													assign node1369 = (inp[0]) ? 4'b1000 : 4'b1010;
									assign node1372 = (inp[7]) ? node1418 : node1373;
										assign node1373 = (inp[8]) ? node1399 : node1374;
											assign node1374 = (inp[2]) ? node1390 : node1375;
												assign node1375 = (inp[14]) ? node1383 : node1376;
													assign node1376 = (inp[0]) ? 4'b1011 : node1377;
														assign node1377 = (inp[15]) ? 4'b1001 : node1378;
															assign node1378 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node1383 = (inp[15]) ? node1385 : 4'b1010;
														assign node1385 = (inp[3]) ? node1387 : 4'b1000;
															assign node1387 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node1390 = (inp[15]) ? node1392 : 4'b1000;
													assign node1392 = (inp[0]) ? node1394 : 4'b1000;
														assign node1394 = (inp[3]) ? node1396 : 4'b1010;
															assign node1396 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node1399 = (inp[14]) ? node1407 : node1400;
												assign node1400 = (inp[2]) ? node1402 : 4'b1000;
													assign node1402 = (inp[5]) ? 4'b0011 : node1403;
														assign node1403 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node1407 = (inp[0]) ? node1409 : 4'b0011;
													assign node1409 = (inp[5]) ? node1411 : 4'b0001;
														assign node1411 = (inp[3]) ? node1415 : node1412;
															assign node1412 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node1415 = (inp[15]) ? 4'b0001 : 4'b0011;
										assign node1418 = (inp[8]) ? node1442 : node1419;
											assign node1419 = (inp[14]) ? node1429 : node1420;
												assign node1420 = (inp[2]) ? node1424 : node1421;
													assign node1421 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node1424 = (inp[5]) ? node1426 : 4'b0001;
														assign node1426 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node1429 = (inp[5]) ? node1437 : node1430;
													assign node1430 = (inp[2]) ? node1434 : node1431;
														assign node1431 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node1434 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node1437 = (inp[0]) ? node1439 : 4'b0011;
														assign node1439 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node1442 = (inp[2]) ? node1450 : node1443;
												assign node1443 = (inp[14]) ? node1447 : node1444;
													assign node1444 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node1447 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node1450 = (inp[5]) ? 4'b0000 : node1451;
													assign node1451 = (inp[3]) ? node1455 : node1452;
														assign node1452 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node1455 = (inp[0]) ? node1457 : 4'b0000;
															assign node1457 = (inp[15]) ? 4'b0010 : 4'b0000;
					assign node1461 = (inp[10]) ? node2143 : node1462;
						assign node1462 = (inp[11]) ? node1794 : node1463;
							assign node1463 = (inp[6]) ? node1627 : node1464;
								assign node1464 = (inp[1]) ? node1546 : node1465;
									assign node1465 = (inp[7]) ? node1507 : node1466;
										assign node1466 = (inp[8]) ? node1490 : node1467;
											assign node1467 = (inp[14]) ? node1477 : node1468;
												assign node1468 = (inp[2]) ? node1474 : node1469;
													assign node1469 = (inp[0]) ? node1471 : 4'b1101;
														assign node1471 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node1474 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node1477 = (inp[3]) ? node1479 : 4'b1100;
													assign node1479 = (inp[15]) ? node1485 : node1480;
														assign node1480 = (inp[2]) ? 4'b1100 : node1481;
															assign node1481 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node1485 = (inp[5]) ? 4'b1100 : node1486;
															assign node1486 = (inp[0]) ? 4'b1110 : 4'b1100;
											assign node1490 = (inp[15]) ? node1498 : node1491;
												assign node1491 = (inp[2]) ? node1493 : 4'b1100;
													assign node1493 = (inp[0]) ? 4'b1101 : node1494;
														assign node1494 = (inp[14]) ? 4'b1101 : 4'b1111;
												assign node1498 = (inp[14]) ? node1502 : node1499;
													assign node1499 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node1502 = (inp[3]) ? node1504 : 4'b1111;
														assign node1504 = (inp[0]) ? 4'b1101 : 4'b1111;
										assign node1507 = (inp[8]) ? node1529 : node1508;
											assign node1508 = (inp[14]) ? node1518 : node1509;
												assign node1509 = (inp[2]) ? node1515 : node1510;
													assign node1510 = (inp[15]) ? node1512 : 4'b1110;
														assign node1512 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node1515 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node1518 = (inp[0]) ? node1522 : node1519;
													assign node1519 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node1522 = (inp[15]) ? 4'b1111 : node1523;
														assign node1523 = (inp[3]) ? node1525 : 4'b1101;
															assign node1525 = (inp[2]) ? 4'b1101 : 4'b1111;
											assign node1529 = (inp[2]) ? node1541 : node1530;
												assign node1530 = (inp[14]) ? 4'b1100 : node1531;
													assign node1531 = (inp[3]) ? 4'b1101 : node1532;
														assign node1532 = (inp[15]) ? node1536 : node1533;
															assign node1533 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node1536 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node1541 = (inp[0]) ? node1543 : 4'b1110;
													assign node1543 = (inp[15]) ? 4'b1110 : 4'b1100;
									assign node1546 = (inp[8]) ? node1592 : node1547;
										assign node1547 = (inp[7]) ? node1571 : node1548;
											assign node1548 = (inp[14]) ? node1562 : node1549;
												assign node1549 = (inp[2]) ? node1557 : node1550;
													assign node1550 = (inp[0]) ? node1552 : 4'b1111;
														assign node1552 = (inp[15]) ? node1554 : 4'b1101;
															assign node1554 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node1557 = (inp[15]) ? 4'b1110 : node1558;
														assign node1558 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node1562 = (inp[2]) ? 4'b1100 : node1563;
													assign node1563 = (inp[0]) ? node1565 : 4'b1110;
														assign node1565 = (inp[3]) ? 4'b1100 : node1566;
															assign node1566 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node1571 = (inp[14]) ? node1581 : node1572;
												assign node1572 = (inp[2]) ? 4'b0101 : node1573;
													assign node1573 = (inp[0]) ? 4'b1110 : node1574;
														assign node1574 = (inp[3]) ? 4'b1110 : node1575;
															assign node1575 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node1581 = (inp[0]) ? 4'b0101 : node1582;
													assign node1582 = (inp[2]) ? node1586 : node1583;
														assign node1583 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node1586 = (inp[5]) ? node1588 : 4'b0101;
															assign node1588 = (inp[15]) ? 4'b0111 : 4'b0101;
										assign node1592 = (inp[7]) ? node1606 : node1593;
											assign node1593 = (inp[15]) ? 4'b0101 : node1594;
												assign node1594 = (inp[3]) ? node1598 : node1595;
													assign node1595 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node1598 = (inp[2]) ? node1600 : 4'b1110;
														assign node1600 = (inp[5]) ? node1602 : 4'b0111;
															assign node1602 = (inp[0]) ? 4'b0111 : 4'b0101;
											assign node1606 = (inp[2]) ? node1618 : node1607;
												assign node1607 = (inp[14]) ? node1611 : node1608;
													assign node1608 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node1611 = (inp[0]) ? 4'b0100 : node1612;
														assign node1612 = (inp[15]) ? node1614 : 4'b0110;
															assign node1614 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node1618 = (inp[15]) ? node1622 : node1619;
													assign node1619 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node1622 = (inp[0]) ? node1624 : 4'b0100;
														assign node1624 = (inp[3]) ? 4'b0100 : 4'b0110;
								assign node1627 = (inp[1]) ? node1723 : node1628;
									assign node1628 = (inp[2]) ? node1678 : node1629;
										assign node1629 = (inp[3]) ? node1661 : node1630;
											assign node1630 = (inp[15]) ? node1646 : node1631;
												assign node1631 = (inp[0]) ? node1641 : node1632;
													assign node1632 = (inp[8]) ? node1636 : node1633;
														assign node1633 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node1636 = (inp[5]) ? node1638 : 4'b0110;
															assign node1638 = (inp[14]) ? 4'b0110 : 4'b0110;
													assign node1641 = (inp[7]) ? 4'b0101 : node1642;
														assign node1642 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node1646 = (inp[0]) ? node1654 : node1647;
													assign node1647 = (inp[7]) ? 4'b0100 : node1648;
														assign node1648 = (inp[5]) ? 4'b0100 : node1649;
															assign node1649 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node1654 = (inp[8]) ? 4'b0111 : node1655;
														assign node1655 = (inp[7]) ? node1657 : 4'b0110;
															assign node1657 = (inp[14]) ? 4'b0111 : 4'b0110;
											assign node1661 = (inp[15]) ? node1671 : node1662;
												assign node1662 = (inp[0]) ? node1668 : node1663;
													assign node1663 = (inp[5]) ? node1665 : 4'b0111;
														assign node1665 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node1668 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node1671 = (inp[0]) ? 4'b0111 : node1672;
													assign node1672 = (inp[8]) ? node1674 : 4'b0111;
														assign node1674 = (inp[5]) ? 4'b0110 : 4'b0100;
										assign node1678 = (inp[8]) ? node1698 : node1679;
											assign node1679 = (inp[7]) ? node1687 : node1680;
												assign node1680 = (inp[5]) ? node1682 : 4'b0100;
													assign node1682 = (inp[3]) ? 4'b0100 : node1683;
														assign node1683 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node1687 = (inp[3]) ? node1693 : node1688;
													assign node1688 = (inp[15]) ? 4'b0101 : node1689;
														assign node1689 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node1693 = (inp[5]) ? 4'b0111 : node1694;
														assign node1694 = (inp[15]) ? 4'b0111 : 4'b0101;
											assign node1698 = (inp[7]) ? node1712 : node1699;
												assign node1699 = (inp[15]) ? node1707 : node1700;
													assign node1700 = (inp[0]) ? node1702 : 4'b0111;
														assign node1702 = (inp[3]) ? node1704 : 4'b0101;
															assign node1704 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node1707 = (inp[0]) ? node1709 : 4'b0101;
														assign node1709 = (inp[14]) ? 4'b0101 : 4'b0111;
												assign node1712 = (inp[3]) ? node1718 : node1713;
													assign node1713 = (inp[0]) ? 4'b0110 : node1714;
														assign node1714 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node1718 = (inp[14]) ? node1720 : 4'b0100;
														assign node1720 = (inp[5]) ? 4'b0100 : 4'b0110;
									assign node1723 = (inp[8]) ? node1761 : node1724;
										assign node1724 = (inp[7]) ? node1742 : node1725;
											assign node1725 = (inp[2]) ? node1735 : node1726;
												assign node1726 = (inp[14]) ? node1732 : node1727;
													assign node1727 = (inp[0]) ? 4'b0111 : node1728;
														assign node1728 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node1732 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node1735 = (inp[0]) ? node1739 : node1736;
													assign node1736 = (inp[14]) ? 4'b0110 : 4'b0100;
													assign node1739 = (inp[14]) ? 4'b0100 : 4'b0110;
											assign node1742 = (inp[2]) ? node1754 : node1743;
												assign node1743 = (inp[14]) ? 4'b1011 : node1744;
													assign node1744 = (inp[5]) ? node1750 : node1745;
														assign node1745 = (inp[0]) ? node1747 : 4'b0110;
															assign node1747 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node1750 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node1754 = (inp[15]) ? node1756 : 4'b1001;
													assign node1756 = (inp[3]) ? 4'b1011 : node1757;
														assign node1757 = (inp[0]) ? 4'b1011 : 4'b1001;
										assign node1761 = (inp[7]) ? node1779 : node1762;
											assign node1762 = (inp[2]) ? node1768 : node1763;
												assign node1763 = (inp[14]) ? 4'b1011 : node1764;
													assign node1764 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node1768 = (inp[15]) ? node1774 : node1769;
													assign node1769 = (inp[5]) ? node1771 : 4'b1011;
														assign node1771 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node1774 = (inp[0]) ? node1776 : 4'b1001;
														assign node1776 = (inp[14]) ? 4'b1001 : 4'b1011;
											assign node1779 = (inp[15]) ? node1789 : node1780;
												assign node1780 = (inp[0]) ? node1784 : node1781;
													assign node1781 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node1784 = (inp[14]) ? 4'b1000 : node1785;
														assign node1785 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node1789 = (inp[0]) ? 4'b1010 : node1790;
													assign node1790 = (inp[14]) ? 4'b1010 : 4'b1000;
							assign node1794 = (inp[6]) ? node1956 : node1795;
								assign node1795 = (inp[1]) ? node1869 : node1796;
									assign node1796 = (inp[8]) ? node1830 : node1797;
										assign node1797 = (inp[7]) ? node1813 : node1798;
											assign node1798 = (inp[14]) ? node1806 : node1799;
												assign node1799 = (inp[2]) ? node1801 : 4'b0101;
													assign node1801 = (inp[5]) ? node1803 : 4'b0100;
														assign node1803 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node1806 = (inp[0]) ? node1808 : 4'b0110;
													assign node1808 = (inp[15]) ? node1810 : 4'b0100;
														assign node1810 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node1813 = (inp[14]) ? node1823 : node1814;
												assign node1814 = (inp[2]) ? 4'b0101 : node1815;
													assign node1815 = (inp[5]) ? node1817 : 4'b0100;
														assign node1817 = (inp[0]) ? node1819 : 4'b0110;
															assign node1819 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node1823 = (inp[5]) ? node1825 : 4'b0101;
													assign node1825 = (inp[0]) ? 4'b0111 : node1826;
														assign node1826 = (inp[3]) ? 4'b0111 : 4'b0101;
										assign node1830 = (inp[7]) ? node1856 : node1831;
											assign node1831 = (inp[2]) ? node1849 : node1832;
												assign node1832 = (inp[14]) ? node1844 : node1833;
													assign node1833 = (inp[5]) ? node1839 : node1834;
														assign node1834 = (inp[3]) ? node1836 : 4'b0110;
															assign node1836 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node1839 = (inp[3]) ? node1841 : 4'b0100;
															assign node1841 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node1844 = (inp[3]) ? node1846 : 4'b0101;
														assign node1846 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node1849 = (inp[15]) ? node1851 : 4'b0111;
													assign node1851 = (inp[0]) ? 4'b0111 : node1852;
														assign node1852 = (inp[3]) ? 4'b0111 : 4'b0101;
											assign node1856 = (inp[14]) ? node1862 : node1857;
												assign node1857 = (inp[2]) ? node1859 : 4'b0111;
													assign node1859 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node1862 = (inp[15]) ? 4'b0110 : node1863;
													assign node1863 = (inp[0]) ? 4'b0100 : node1864;
														assign node1864 = (inp[3]) ? 4'b0100 : 4'b0110;
									assign node1869 = (inp[8]) ? node1913 : node1870;
										assign node1870 = (inp[7]) ? node1892 : node1871;
											assign node1871 = (inp[14]) ? node1883 : node1872;
												assign node1872 = (inp[2]) ? node1878 : node1873;
													assign node1873 = (inp[15]) ? 4'b0101 : node1874;
														assign node1874 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node1878 = (inp[0]) ? node1880 : 4'b0110;
														assign node1880 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node1883 = (inp[5]) ? 4'b0100 : node1884;
													assign node1884 = (inp[0]) ? node1888 : node1885;
														assign node1885 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node1888 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node1892 = (inp[2]) ? node1904 : node1893;
												assign node1893 = (inp[14]) ? 4'b1011 : node1894;
													assign node1894 = (inp[5]) ? node1900 : node1895;
														assign node1895 = (inp[3]) ? node1897 : 4'b0100;
															assign node1897 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node1900 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node1904 = (inp[0]) ? 4'b1001 : node1905;
													assign node1905 = (inp[15]) ? 4'b1001 : node1906;
														assign node1906 = (inp[3]) ? node1908 : 4'b1011;
															assign node1908 = (inp[14]) ? 4'b1001 : 4'b1011;
										assign node1913 = (inp[7]) ? node1927 : node1914;
											assign node1914 = (inp[14]) ? 4'b1001 : node1915;
												assign node1915 = (inp[2]) ? node1919 : node1916;
													assign node1916 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node1919 = (inp[15]) ? node1921 : 4'b1001;
														assign node1921 = (inp[5]) ? node1923 : 4'b1011;
															assign node1923 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node1927 = (inp[14]) ? node1941 : node1928;
												assign node1928 = (inp[2]) ? node1936 : node1929;
													assign node1929 = (inp[15]) ? node1931 : 4'b1001;
														assign node1931 = (inp[5]) ? node1933 : 4'b1011;
															assign node1933 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node1936 = (inp[15]) ? node1938 : 4'b1010;
														assign node1938 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node1941 = (inp[5]) ? node1949 : node1942;
													assign node1942 = (inp[2]) ? node1944 : 4'b1010;
														assign node1944 = (inp[3]) ? 4'b1010 : node1945;
															assign node1945 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node1949 = (inp[2]) ? node1951 : 4'b1000;
														assign node1951 = (inp[3]) ? node1953 : 4'b1010;
															assign node1953 = (inp[0]) ? 4'b1000 : 4'b1000;
								assign node1956 = (inp[1]) ? node2054 : node1957;
									assign node1957 = (inp[3]) ? node2009 : node1958;
										assign node1958 = (inp[7]) ? node1978 : node1959;
											assign node1959 = (inp[8]) ? node1969 : node1960;
												assign node1960 = (inp[14]) ? node1964 : node1961;
													assign node1961 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node1964 = (inp[2]) ? 4'b1000 : node1965;
														assign node1965 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node1969 = (inp[2]) ? node1975 : node1970;
													assign node1970 = (inp[14]) ? node1972 : 4'b1000;
														assign node1972 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node1975 = (inp[14]) ? 4'b1001 : 4'b1011;
											assign node1978 = (inp[8]) ? node1994 : node1979;
												assign node1979 = (inp[14]) ? node1985 : node1980;
													assign node1980 = (inp[15]) ? 4'b1000 : node1981;
														assign node1981 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node1985 = (inp[2]) ? 4'b1011 : node1986;
														assign node1986 = (inp[15]) ? node1990 : node1987;
															assign node1987 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node1990 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node1994 = (inp[2]) ? node2002 : node1995;
													assign node1995 = (inp[14]) ? node1997 : 4'b1001;
														assign node1997 = (inp[15]) ? 4'b1000 : node1998;
															assign node1998 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node2002 = (inp[0]) ? node2006 : node2003;
														assign node2003 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node2006 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node2009 = (inp[15]) ? node2033 : node2010;
											assign node2010 = (inp[7]) ? node2022 : node2011;
												assign node2011 = (inp[8]) ? node2019 : node2012;
													assign node2012 = (inp[14]) ? node2016 : node2013;
														assign node2013 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node2016 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node2019 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node2022 = (inp[5]) ? 4'b1011 : node2023;
													assign node2023 = (inp[0]) ? node2029 : node2024;
														assign node2024 = (inp[14]) ? 4'b1011 : node2025;
															assign node2025 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node2029 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node2033 = (inp[7]) ? node2045 : node2034;
												assign node2034 = (inp[5]) ? 4'b1010 : node2035;
													assign node2035 = (inp[0]) ? node2039 : node2036;
														assign node2036 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node2039 = (inp[14]) ? 4'b1010 : node2040;
															assign node2040 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node2045 = (inp[5]) ? node2047 : 4'b1010;
													assign node2047 = (inp[0]) ? 4'b1001 : node2048;
														assign node2048 = (inp[8]) ? node2050 : 4'b1011;
															assign node2050 = (inp[14]) ? 4'b1010 : 4'b1011;
									assign node2054 = (inp[8]) ? node2090 : node2055;
										assign node2055 = (inp[7]) ? node2069 : node2056;
											assign node2056 = (inp[2]) ? 4'b1010 : node2057;
												assign node2057 = (inp[14]) ? node2065 : node2058;
													assign node2058 = (inp[0]) ? node2060 : 4'b1011;
														assign node2060 = (inp[15]) ? node2062 : 4'b1001;
															assign node2062 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node2065 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node2069 = (inp[2]) ? node2081 : node2070;
												assign node2070 = (inp[14]) ? node2078 : node2071;
													assign node2071 = (inp[15]) ? node2073 : 4'b1000;
														assign node2073 = (inp[5]) ? 4'b1010 : node2074;
															assign node2074 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node2078 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node2081 = (inp[3]) ? node2083 : 4'b0011;
													assign node2083 = (inp[15]) ? node2085 : 4'b0001;
														assign node2085 = (inp[14]) ? 4'b0011 : node2086;
															assign node2086 = (inp[0]) ? 4'b0001 : 4'b0001;
										assign node2090 = (inp[7]) ? node2114 : node2091;
											assign node2091 = (inp[14]) ? node2099 : node2092;
												assign node2092 = (inp[2]) ? node2096 : node2093;
													assign node2093 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node2096 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node2099 = (inp[2]) ? node2109 : node2100;
													assign node2100 = (inp[5]) ? 4'b0011 : node2101;
														assign node2101 = (inp[15]) ? node2105 : node2102;
															assign node2102 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node2105 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node2109 = (inp[15]) ? node2111 : 4'b0001;
														assign node2111 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node2114 = (inp[2]) ? node2128 : node2115;
												assign node2115 = (inp[14]) ? node2125 : node2116;
													assign node2116 = (inp[0]) ? node2122 : node2117;
														assign node2117 = (inp[15]) ? node2119 : 4'b0011;
															assign node2119 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node2122 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node2125 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node2128 = (inp[5]) ? node2138 : node2129;
													assign node2129 = (inp[3]) ? node2131 : 4'b0010;
														assign node2131 = (inp[15]) ? node2135 : node2132;
															assign node2132 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node2135 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node2138 = (inp[3]) ? node2140 : 4'b0000;
														assign node2140 = (inp[15]) ? 4'b0000 : 4'b0010;
						assign node2143 = (inp[14]) ? node2527 : node2144;
							assign node2144 = (inp[15]) ? node2348 : node2145;
								assign node2145 = (inp[0]) ? node2247 : node2146;
									assign node2146 = (inp[5]) ? node2196 : node2147;
										assign node2147 = (inp[8]) ? node2171 : node2148;
											assign node2148 = (inp[6]) ? node2160 : node2149;
												assign node2149 = (inp[11]) ? node2153 : node2150;
													assign node2150 = (inp[3]) ? 4'b1011 : 4'b0011;
													assign node2153 = (inp[1]) ? 4'b0010 : node2154;
														assign node2154 = (inp[2]) ? node2156 : 4'b0011;
															assign node2156 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node2160 = (inp[11]) ? node2164 : node2161;
													assign node2161 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node2164 = (inp[2]) ? node2166 : 4'b1010;
														assign node2166 = (inp[7]) ? node2168 : 4'b1010;
															assign node2168 = (inp[3]) ? 4'b1011 : 4'b0011;
											assign node2171 = (inp[1]) ? node2187 : node2172;
												assign node2172 = (inp[3]) ? node2180 : node2173;
													assign node2173 = (inp[2]) ? node2175 : 4'b1011;
														assign node2175 = (inp[11]) ? 4'b0010 : node2176;
															assign node2176 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node2180 = (inp[7]) ? 4'b1011 : node2181;
														assign node2181 = (inp[6]) ? 4'b1011 : node2182;
															assign node2182 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node2187 = (inp[6]) ? node2189 : 4'b1011;
													assign node2189 = (inp[11]) ? 4'b1010 : node2190;
														assign node2190 = (inp[3]) ? node2192 : 4'b1011;
															assign node2192 = (inp[2]) ? 4'b1010 : 4'b0010;
										assign node2196 = (inp[3]) ? node2222 : node2197;
											assign node2197 = (inp[1]) ? node2207 : node2198;
												assign node2198 = (inp[2]) ? 4'b1010 : node2199;
													assign node2199 = (inp[8]) ? node2203 : node2200;
														assign node2200 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node2203 = (inp[6]) ? 4'b1011 : 4'b1010;
												assign node2207 = (inp[6]) ? node2213 : node2208;
													assign node2208 = (inp[2]) ? node2210 : 4'b1010;
														assign node2210 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node2213 = (inp[2]) ? 4'b1011 : node2214;
														assign node2214 = (inp[7]) ? node2218 : node2215;
															assign node2215 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node2218 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node2222 = (inp[1]) ? node2234 : node2223;
												assign node2223 = (inp[7]) ? 4'b1000 : node2224;
													assign node2224 = (inp[8]) ? node2228 : node2225;
														assign node2225 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node2228 = (inp[2]) ? node2230 : 4'b0000;
															assign node2230 = (inp[6]) ? 4'b1001 : 4'b0001;
												assign node2234 = (inp[6]) ? node2238 : node2235;
													assign node2235 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node2238 = (inp[2]) ? node2240 : 4'b1000;
														assign node2240 = (inp[11]) ? node2244 : node2241;
															assign node2241 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node2244 = (inp[8]) ? 4'b0000 : 4'b1000;
									assign node2247 = (inp[3]) ? node2299 : node2248;
										assign node2248 = (inp[1]) ? node2282 : node2249;
											assign node2249 = (inp[2]) ? node2267 : node2250;
												assign node2250 = (inp[5]) ? node2256 : node2251;
													assign node2251 = (inp[7]) ? node2253 : 4'b1000;
														assign node2253 = (inp[11]) ? 4'b1000 : 4'b0001;
													assign node2256 = (inp[11]) ? node2262 : node2257;
														assign node2257 = (inp[6]) ? 4'b0001 : node2258;
															assign node2258 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node2262 = (inp[8]) ? node2264 : 4'b0000;
															assign node2264 = (inp[6]) ? 4'b1001 : 4'b0001;
												assign node2267 = (inp[7]) ? node2275 : node2268;
													assign node2268 = (inp[8]) ? node2270 : 4'b0000;
														assign node2270 = (inp[5]) ? 4'b0001 : node2271;
															assign node2271 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node2275 = (inp[8]) ? 4'b1000 : node2276;
														assign node2276 = (inp[5]) ? node2278 : 4'b0001;
															assign node2278 = (inp[11]) ? 4'b1001 : 4'b0001;
											assign node2282 = (inp[11]) ? node2288 : node2283;
												assign node2283 = (inp[6]) ? 4'b0000 : node2284;
													assign node2284 = (inp[8]) ? 4'b0000 : 4'b1000;
												assign node2288 = (inp[7]) ? node2296 : node2289;
													assign node2289 = (inp[2]) ? node2293 : node2290;
														assign node2290 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node2293 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node2296 = (inp[8]) ? 4'b0000 : 4'b1000;
										assign node2299 = (inp[5]) ? node2325 : node2300;
											assign node2300 = (inp[6]) ? node2308 : node2301;
												assign node2301 = (inp[2]) ? node2303 : 4'b1000;
													assign node2303 = (inp[7]) ? node2305 : 4'b0001;
														assign node2305 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node2308 = (inp[1]) ? node2316 : node2309;
													assign node2309 = (inp[11]) ? node2311 : 4'b0001;
														assign node2311 = (inp[8]) ? node2313 : 4'b1001;
															assign node2313 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node2316 = (inp[2]) ? node2318 : 4'b0000;
														assign node2318 = (inp[11]) ? node2322 : node2319;
															assign node2319 = (inp[7]) ? 4'b1001 : 4'b0000;
															assign node2322 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node2325 = (inp[1]) ? node2337 : node2326;
												assign node2326 = (inp[11]) ? node2330 : node2327;
													assign node2327 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node2330 = (inp[6]) ? node2332 : 4'b0010;
														assign node2332 = (inp[7]) ? node2334 : 4'b1010;
															assign node2334 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node2337 = (inp[11]) ? 4'b0011 : node2338;
													assign node2338 = (inp[6]) ? node2344 : node2339;
														assign node2339 = (inp[7]) ? node2341 : 4'b0011;
															assign node2341 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node2344 = (inp[7]) ? 4'b1011 : 4'b0010;
								assign node2348 = (inp[0]) ? node2420 : node2349;
									assign node2349 = (inp[3]) ? node2381 : node2350;
										assign node2350 = (inp[6]) ? node2362 : node2351;
											assign node2351 = (inp[11]) ? node2355 : node2352;
												assign node2352 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node2355 = (inp[1]) ? node2357 : 4'b0000;
													assign node2357 = (inp[5]) ? 4'b1001 : node2358;
														assign node2358 = (inp[8]) ? 4'b1000 : 4'b0000;
											assign node2362 = (inp[7]) ? node2372 : node2363;
												assign node2363 = (inp[8]) ? node2367 : node2364;
													assign node2364 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node2367 = (inp[2]) ? 4'b1001 : node2368;
														assign node2368 = (inp[11]) ? 4'b1000 : 4'b0000;
												assign node2372 = (inp[2]) ? node2378 : node2373;
													assign node2373 = (inp[11]) ? node2375 : 4'b0001;
														assign node2375 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node2378 = (inp[11]) ? 4'b0001 : 4'b1001;
										assign node2381 = (inp[5]) ? node2399 : node2382;
											assign node2382 = (inp[11]) ? node2390 : node2383;
												assign node2383 = (inp[7]) ? node2387 : node2384;
													assign node2384 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node2387 = (inp[6]) ? 4'b0001 : 4'b0000;
												assign node2390 = (inp[2]) ? node2394 : node2391;
													assign node2391 = (inp[6]) ? 4'b1001 : 4'b0001;
													assign node2394 = (inp[1]) ? node2396 : 4'b1001;
														assign node2396 = (inp[6]) ? 4'b0001 : 4'b1001;
											assign node2399 = (inp[6]) ? node2409 : node2400;
												assign node2400 = (inp[8]) ? node2402 : 4'b0011;
													assign node2402 = (inp[7]) ? node2406 : node2403;
														assign node2403 = (inp[1]) ? 4'b1010 : 4'b0010;
														assign node2406 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node2409 = (inp[11]) ? node2413 : node2410;
													assign node2410 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node2413 = (inp[7]) ? 4'b1010 : node2414;
														assign node2414 = (inp[2]) ? 4'b1010 : node2415;
															assign node2415 = (inp[8]) ? 4'b1010 : 4'b1011;
									assign node2420 = (inp[5]) ? node2480 : node2421;
										assign node2421 = (inp[1]) ? node2443 : node2422;
											assign node2422 = (inp[11]) ? node2434 : node2423;
												assign node2423 = (inp[6]) ? 4'b0010 : node2424;
													assign node2424 = (inp[2]) ? node2428 : node2425;
														assign node2425 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node2428 = (inp[7]) ? node2430 : 4'b1011;
															assign node2430 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node2434 = (inp[6]) ? node2436 : 4'b0011;
													assign node2436 = (inp[7]) ? 4'b1011 : node2437;
														assign node2437 = (inp[2]) ? node2439 : 4'b1010;
															assign node2439 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node2443 = (inp[3]) ? node2463 : node2444;
												assign node2444 = (inp[6]) ? node2450 : node2445;
													assign node2445 = (inp[2]) ? 4'b0010 : node2446;
														assign node2446 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node2450 = (inp[2]) ? node2456 : node2451;
														assign node2451 = (inp[11]) ? node2453 : 4'b0011;
															assign node2453 = (inp[7]) ? 4'b0010 : 4'b1010;
														assign node2456 = (inp[11]) ? node2460 : node2457;
															assign node2457 = (inp[7]) ? 4'b1010 : 4'b0010;
															assign node2460 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node2463 = (inp[8]) ? node2471 : node2464;
													assign node2464 = (inp[6]) ? node2466 : 4'b1010;
														assign node2466 = (inp[2]) ? node2468 : 4'b1011;
															assign node2468 = (inp[7]) ? 4'b1011 : 4'b0010;
													assign node2471 = (inp[6]) ? node2475 : node2472;
														assign node2472 = (inp[2]) ? 4'b1011 : 4'b0011;
														assign node2475 = (inp[11]) ? node2477 : 4'b0010;
															assign node2477 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node2480 = (inp[3]) ? node2504 : node2481;
											assign node2481 = (inp[8]) ? node2489 : node2482;
												assign node2482 = (inp[6]) ? node2486 : node2483;
													assign node2483 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node2486 = (inp[1]) ? 4'b1011 : 4'b0011;
												assign node2489 = (inp[11]) ? node2499 : node2490;
													assign node2490 = (inp[2]) ? node2494 : node2491;
														assign node2491 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node2494 = (inp[6]) ? node2496 : 4'b0011;
															assign node2496 = (inp[1]) ? 4'b1011 : 4'b0011;
													assign node2499 = (inp[7]) ? 4'b1010 : node2500;
														assign node2500 = (inp[1]) ? 4'b1010 : 4'b1011;
											assign node2504 = (inp[7]) ? node2520 : node2505;
												assign node2505 = (inp[6]) ? node2509 : node2506;
													assign node2506 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node2509 = (inp[11]) ? node2517 : node2510;
														assign node2510 = (inp[1]) ? node2514 : node2511;
															assign node2511 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node2514 = (inp[2]) ? 4'b1001 : 4'b0000;
														assign node2517 = (inp[1]) ? 4'b1000 : 4'b1001;
												assign node2520 = (inp[1]) ? node2522 : 4'b1001;
													assign node2522 = (inp[8]) ? node2524 : 4'b0001;
														assign node2524 = (inp[2]) ? 4'b0000 : 4'b0001;
							assign node2527 = (inp[0]) ? node2747 : node2528;
								assign node2528 = (inp[15]) ? node2638 : node2529;
									assign node2529 = (inp[3]) ? node2577 : node2530;
										assign node2530 = (inp[2]) ? node2552 : node2531;
											assign node2531 = (inp[7]) ? node2545 : node2532;
												assign node2532 = (inp[8]) ? node2540 : node2533;
													assign node2533 = (inp[5]) ? 4'b0010 : node2534;
														assign node2534 = (inp[6]) ? 4'b1010 : node2535;
															assign node2535 = (inp[11]) ? 4'b0010 : 4'b1010;
													assign node2540 = (inp[6]) ? node2542 : 4'b1011;
														assign node2542 = (inp[1]) ? 4'b0011 : 4'b1011;
												assign node2545 = (inp[8]) ? 4'b0010 : node2546;
													assign node2546 = (inp[11]) ? 4'b0011 : node2547;
														assign node2547 = (inp[5]) ? 4'b1011 : 4'b0011;
											assign node2552 = (inp[5]) ? node2560 : node2553;
												assign node2553 = (inp[8]) ? node2557 : node2554;
													assign node2554 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node2557 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node2560 = (inp[1]) ? node2574 : node2561;
													assign node2561 = (inp[11]) ? node2567 : node2562;
														assign node2562 = (inp[7]) ? node2564 : 4'b1010;
															assign node2564 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node2567 = (inp[6]) ? node2571 : node2568;
															assign node2568 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node2571 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node2574 = (inp[11]) ? 4'b0011 : 4'b1011;
										assign node2577 = (inp[5]) ? node2605 : node2578;
											assign node2578 = (inp[2]) ? node2594 : node2579;
												assign node2579 = (inp[7]) ? node2587 : node2580;
													assign node2580 = (inp[8]) ? node2582 : 4'b0010;
														assign node2582 = (inp[6]) ? node2584 : 4'b0011;
															assign node2584 = (inp[11]) ? 4'b1011 : 4'b0011;
													assign node2587 = (inp[8]) ? node2589 : 4'b1011;
														assign node2589 = (inp[11]) ? node2591 : 4'b0010;
															assign node2591 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node2594 = (inp[1]) ? node2598 : node2595;
													assign node2595 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node2598 = (inp[8]) ? 4'b0011 : node2599;
														assign node2599 = (inp[7]) ? node2601 : 4'b1010;
															assign node2601 = (inp[6]) ? 4'b0011 : 4'b1011;
											assign node2605 = (inp[6]) ? node2625 : node2606;
												assign node2606 = (inp[2]) ? node2614 : node2607;
													assign node2607 = (inp[7]) ? node2609 : 4'b0000;
														assign node2609 = (inp[11]) ? 4'b1001 : node2610;
															assign node2610 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node2614 = (inp[1]) ? node2620 : node2615;
														assign node2615 = (inp[11]) ? node2617 : 4'b1001;
															assign node2617 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node2620 = (inp[11]) ? 4'b0000 : node2621;
															assign node2621 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node2625 = (inp[2]) ? node2629 : node2626;
													assign node2626 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node2629 = (inp[7]) ? node2633 : node2630;
														assign node2630 = (inp[8]) ? 4'b0001 : 4'b1000;
														assign node2633 = (inp[8]) ? node2635 : 4'b0001;
															assign node2635 = (inp[11]) ? 4'b0000 : 4'b0000;
									assign node2638 = (inp[3]) ? node2694 : node2639;
										assign node2639 = (inp[2]) ? node2665 : node2640;
											assign node2640 = (inp[5]) ? node2660 : node2641;
												assign node2641 = (inp[7]) ? node2653 : node2642;
													assign node2642 = (inp[8]) ? node2648 : node2643;
														assign node2643 = (inp[11]) ? node2645 : 4'b0000;
															assign node2645 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node2648 = (inp[6]) ? node2650 : 4'b0001;
															assign node2650 = (inp[1]) ? 4'b0001 : 4'b0001;
													assign node2653 = (inp[8]) ? node2655 : 4'b1001;
														assign node2655 = (inp[1]) ? 4'b1000 : node2656;
															assign node2656 = (inp[6]) ? 4'b0000 : 4'b1000;
												assign node2660 = (inp[7]) ? 4'b0001 : node2661;
													assign node2661 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node2665 = (inp[11]) ? node2683 : node2666;
												assign node2666 = (inp[6]) ? node2676 : node2667;
													assign node2667 = (inp[1]) ? node2673 : node2668;
														assign node2668 = (inp[7]) ? node2670 : 4'b1001;
															assign node2670 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node2673 = (inp[8]) ? 4'b0001 : 4'b1000;
													assign node2676 = (inp[1]) ? 4'b1001 : node2677;
														assign node2677 = (inp[7]) ? node2679 : 4'b0000;
															assign node2679 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node2683 = (inp[8]) ? node2687 : node2684;
													assign node2684 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node2687 = (inp[7]) ? 4'b0000 : node2688;
														assign node2688 = (inp[5]) ? node2690 : 4'b1001;
															assign node2690 = (inp[6]) ? 4'b1001 : 4'b0001;
										assign node2694 = (inp[5]) ? node2720 : node2695;
											assign node2695 = (inp[1]) ? node2707 : node2696;
												assign node2696 = (inp[11]) ? node2702 : node2697;
													assign node2697 = (inp[6]) ? 4'b0000 : node2698;
														assign node2698 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node2702 = (inp[6]) ? 4'b1001 : node2703;
														assign node2703 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node2707 = (inp[6]) ? node2713 : node2708;
													assign node2708 = (inp[2]) ? 4'b0000 : node2709;
														assign node2709 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node2713 = (inp[8]) ? 4'b1000 : node2714;
														assign node2714 = (inp[7]) ? node2716 : 4'b0000;
															assign node2716 = (inp[11]) ? 4'b0001 : 4'b1001;
											assign node2720 = (inp[1]) ? node2734 : node2721;
												assign node2721 = (inp[7]) ? node2729 : node2722;
													assign node2722 = (inp[8]) ? node2724 : 4'b1010;
														assign node2724 = (inp[6]) ? node2726 : 4'b0011;
															assign node2726 = (inp[11]) ? 4'b1011 : 4'b0011;
													assign node2729 = (inp[11]) ? node2731 : 4'b0010;
														assign node2731 = (inp[6]) ? 4'b1010 : 4'b0010;
												assign node2734 = (inp[2]) ? node2742 : node2735;
													assign node2735 = (inp[7]) ? node2739 : node2736;
														assign node2736 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node2739 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node2742 = (inp[11]) ? 4'b0011 : node2743;
														assign node2743 = (inp[8]) ? 4'b0011 : 4'b1011;
								assign node2747 = (inp[15]) ? node2815 : node2748;
									assign node2748 = (inp[3]) ? node2778 : node2749;
										assign node2749 = (inp[7]) ? node2763 : node2750;
											assign node2750 = (inp[8]) ? node2754 : node2751;
												assign node2751 = (inp[2]) ? 4'b1000 : 4'b0000;
												assign node2754 = (inp[11]) ? node2756 : 4'b0001;
													assign node2756 = (inp[1]) ? node2760 : node2757;
														assign node2757 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node2760 = (inp[6]) ? 4'b0001 : 4'b1001;
											assign node2763 = (inp[8]) ? node2769 : node2764;
												assign node2764 = (inp[6]) ? 4'b1001 : node2765;
													assign node2765 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node2769 = (inp[2]) ? node2771 : 4'b0000;
													assign node2771 = (inp[1]) ? 4'b0000 : node2772;
														assign node2772 = (inp[5]) ? node2774 : 4'b1000;
															assign node2774 = (inp[6]) ? 4'b1000 : 4'b0000;
										assign node2778 = (inp[5]) ? node2794 : node2779;
											assign node2779 = (inp[8]) ? node2789 : node2780;
												assign node2780 = (inp[7]) ? 4'b0001 : node2781;
													assign node2781 = (inp[2]) ? node2785 : node2782;
														assign node2782 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node2785 = (inp[6]) ? 4'b0000 : 4'b1000;
												assign node2789 = (inp[7]) ? node2791 : 4'b0001;
													assign node2791 = (inp[1]) ? 4'b1000 : 4'b0000;
											assign node2794 = (inp[11]) ? node2800 : node2795;
												assign node2795 = (inp[8]) ? 4'b0010 : node2796;
													assign node2796 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node2800 = (inp[1]) ? node2810 : node2801;
													assign node2801 = (inp[6]) ? node2807 : node2802;
														assign node2802 = (inp[7]) ? 4'b0010 : node2803;
															assign node2803 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node2807 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node2810 = (inp[6]) ? node2812 : 4'b1011;
														assign node2812 = (inp[2]) ? 4'b0011 : 4'b0010;
									assign node2815 = (inp[3]) ? node2869 : node2816;
										assign node2816 = (inp[6]) ? node2840 : node2817;
											assign node2817 = (inp[11]) ? node2827 : node2818;
												assign node2818 = (inp[1]) ? node2824 : node2819;
													assign node2819 = (inp[2]) ? 4'b1011 : node2820;
														assign node2820 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node2824 = (inp[8]) ? 4'b0010 : 4'b1010;
												assign node2827 = (inp[1]) ? node2835 : node2828;
													assign node2828 = (inp[5]) ? node2830 : 4'b0010;
														assign node2830 = (inp[7]) ? 4'b0011 : node2831;
															assign node2831 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node2835 = (inp[5]) ? 4'b1011 : node2836;
														assign node2836 = (inp[7]) ? 4'b1011 : 4'b0010;
											assign node2840 = (inp[11]) ? node2854 : node2841;
												assign node2841 = (inp[1]) ? 4'b0010 : node2842;
													assign node2842 = (inp[2]) ? node2848 : node2843;
														assign node2843 = (inp[7]) ? 4'b0011 : node2844;
															assign node2844 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node2848 = (inp[7]) ? 4'b0010 : node2849;
															assign node2849 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node2854 = (inp[1]) ? node2864 : node2855;
													assign node2855 = (inp[2]) ? node2857 : 4'b1011;
														assign node2857 = (inp[7]) ? node2861 : node2858;
															assign node2858 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node2861 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node2864 = (inp[5]) ? 4'b0011 : node2865;
														assign node2865 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node2869 = (inp[5]) ? node2897 : node2870;
											assign node2870 = (inp[2]) ? node2884 : node2871;
												assign node2871 = (inp[1]) ? node2877 : node2872;
													assign node2872 = (inp[11]) ? node2874 : 4'b0011;
														assign node2874 = (inp[6]) ? 4'b1011 : 4'b0011;
													assign node2877 = (inp[6]) ? node2879 : 4'b1011;
														assign node2879 = (inp[11]) ? 4'b1010 : node2880;
															assign node2880 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node2884 = (inp[6]) ? node2892 : node2885;
													assign node2885 = (inp[11]) ? 4'b0010 : node2886;
														assign node2886 = (inp[7]) ? node2888 : 4'b0011;
															assign node2888 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node2892 = (inp[11]) ? 4'b0010 : node2893;
														assign node2893 = (inp[8]) ? 4'b1010 : 4'b0010;
											assign node2897 = (inp[1]) ? node2911 : node2898;
												assign node2898 = (inp[6]) ? 4'b0001 : node2899;
													assign node2899 = (inp[11]) ? node2907 : node2900;
														assign node2900 = (inp[2]) ? node2904 : node2901;
															assign node2901 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node2904 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node2907 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node2911 = (inp[7]) ? node2917 : node2912;
													assign node2912 = (inp[8]) ? 4'b0001 : node2913;
														assign node2913 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node2917 = (inp[8]) ? 4'b0000 : 4'b0001;
				assign node2920 = (inp[12]) ? node4242 : node2921;
					assign node2921 = (inp[10]) ? node3621 : node2922;
						assign node2922 = (inp[0]) ? node3240 : node2923;
							assign node2923 = (inp[15]) ? node3089 : node2924;
								assign node2924 = (inp[5]) ? node3016 : node2925;
									assign node2925 = (inp[1]) ? node2967 : node2926;
										assign node2926 = (inp[11]) ? node2946 : node2927;
											assign node2927 = (inp[6]) ? node2941 : node2928;
												assign node2928 = (inp[8]) ? node2938 : node2929;
													assign node2929 = (inp[14]) ? node2935 : node2930;
														assign node2930 = (inp[2]) ? 4'b1011 : node2931;
															assign node2931 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node2935 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node2938 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node2941 = (inp[14]) ? node2943 : 4'b0010;
													assign node2943 = (inp[8]) ? 4'b0011 : 4'b0010;
											assign node2946 = (inp[6]) ? node2956 : node2947;
												assign node2947 = (inp[8]) ? node2949 : 4'b0011;
													assign node2949 = (inp[3]) ? node2951 : 4'b0010;
														assign node2951 = (inp[7]) ? node2953 : 4'b0011;
															assign node2953 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node2956 = (inp[14]) ? node2962 : node2957;
													assign node2957 = (inp[8]) ? node2959 : 4'b1010;
														assign node2959 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node2962 = (inp[3]) ? node2964 : 4'b1011;
														assign node2964 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node2967 = (inp[2]) ? node2991 : node2968;
											assign node2968 = (inp[3]) ? node2974 : node2969;
												assign node2969 = (inp[6]) ? node2971 : 4'b0010;
													assign node2971 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node2974 = (inp[14]) ? node2986 : node2975;
													assign node2975 = (inp[6]) ? node2983 : node2976;
														assign node2976 = (inp[7]) ? node2980 : node2977;
															assign node2977 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node2980 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node2983 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node2986 = (inp[6]) ? node2988 : 4'b0011;
														assign node2988 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node2991 = (inp[11]) ? node3003 : node2992;
												assign node2992 = (inp[6]) ? node2998 : node2993;
													assign node2993 = (inp[3]) ? 4'b0011 : node2994;
														assign node2994 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node2998 = (inp[8]) ? 4'b1011 : node2999;
														assign node2999 = (inp[7]) ? 4'b1011 : 4'b0010;
												assign node3003 = (inp[6]) ? node3009 : node3004;
													assign node3004 = (inp[8]) ? node3006 : 4'b0010;
														assign node3006 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node3009 = (inp[8]) ? node3013 : node3010;
														assign node3010 = (inp[7]) ? 4'b0011 : 4'b1010;
														assign node3013 = (inp[7]) ? 4'b0010 : 4'b0011;
									assign node3016 = (inp[3]) ? node3058 : node3017;
										assign node3017 = (inp[2]) ? node3043 : node3018;
											assign node3018 = (inp[8]) ? node3038 : node3019;
												assign node3019 = (inp[6]) ? node3027 : node3020;
													assign node3020 = (inp[14]) ? node3024 : node3021;
														assign node3021 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node3024 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node3027 = (inp[11]) ? node3035 : node3028;
														assign node3028 = (inp[14]) ? node3032 : node3029;
															assign node3029 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node3032 = (inp[1]) ? 4'b1011 : 4'b0011;
														assign node3035 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node3038 = (inp[7]) ? 4'b0010 : node3039;
													assign node3039 = (inp[14]) ? 4'b0011 : 4'b0010;
											assign node3043 = (inp[6]) ? node3053 : node3044;
												assign node3044 = (inp[8]) ? node3048 : node3045;
													assign node3045 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node3048 = (inp[14]) ? node3050 : 4'b0010;
														assign node3050 = (inp[1]) ? 4'b0011 : 4'b1011;
												assign node3053 = (inp[1]) ? 4'b1010 : node3054;
													assign node3054 = (inp[11]) ? 4'b1010 : 4'b0010;
										assign node3058 = (inp[7]) ? node3080 : node3059;
											assign node3059 = (inp[8]) ? node3069 : node3060;
												assign node3060 = (inp[1]) ? node3066 : node3061;
													assign node3061 = (inp[11]) ? 4'b0000 : node3062;
														assign node3062 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node3066 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node3069 = (inp[11]) ? node3073 : node3070;
													assign node3070 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node3073 = (inp[1]) ? node3077 : node3074;
														assign node3074 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node3077 = (inp[6]) ? 4'b1000 : 4'b1001;
											assign node3080 = (inp[8]) ? node3082 : 4'b1001;
												assign node3082 = (inp[14]) ? 4'b1000 : node3083;
													assign node3083 = (inp[1]) ? 4'b0001 : node3084;
														assign node3084 = (inp[2]) ? 4'b1000 : 4'b1001;
								assign node3089 = (inp[5]) ? node3163 : node3090;
									assign node3090 = (inp[1]) ? node3132 : node3091;
										assign node3091 = (inp[8]) ? node3111 : node3092;
											assign node3092 = (inp[7]) ? node3102 : node3093;
												assign node3093 = (inp[14]) ? node3097 : node3094;
													assign node3094 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node3097 = (inp[3]) ? 4'b1000 : node3098;
														assign node3098 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node3102 = (inp[2]) ? node3108 : node3103;
													assign node3103 = (inp[14]) ? node3105 : 4'b0000;
														assign node3105 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node3108 = (inp[11]) ? 4'b1001 : 4'b0001;
											assign node3111 = (inp[7]) ? node3117 : node3112;
												assign node3112 = (inp[2]) ? node3114 : 4'b0000;
													assign node3114 = (inp[3]) ? 4'b0001 : 4'b1001;
												assign node3117 = (inp[3]) ? node3127 : node3118;
													assign node3118 = (inp[2]) ? node3120 : 4'b1000;
														assign node3120 = (inp[14]) ? node3124 : node3121;
															assign node3121 = (inp[11]) ? 4'b1000 : 4'b0000;
															assign node3124 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node3127 = (inp[11]) ? node3129 : 4'b0000;
														assign node3129 = (inp[6]) ? 4'b1000 : 4'b0000;
										assign node3132 = (inp[11]) ? node3148 : node3133;
											assign node3133 = (inp[6]) ? node3141 : node3134;
												assign node3134 = (inp[8]) ? 4'b0001 : node3135;
													assign node3135 = (inp[2]) ? node3137 : 4'b1000;
														assign node3137 = (inp[7]) ? 4'b0001 : 4'b1000;
												assign node3141 = (inp[3]) ? node3143 : 4'b1001;
													assign node3143 = (inp[8]) ? node3145 : 4'b1001;
														assign node3145 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node3148 = (inp[6]) ? node3154 : node3149;
												assign node3149 = (inp[7]) ? node3151 : 4'b0000;
													assign node3151 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node3154 = (inp[8]) ? node3156 : 4'b1000;
													assign node3156 = (inp[7]) ? 4'b0000 : node3157;
														assign node3157 = (inp[3]) ? 4'b0001 : node3158;
															assign node3158 = (inp[2]) ? 4'b0001 : 4'b1000;
									assign node3163 = (inp[3]) ? node3203 : node3164;
										assign node3164 = (inp[1]) ? node3182 : node3165;
											assign node3165 = (inp[6]) ? node3175 : node3166;
												assign node3166 = (inp[11]) ? node3168 : 4'b1001;
													assign node3168 = (inp[14]) ? node3170 : 4'b0001;
														assign node3170 = (inp[2]) ? node3172 : 4'b0001;
															assign node3172 = (inp[7]) ? 4'b0000 : 4'b0000;
												assign node3175 = (inp[2]) ? node3177 : 4'b0000;
													assign node3177 = (inp[8]) ? node3179 : 4'b1000;
														assign node3179 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node3182 = (inp[6]) ? node3198 : node3183;
												assign node3183 = (inp[2]) ? node3193 : node3184;
													assign node3184 = (inp[8]) ? node3188 : node3185;
														assign node3185 = (inp[14]) ? 4'b1001 : 4'b0001;
														assign node3188 = (inp[11]) ? 4'b1000 : node3189;
															assign node3189 = (inp[14]) ? 4'b0000 : 4'b1000;
													assign node3193 = (inp[8]) ? 4'b1000 : node3194;
														assign node3194 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node3198 = (inp[2]) ? node3200 : 4'b1000;
													assign node3200 = (inp[14]) ? 4'b0001 : 4'b1001;
										assign node3203 = (inp[6]) ? node3217 : node3204;
											assign node3204 = (inp[7]) ? node3210 : node3205;
												assign node3205 = (inp[14]) ? node3207 : 4'b1011;
													assign node3207 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node3210 = (inp[11]) ? node3214 : node3211;
													assign node3211 = (inp[1]) ? 4'b0010 : 4'b1010;
													assign node3214 = (inp[14]) ? 4'b1010 : 4'b1011;
											assign node3217 = (inp[11]) ? node3227 : node3218;
												assign node3218 = (inp[1]) ? node3224 : node3219;
													assign node3219 = (inp[8]) ? node3221 : 4'b0011;
														assign node3221 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node3224 = (inp[7]) ? 4'b1010 : 4'b0010;
												assign node3227 = (inp[1]) ? node3235 : node3228;
													assign node3228 = (inp[14]) ? 4'b1011 : node3229;
														assign node3229 = (inp[8]) ? node3231 : 4'b1010;
															assign node3231 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node3235 = (inp[2]) ? node3237 : 4'b1010;
														assign node3237 = (inp[8]) ? 4'b0010 : 4'b0011;
							assign node3240 = (inp[15]) ? node3434 : node3241;
								assign node3241 = (inp[5]) ? node3335 : node3242;
									assign node3242 = (inp[14]) ? node3296 : node3243;
										assign node3243 = (inp[1]) ? node3275 : node3244;
											assign node3244 = (inp[11]) ? node3260 : node3245;
												assign node3245 = (inp[6]) ? node3253 : node3246;
													assign node3246 = (inp[2]) ? node3248 : 4'b1000;
														assign node3248 = (inp[7]) ? node3250 : 4'b1001;
															assign node3250 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node3253 = (inp[2]) ? 4'b0001 : node3254;
														assign node3254 = (inp[8]) ? node3256 : 4'b0000;
															assign node3256 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node3260 = (inp[6]) ? node3272 : node3261;
													assign node3261 = (inp[8]) ? node3267 : node3262;
														assign node3262 = (inp[7]) ? 4'b0000 : node3263;
															assign node3263 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node3267 = (inp[2]) ? node3269 : 4'b0001;
															assign node3269 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node3272 = (inp[3]) ? 4'b1000 : 4'b1001;
											assign node3275 = (inp[7]) ? node3289 : node3276;
												assign node3276 = (inp[11]) ? node3286 : node3277;
													assign node3277 = (inp[8]) ? node3281 : node3278;
														assign node3278 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node3281 = (inp[2]) ? node3283 : 4'b1000;
															assign node3283 = (inp[3]) ? 4'b1001 : 4'b0001;
													assign node3286 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node3289 = (inp[6]) ? node3293 : node3290;
													assign node3290 = (inp[11]) ? 4'b1001 : 4'b0001;
													assign node3293 = (inp[11]) ? 4'b0001 : 4'b1001;
										assign node3296 = (inp[2]) ? node3308 : node3297;
											assign node3297 = (inp[11]) ? node3303 : node3298;
												assign node3298 = (inp[7]) ? node3300 : 4'b1001;
													assign node3300 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node3303 = (inp[7]) ? 4'b0000 : node3304;
													assign node3304 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node3308 = (inp[11]) ? node3328 : node3309;
												assign node3309 = (inp[3]) ? node3319 : node3310;
													assign node3310 = (inp[7]) ? node3314 : node3311;
														assign node3311 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node3314 = (inp[6]) ? 4'b1000 : node3315;
															assign node3315 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node3319 = (inp[1]) ? node3325 : node3320;
														assign node3320 = (inp[7]) ? 4'b1000 : node3321;
															assign node3321 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node3325 = (inp[6]) ? 4'b1000 : 4'b0000;
												assign node3328 = (inp[3]) ? 4'b1001 : node3329;
													assign node3329 = (inp[6]) ? node3331 : 4'b1000;
														assign node3331 = (inp[7]) ? 4'b0001 : 4'b1000;
									assign node3335 = (inp[3]) ? node3379 : node3336;
										assign node3336 = (inp[8]) ? node3354 : node3337;
											assign node3337 = (inp[7]) ? node3339 : 4'b0000;
												assign node3339 = (inp[2]) ? node3347 : node3340;
													assign node3340 = (inp[14]) ? node3344 : node3341;
														assign node3341 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node3344 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node3347 = (inp[14]) ? 4'b0001 : node3348;
														assign node3348 = (inp[11]) ? node3350 : 4'b1001;
															assign node3350 = (inp[1]) ? 4'b1001 : 4'b0001;
											assign node3354 = (inp[7]) ? node3368 : node3355;
												assign node3355 = (inp[11]) ? node3363 : node3356;
													assign node3356 = (inp[14]) ? node3358 : 4'b1001;
														assign node3358 = (inp[6]) ? 4'b0001 : node3359;
															assign node3359 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node3363 = (inp[14]) ? 4'b1001 : node3364;
														assign node3364 = (inp[1]) ? 4'b0001 : 4'b1000;
												assign node3368 = (inp[11]) ? node3376 : node3369;
													assign node3369 = (inp[6]) ? 4'b1001 : node3370;
														assign node3370 = (inp[2]) ? 4'b1000 : node3371;
															assign node3371 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node3376 = (inp[1]) ? 4'b1000 : 4'b0000;
										assign node3379 = (inp[14]) ? node3419 : node3380;
											assign node3380 = (inp[8]) ? node3404 : node3381;
												assign node3381 = (inp[1]) ? node3391 : node3382;
													assign node3382 = (inp[6]) ? node3388 : node3383;
														assign node3383 = (inp[11]) ? 4'b0010 : node3384;
															assign node3384 = (inp[2]) ? 4'b1010 : 4'b1010;
														assign node3388 = (inp[7]) ? 4'b0010 : 4'b1010;
													assign node3391 = (inp[7]) ? node3399 : node3392;
														assign node3392 = (inp[2]) ? node3396 : node3393;
															assign node3393 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node3396 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node3399 = (inp[6]) ? node3401 : 4'b1011;
															assign node3401 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node3404 = (inp[7]) ? node3412 : node3405;
													assign node3405 = (inp[2]) ? node3409 : node3406;
														assign node3406 = (inp[6]) ? 4'b0010 : 4'b1010;
														assign node3409 = (inp[6]) ? 4'b1011 : 4'b0011;
													assign node3412 = (inp[2]) ? node3414 : 4'b1011;
														assign node3414 = (inp[6]) ? 4'b1010 : node3415;
															assign node3415 = (inp[11]) ? 4'b0010 : 4'b0010;
											assign node3419 = (inp[1]) ? node3425 : node3420;
												assign node3420 = (inp[2]) ? 4'b0011 : node3421;
													assign node3421 = (inp[8]) ? 4'b1011 : 4'b0011;
												assign node3425 = (inp[6]) ? node3431 : node3426;
													assign node3426 = (inp[7]) ? 4'b0010 : node3427;
														assign node3427 = (inp[11]) ? 4'b0010 : 4'b1010;
													assign node3431 = (inp[11]) ? 4'b1010 : 4'b1011;
								assign node3434 = (inp[3]) ? node3520 : node3435;
									assign node3435 = (inp[8]) ? node3477 : node3436;
										assign node3436 = (inp[7]) ? node3462 : node3437;
											assign node3437 = (inp[14]) ? node3449 : node3438;
												assign node3438 = (inp[2]) ? node3446 : node3439;
													assign node3439 = (inp[5]) ? node3441 : 4'b1011;
														assign node3441 = (inp[11]) ? node3443 : 4'b0011;
															assign node3443 = (inp[6]) ? 4'b1011 : 4'b0011;
													assign node3446 = (inp[1]) ? 4'b1010 : 4'b0010;
												assign node3449 = (inp[1]) ? node3451 : 4'b1010;
													assign node3451 = (inp[5]) ? node3457 : node3452;
														assign node3452 = (inp[6]) ? 4'b0010 : node3453;
															assign node3453 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node3457 = (inp[6]) ? node3459 : 4'b1010;
															assign node3459 = (inp[11]) ? 4'b1010 : 4'b0010;
											assign node3462 = (inp[2]) ? node3472 : node3463;
												assign node3463 = (inp[14]) ? 4'b0011 : node3464;
													assign node3464 = (inp[1]) ? node3466 : 4'b1010;
														assign node3466 = (inp[11]) ? 4'b0010 : node3467;
															assign node3467 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node3472 = (inp[5]) ? node3474 : 4'b1011;
													assign node3474 = (inp[6]) ? 4'b0011 : 4'b1011;
										assign node3477 = (inp[7]) ? node3499 : node3478;
											assign node3478 = (inp[2]) ? node3486 : node3479;
												assign node3479 = (inp[14]) ? 4'b0011 : node3480;
													assign node3480 = (inp[11]) ? node3482 : 4'b0010;
														assign node3482 = (inp[6]) ? 4'b1010 : 4'b0010;
												assign node3486 = (inp[1]) ? node3494 : node3487;
													assign node3487 = (inp[14]) ? node3489 : 4'b0011;
														assign node3489 = (inp[6]) ? 4'b1011 : node3490;
															assign node3490 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node3494 = (inp[11]) ? 4'b0011 : node3495;
														assign node3495 = (inp[6]) ? 4'b1011 : 4'b0011;
											assign node3499 = (inp[2]) ? node3511 : node3500;
												assign node3500 = (inp[14]) ? node3508 : node3501;
													assign node3501 = (inp[6]) ? 4'b1011 : node3502;
														assign node3502 = (inp[11]) ? node3504 : 4'b1011;
															assign node3504 = (inp[1]) ? 4'b1011 : 4'b0011;
													assign node3508 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node3511 = (inp[6]) ? node3513 : 4'b1010;
													assign node3513 = (inp[14]) ? node3517 : node3514;
														assign node3514 = (inp[1]) ? 4'b0010 : 4'b1010;
														assign node3517 = (inp[1]) ? 4'b1010 : 4'b0010;
									assign node3520 = (inp[5]) ? node3564 : node3521;
										assign node3521 = (inp[8]) ? node3535 : node3522;
											assign node3522 = (inp[7]) ? node3526 : node3523;
												assign node3523 = (inp[11]) ? 4'b0010 : 4'b1010;
												assign node3526 = (inp[6]) ? node3532 : node3527;
													assign node3527 = (inp[14]) ? 4'b0011 : node3528;
														assign node3528 = (inp[1]) ? 4'b1011 : 4'b0010;
													assign node3532 = (inp[14]) ? 4'b1011 : 4'b0011;
											assign node3535 = (inp[7]) ? node3547 : node3536;
												assign node3536 = (inp[14]) ? node3538 : 4'b0011;
													assign node3538 = (inp[6]) ? 4'b1011 : node3539;
														assign node3539 = (inp[2]) ? node3543 : node3540;
															assign node3540 = (inp[11]) ? 4'b0011 : 4'b1011;
															assign node3543 = (inp[1]) ? 4'b0011 : 4'b1011;
												assign node3547 = (inp[2]) ? node3557 : node3548;
													assign node3548 = (inp[14]) ? node3554 : node3549;
														assign node3549 = (inp[1]) ? node3551 : 4'b1011;
															assign node3551 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node3554 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node3557 = (inp[6]) ? node3559 : 4'b1010;
														assign node3559 = (inp[11]) ? 4'b0010 : node3560;
															assign node3560 = (inp[1]) ? 4'b1010 : 4'b0010;
										assign node3564 = (inp[2]) ? node3598 : node3565;
											assign node3565 = (inp[1]) ? node3583 : node3566;
												assign node3566 = (inp[11]) ? node3580 : node3567;
													assign node3567 = (inp[6]) ? node3573 : node3568;
														assign node3568 = (inp[8]) ? 4'b1000 : node3569;
															assign node3569 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node3573 = (inp[7]) ? node3577 : node3574;
															assign node3574 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node3577 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node3580 = (inp[6]) ? 4'b1000 : 4'b0000;
												assign node3583 = (inp[14]) ? node3591 : node3584;
													assign node3584 = (inp[6]) ? 4'b1000 : node3585;
														assign node3585 = (inp[11]) ? 4'b1001 : node3586;
															assign node3586 = (inp[8]) ? 4'b0000 : 4'b1000;
													assign node3591 = (inp[11]) ? node3593 : 4'b1000;
														assign node3593 = (inp[8]) ? 4'b0001 : node3594;
															assign node3594 = (inp[6]) ? 4'b1000 : 4'b0000;
											assign node3598 = (inp[8]) ? node3614 : node3599;
												assign node3599 = (inp[7]) ? node3607 : node3600;
													assign node3600 = (inp[1]) ? node3602 : 4'b0000;
														assign node3602 = (inp[14]) ? 4'b1000 : node3603;
															assign node3603 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node3607 = (inp[14]) ? node3609 : 4'b0001;
														assign node3609 = (inp[11]) ? 4'b1001 : node3610;
															assign node3610 = (inp[6]) ? 4'b1001 : 4'b0001;
												assign node3614 = (inp[1]) ? 4'b0001 : node3615;
													assign node3615 = (inp[14]) ? 4'b1001 : node3616;
														assign node3616 = (inp[6]) ? 4'b0001 : 4'b1001;
						assign node3621 = (inp[6]) ? node3933 : node3622;
							assign node3622 = (inp[11]) ? node3788 : node3623;
								assign node3623 = (inp[1]) ? node3719 : node3624;
									assign node3624 = (inp[5]) ? node3670 : node3625;
										assign node3625 = (inp[14]) ? node3651 : node3626;
											assign node3626 = (inp[15]) ? node3638 : node3627;
												assign node3627 = (inp[3]) ? node3633 : node3628;
													assign node3628 = (inp[7]) ? 4'b1011 : node3629;
														assign node3629 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node3633 = (inp[8]) ? node3635 : 4'b1010;
														assign node3635 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node3638 = (inp[0]) ? node3646 : node3639;
													assign node3639 = (inp[8]) ? 4'b1000 : node3640;
														assign node3640 = (inp[2]) ? node3642 : 4'b1001;
															assign node3642 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node3646 = (inp[3]) ? 4'b1011 : node3647;
														assign node3647 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node3651 = (inp[15]) ? node3659 : node3652;
												assign node3652 = (inp[0]) ? node3654 : 4'b1010;
													assign node3654 = (inp[7]) ? node3656 : 4'b1000;
														assign node3656 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node3659 = (inp[0]) ? node3665 : node3660;
													assign node3660 = (inp[8]) ? node3662 : 4'b1001;
														assign node3662 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node3665 = (inp[7]) ? 4'b1010 : node3666;
														assign node3666 = (inp[8]) ? 4'b1011 : 4'b1010;
										assign node3670 = (inp[8]) ? node3700 : node3671;
											assign node3671 = (inp[7]) ? node3685 : node3672;
												assign node3672 = (inp[0]) ? node3678 : node3673;
													assign node3673 = (inp[15]) ? 4'b1010 : node3674;
														assign node3674 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node3678 = (inp[14]) ? node3682 : node3679;
														assign node3679 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node3682 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node3685 = (inp[2]) ? node3691 : node3686;
													assign node3686 = (inp[14]) ? 4'b1011 : node3687;
														assign node3687 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node3691 = (inp[15]) ? node3693 : 4'b1011;
														assign node3693 = (inp[0]) ? node3697 : node3694;
															assign node3694 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node3697 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node3700 = (inp[7]) ? node3712 : node3701;
												assign node3701 = (inp[3]) ? node3707 : node3702;
													assign node3702 = (inp[2]) ? 4'b1001 : node3703;
														assign node3703 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node3707 = (inp[0]) ? node3709 : 4'b1010;
														assign node3709 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node3712 = (inp[0]) ? 4'b1010 : node3713;
													assign node3713 = (inp[3]) ? node3715 : 4'b1000;
														assign node3715 = (inp[14]) ? 4'b1000 : 4'b1001;
									assign node3719 = (inp[7]) ? node3753 : node3720;
										assign node3720 = (inp[8]) ? node3738 : node3721;
											assign node3721 = (inp[2]) ? node3729 : node3722;
												assign node3722 = (inp[14]) ? 4'b1000 : node3723;
													assign node3723 = (inp[15]) ? 4'b1011 : node3724;
														assign node3724 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node3729 = (inp[15]) ? node3735 : node3730;
													assign node3730 = (inp[0]) ? 4'b1000 : node3731;
														assign node3731 = (inp[14]) ? 4'b1010 : 4'b1000;
													assign node3735 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node3738 = (inp[14]) ? node3748 : node3739;
												assign node3739 = (inp[2]) ? node3745 : node3740;
													assign node3740 = (inp[0]) ? node3742 : 4'b1010;
														assign node3742 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node3745 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node3748 = (inp[2]) ? 4'b0011 : node3749;
													assign node3749 = (inp[15]) ? 4'b0011 : 4'b0001;
										assign node3753 = (inp[8]) ? node3775 : node3754;
											assign node3754 = (inp[2]) ? node3760 : node3755;
												assign node3755 = (inp[3]) ? node3757 : 4'b1010;
													assign node3757 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node3760 = (inp[5]) ? node3762 : 4'b0001;
													assign node3762 = (inp[15]) ? node3768 : node3763;
														assign node3763 = (inp[0]) ? 4'b0001 : node3764;
															assign node3764 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node3768 = (inp[14]) ? node3772 : node3769;
															assign node3769 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node3772 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node3775 = (inp[14]) ? node3781 : node3776;
												assign node3776 = (inp[2]) ? 4'b0000 : node3777;
													assign node3777 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node3781 = (inp[3]) ? 4'b0010 : node3782;
													assign node3782 = (inp[2]) ? node3784 : 4'b0000;
														assign node3784 = (inp[15]) ? 4'b0010 : 4'b0000;
								assign node3788 = (inp[1]) ? node3874 : node3789;
									assign node3789 = (inp[15]) ? node3827 : node3790;
										assign node3790 = (inp[0]) ? node3808 : node3791;
											assign node3791 = (inp[3]) ? node3799 : node3792;
												assign node3792 = (inp[7]) ? 4'b0011 : node3793;
													assign node3793 = (inp[8]) ? node3795 : 4'b0010;
														assign node3795 = (inp[14]) ? 4'b0011 : 4'b0010;
												assign node3799 = (inp[5]) ? 4'b0000 : node3800;
													assign node3800 = (inp[7]) ? 4'b0010 : node3801;
														assign node3801 = (inp[8]) ? 4'b0011 : node3802;
															assign node3802 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node3808 = (inp[5]) ? node3816 : node3809;
												assign node3809 = (inp[3]) ? 4'b0000 : node3810;
													assign node3810 = (inp[7]) ? node3812 : 4'b0000;
														assign node3812 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node3816 = (inp[3]) ? node3818 : 4'b0000;
													assign node3818 = (inp[8]) ? node3820 : 4'b0010;
														assign node3820 = (inp[2]) ? node3824 : node3821;
															assign node3821 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node3824 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node3827 = (inp[0]) ? node3857 : node3828;
											assign node3828 = (inp[5]) ? node3842 : node3829;
												assign node3829 = (inp[8]) ? node3837 : node3830;
													assign node3830 = (inp[7]) ? node3832 : 4'b0000;
														assign node3832 = (inp[14]) ? 4'b0001 : node3833;
															assign node3833 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node3837 = (inp[2]) ? node3839 : 4'b0001;
														assign node3839 = (inp[3]) ? 4'b0000 : 4'b0001;
												assign node3842 = (inp[3]) ? node3850 : node3843;
													assign node3843 = (inp[8]) ? 4'b0000 : node3844;
														assign node3844 = (inp[7]) ? node3846 : 4'b0001;
															assign node3846 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node3850 = (inp[8]) ? node3854 : node3851;
														assign node3851 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node3854 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node3857 = (inp[3]) ? node3867 : node3858;
												assign node3858 = (inp[8]) ? node3864 : node3859;
													assign node3859 = (inp[7]) ? 4'b0011 : node3860;
														assign node3860 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node3864 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node3867 = (inp[5]) ? node3871 : node3868;
													assign node3868 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node3871 = (inp[8]) ? 4'b0001 : 4'b0000;
									assign node3874 = (inp[8]) ? node3908 : node3875;
										assign node3875 = (inp[7]) ? node3897 : node3876;
											assign node3876 = (inp[2]) ? node3884 : node3877;
												assign node3877 = (inp[14]) ? node3879 : 4'b0011;
													assign node3879 = (inp[5]) ? node3881 : 4'b0000;
														assign node3881 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node3884 = (inp[15]) ? node3888 : node3885;
													assign node3885 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node3888 = (inp[0]) ? node3894 : node3889;
														assign node3889 = (inp[14]) ? 4'b0000 : node3890;
															assign node3890 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node3894 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node3897 = (inp[2]) ? node3901 : node3898;
												assign node3898 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node3901 = (inp[3]) ? node3903 : 4'b1111;
													assign node3903 = (inp[5]) ? node3905 : 4'b1101;
														assign node3905 = (inp[15]) ? 4'b1111 : 4'b1101;
										assign node3908 = (inp[2]) ? node3918 : node3909;
											assign node3909 = (inp[7]) ? node3913 : node3910;
												assign node3910 = (inp[14]) ? 4'b1111 : 4'b0010;
												assign node3913 = (inp[14]) ? 4'b1100 : node3914;
													assign node3914 = (inp[15]) ? 4'b1111 : 4'b1101;
											assign node3918 = (inp[7]) ? node3928 : node3919;
												assign node3919 = (inp[3]) ? node3921 : 4'b1101;
													assign node3921 = (inp[0]) ? node3925 : node3922;
														assign node3922 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node3925 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node3928 = (inp[3]) ? node3930 : 4'b1100;
													assign node3930 = (inp[15]) ? 4'b1100 : 4'b1110;
							assign node3933 = (inp[11]) ? node4085 : node3934;
								assign node3934 = (inp[1]) ? node4024 : node3935;
									assign node3935 = (inp[15]) ? node3983 : node3936;
										assign node3936 = (inp[0]) ? node3968 : node3937;
											assign node3937 = (inp[3]) ? node3955 : node3938;
												assign node3938 = (inp[8]) ? node3950 : node3939;
													assign node3939 = (inp[7]) ? node3945 : node3940;
														assign node3940 = (inp[14]) ? 4'b0010 : node3941;
															assign node3941 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node3945 = (inp[14]) ? 4'b0011 : node3946;
															assign node3946 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node3950 = (inp[7]) ? 4'b0010 : node3951;
														assign node3951 = (inp[14]) ? 4'b0011 : 4'b0010;
												assign node3955 = (inp[5]) ? node3961 : node3956;
													assign node3956 = (inp[14]) ? 4'b0010 : node3957;
														assign node3957 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node3961 = (inp[7]) ? node3963 : 4'b0001;
														assign node3963 = (inp[14]) ? node3965 : 4'b0000;
															assign node3965 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node3968 = (inp[5]) ? node3972 : node3969;
												assign node3969 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node3972 = (inp[3]) ? node3978 : node3973;
													assign node3973 = (inp[7]) ? 4'b0000 : node3974;
														assign node3974 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node3978 = (inp[14]) ? node3980 : 4'b0011;
														assign node3980 = (inp[2]) ? 4'b0011 : 4'b0010;
										assign node3983 = (inp[5]) ? node3999 : node3984;
											assign node3984 = (inp[0]) ? 4'b0011 : node3985;
												assign node3985 = (inp[7]) ? node3993 : node3986;
													assign node3986 = (inp[3]) ? node3988 : 4'b0001;
														assign node3988 = (inp[2]) ? 4'b0001 : node3989;
															assign node3989 = (inp[14]) ? 4'b0000 : 4'b0000;
													assign node3993 = (inp[14]) ? 4'b0000 : node3994;
														assign node3994 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node3999 = (inp[2]) ? node4011 : node4000;
												assign node4000 = (inp[14]) ? node4002 : 4'b0010;
													assign node4002 = (inp[8]) ? node4006 : node4003;
														assign node4003 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node4006 = (inp[0]) ? 4'b0000 : node4007;
															assign node4007 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node4011 = (inp[8]) ? node4017 : node4012;
													assign node4012 = (inp[3]) ? node4014 : 4'b0000;
														assign node4014 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node4017 = (inp[7]) ? node4019 : 4'b0001;
														assign node4019 = (inp[3]) ? 4'b0000 : node4020;
															assign node4020 = (inp[0]) ? 4'b0010 : 4'b0000;
									assign node4024 = (inp[7]) ? node4052 : node4025;
										assign node4025 = (inp[8]) ? node4035 : node4026;
											assign node4026 = (inp[2]) ? node4030 : node4027;
												assign node4027 = (inp[0]) ? 4'b0011 : 4'b0000;
												assign node4030 = (inp[0]) ? 4'b0000 : node4031;
													assign node4031 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node4035 = (inp[2]) ? node4045 : node4036;
												assign node4036 = (inp[14]) ? 4'b1101 : node4037;
													assign node4037 = (inp[15]) ? node4041 : node4038;
														assign node4038 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node4041 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node4045 = (inp[0]) ? 4'b1111 : node4046;
													assign node4046 = (inp[3]) ? node4048 : 4'b1101;
														assign node4048 = (inp[15]) ? 4'b1111 : 4'b1101;
										assign node4052 = (inp[8]) ? node4064 : node4053;
											assign node4053 = (inp[14]) ? node4059 : node4054;
												assign node4054 = (inp[2]) ? node4056 : 4'b0000;
													assign node4056 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node4059 = (inp[5]) ? node4061 : 4'b1111;
													assign node4061 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node4064 = (inp[14]) ? node4072 : node4065;
												assign node4065 = (inp[2]) ? node4067 : 4'b1111;
													assign node4067 = (inp[3]) ? 4'b1100 : node4068;
														assign node4068 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node4072 = (inp[5]) ? 4'b1100 : node4073;
													assign node4073 = (inp[0]) ? node4079 : node4074;
														assign node4074 = (inp[15]) ? 4'b1100 : node4075;
															assign node4075 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node4079 = (inp[2]) ? 4'b1110 : node4080;
															assign node4080 = (inp[15]) ? 4'b1100 : 4'b1110;
								assign node4085 = (inp[1]) ? node4155 : node4086;
									assign node4086 = (inp[7]) ? node4116 : node4087;
										assign node4087 = (inp[8]) ? node4099 : node4088;
											assign node4088 = (inp[2]) ? node4092 : node4089;
												assign node4089 = (inp[3]) ? 4'b1101 : 4'b1100;
												assign node4092 = (inp[0]) ? node4094 : 4'b1110;
													assign node4094 = (inp[3]) ? 4'b1110 : node4095;
														assign node4095 = (inp[14]) ? 4'b1100 : 4'b1110;
											assign node4099 = (inp[14]) ? node4111 : node4100;
												assign node4100 = (inp[0]) ? node4102 : 4'b1101;
													assign node4102 = (inp[15]) ? node4106 : node4103;
														assign node4103 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node4106 = (inp[5]) ? 4'b1100 : node4107;
															assign node4107 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node4111 = (inp[3]) ? node4113 : 4'b1111;
													assign node4113 = (inp[0]) ? 4'b1101 : 4'b1111;
										assign node4116 = (inp[3]) ? node4138 : node4117;
											assign node4117 = (inp[8]) ? node4131 : node4118;
												assign node4118 = (inp[14]) ? node4124 : node4119;
													assign node4119 = (inp[2]) ? 4'b1101 : node4120;
														assign node4120 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node4124 = (inp[15]) ? node4126 : 4'b1101;
														assign node4126 = (inp[5]) ? 4'b1111 : node4127;
															assign node4127 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node4131 = (inp[15]) ? node4135 : node4132;
													assign node4132 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node4135 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node4138 = (inp[14]) ? node4152 : node4139;
												assign node4139 = (inp[5]) ? node4147 : node4140;
													assign node4140 = (inp[2]) ? 4'b1100 : node4141;
														assign node4141 = (inp[0]) ? node4143 : 4'b1101;
															assign node4143 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node4147 = (inp[2]) ? 4'b1111 : node4148;
														assign node4148 = (inp[8]) ? 4'b1111 : 4'b1110;
												assign node4152 = (inp[8]) ? 4'b1110 : 4'b1111;
									assign node4155 = (inp[8]) ? node4199 : node4156;
										assign node4156 = (inp[7]) ? node4180 : node4157;
											assign node4157 = (inp[2]) ? node4169 : node4158;
												assign node4158 = (inp[14]) ? node4166 : node4159;
													assign node4159 = (inp[0]) ? node4161 : 4'b1101;
														assign node4161 = (inp[3]) ? 4'b1111 : node4162;
															assign node4162 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node4166 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node4169 = (inp[3]) ? node4175 : node4170;
													assign node4170 = (inp[14]) ? node4172 : 4'b1110;
														assign node4172 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node4175 = (inp[0]) ? node4177 : 4'b1100;
														assign node4177 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node4180 = (inp[2]) ? node4190 : node4181;
												assign node4181 = (inp[14]) ? node4185 : node4182;
													assign node4182 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node4185 = (inp[5]) ? node4187 : 4'b0111;
														assign node4187 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node4190 = (inp[3]) ? node4196 : node4191;
													assign node4191 = (inp[14]) ? 4'b0101 : node4192;
														assign node4192 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node4196 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node4199 = (inp[7]) ? node4223 : node4200;
											assign node4200 = (inp[2]) ? node4214 : node4201;
												assign node4201 = (inp[14]) ? node4209 : node4202;
													assign node4202 = (inp[5]) ? node4204 : 4'b1100;
														assign node4204 = (inp[3]) ? node4206 : 4'b1100;
															assign node4206 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node4209 = (inp[5]) ? 4'b0101 : node4210;
														assign node4210 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node4214 = (inp[0]) ? node4218 : node4215;
													assign node4215 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node4218 = (inp[14]) ? node4220 : 4'b0101;
														assign node4220 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node4223 = (inp[2]) ? node4231 : node4224;
												assign node4224 = (inp[14]) ? 4'b0110 : node4225;
													assign node4225 = (inp[15]) ? 4'b0101 : node4226;
														assign node4226 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node4231 = (inp[5]) ? 4'b0100 : node4232;
													assign node4232 = (inp[15]) ? node4238 : node4233;
														assign node4233 = (inp[14]) ? node4235 : 4'b0100;
															assign node4235 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node4238 = (inp[14]) ? 4'b0100 : 4'b0110;
					assign node4242 = (inp[10]) ? node4916 : node4243;
						assign node4243 = (inp[6]) ? node4571 : node4244;
							assign node4244 = (inp[11]) ? node4402 : node4245;
								assign node4245 = (inp[1]) ? node4323 : node4246;
									assign node4246 = (inp[5]) ? node4278 : node4247;
										assign node4247 = (inp[8]) ? node4265 : node4248;
											assign node4248 = (inp[7]) ? node4260 : node4249;
												assign node4249 = (inp[14]) ? node4255 : node4250;
													assign node4250 = (inp[2]) ? 4'b1000 : node4251;
														assign node4251 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node4255 = (inp[3]) ? node4257 : 4'b1000;
														assign node4257 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node4260 = (inp[14]) ? 4'b1001 : node4261;
													assign node4261 = (inp[0]) ? 4'b1000 : 4'b1011;
											assign node4265 = (inp[7]) ? node4275 : node4266;
												assign node4266 = (inp[0]) ? node4270 : node4267;
													assign node4267 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node4270 = (inp[15]) ? 4'b1011 : node4271;
														assign node4271 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node4275 = (inp[14]) ? 4'b1010 : 4'b1001;
										assign node4278 = (inp[8]) ? node4296 : node4279;
											assign node4279 = (inp[7]) ? node4283 : node4280;
												assign node4280 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node4283 = (inp[2]) ? node4289 : node4284;
													assign node4284 = (inp[14]) ? 4'b1011 : node4285;
														assign node4285 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node4289 = (inp[3]) ? node4291 : 4'b1011;
														assign node4291 = (inp[0]) ? 4'b1001 : node4292;
															assign node4292 = (inp[15]) ? 4'b1011 : 4'b1001;
											assign node4296 = (inp[7]) ? node4314 : node4297;
												assign node4297 = (inp[2]) ? node4307 : node4298;
													assign node4298 = (inp[14]) ? node4304 : node4299;
														assign node4299 = (inp[3]) ? 4'b1010 : node4300;
															assign node4300 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node4304 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node4307 = (inp[0]) ? node4309 : 4'b1001;
														assign node4309 = (inp[14]) ? 4'b1011 : node4310;
															assign node4310 = (inp[3]) ? 4'b1001 : 4'b1001;
												assign node4314 = (inp[14]) ? 4'b1000 : node4315;
													assign node4315 = (inp[3]) ? node4317 : 4'b1010;
														assign node4317 = (inp[15]) ? node4319 : 4'b1000;
															assign node4319 = (inp[0]) ? 4'b1000 : 4'b1010;
									assign node4323 = (inp[7]) ? node4363 : node4324;
										assign node4324 = (inp[8]) ? node4354 : node4325;
											assign node4325 = (inp[2]) ? node4341 : node4326;
												assign node4326 = (inp[14]) ? node4336 : node4327;
													assign node4327 = (inp[3]) ? node4333 : node4328;
														assign node4328 = (inp[5]) ? 4'b1011 : node4329;
															assign node4329 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node4333 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node4336 = (inp[3]) ? 4'b1000 : node4337;
														assign node4337 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node4341 = (inp[0]) ? node4349 : node4342;
													assign node4342 = (inp[15]) ? node4346 : node4343;
														assign node4343 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node4346 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node4349 = (inp[3]) ? node4351 : 4'b1000;
														assign node4351 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node4354 = (inp[14]) ? node4360 : node4355;
												assign node4355 = (inp[2]) ? 4'b0011 : node4356;
													assign node4356 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node4360 = (inp[3]) ? 4'b0011 : 4'b0001;
										assign node4363 = (inp[8]) ? node4385 : node4364;
											assign node4364 = (inp[14]) ? node4376 : node4365;
												assign node4365 = (inp[2]) ? node4371 : node4366;
													assign node4366 = (inp[15]) ? node4368 : 4'b1010;
														assign node4368 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node4371 = (inp[15]) ? 4'b0001 : node4372;
														assign node4372 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node4376 = (inp[3]) ? node4378 : 4'b0011;
													assign node4378 = (inp[2]) ? node4380 : 4'b0011;
														assign node4380 = (inp[5]) ? node4382 : 4'b0011;
															assign node4382 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node4385 = (inp[14]) ? node4393 : node4386;
												assign node4386 = (inp[2]) ? 4'b0000 : node4387;
													assign node4387 = (inp[15]) ? node4389 : 4'b0001;
														assign node4389 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node4393 = (inp[0]) ? node4399 : node4394;
													assign node4394 = (inp[2]) ? 4'b0010 : node4395;
														assign node4395 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node4399 = (inp[15]) ? 4'b0010 : 4'b0000;
								assign node4402 = (inp[1]) ? node4488 : node4403;
									assign node4403 = (inp[8]) ? node4433 : node4404;
										assign node4404 = (inp[7]) ? node4416 : node4405;
											assign node4405 = (inp[2]) ? node4413 : node4406;
												assign node4406 = (inp[14]) ? 4'b0000 : node4407;
													assign node4407 = (inp[0]) ? 4'b0001 : node4408;
														assign node4408 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node4413 = (inp[5]) ? 4'b0010 : 4'b0000;
											assign node4416 = (inp[3]) ? node4424 : node4417;
												assign node4417 = (inp[15]) ? node4421 : node4418;
													assign node4418 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node4421 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node4424 = (inp[14]) ? 4'b0011 : node4425;
													assign node4425 = (inp[2]) ? 4'b0011 : node4426;
														assign node4426 = (inp[0]) ? node4428 : 4'b0000;
															assign node4428 = (inp[5]) ? 4'b0000 : 4'b0010;
										assign node4433 = (inp[7]) ? node4459 : node4434;
											assign node4434 = (inp[14]) ? node4442 : node4435;
												assign node4435 = (inp[2]) ? 4'b0011 : node4436;
													assign node4436 = (inp[15]) ? node4438 : 4'b0010;
														assign node4438 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node4442 = (inp[2]) ? node4448 : node4443;
													assign node4443 = (inp[5]) ? 4'b0001 : node4444;
														assign node4444 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node4448 = (inp[3]) ? node4454 : node4449;
														assign node4449 = (inp[15]) ? 4'b0011 : node4450;
															assign node4450 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node4454 = (inp[15]) ? node4456 : 4'b0011;
															assign node4456 = (inp[5]) ? 4'b0011 : 4'b0001;
											assign node4459 = (inp[14]) ? node4471 : node4460;
												assign node4460 = (inp[2]) ? 4'b0010 : node4461;
													assign node4461 = (inp[0]) ? node4465 : node4462;
														assign node4462 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node4465 = (inp[3]) ? node4467 : 4'b0011;
															assign node4467 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node4471 = (inp[2]) ? node4481 : node4472;
													assign node4472 = (inp[5]) ? 4'b0010 : node4473;
														assign node4473 = (inp[3]) ? node4477 : node4474;
															assign node4474 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node4477 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node4481 = (inp[15]) ? node4485 : node4482;
														assign node4482 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node4485 = (inp[0]) ? 4'b0010 : 4'b0000;
									assign node4488 = (inp[8]) ? node4524 : node4489;
										assign node4489 = (inp[7]) ? node4509 : node4490;
											assign node4490 = (inp[14]) ? node4500 : node4491;
												assign node4491 = (inp[2]) ? node4495 : node4492;
													assign node4492 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node4495 = (inp[0]) ? 4'b0010 : node4496;
														assign node4496 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node4500 = (inp[3]) ? 4'b0010 : node4501;
													assign node4501 = (inp[5]) ? node4505 : node4502;
														assign node4502 = (inp[2]) ? 4'b0010 : 4'b0000;
														assign node4505 = (inp[0]) ? 4'b0000 : 4'b0010;
											assign node4509 = (inp[14]) ? node4517 : node4510;
												assign node4510 = (inp[2]) ? 4'b1101 : node4511;
													assign node4511 = (inp[3]) ? node4513 : 4'b0010;
														assign node4513 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node4517 = (inp[2]) ? node4519 : 4'b1101;
													assign node4519 = (inp[15]) ? node4521 : 4'b1111;
														assign node4521 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node4524 = (inp[7]) ? node4552 : node4525;
											assign node4525 = (inp[2]) ? node4535 : node4526;
												assign node4526 = (inp[14]) ? node4532 : node4527;
													assign node4527 = (inp[15]) ? node4529 : 4'b0010;
														assign node4529 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node4532 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node4535 = (inp[0]) ? node4543 : node4536;
													assign node4536 = (inp[3]) ? 4'b1111 : node4537;
														assign node4537 = (inp[14]) ? node4539 : 4'b1101;
															assign node4539 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node4543 = (inp[3]) ? node4549 : node4544;
														assign node4544 = (inp[15]) ? 4'b1111 : node4545;
															assign node4545 = (inp[14]) ? 4'b1101 : 4'b1111;
														assign node4549 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node4552 = (inp[2]) ? node4564 : node4553;
												assign node4553 = (inp[14]) ? node4559 : node4554;
													assign node4554 = (inp[5]) ? 4'b1101 : node4555;
														assign node4555 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node4559 = (inp[3]) ? node4561 : 4'b1100;
														assign node4561 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node4564 = (inp[5]) ? node4566 : 4'b1100;
													assign node4566 = (inp[15]) ? 4'b1110 : node4567;
														assign node4567 = (inp[14]) ? 4'b1100 : 4'b1110;
							assign node4571 = (inp[11]) ? node4747 : node4572;
								assign node4572 = (inp[1]) ? node4658 : node4573;
									assign node4573 = (inp[14]) ? node4617 : node4574;
										assign node4574 = (inp[3]) ? node4600 : node4575;
											assign node4575 = (inp[2]) ? node4589 : node4576;
												assign node4576 = (inp[0]) ? node4584 : node4577;
													assign node4577 = (inp[15]) ? 4'b0000 : node4578;
														assign node4578 = (inp[5]) ? node4580 : 4'b0010;
															assign node4580 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node4584 = (inp[15]) ? node4586 : 4'b0000;
														assign node4586 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node4589 = (inp[0]) ? node4597 : node4590;
													assign node4590 = (inp[15]) ? node4594 : node4591;
														assign node4591 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node4594 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node4597 = (inp[15]) ? 4'b0011 : 4'b0001;
											assign node4600 = (inp[0]) ? node4614 : node4601;
												assign node4601 = (inp[8]) ? node4605 : node4602;
													assign node4602 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node4605 = (inp[5]) ? node4611 : node4606;
														assign node4606 = (inp[15]) ? 4'b0000 : node4607;
															assign node4607 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node4611 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node4614 = (inp[8]) ? 4'b0001 : 4'b0011;
										assign node4617 = (inp[5]) ? node4631 : node4618;
											assign node4618 = (inp[3]) ? node4626 : node4619;
												assign node4619 = (inp[15]) ? 4'b0011 : node4620;
													assign node4620 = (inp[0]) ? node4622 : 4'b0010;
														assign node4622 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node4626 = (inp[15]) ? node4628 : 4'b0010;
													assign node4628 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node4631 = (inp[2]) ? node4645 : node4632;
												assign node4632 = (inp[0]) ? node4642 : node4633;
													assign node4633 = (inp[7]) ? node4639 : node4634;
														assign node4634 = (inp[15]) ? node4636 : 4'b0001;
															assign node4636 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node4639 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node4642 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node4645 = (inp[7]) ? node4651 : node4646;
													assign node4646 = (inp[8]) ? 4'b0011 : node4647;
														assign node4647 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node4651 = (inp[8]) ? node4653 : 4'b0001;
														assign node4653 = (inp[3]) ? 4'b0000 : node4654;
															assign node4654 = (inp[15]) ? 4'b0010 : 4'b0000;
									assign node4658 = (inp[8]) ? node4712 : node4659;
										assign node4659 = (inp[7]) ? node4687 : node4660;
											assign node4660 = (inp[14]) ? node4674 : node4661;
												assign node4661 = (inp[2]) ? node4669 : node4662;
													assign node4662 = (inp[3]) ? node4664 : 4'b0001;
														assign node4664 = (inp[0]) ? node4666 : 4'b0011;
															assign node4666 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node4669 = (inp[3]) ? node4671 : 4'b0000;
														assign node4671 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node4674 = (inp[0]) ? node4678 : node4675;
													assign node4675 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node4678 = (inp[3]) ? node4682 : node4679;
														assign node4679 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node4682 = (inp[15]) ? node4684 : 4'b0010;
															assign node4684 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node4687 = (inp[14]) ? node4699 : node4688;
												assign node4688 = (inp[2]) ? node4692 : node4689;
													assign node4689 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node4692 = (inp[5]) ? node4694 : 4'b1101;
														assign node4694 = (inp[15]) ? 4'b1111 : node4695;
															assign node4695 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node4699 = (inp[5]) ? node4705 : node4700;
													assign node4700 = (inp[2]) ? node4702 : 4'b1101;
														assign node4702 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node4705 = (inp[3]) ? node4707 : 4'b1111;
														assign node4707 = (inp[0]) ? 4'b1101 : node4708;
															assign node4708 = (inp[15]) ? 4'b1111 : 4'b1101;
										assign node4712 = (inp[7]) ? node4728 : node4713;
											assign node4713 = (inp[15]) ? node4719 : node4714;
												assign node4714 = (inp[0]) ? node4716 : 4'b1101;
													assign node4716 = (inp[14]) ? 4'b1111 : 4'b1101;
												assign node4719 = (inp[14]) ? node4723 : node4720;
													assign node4720 = (inp[2]) ? 4'b1111 : 4'b0010;
													assign node4723 = (inp[0]) ? node4725 : 4'b1111;
														assign node4725 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node4728 = (inp[14]) ? node4734 : node4729;
												assign node4729 = (inp[2]) ? 4'b1100 : node4730;
													assign node4730 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node4734 = (inp[15]) ? node4736 : 4'b1100;
													assign node4736 = (inp[0]) ? node4742 : node4737;
														assign node4737 = (inp[5]) ? 4'b1110 : node4738;
															assign node4738 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node4742 = (inp[5]) ? 4'b1100 : node4743;
															assign node4743 = (inp[3]) ? 4'b1100 : 4'b1110;
								assign node4747 = (inp[1]) ? node4837 : node4748;
									assign node4748 = (inp[2]) ? node4802 : node4749;
										assign node4749 = (inp[0]) ? node4779 : node4750;
											assign node4750 = (inp[15]) ? node4760 : node4751;
												assign node4751 = (inp[5]) ? node4753 : 4'b1110;
													assign node4753 = (inp[14]) ? node4755 : 4'b1100;
														assign node4755 = (inp[7]) ? 4'b1101 : node4756;
															assign node4756 = (inp[3]) ? 4'b1101 : 4'b1100;
												assign node4760 = (inp[5]) ? node4768 : node4761;
													assign node4761 = (inp[3]) ? node4763 : 4'b1100;
														assign node4763 = (inp[7]) ? 4'b1110 : node4764;
															assign node4764 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node4768 = (inp[14]) ? node4774 : node4769;
														assign node4769 = (inp[7]) ? node4771 : 4'b1111;
															assign node4771 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node4774 = (inp[8]) ? 4'b1110 : node4775;
															assign node4775 = (inp[7]) ? 4'b1111 : 4'b1110;
											assign node4779 = (inp[14]) ? node4795 : node4780;
												assign node4780 = (inp[15]) ? node4786 : node4781;
													assign node4781 = (inp[3]) ? node4783 : 4'b1100;
														assign node4783 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node4786 = (inp[5]) ? node4790 : node4787;
														assign node4787 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node4790 = (inp[8]) ? 4'b1100 : node4791;
															assign node4791 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node4795 = (inp[3]) ? 4'b1100 : node4796;
													assign node4796 = (inp[5]) ? node4798 : 4'b1110;
														assign node4798 = (inp[7]) ? 4'b1110 : 4'b1111;
										assign node4802 = (inp[5]) ? node4828 : node4803;
											assign node4803 = (inp[7]) ? node4815 : node4804;
												assign node4804 = (inp[8]) ? node4806 : 4'b1110;
													assign node4806 = (inp[15]) ? node4808 : 4'b1111;
														assign node4808 = (inp[14]) ? node4812 : node4809;
															assign node4809 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node4812 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node4815 = (inp[8]) ? node4823 : node4816;
													assign node4816 = (inp[14]) ? 4'b1101 : node4817;
														assign node4817 = (inp[3]) ? node4819 : 4'b1111;
															assign node4819 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node4823 = (inp[15]) ? 4'b1100 : node4824;
														assign node4824 = (inp[3]) ? 4'b1100 : 4'b1110;
											assign node4828 = (inp[0]) ? node4832 : node4829;
												assign node4829 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node4832 = (inp[15]) ? node4834 : 4'b1111;
													assign node4834 = (inp[7]) ? 4'b1101 : 4'b1100;
									assign node4837 = (inp[7]) ? node4871 : node4838;
										assign node4838 = (inp[8]) ? node4856 : node4839;
											assign node4839 = (inp[14]) ? node4845 : node4840;
												assign node4840 = (inp[2]) ? 4'b1110 : node4841;
													assign node4841 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node4845 = (inp[0]) ? node4849 : node4846;
													assign node4846 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node4849 = (inp[3]) ? 4'b1100 : node4850;
														assign node4850 = (inp[2]) ? 4'b1110 : node4851;
															assign node4851 = (inp[15]) ? 4'b1100 : 4'b1100;
											assign node4856 = (inp[2]) ? node4864 : node4857;
												assign node4857 = (inp[14]) ? 4'b0111 : node4858;
													assign node4858 = (inp[3]) ? 4'b1110 : node4859;
														assign node4859 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node4864 = (inp[14]) ? node4866 : 4'b0101;
													assign node4866 = (inp[5]) ? node4868 : 4'b0111;
														assign node4868 = (inp[3]) ? 4'b0111 : 4'b0101;
										assign node4871 = (inp[8]) ? node4897 : node4872;
											assign node4872 = (inp[2]) ? node4886 : node4873;
												assign node4873 = (inp[14]) ? node4883 : node4874;
													assign node4874 = (inp[0]) ? node4878 : node4875;
														assign node4875 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node4878 = (inp[5]) ? node4880 : 4'b1110;
															assign node4880 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node4883 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node4886 = (inp[0]) ? node4888 : 4'b0111;
													assign node4888 = (inp[3]) ? 4'b0101 : node4889;
														assign node4889 = (inp[5]) ? node4893 : node4890;
															assign node4890 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node4893 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node4897 = (inp[14]) ? node4905 : node4898;
												assign node4898 = (inp[2]) ? node4900 : 4'b0101;
													assign node4900 = (inp[0]) ? 4'b0100 : node4901;
														assign node4901 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node4905 = (inp[15]) ? node4911 : node4906;
													assign node4906 = (inp[2]) ? 4'b0100 : node4907;
														assign node4907 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node4911 = (inp[3]) ? 4'b0110 : node4912;
														assign node4912 = (inp[2]) ? 4'b0110 : 4'b0100;
						assign node4916 = (inp[0]) ? node5276 : node4917;
							assign node4917 = (inp[15]) ? node5091 : node4918;
								assign node4918 = (inp[5]) ? node5000 : node4919;
									assign node4919 = (inp[3]) ? node4963 : node4920;
										assign node4920 = (inp[2]) ? node4944 : node4921;
											assign node4921 = (inp[8]) ? node4935 : node4922;
												assign node4922 = (inp[11]) ? node4926 : node4923;
													assign node4923 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node4926 = (inp[6]) ? node4930 : node4927;
														assign node4927 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node4930 = (inp[7]) ? node4932 : 4'b1110;
															assign node4932 = (inp[14]) ? 4'b0111 : 4'b1110;
												assign node4935 = (inp[7]) ? node4941 : node4936;
													assign node4936 = (inp[6]) ? 4'b1111 : node4937;
														assign node4937 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node4941 = (inp[14]) ? 4'b1110 : 4'b1111;
											assign node4944 = (inp[11]) ? node4952 : node4945;
												assign node4945 = (inp[7]) ? node4949 : node4946;
													assign node4946 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node4949 = (inp[1]) ? 4'b1111 : 4'b1110;
												assign node4952 = (inp[8]) ? node4960 : node4953;
													assign node4953 = (inp[7]) ? node4955 : 4'b1110;
														assign node4955 = (inp[6]) ? 4'b1111 : node4956;
															assign node4956 = (inp[1]) ? 4'b1111 : 4'b0111;
													assign node4960 = (inp[7]) ? 4'b1110 : 4'b1111;
										assign node4963 = (inp[7]) ? node4983 : node4964;
											assign node4964 = (inp[8]) ? node4972 : node4965;
												assign node4965 = (inp[14]) ? node4967 : 4'b1101;
													assign node4967 = (inp[1]) ? 4'b0100 : node4968;
														assign node4968 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node4972 = (inp[1]) ? 4'b1101 : node4973;
													assign node4973 = (inp[14]) ? node4975 : 4'b0101;
														assign node4975 = (inp[2]) ? node4979 : node4976;
															assign node4976 = (inp[11]) ? 4'b0101 : 4'b1101;
															assign node4979 = (inp[6]) ? 4'b0101 : 4'b0101;
											assign node4983 = (inp[14]) ? node4993 : node4984;
												assign node4984 = (inp[8]) ? node4990 : node4985;
													assign node4985 = (inp[6]) ? node4987 : 4'b0100;
														assign node4987 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node4990 = (inp[2]) ? 4'b1100 : 4'b0101;
												assign node4993 = (inp[8]) ? node4995 : 4'b0101;
													assign node4995 = (inp[6]) ? 4'b0100 : node4996;
														assign node4996 = (inp[11]) ? 4'b0100 : 4'b1100;
									assign node5000 = (inp[1]) ? node5048 : node5001;
										assign node5001 = (inp[8]) ? node5025 : node5002;
											assign node5002 = (inp[7]) ? node5014 : node5003;
												assign node5003 = (inp[14]) ? node5009 : node5004;
													assign node5004 = (inp[2]) ? node5006 : 4'b1101;
														assign node5006 = (inp[3]) ? 4'b0100 : 4'b1100;
													assign node5009 = (inp[11]) ? node5011 : 4'b1100;
														assign node5011 = (inp[6]) ? 4'b1100 : 4'b0100;
												assign node5014 = (inp[14]) ? node5018 : node5015;
													assign node5015 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node5018 = (inp[2]) ? 4'b1101 : node5019;
														assign node5019 = (inp[6]) ? 4'b0101 : node5020;
															assign node5020 = (inp[11]) ? 4'b0101 : 4'b1101;
											assign node5025 = (inp[3]) ? node5039 : node5026;
												assign node5026 = (inp[6]) ? node5032 : node5027;
													assign node5027 = (inp[7]) ? 4'b1100 : node5028;
														assign node5028 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node5032 = (inp[11]) ? 4'b1100 : node5033;
														assign node5033 = (inp[2]) ? 4'b0100 : node5034;
															assign node5034 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node5039 = (inp[7]) ? node5045 : node5040;
													assign node5040 = (inp[11]) ? node5042 : 4'b0101;
														assign node5042 = (inp[2]) ? 4'b1101 : 4'b0101;
													assign node5045 = (inp[11]) ? 4'b0101 : 4'b1101;
										assign node5048 = (inp[14]) ? node5068 : node5049;
											assign node5049 = (inp[6]) ? node5055 : node5050;
												assign node5050 = (inp[7]) ? 4'b1100 : node5051;
													assign node5051 = (inp[2]) ? 4'b1100 : 4'b0100;
												assign node5055 = (inp[7]) ? node5063 : node5056;
													assign node5056 = (inp[11]) ? node5058 : 4'b0100;
														assign node5058 = (inp[2]) ? node5060 : 4'b1100;
															assign node5060 = (inp[8]) ? 4'b0101 : 4'b1100;
													assign node5063 = (inp[11]) ? node5065 : 4'b0100;
														assign node5065 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node5068 = (inp[8]) ? node5082 : node5069;
												assign node5069 = (inp[7]) ? node5075 : node5070;
													assign node5070 = (inp[11]) ? 4'b1100 : node5071;
														assign node5071 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node5075 = (inp[2]) ? node5077 : 4'b1101;
														assign node5077 = (inp[11]) ? node5079 : 4'b0101;
															assign node5079 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node5082 = (inp[7]) ? node5086 : node5083;
													assign node5083 = (inp[2]) ? 4'b0101 : 4'b1101;
													assign node5086 = (inp[3]) ? 4'b1100 : node5087;
														assign node5087 = (inp[2]) ? 4'b1100 : 4'b0100;
								assign node5091 = (inp[5]) ? node5193 : node5092;
									assign node5092 = (inp[3]) ? node5156 : node5093;
										assign node5093 = (inp[8]) ? node5125 : node5094;
											assign node5094 = (inp[7]) ? node5106 : node5095;
												assign node5095 = (inp[14]) ? node5101 : node5096;
													assign node5096 = (inp[11]) ? node5098 : 4'b1101;
														assign node5098 = (inp[6]) ? 4'b1101 : 4'b0101;
													assign node5101 = (inp[11]) ? node5103 : 4'b0100;
														assign node5103 = (inp[6]) ? 4'b1100 : 4'b0100;
												assign node5106 = (inp[14]) ? node5112 : node5107;
													assign node5107 = (inp[2]) ? 4'b1101 : node5108;
														assign node5108 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node5112 = (inp[1]) ? node5118 : node5113;
														assign node5113 = (inp[6]) ? 4'b0101 : node5114;
															assign node5114 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node5118 = (inp[11]) ? node5122 : node5119;
															assign node5119 = (inp[2]) ? 4'b1101 : 4'b0101;
															assign node5122 = (inp[6]) ? 4'b0101 : 4'b1101;
											assign node5125 = (inp[14]) ? node5145 : node5126;
												assign node5126 = (inp[2]) ? node5138 : node5127;
													assign node5127 = (inp[7]) ? node5133 : node5128;
														assign node5128 = (inp[11]) ? 4'b0100 : node5129;
															assign node5129 = (inp[6]) ? 4'b0100 : 4'b1100;
														assign node5133 = (inp[1]) ? 4'b1101 : node5134;
															assign node5134 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node5138 = (inp[7]) ? node5140 : 4'b0101;
														assign node5140 = (inp[6]) ? node5142 : 4'b0100;
															assign node5142 = (inp[11]) ? 4'b1100 : 4'b0100;
												assign node5145 = (inp[7]) ? node5153 : node5146;
													assign node5146 = (inp[11]) ? node5150 : node5147;
														assign node5147 = (inp[1]) ? 4'b0101 : 4'b1101;
														assign node5150 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node5153 = (inp[2]) ? 4'b1100 : 4'b0100;
										assign node5156 = (inp[11]) ? node5182 : node5157;
											assign node5157 = (inp[6]) ? node5169 : node5158;
												assign node5158 = (inp[1]) ? node5164 : node5159;
													assign node5159 = (inp[14]) ? node5161 : 4'b1111;
														assign node5161 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node5164 = (inp[14]) ? node5166 : 4'b1110;
														assign node5166 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node5169 = (inp[1]) ? node5175 : node5170;
													assign node5170 = (inp[14]) ? node5172 : 4'b0110;
														assign node5172 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node5175 = (inp[14]) ? node5177 : 4'b0111;
														assign node5177 = (inp[2]) ? 4'b1111 : node5178;
															assign node5178 = (inp[7]) ? 4'b1110 : 4'b0110;
											assign node5182 = (inp[1]) ? node5186 : node5183;
												assign node5183 = (inp[6]) ? 4'b1110 : 4'b0110;
												assign node5186 = (inp[14]) ? 4'b0110 : node5187;
													assign node5187 = (inp[8]) ? node5189 : 4'b0111;
														assign node5189 = (inp[7]) ? 4'b0110 : 4'b0111;
									assign node5193 = (inp[1]) ? node5229 : node5194;
										assign node5194 = (inp[8]) ? node5208 : node5195;
											assign node5195 = (inp[7]) ? node5203 : node5196;
												assign node5196 = (inp[2]) ? node5198 : 4'b0111;
													assign node5198 = (inp[14]) ? node5200 : 4'b1110;
														assign node5200 = (inp[3]) ? 4'b0110 : 4'b1110;
												assign node5203 = (inp[11]) ? 4'b0111 : node5204;
													assign node5204 = (inp[6]) ? 4'b0111 : 4'b1111;
											assign node5208 = (inp[7]) ? node5222 : node5209;
												assign node5209 = (inp[2]) ? node5217 : node5210;
													assign node5210 = (inp[14]) ? 4'b1111 : node5211;
														assign node5211 = (inp[11]) ? 4'b1110 : node5212;
															assign node5212 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node5217 = (inp[6]) ? node5219 : 4'b1111;
														assign node5219 = (inp[11]) ? 4'b1111 : 4'b0111;
												assign node5222 = (inp[6]) ? node5226 : node5223;
													assign node5223 = (inp[11]) ? 4'b0110 : 4'b1110;
													assign node5226 = (inp[11]) ? 4'b1110 : 4'b0110;
										assign node5229 = (inp[11]) ? node5251 : node5230;
											assign node5230 = (inp[14]) ? node5242 : node5231;
												assign node5231 = (inp[6]) ? node5237 : node5232;
													assign node5232 = (inp[3]) ? 4'b1110 : node5233;
														assign node5233 = (inp[8]) ? 4'b0111 : 4'b1110;
													assign node5237 = (inp[8]) ? 4'b1111 : node5238;
														assign node5238 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node5242 = (inp[8]) ? node5248 : node5243;
													assign node5243 = (inp[3]) ? node5245 : 4'b1111;
														assign node5245 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node5248 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node5251 = (inp[7]) ? node5269 : node5252;
												assign node5252 = (inp[2]) ? node5264 : node5253;
													assign node5253 = (inp[6]) ? node5259 : node5254;
														assign node5254 = (inp[14]) ? 4'b0110 : node5255;
															assign node5255 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node5259 = (inp[8]) ? 4'b0111 : node5260;
															assign node5260 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node5264 = (inp[8]) ? node5266 : 4'b0110;
														assign node5266 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node5269 = (inp[6]) ? 4'b0111 : node5270;
													assign node5270 = (inp[14]) ? node5272 : 4'b1111;
														assign node5272 = (inp[2]) ? 4'b1111 : 4'b1110;
							assign node5276 = (inp[15]) ? node5454 : node5277;
								assign node5277 = (inp[3]) ? node5367 : node5278;
									assign node5278 = (inp[5]) ? node5314 : node5279;
										assign node5279 = (inp[2]) ? node5303 : node5280;
											assign node5280 = (inp[1]) ? node5292 : node5281;
												assign node5281 = (inp[6]) ? node5285 : node5282;
													assign node5282 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node5285 = (inp[11]) ? node5289 : node5286;
														assign node5286 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node5289 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node5292 = (inp[14]) ? node5298 : node5293;
													assign node5293 = (inp[11]) ? node5295 : 4'b0101;
														assign node5295 = (inp[6]) ? 4'b0101 : 4'b0100;
													assign node5298 = (inp[6]) ? node5300 : 4'b0100;
														assign node5300 = (inp[11]) ? 4'b0100 : 4'b1100;
											assign node5303 = (inp[6]) ? node5307 : node5304;
												assign node5304 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node5307 = (inp[1]) ? 4'b1101 : node5308;
													assign node5308 = (inp[11]) ? node5310 : 4'b0100;
														assign node5310 = (inp[7]) ? 4'b1101 : 4'b1100;
										assign node5314 = (inp[6]) ? node5340 : node5315;
											assign node5315 = (inp[2]) ? node5331 : node5316;
												assign node5316 = (inp[11]) ? node5318 : 4'b0111;
													assign node5318 = (inp[1]) ? node5324 : node5319;
														assign node5319 = (inp[8]) ? node5321 : 4'b0111;
															assign node5321 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node5324 = (inp[14]) ? node5328 : node5325;
															assign node5325 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node5328 = (inp[7]) ? 4'b1110 : 4'b0110;
												assign node5331 = (inp[7]) ? node5333 : 4'b1111;
													assign node5333 = (inp[8]) ? 4'b0110 : node5334;
														assign node5334 = (inp[1]) ? node5336 : 4'b0111;
															assign node5336 = (inp[11]) ? 4'b1111 : 4'b0111;
											assign node5340 = (inp[11]) ? node5354 : node5341;
												assign node5341 = (inp[1]) ? node5349 : node5342;
													assign node5342 = (inp[2]) ? 4'b0111 : node5343;
														assign node5343 = (inp[14]) ? node5345 : 4'b0110;
															assign node5345 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node5349 = (inp[14]) ? node5351 : 4'b1111;
														assign node5351 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node5354 = (inp[1]) ? node5364 : node5355;
													assign node5355 = (inp[14]) ? 4'b1111 : node5356;
														assign node5356 = (inp[8]) ? node5360 : node5357;
															assign node5357 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node5360 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node5364 = (inp[7]) ? 4'b0110 : 4'b1110;
									assign node5367 = (inp[8]) ? node5419 : node5368;
										assign node5368 = (inp[7]) ? node5392 : node5369;
											assign node5369 = (inp[2]) ? node5379 : node5370;
												assign node5370 = (inp[14]) ? node5374 : node5371;
													assign node5371 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node5374 = (inp[11]) ? 4'b1110 : node5375;
														assign node5375 = (inp[6]) ? 4'b0110 : 4'b1110;
												assign node5379 = (inp[5]) ? node5385 : node5380;
													assign node5380 = (inp[6]) ? 4'b0110 : node5381;
														assign node5381 = (inp[11]) ? 4'b0110 : 4'b1110;
													assign node5385 = (inp[14]) ? node5389 : node5386;
														assign node5386 = (inp[1]) ? 4'b0110 : 4'b1110;
														assign node5389 = (inp[11]) ? 4'b1110 : 4'b0110;
											assign node5392 = (inp[2]) ? node5406 : node5393;
												assign node5393 = (inp[14]) ? node5399 : node5394;
													assign node5394 = (inp[11]) ? 4'b1110 : node5395;
														assign node5395 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node5399 = (inp[1]) ? node5401 : 4'b0111;
														assign node5401 = (inp[11]) ? 4'b1111 : node5402;
															assign node5402 = (inp[6]) ? 4'b1111 : 4'b0111;
												assign node5406 = (inp[6]) ? node5412 : node5407;
													assign node5407 = (inp[14]) ? node5409 : 4'b0111;
														assign node5409 = (inp[1]) ? 4'b1111 : 4'b0111;
													assign node5412 = (inp[11]) ? node5416 : node5413;
														assign node5413 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node5416 = (inp[5]) ? 4'b1111 : 4'b0111;
										assign node5419 = (inp[7]) ? node5443 : node5420;
											assign node5420 = (inp[2]) ? node5430 : node5421;
												assign node5421 = (inp[14]) ? node5427 : node5422;
													assign node5422 = (inp[5]) ? node5424 : 4'b0110;
														assign node5424 = (inp[11]) ? 4'b0110 : 4'b1110;
													assign node5427 = (inp[5]) ? 4'b1111 : 4'b0111;
												assign node5430 = (inp[14]) ? node5436 : node5431;
													assign node5431 = (inp[6]) ? node5433 : 4'b0111;
														assign node5433 = (inp[11]) ? 4'b1111 : 4'b0111;
													assign node5436 = (inp[1]) ? node5438 : 4'b0111;
														assign node5438 = (inp[6]) ? node5440 : 4'b1111;
															assign node5440 = (inp[11]) ? 4'b0111 : 4'b1111;
											assign node5443 = (inp[1]) ? node5451 : node5444;
												assign node5444 = (inp[14]) ? node5446 : 4'b1111;
													assign node5446 = (inp[6]) ? node5448 : 4'b1110;
														assign node5448 = (inp[11]) ? 4'b1110 : 4'b0110;
												assign node5451 = (inp[2]) ? 4'b0110 : 4'b0111;
								assign node5454 = (inp[5]) ? node5546 : node5455;
									assign node5455 = (inp[3]) ? node5499 : node5456;
										assign node5456 = (inp[8]) ? node5480 : node5457;
											assign node5457 = (inp[7]) ? node5473 : node5458;
												assign node5458 = (inp[1]) ? node5464 : node5459;
													assign node5459 = (inp[14]) ? 4'b0110 : node5460;
														assign node5460 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node5464 = (inp[2]) ? node5468 : node5465;
														assign node5465 = (inp[14]) ? 4'b0110 : 4'b1111;
														assign node5468 = (inp[14]) ? 4'b1110 : node5469;
															assign node5469 = (inp[6]) ? 4'b1110 : 4'b0110;
												assign node5473 = (inp[14]) ? node5475 : 4'b0110;
													assign node5475 = (inp[1]) ? 4'b0111 : node5476;
														assign node5476 = (inp[6]) ? 4'b0111 : 4'b1111;
											assign node5480 = (inp[7]) ? node5494 : node5481;
												assign node5481 = (inp[1]) ? node5489 : node5482;
													assign node5482 = (inp[2]) ? node5484 : 4'b1110;
														assign node5484 = (inp[14]) ? 4'b1111 : node5485;
															assign node5485 = (inp[11]) ? 4'b1111 : 4'b0111;
													assign node5489 = (inp[14]) ? 4'b0111 : node5490;
														assign node5490 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node5494 = (inp[2]) ? 4'b0110 : node5495;
													assign node5495 = (inp[14]) ? 4'b1110 : 4'b1111;
										assign node5499 = (inp[2]) ? node5527 : node5500;
											assign node5500 = (inp[1]) ? node5518 : node5501;
												assign node5501 = (inp[6]) ? node5509 : node5502;
													assign node5502 = (inp[11]) ? 4'b0101 : node5503;
														assign node5503 = (inp[7]) ? 4'b1100 : node5504;
															assign node5504 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node5509 = (inp[11]) ? node5513 : node5510;
														assign node5510 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node5513 = (inp[8]) ? node5515 : 4'b1100;
															assign node5515 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node5518 = (inp[11]) ? node5524 : node5519;
													assign node5519 = (inp[6]) ? 4'b0100 : node5520;
														assign node5520 = (inp[8]) ? 4'b0100 : 4'b1100;
													assign node5524 = (inp[8]) ? 4'b1101 : 4'b1100;
											assign node5527 = (inp[11]) ? node5529 : 4'b1100;
												assign node5529 = (inp[14]) ? node5539 : node5530;
													assign node5530 = (inp[1]) ? node5534 : node5531;
														assign node5531 = (inp[8]) ? 4'b0101 : 4'b1100;
														assign node5534 = (inp[6]) ? node5536 : 4'b0100;
															assign node5536 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node5539 = (inp[1]) ? 4'b1101 : node5540;
														assign node5540 = (inp[8]) ? node5542 : 4'b0101;
															assign node5542 = (inp[7]) ? 4'b0100 : 4'b0101;
									assign node5546 = (inp[3]) ? node5600 : node5547;
										assign node5547 = (inp[2]) ? node5567 : node5548;
											assign node5548 = (inp[1]) ? node5562 : node5549;
												assign node5549 = (inp[8]) ? node5557 : node5550;
													assign node5550 = (inp[6]) ? node5554 : node5551;
														assign node5551 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node5554 = (inp[14]) ? 4'b0100 : 4'b1100;
													assign node5557 = (inp[6]) ? node5559 : 4'b0101;
														assign node5559 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node5562 = (inp[11]) ? 4'b1100 : node5563;
													assign node5563 = (inp[6]) ? 4'b0101 : 4'b1100;
											assign node5567 = (inp[14]) ? node5585 : node5568;
												assign node5568 = (inp[6]) ? node5576 : node5569;
													assign node5569 = (inp[11]) ? 4'b0100 : node5570;
														assign node5570 = (inp[8]) ? node5572 : 4'b0101;
															assign node5572 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node5576 = (inp[7]) ? node5578 : 4'b0101;
														assign node5578 = (inp[8]) ? node5582 : node5579;
															assign node5579 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node5582 = (inp[1]) ? 4'b1100 : 4'b0100;
												assign node5585 = (inp[7]) ? node5593 : node5586;
													assign node5586 = (inp[6]) ? node5590 : node5587;
														assign node5587 = (inp[11]) ? 4'b0100 : 4'b1100;
														assign node5590 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node5593 = (inp[8]) ? 4'b0100 : node5594;
														assign node5594 = (inp[11]) ? 4'b0101 : node5595;
															assign node5595 = (inp[6]) ? 4'b0101 : 4'b1101;
										assign node5600 = (inp[14]) ? node5624 : node5601;
											assign node5601 = (inp[1]) ? node5619 : node5602;
												assign node5602 = (inp[6]) ? node5610 : node5603;
													assign node5603 = (inp[11]) ? 4'b0101 : node5604;
														assign node5604 = (inp[2]) ? 4'b1101 : node5605;
															assign node5605 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node5610 = (inp[11]) ? node5616 : node5611;
														assign node5611 = (inp[7]) ? 4'b0100 : node5612;
															assign node5612 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node5616 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node5619 = (inp[6]) ? node5621 : 4'b0100;
													assign node5621 = (inp[11]) ? 4'b0101 : 4'b1101;
											assign node5624 = (inp[1]) ? node5636 : node5625;
												assign node5625 = (inp[2]) ? node5631 : node5626;
													assign node5626 = (inp[8]) ? node5628 : 4'b0100;
														assign node5628 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node5631 = (inp[6]) ? node5633 : 4'b0101;
														assign node5633 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node5636 = (inp[8]) ? node5642 : node5637;
													assign node5637 = (inp[11]) ? node5639 : 4'b0101;
														assign node5639 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node5642 = (inp[7]) ? 4'b1100 : node5643;
														assign node5643 = (inp[6]) ? 4'b1101 : node5644;
															assign node5644 = (inp[11]) ? 4'b1101 : 4'b0101;
			assign node5649 = (inp[4]) ? node8381 : node5650;
				assign node5650 = (inp[10]) ? node7052 : node5651;
					assign node5651 = (inp[12]) ? node6383 : node5652;
						assign node5652 = (inp[0]) ? node6000 : node5653;
							assign node5653 = (inp[15]) ? node5823 : node5654;
								assign node5654 = (inp[3]) ? node5726 : node5655;
									assign node5655 = (inp[11]) ? node5687 : node5656;
										assign node5656 = (inp[2]) ? node5668 : node5657;
											assign node5657 = (inp[6]) ? node5661 : node5658;
												assign node5658 = (inp[1]) ? 4'b1010 : 4'b1011;
												assign node5661 = (inp[14]) ? node5665 : node5662;
													assign node5662 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node5665 = (inp[1]) ? 4'b1011 : 4'b0010;
											assign node5668 = (inp[8]) ? node5676 : node5669;
												assign node5669 = (inp[14]) ? node5673 : node5670;
													assign node5670 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node5673 = (inp[6]) ? 4'b1011 : 4'b0011;
												assign node5676 = (inp[7]) ? node5682 : node5677;
													assign node5677 = (inp[6]) ? 4'b0011 : node5678;
														assign node5678 = (inp[5]) ? 4'b0011 : 4'b1011;
													assign node5682 = (inp[1]) ? node5684 : 4'b0010;
														assign node5684 = (inp[6]) ? 4'b1010 : 4'b0010;
										assign node5687 = (inp[6]) ? node5697 : node5688;
											assign node5688 = (inp[8]) ? 4'b1011 : node5689;
												assign node5689 = (inp[7]) ? node5691 : 4'b0010;
													assign node5691 = (inp[1]) ? 4'b1011 : node5692;
														assign node5692 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node5697 = (inp[1]) ? node5715 : node5698;
												assign node5698 = (inp[2]) ? node5708 : node5699;
													assign node5699 = (inp[8]) ? node5701 : 4'b1010;
														assign node5701 = (inp[7]) ? node5705 : node5702;
															assign node5702 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node5705 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node5708 = (inp[5]) ? 4'b1011 : node5709;
														assign node5709 = (inp[14]) ? 4'b1011 : node5710;
															assign node5710 = (inp[8]) ? 4'b1010 : 4'b1010;
												assign node5715 = (inp[7]) ? 4'b0010 : node5716;
													assign node5716 = (inp[5]) ? 4'b1010 : node5717;
														assign node5717 = (inp[8]) ? node5721 : node5718;
															assign node5718 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node5721 = (inp[2]) ? 4'b0011 : 4'b1010;
									assign node5726 = (inp[5]) ? node5764 : node5727;
										assign node5727 = (inp[8]) ? node5745 : node5728;
											assign node5728 = (inp[2]) ? node5734 : node5729;
												assign node5729 = (inp[14]) ? 4'b1011 : node5730;
													assign node5730 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node5734 = (inp[7]) ? node5740 : node5735;
													assign node5735 = (inp[14]) ? node5737 : 4'b1010;
														assign node5737 = (inp[11]) ? 4'b0010 : 4'b1010;
													assign node5740 = (inp[6]) ? 4'b0011 : node5741;
														assign node5741 = (inp[1]) ? 4'b0011 : 4'b1011;
											assign node5745 = (inp[7]) ? node5751 : node5746;
												assign node5746 = (inp[11]) ? 4'b1011 : node5747;
													assign node5747 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node5751 = (inp[2]) ? node5755 : node5752;
													assign node5752 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node5755 = (inp[11]) ? node5757 : 4'b1010;
														assign node5757 = (inp[6]) ? node5761 : node5758;
															assign node5758 = (inp[1]) ? 4'b1010 : 4'b0010;
															assign node5761 = (inp[1]) ? 4'b0010 : 4'b1010;
										assign node5764 = (inp[8]) ? node5794 : node5765;
											assign node5765 = (inp[7]) ? node5779 : node5766;
												assign node5766 = (inp[11]) ? node5772 : node5767;
													assign node5767 = (inp[6]) ? node5769 : 4'b1000;
														assign node5769 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node5772 = (inp[6]) ? node5774 : 4'b0000;
														assign node5774 = (inp[14]) ? 4'b1000 : node5775;
															assign node5775 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node5779 = (inp[2]) ? node5787 : node5780;
													assign node5780 = (inp[14]) ? 4'b1001 : node5781;
														assign node5781 = (inp[1]) ? 4'b1000 : node5782;
															assign node5782 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node5787 = (inp[6]) ? node5789 : 4'b0001;
														assign node5789 = (inp[14]) ? node5791 : 4'b0001;
															assign node5791 = (inp[11]) ? 4'b1001 : 4'b0001;
											assign node5794 = (inp[6]) ? node5808 : node5795;
												assign node5795 = (inp[7]) ? node5801 : node5796;
													assign node5796 = (inp[14]) ? 4'b1001 : node5797;
														assign node5797 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node5801 = (inp[14]) ? 4'b1000 : node5802;
														assign node5802 = (inp[2]) ? 4'b1000 : node5803;
															assign node5803 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node5808 = (inp[2]) ? node5814 : node5809;
													assign node5809 = (inp[11]) ? 4'b1000 : node5810;
														assign node5810 = (inp[7]) ? 4'b1001 : 4'b0000;
													assign node5814 = (inp[7]) ? 4'b0000 : node5815;
														assign node5815 = (inp[14]) ? node5819 : node5816;
															assign node5816 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node5819 = (inp[1]) ? 4'b0001 : 4'b0001;
								assign node5823 = (inp[5]) ? node5921 : node5824;
									assign node5824 = (inp[1]) ? node5880 : node5825;
										assign node5825 = (inp[8]) ? node5847 : node5826;
											assign node5826 = (inp[7]) ? node5838 : node5827;
												assign node5827 = (inp[14]) ? 4'b1000 : node5828;
													assign node5828 = (inp[2]) ? node5832 : node5829;
														assign node5829 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node5832 = (inp[3]) ? node5834 : 4'b1000;
															assign node5834 = (inp[11]) ? 4'b1000 : 4'b0000;
												assign node5838 = (inp[14]) ? node5844 : node5839;
													assign node5839 = (inp[2]) ? 4'b0001 : node5840;
														assign node5840 = (inp[3]) ? 4'b0000 : 4'b1000;
													assign node5844 = (inp[3]) ? 4'b0001 : 4'b1001;
											assign node5847 = (inp[7]) ? node5869 : node5848;
												assign node5848 = (inp[2]) ? node5856 : node5849;
													assign node5849 = (inp[14]) ? node5853 : node5850;
														assign node5850 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node5853 = (inp[6]) ? 4'b1001 : 4'b0001;
													assign node5856 = (inp[14]) ? node5862 : node5857;
														assign node5857 = (inp[3]) ? 4'b1001 : node5858;
															assign node5858 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node5862 = (inp[6]) ? node5866 : node5863;
															assign node5863 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node5866 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node5869 = (inp[2]) ? node5877 : node5870;
													assign node5870 = (inp[14]) ? 4'b1000 : node5871;
														assign node5871 = (inp[3]) ? 4'b0001 : node5872;
															assign node5872 = (inp[6]) ? 4'b1001 : 4'b0001;
													assign node5877 = (inp[11]) ? 4'b1000 : 4'b0000;
										assign node5880 = (inp[7]) ? node5898 : node5881;
											assign node5881 = (inp[8]) ? node5891 : node5882;
												assign node5882 = (inp[3]) ? 4'b1000 : node5883;
													assign node5883 = (inp[14]) ? node5885 : 4'b1001;
														assign node5885 = (inp[2]) ? node5887 : 4'b0000;
															assign node5887 = (inp[6]) ? 4'b0000 : 4'b1000;
												assign node5891 = (inp[14]) ? node5895 : node5892;
													assign node5892 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node5895 = (inp[6]) ? 4'b1001 : 4'b0001;
											assign node5898 = (inp[8]) ? node5912 : node5899;
												assign node5899 = (inp[2]) ? node5907 : node5900;
													assign node5900 = (inp[14]) ? 4'b1001 : node5901;
														assign node5901 = (inp[11]) ? 4'b1000 : node5902;
															assign node5902 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node5907 = (inp[3]) ? node5909 : 4'b0001;
														assign node5909 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node5912 = (inp[14]) ? node5914 : 4'b0001;
													assign node5914 = (inp[2]) ? 4'b1000 : node5915;
														assign node5915 = (inp[11]) ? node5917 : 4'b0000;
															assign node5917 = (inp[6]) ? 4'b0000 : 4'b1000;
									assign node5921 = (inp[3]) ? node5961 : node5922;
										assign node5922 = (inp[2]) ? node5940 : node5923;
											assign node5923 = (inp[11]) ? node5927 : node5924;
												assign node5924 = (inp[6]) ? 4'b0000 : 4'b1000;
												assign node5927 = (inp[6]) ? node5937 : node5928;
													assign node5928 = (inp[7]) ? node5932 : node5929;
														assign node5929 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node5932 = (inp[1]) ? 4'b1001 : node5933;
															assign node5933 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node5937 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node5940 = (inp[8]) ? node5950 : node5941;
												assign node5941 = (inp[7]) ? node5943 : 4'b1000;
													assign node5943 = (inp[11]) ? 4'b1001 : node5944;
														assign node5944 = (inp[6]) ? node5946 : 4'b0001;
															assign node5946 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node5950 = (inp[7]) ? node5954 : node5951;
													assign node5951 = (inp[14]) ? 4'b0001 : 4'b1001;
													assign node5954 = (inp[14]) ? node5958 : node5955;
														assign node5955 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node5958 = (inp[1]) ? 4'b1000 : 4'b0000;
										assign node5961 = (inp[7]) ? node5977 : node5962;
											assign node5962 = (inp[8]) ? 4'b1011 : node5963;
												assign node5963 = (inp[2]) ? node5971 : node5964;
													assign node5964 = (inp[14]) ? 4'b1010 : node5965;
														assign node5965 = (inp[6]) ? 4'b1011 : node5966;
															assign node5966 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node5971 = (inp[6]) ? 4'b1010 : node5972;
														assign node5972 = (inp[11]) ? 4'b0010 : 4'b1010;
											assign node5977 = (inp[8]) ? node5989 : node5978;
												assign node5978 = (inp[14]) ? node5982 : node5979;
													assign node5979 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node5982 = (inp[1]) ? node5986 : node5983;
														assign node5983 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node5986 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node5989 = (inp[2]) ? node5993 : node5990;
													assign node5990 = (inp[6]) ? 4'b1010 : 4'b1011;
													assign node5993 = (inp[6]) ? node5995 : 4'b0010;
														assign node5995 = (inp[14]) ? 4'b1010 : node5996;
															assign node5996 = (inp[1]) ? 4'b1010 : 4'b0010;
							assign node6000 = (inp[15]) ? node6204 : node6001;
								assign node6001 = (inp[5]) ? node6099 : node6002;
									assign node6002 = (inp[3]) ? node6052 : node6003;
										assign node6003 = (inp[8]) ? node6023 : node6004;
											assign node6004 = (inp[7]) ? node6010 : node6005;
												assign node6005 = (inp[11]) ? node6007 : 4'b1000;
													assign node6007 = (inp[6]) ? 4'b1000 : 4'b0000;
												assign node6010 = (inp[2]) ? node6018 : node6011;
													assign node6011 = (inp[14]) ? 4'b1001 : node6012;
														assign node6012 = (inp[6]) ? 4'b0000 : node6013;
															assign node6013 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node6018 = (inp[6]) ? 4'b0001 : node6019;
														assign node6019 = (inp[11]) ? 4'b1001 : 4'b0001;
											assign node6023 = (inp[2]) ? node6041 : node6024;
												assign node6024 = (inp[6]) ? node6032 : node6025;
													assign node6025 = (inp[7]) ? node6029 : node6026;
														assign node6026 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node6029 = (inp[11]) ? 4'b1001 : 4'b0001;
													assign node6032 = (inp[7]) ? node6036 : node6033;
														assign node6033 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node6036 = (inp[11]) ? 4'b1000 : node6037;
															assign node6037 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node6041 = (inp[7]) ? node6045 : node6042;
													assign node6042 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node6045 = (inp[1]) ? 4'b1000 : node6046;
														assign node6046 = (inp[6]) ? node6048 : 4'b1000;
															assign node6048 = (inp[11]) ? 4'b1000 : 4'b0000;
										assign node6052 = (inp[11]) ? node6082 : node6053;
											assign node6053 = (inp[6]) ? node6065 : node6054;
												assign node6054 = (inp[7]) ? node6062 : node6055;
													assign node6055 = (inp[8]) ? node6057 : 4'b1000;
														assign node6057 = (inp[14]) ? 4'b0001 : node6058;
															assign node6058 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node6062 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node6065 = (inp[7]) ? node6073 : node6066;
													assign node6066 = (inp[8]) ? 4'b0001 : node6067;
														assign node6067 = (inp[2]) ? 4'b0000 : node6068;
															assign node6068 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node6073 = (inp[1]) ? node6075 : 4'b0000;
														assign node6075 = (inp[14]) ? node6079 : node6076;
															assign node6076 = (inp[8]) ? 4'b1001 : 4'b0000;
															assign node6079 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node6082 = (inp[6]) ? node6092 : node6083;
												assign node6083 = (inp[1]) ? 4'b1001 : node6084;
													assign node6084 = (inp[7]) ? node6086 : 4'b0001;
														assign node6086 = (inp[8]) ? node6088 : 4'b0001;
															assign node6088 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node6092 = (inp[2]) ? node6094 : 4'b1000;
													assign node6094 = (inp[1]) ? 4'b0001 : node6095;
														assign node6095 = (inp[7]) ? 4'b1001 : 4'b1000;
									assign node6099 = (inp[3]) ? node6143 : node6100;
										assign node6100 = (inp[1]) ? node6118 : node6101;
											assign node6101 = (inp[6]) ? node6113 : node6102;
												assign node6102 = (inp[11]) ? node6110 : node6103;
													assign node6103 = (inp[8]) ? node6105 : 4'b1001;
														assign node6105 = (inp[7]) ? node6107 : 4'b1000;
															assign node6107 = (inp[14]) ? 4'b1000 : 4'b1000;
													assign node6110 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node6113 = (inp[8]) ? 4'b0001 : node6114;
													assign node6114 = (inp[11]) ? 4'b1000 : 4'b0000;
											assign node6118 = (inp[6]) ? node6128 : node6119;
												assign node6119 = (inp[11]) ? node6125 : node6120;
													assign node6120 = (inp[8]) ? node6122 : 4'b1000;
														assign node6122 = (inp[2]) ? 4'b0000 : 4'b1000;
													assign node6125 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node6128 = (inp[11]) ? node6136 : node6129;
													assign node6129 = (inp[7]) ? node6133 : node6130;
														assign node6130 = (inp[2]) ? 4'b1001 : 4'b0000;
														assign node6133 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node6136 = (inp[7]) ? 4'b0000 : node6137;
														assign node6137 = (inp[14]) ? 4'b1000 : node6138;
															assign node6138 = (inp[2]) ? 4'b0001 : 4'b1000;
										assign node6143 = (inp[11]) ? node6175 : node6144;
											assign node6144 = (inp[6]) ? node6162 : node6145;
												assign node6145 = (inp[1]) ? node6153 : node6146;
													assign node6146 = (inp[7]) ? 4'b1010 : node6147;
														assign node6147 = (inp[14]) ? 4'b1010 : node6148;
															assign node6148 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node6153 = (inp[7]) ? node6159 : node6154;
														assign node6154 = (inp[14]) ? 4'b0011 : node6155;
															assign node6155 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node6159 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node6162 = (inp[1]) ? node6170 : node6163;
													assign node6163 = (inp[8]) ? node6165 : 4'b0010;
														assign node6165 = (inp[2]) ? 4'b0010 : node6166;
															assign node6166 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node6170 = (inp[14]) ? node6172 : 4'b0010;
														assign node6172 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node6175 = (inp[2]) ? node6191 : node6176;
												assign node6176 = (inp[8]) ? node6186 : node6177;
													assign node6177 = (inp[1]) ? node6179 : 4'b1011;
														assign node6179 = (inp[14]) ? node6183 : node6180;
															assign node6180 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node6183 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node6186 = (inp[14]) ? 4'b0011 : node6187;
														assign node6187 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node6191 = (inp[8]) ? 4'b1010 : node6192;
													assign node6192 = (inp[7]) ? node6196 : node6193;
														assign node6193 = (inp[1]) ? 4'b1010 : 4'b0010;
														assign node6196 = (inp[1]) ? node6200 : node6197;
															assign node6197 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node6200 = (inp[14]) ? 4'b0011 : 4'b1011;
								assign node6204 = (inp[3]) ? node6292 : node6205;
									assign node6205 = (inp[8]) ? node6239 : node6206;
										assign node6206 = (inp[7]) ? node6218 : node6207;
											assign node6207 = (inp[14]) ? node6213 : node6208;
												assign node6208 = (inp[2]) ? node6210 : 4'b0011;
													assign node6210 = (inp[11]) ? 4'b1010 : 4'b0010;
												assign node6213 = (inp[6]) ? node6215 : 4'b1010;
													assign node6215 = (inp[11]) ? 4'b1010 : 4'b0010;
											assign node6218 = (inp[14]) ? node6222 : node6219;
												assign node6219 = (inp[2]) ? 4'b1011 : 4'b0010;
												assign node6222 = (inp[2]) ? node6230 : node6223;
													assign node6223 = (inp[11]) ? node6225 : 4'b0011;
														assign node6225 = (inp[6]) ? 4'b0011 : node6226;
															assign node6226 = (inp[1]) ? 4'b1011 : 4'b0011;
													assign node6230 = (inp[1]) ? 4'b0011 : node6231;
														assign node6231 = (inp[5]) ? node6235 : node6232;
															assign node6232 = (inp[11]) ? 4'b0011 : 4'b1011;
															assign node6235 = (inp[11]) ? 4'b1011 : 4'b0011;
										assign node6239 = (inp[7]) ? node6275 : node6240;
											assign node6240 = (inp[2]) ? node6256 : node6241;
												assign node6241 = (inp[14]) ? node6247 : node6242;
													assign node6242 = (inp[11]) ? 4'b1010 : node6243;
														assign node6243 = (inp[1]) ? 4'b0010 : 4'b1010;
													assign node6247 = (inp[5]) ? node6249 : 4'b1011;
														assign node6249 = (inp[11]) ? node6253 : node6250;
															assign node6250 = (inp[6]) ? 4'b0011 : 4'b1011;
															assign node6253 = (inp[6]) ? 4'b1011 : 4'b0011;
												assign node6256 = (inp[5]) ? node6266 : node6257;
													assign node6257 = (inp[6]) ? node6259 : 4'b1011;
														assign node6259 = (inp[11]) ? node6263 : node6260;
															assign node6260 = (inp[1]) ? 4'b1011 : 4'b0011;
															assign node6263 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node6266 = (inp[11]) ? 4'b0011 : node6267;
														assign node6267 = (inp[1]) ? node6271 : node6268;
															assign node6268 = (inp[6]) ? 4'b0011 : 4'b1011;
															assign node6271 = (inp[6]) ? 4'b1011 : 4'b0011;
											assign node6275 = (inp[14]) ? node6285 : node6276;
												assign node6276 = (inp[2]) ? 4'b0010 : node6277;
													assign node6277 = (inp[1]) ? node6279 : 4'b1011;
														assign node6279 = (inp[6]) ? node6281 : 4'b0011;
															assign node6281 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node6285 = (inp[6]) ? node6287 : 4'b1010;
													assign node6287 = (inp[2]) ? node6289 : 4'b1010;
														assign node6289 = (inp[5]) ? 4'b0010 : 4'b1010;
									assign node6292 = (inp[5]) ? node6340 : node6293;
										assign node6293 = (inp[2]) ? node6317 : node6294;
											assign node6294 = (inp[11]) ? node6302 : node6295;
												assign node6295 = (inp[6]) ? node6297 : 4'b1010;
													assign node6297 = (inp[7]) ? node6299 : 4'b0010;
														assign node6299 = (inp[8]) ? 4'b1011 : 4'b0010;
												assign node6302 = (inp[1]) ? node6310 : node6303;
													assign node6303 = (inp[6]) ? 4'b1010 : node6304;
														assign node6304 = (inp[8]) ? node6306 : 4'b0011;
															assign node6306 = (inp[7]) ? 4'b0010 : 4'b0010;
													assign node6310 = (inp[6]) ? 4'b0011 : node6311;
														assign node6311 = (inp[7]) ? node6313 : 4'b1011;
															assign node6313 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node6317 = (inp[8]) ? node6327 : node6318;
												assign node6318 = (inp[7]) ? node6320 : 4'b1010;
													assign node6320 = (inp[6]) ? 4'b1011 : node6321;
														assign node6321 = (inp[1]) ? node6323 : 4'b1011;
															assign node6323 = (inp[11]) ? 4'b1011 : 4'b0011;
												assign node6327 = (inp[7]) ? node6337 : node6328;
													assign node6328 = (inp[11]) ? node6332 : node6329;
														assign node6329 = (inp[14]) ? 4'b0011 : 4'b1011;
														assign node6332 = (inp[6]) ? 4'b0011 : node6333;
															assign node6333 = (inp[1]) ? 4'b1011 : 4'b0011;
													assign node6337 = (inp[11]) ? 4'b1010 : 4'b0010;
										assign node6340 = (inp[11]) ? node6364 : node6341;
											assign node6341 = (inp[8]) ? node6349 : node6342;
												assign node6342 = (inp[6]) ? node6346 : node6343;
													assign node6343 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node6346 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node6349 = (inp[7]) ? node6353 : node6350;
													assign node6350 = (inp[6]) ? 4'b1001 : 4'b0001;
													assign node6353 = (inp[14]) ? node6357 : node6354;
														assign node6354 = (inp[2]) ? 4'b0000 : 4'b1001;
														assign node6357 = (inp[2]) ? node6361 : node6358;
															assign node6358 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node6361 = (inp[6]) ? 4'b0000 : 4'b1000;
											assign node6364 = (inp[6]) ? node6378 : node6365;
												assign node6365 = (inp[8]) ? node6373 : node6366;
													assign node6366 = (inp[14]) ? 4'b0000 : node6367;
														assign node6367 = (inp[2]) ? 4'b0000 : node6368;
															assign node6368 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node6373 = (inp[2]) ? node6375 : 4'b0001;
														assign node6375 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node6378 = (inp[14]) ? 4'b1000 : node6379;
													assign node6379 = (inp[2]) ? 4'b0001 : 4'b1001;
						assign node6383 = (inp[11]) ? node6701 : node6384;
							assign node6384 = (inp[6]) ? node6548 : node6385;
								assign node6385 = (inp[1]) ? node6459 : node6386;
									assign node6386 = (inp[2]) ? node6418 : node6387;
										assign node6387 = (inp[15]) ? node6403 : node6388;
											assign node6388 = (inp[0]) ? node6398 : node6389;
												assign node6389 = (inp[3]) ? node6393 : node6390;
													assign node6390 = (inp[5]) ? 4'b1010 : 4'b1011;
													assign node6393 = (inp[5]) ? node6395 : 4'b1011;
														assign node6395 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node6398 = (inp[3]) ? node6400 : 4'b1001;
													assign node6400 = (inp[5]) ? 4'b1011 : 4'b1001;
											assign node6403 = (inp[0]) ? node6411 : node6404;
												assign node6404 = (inp[5]) ? node6408 : node6405;
													assign node6405 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node6408 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node6411 = (inp[5]) ? node6415 : node6412;
													assign node6412 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node6415 = (inp[3]) ? 4'b1000 : 4'b1010;
										assign node6418 = (inp[5]) ? node6428 : node6419;
											assign node6419 = (inp[7]) ? node6421 : 4'b1011;
												assign node6421 = (inp[8]) ? node6423 : 4'b1011;
													assign node6423 = (inp[0]) ? 4'b1010 : node6424;
														assign node6424 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node6428 = (inp[3]) ? node6446 : node6429;
												assign node6429 = (inp[14]) ? node6437 : node6430;
													assign node6430 = (inp[8]) ? 4'b1010 : node6431;
														assign node6431 = (inp[15]) ? 4'b1000 : node6432;
															assign node6432 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node6437 = (inp[15]) ? node6441 : node6438;
														assign node6438 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node6441 = (inp[8]) ? node6443 : 4'b1010;
															assign node6443 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node6446 = (inp[8]) ? node6454 : node6447;
													assign node6447 = (inp[7]) ? node6449 : 4'b1010;
														assign node6449 = (inp[14]) ? 4'b1001 : node6450;
															assign node6450 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node6454 = (inp[0]) ? node6456 : 4'b1010;
														assign node6456 = (inp[7]) ? 4'b1000 : 4'b1001;
									assign node6459 = (inp[7]) ? node6495 : node6460;
										assign node6460 = (inp[8]) ? node6472 : node6461;
											assign node6461 = (inp[15]) ? node6465 : node6462;
												assign node6462 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node6465 = (inp[0]) ? node6469 : node6466;
													assign node6466 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node6469 = (inp[14]) ? 4'b1010 : 4'b1011;
											assign node6472 = (inp[2]) ? node6484 : node6473;
												assign node6473 = (inp[14]) ? node6481 : node6474;
													assign node6474 = (inp[15]) ? 4'b1000 : node6475;
														assign node6475 = (inp[3]) ? 4'b1000 : node6476;
															assign node6476 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node6481 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node6484 = (inp[14]) ? 4'b0001 : node6485;
													assign node6485 = (inp[5]) ? node6491 : node6486;
														assign node6486 = (inp[15]) ? node6488 : 4'b0001;
															assign node6488 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node6491 = (inp[15]) ? 4'b0001 : 4'b0011;
										assign node6495 = (inp[8]) ? node6519 : node6496;
											assign node6496 = (inp[2]) ? node6512 : node6497;
												assign node6497 = (inp[14]) ? node6505 : node6498;
													assign node6498 = (inp[0]) ? node6500 : 4'b1000;
														assign node6500 = (inp[3]) ? node6502 : 4'b1010;
															assign node6502 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node6505 = (inp[5]) ? node6507 : 4'b0011;
														assign node6507 = (inp[3]) ? 4'b0011 : node6508;
															assign node6508 = (inp[15]) ? 4'b0001 : 4'b0001;
												assign node6512 = (inp[15]) ? node6514 : 4'b0001;
													assign node6514 = (inp[3]) ? 4'b0011 : node6515;
														assign node6515 = (inp[0]) ? 4'b0011 : 4'b0001;
											assign node6519 = (inp[2]) ? node6533 : node6520;
												assign node6520 = (inp[14]) ? node6528 : node6521;
													assign node6521 = (inp[5]) ? 4'b0011 : node6522;
														assign node6522 = (inp[3]) ? node6524 : 4'b0001;
															assign node6524 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node6528 = (inp[0]) ? 4'b0010 : node6529;
														assign node6529 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node6533 = (inp[3]) ? node6541 : node6534;
													assign node6534 = (inp[15]) ? node6538 : node6535;
														assign node6535 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node6538 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node6541 = (inp[5]) ? 4'b0010 : node6542;
														assign node6542 = (inp[14]) ? 4'b0010 : node6543;
															assign node6543 = (inp[15]) ? 4'b0010 : 4'b0000;
								assign node6548 = (inp[1]) ? node6636 : node6549;
									assign node6549 = (inp[14]) ? node6591 : node6550;
										assign node6550 = (inp[5]) ? node6564 : node6551;
											assign node6551 = (inp[15]) ? node6555 : node6552;
												assign node6552 = (inp[0]) ? 4'b0001 : 4'b0010;
												assign node6555 = (inp[0]) ? node6557 : 4'b0001;
													assign node6557 = (inp[2]) ? node6559 : 4'b0011;
														assign node6559 = (inp[3]) ? node6561 : 4'b0010;
															assign node6561 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node6564 = (inp[8]) ? node6580 : node6565;
												assign node6565 = (inp[0]) ? node6573 : node6566;
													assign node6566 = (inp[3]) ? node6570 : node6567;
														assign node6567 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node6570 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node6573 = (inp[7]) ? node6577 : node6574;
														assign node6574 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node6577 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node6580 = (inp[3]) ? 4'b0000 : node6581;
													assign node6581 = (inp[0]) ? node6585 : node6582;
														assign node6582 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node6585 = (inp[7]) ? node6587 : 4'b0001;
															assign node6587 = (inp[15]) ? 4'b0010 : 4'b0000;
										assign node6591 = (inp[5]) ? node6617 : node6592;
											assign node6592 = (inp[2]) ? node6604 : node6593;
												assign node6593 = (inp[3]) ? node6595 : 4'b0010;
													assign node6595 = (inp[15]) ? node6601 : node6596;
														assign node6596 = (inp[0]) ? 4'b0000 : node6597;
															assign node6597 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node6601 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node6604 = (inp[0]) ? node6612 : node6605;
													assign node6605 = (inp[15]) ? node6607 : 4'b0010;
														assign node6607 = (inp[3]) ? node6609 : 4'b0001;
															assign node6609 = (inp[8]) ? 4'b0000 : 4'b0000;
													assign node6612 = (inp[15]) ? node6614 : 4'b0001;
														assign node6614 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node6617 = (inp[15]) ? node6625 : node6618;
												assign node6618 = (inp[2]) ? 4'b0000 : node6619;
													assign node6619 = (inp[0]) ? 4'b0011 : node6620;
														assign node6620 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node6625 = (inp[8]) ? node6629 : node6626;
													assign node6626 = (inp[3]) ? 4'b0010 : 4'b0011;
													assign node6629 = (inp[7]) ? 4'b0010 : node6630;
														assign node6630 = (inp[0]) ? 4'b0011 : node6631;
															assign node6631 = (inp[3]) ? 4'b0011 : 4'b0001;
									assign node6636 = (inp[8]) ? node6672 : node6637;
										assign node6637 = (inp[7]) ? node6659 : node6638;
											assign node6638 = (inp[14]) ? node6650 : node6639;
												assign node6639 = (inp[2]) ? node6647 : node6640;
													assign node6640 = (inp[0]) ? node6642 : 4'b0011;
														assign node6642 = (inp[5]) ? node6644 : 4'b0011;
															assign node6644 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node6647 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node6650 = (inp[15]) ? 4'b0010 : node6651;
													assign node6651 = (inp[0]) ? 4'b0000 : node6652;
														assign node6652 = (inp[3]) ? node6654 : 4'b0010;
															assign node6654 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node6659 = (inp[14]) ? node6667 : node6660;
												assign node6660 = (inp[2]) ? 4'b1111 : node6661;
													assign node6661 = (inp[3]) ? 4'b0010 : node6662;
														assign node6662 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node6667 = (inp[15]) ? 4'b1111 : node6668;
													assign node6668 = (inp[3]) ? 4'b1111 : 4'b1101;
										assign node6672 = (inp[7]) ? node6688 : node6673;
											assign node6673 = (inp[2]) ? node6679 : node6674;
												assign node6674 = (inp[14]) ? 4'b1111 : node6675;
													assign node6675 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node6679 = (inp[0]) ? node6681 : 4'b1111;
													assign node6681 = (inp[14]) ? node6683 : 4'b1101;
														assign node6683 = (inp[3]) ? node6685 : 4'b1111;
															assign node6685 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node6688 = (inp[2]) ? node6694 : node6689;
												assign node6689 = (inp[14]) ? node6691 : 4'b1101;
													assign node6691 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node6694 = (inp[3]) ? node6696 : 4'b1100;
													assign node6696 = (inp[15]) ? node6698 : 4'b1100;
														assign node6698 = (inp[0]) ? 4'b1100 : 4'b1110;
							assign node6701 = (inp[6]) ? node6871 : node6702;
								assign node6702 = (inp[1]) ? node6776 : node6703;
									assign node6703 = (inp[15]) ? node6735 : node6704;
										assign node6704 = (inp[0]) ? node6712 : node6705;
											assign node6705 = (inp[5]) ? node6707 : 4'b0010;
												assign node6707 = (inp[3]) ? node6709 : 4'b0011;
													assign node6709 = (inp[14]) ? 4'b0001 : 4'b0000;
											assign node6712 = (inp[5]) ? node6726 : node6713;
												assign node6713 = (inp[2]) ? node6715 : 4'b0000;
													assign node6715 = (inp[3]) ? node6721 : node6716;
														assign node6716 = (inp[8]) ? 4'b0000 : node6717;
															assign node6717 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node6721 = (inp[7]) ? 4'b0001 : node6722;
															assign node6722 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node6726 = (inp[3]) ? node6728 : 4'b0000;
													assign node6728 = (inp[8]) ? node6730 : 4'b0010;
														assign node6730 = (inp[2]) ? 4'b0010 : node6731;
															assign node6731 = (inp[7]) ? 4'b0011 : 4'b0010;
										assign node6735 = (inp[0]) ? node6765 : node6736;
											assign node6736 = (inp[5]) ? node6750 : node6737;
												assign node6737 = (inp[2]) ? node6743 : node6738;
													assign node6738 = (inp[3]) ? 4'b0001 : node6739;
														assign node6739 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node6743 = (inp[3]) ? 4'b0000 : node6744;
														assign node6744 = (inp[7]) ? 4'b0001 : node6745;
															assign node6745 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node6750 = (inp[3]) ? node6758 : node6751;
													assign node6751 = (inp[2]) ? 4'b0000 : node6752;
														assign node6752 = (inp[7]) ? 4'b0001 : node6753;
															assign node6753 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node6758 = (inp[8]) ? node6760 : 4'b0011;
														assign node6760 = (inp[7]) ? 4'b0010 : node6761;
															assign node6761 = (inp[14]) ? 4'b0011 : 4'b0010;
											assign node6765 = (inp[5]) ? node6771 : node6766;
												assign node6766 = (inp[7]) ? node6768 : 4'b0011;
													assign node6768 = (inp[14]) ? 4'b0011 : 4'b0010;
												assign node6771 = (inp[3]) ? 4'b0000 : node6772;
													assign node6772 = (inp[14]) ? 4'b0010 : 4'b0011;
									assign node6776 = (inp[8]) ? node6820 : node6777;
										assign node6777 = (inp[7]) ? node6799 : node6778;
											assign node6778 = (inp[14]) ? node6788 : node6779;
												assign node6779 = (inp[2]) ? node6785 : node6780;
													assign node6780 = (inp[5]) ? 4'b0011 : node6781;
														assign node6781 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node6785 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node6788 = (inp[0]) ? node6792 : node6789;
													assign node6789 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node6792 = (inp[3]) ? node6794 : 4'b0010;
														assign node6794 = (inp[5]) ? node6796 : 4'b0010;
															assign node6796 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node6799 = (inp[2]) ? node6811 : node6800;
												assign node6800 = (inp[14]) ? node6804 : node6801;
													assign node6801 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node6804 = (inp[15]) ? 4'b1101 : node6805;
														assign node6805 = (inp[0]) ? node6807 : 4'b1111;
															assign node6807 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node6811 = (inp[3]) ? node6817 : node6812;
													assign node6812 = (inp[5]) ? 4'b1101 : node6813;
														assign node6813 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node6817 = (inp[5]) ? 4'b1111 : 4'b1101;
										assign node6820 = (inp[7]) ? node6844 : node6821;
											assign node6821 = (inp[2]) ? node6835 : node6822;
												assign node6822 = (inp[14]) ? node6828 : node6823;
													assign node6823 = (inp[5]) ? node6825 : 4'b0000;
														assign node6825 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node6828 = (inp[15]) ? 4'b1101 : node6829;
														assign node6829 = (inp[3]) ? 4'b1111 : node6830;
															assign node6830 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node6835 = (inp[3]) ? node6837 : 4'b1111;
													assign node6837 = (inp[5]) ? 4'b1101 : node6838;
														assign node6838 = (inp[15]) ? 4'b1111 : node6839;
															assign node6839 = (inp[0]) ? 4'b1111 : 4'b1101;
											assign node6844 = (inp[14]) ? node6854 : node6845;
												assign node6845 = (inp[2]) ? 4'b1110 : node6846;
													assign node6846 = (inp[3]) ? node6848 : 4'b1101;
														assign node6848 = (inp[5]) ? 4'b1111 : node6849;
															assign node6849 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node6854 = (inp[15]) ? node6860 : node6855;
													assign node6855 = (inp[0]) ? 4'b1110 : node6856;
														assign node6856 = (inp[2]) ? 4'b1110 : 4'b1100;
													assign node6860 = (inp[2]) ? node6866 : node6861;
														assign node6861 = (inp[5]) ? node6863 : 4'b1110;
															assign node6863 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node6866 = (inp[0]) ? 4'b1100 : node6867;
															assign node6867 = (inp[5]) ? 4'b1110 : 4'b1100;
								assign node6871 = (inp[1]) ? node6963 : node6872;
									assign node6872 = (inp[3]) ? node6912 : node6873;
										assign node6873 = (inp[14]) ? node6891 : node6874;
											assign node6874 = (inp[5]) ? node6886 : node6875;
												assign node6875 = (inp[8]) ? node6881 : node6876;
													assign node6876 = (inp[7]) ? node6878 : 4'b1110;
														assign node6878 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node6881 = (inp[2]) ? node6883 : 4'b1100;
														assign node6883 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node6886 = (inp[8]) ? node6888 : 4'b1100;
													assign node6888 = (inp[2]) ? 4'b1110 : 4'b1100;
											assign node6891 = (inp[2]) ? node6901 : node6892;
												assign node6892 = (inp[5]) ? node6896 : node6893;
													assign node6893 = (inp[8]) ? 4'b1100 : 4'b1111;
													assign node6896 = (inp[0]) ? 4'b1111 : node6897;
														assign node6897 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node6901 = (inp[5]) ? 4'b1100 : node6902;
													assign node6902 = (inp[15]) ? node6906 : node6903;
														assign node6903 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node6906 = (inp[0]) ? 4'b1111 : node6907;
															assign node6907 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node6912 = (inp[5]) ? node6946 : node6913;
											assign node6913 = (inp[2]) ? node6929 : node6914;
												assign node6914 = (inp[8]) ? node6916 : 4'b1101;
													assign node6916 = (inp[7]) ? node6922 : node6917;
														assign node6917 = (inp[0]) ? 4'b1101 : node6918;
															assign node6918 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node6922 = (inp[0]) ? node6926 : node6923;
															assign node6923 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node6926 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node6929 = (inp[0]) ? node6937 : node6930;
													assign node6930 = (inp[15]) ? 4'b1111 : node6931;
														assign node6931 = (inp[8]) ? 4'b1101 : node6932;
															assign node6932 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node6937 = (inp[15]) ? node6943 : node6938;
														assign node6938 = (inp[14]) ? 4'b1110 : node6939;
															assign node6939 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node6943 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node6946 = (inp[0]) ? node6954 : node6947;
												assign node6947 = (inp[15]) ? node6951 : node6948;
													assign node6948 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node6951 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node6954 = (inp[15]) ? 4'b1101 : node6955;
													assign node6955 = (inp[8]) ? 4'b1111 : node6956;
														assign node6956 = (inp[14]) ? 4'b1111 : node6957;
															assign node6957 = (inp[7]) ? 4'b1110 : 4'b1111;
									assign node6963 = (inp[7]) ? node7015 : node6964;
										assign node6964 = (inp[8]) ? node6982 : node6965;
											assign node6965 = (inp[15]) ? node6979 : node6966;
												assign node6966 = (inp[2]) ? node6970 : node6967;
													assign node6967 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node6970 = (inp[14]) ? node6976 : node6971;
														assign node6971 = (inp[0]) ? node6973 : 4'b1100;
															assign node6973 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node6976 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node6979 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node6982 = (inp[2]) ? node7004 : node6983;
												assign node6983 = (inp[14]) ? node6997 : node6984;
													assign node6984 = (inp[0]) ? node6990 : node6985;
														assign node6985 = (inp[15]) ? 4'b1110 : node6986;
															assign node6986 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node6990 = (inp[5]) ? node6994 : node6991;
															assign node6991 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node6994 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node6997 = (inp[0]) ? 4'b0101 : node6998;
														assign node6998 = (inp[3]) ? node7000 : 4'b0101;
															assign node7000 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node7004 = (inp[0]) ? node7010 : node7005;
													assign node7005 = (inp[15]) ? node7007 : 4'b0101;
														assign node7007 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node7010 = (inp[15]) ? node7012 : 4'b0111;
														assign node7012 = (inp[3]) ? 4'b0101 : 4'b0111;
										assign node7015 = (inp[8]) ? node7029 : node7016;
											assign node7016 = (inp[14]) ? node7020 : node7017;
												assign node7017 = (inp[2]) ? 4'b0101 : 4'b1100;
												assign node7020 = (inp[3]) ? node7022 : 4'b0101;
													assign node7022 = (inp[0]) ? node7026 : node7023;
														assign node7023 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node7026 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node7029 = (inp[14]) ? node7043 : node7030;
												assign node7030 = (inp[2]) ? node7038 : node7031;
													assign node7031 = (inp[3]) ? 4'b0101 : node7032;
														assign node7032 = (inp[5]) ? node7034 : 4'b0111;
															assign node7034 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node7038 = (inp[5]) ? node7040 : 4'b0100;
														assign node7040 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node7043 = (inp[5]) ? node7047 : node7044;
													assign node7044 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node7047 = (inp[15]) ? 4'b0110 : node7048;
														assign node7048 = (inp[0]) ? 4'b0110 : 4'b0100;
					assign node7052 = (inp[12]) ? node7694 : node7053;
						assign node7053 = (inp[11]) ? node7375 : node7054;
							assign node7054 = (inp[6]) ? node7210 : node7055;
								assign node7055 = (inp[1]) ? node7133 : node7056;
									assign node7056 = (inp[2]) ? node7090 : node7057;
										assign node7057 = (inp[14]) ? node7075 : node7058;
											assign node7058 = (inp[3]) ? node7068 : node7059;
												assign node7059 = (inp[8]) ? node7065 : node7060;
													assign node7060 = (inp[15]) ? node7062 : 4'b1001;
														assign node7062 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node7065 = (inp[5]) ? 4'b1000 : 4'b1001;
												assign node7068 = (inp[0]) ? 4'b1011 : node7069;
													assign node7069 = (inp[5]) ? 4'b1001 : node7070;
														assign node7070 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node7075 = (inp[0]) ? node7083 : node7076;
												assign node7076 = (inp[8]) ? node7080 : node7077;
													assign node7077 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node7080 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node7083 = (inp[7]) ? node7087 : node7084;
													assign node7084 = (inp[3]) ? 4'b1001 : 4'b1000;
													assign node7087 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node7090 = (inp[0]) ? node7114 : node7091;
											assign node7091 = (inp[15]) ? node7101 : node7092;
												assign node7092 = (inp[3]) ? node7098 : node7093;
													assign node7093 = (inp[8]) ? node7095 : 4'b1010;
														assign node7095 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node7098 = (inp[8]) ? 4'b1010 : 4'b1000;
												assign node7101 = (inp[3]) ? node7105 : node7102;
													assign node7102 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node7105 = (inp[5]) ? node7107 : 4'b1001;
														assign node7107 = (inp[8]) ? node7111 : node7108;
															assign node7108 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node7111 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node7114 = (inp[14]) ? node7126 : node7115;
												assign node7115 = (inp[8]) ? node7123 : node7116;
													assign node7116 = (inp[7]) ? 4'b1001 : node7117;
														assign node7117 = (inp[3]) ? node7119 : 4'b1010;
															assign node7119 = (inp[5]) ? 4'b1000 : 4'b1000;
													assign node7123 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node7126 = (inp[15]) ? node7128 : 4'b1001;
													assign node7128 = (inp[8]) ? node7130 : 4'b1001;
														assign node7130 = (inp[7]) ? 4'b1010 : 4'b1011;
									assign node7133 = (inp[8]) ? node7177 : node7134;
										assign node7134 = (inp[7]) ? node7156 : node7135;
											assign node7135 = (inp[15]) ? node7141 : node7136;
												assign node7136 = (inp[5]) ? node7138 : 4'b1010;
													assign node7138 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node7141 = (inp[14]) ? node7151 : node7142;
													assign node7142 = (inp[2]) ? node7148 : node7143;
														assign node7143 = (inp[3]) ? node7145 : 4'b1001;
															assign node7145 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node7148 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node7151 = (inp[3]) ? 4'b1000 : node7152;
														assign node7152 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node7156 = (inp[2]) ? node7166 : node7157;
												assign node7157 = (inp[14]) ? node7159 : 4'b1010;
													assign node7159 = (inp[0]) ? 4'b0011 : node7160;
														assign node7160 = (inp[15]) ? node7162 : 4'b0011;
															assign node7162 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node7166 = (inp[14]) ? node7172 : node7167;
													assign node7167 = (inp[3]) ? 4'b0001 : node7168;
														assign node7168 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node7172 = (inp[15]) ? 4'b0001 : node7173;
														assign node7173 = (inp[3]) ? 4'b0011 : 4'b0001;
										assign node7177 = (inp[7]) ? node7189 : node7178;
											assign node7178 = (inp[0]) ? node7184 : node7179;
												assign node7179 = (inp[15]) ? node7181 : 4'b0011;
													assign node7181 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node7184 = (inp[2]) ? node7186 : 4'b1000;
													assign node7186 = (inp[15]) ? 4'b0011 : 4'b0001;
											assign node7189 = (inp[2]) ? node7201 : node7190;
												assign node7190 = (inp[14]) ? node7198 : node7191;
													assign node7191 = (inp[0]) ? node7193 : 4'b0011;
														assign node7193 = (inp[15]) ? node7195 : 4'b0001;
															assign node7195 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node7198 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node7201 = (inp[0]) ? node7203 : 4'b0000;
													assign node7203 = (inp[5]) ? node7205 : 4'b0010;
														assign node7205 = (inp[14]) ? node7207 : 4'b0000;
															assign node7207 = (inp[3]) ? 4'b0010 : 4'b0000;
								assign node7210 = (inp[1]) ? node7292 : node7211;
									assign node7211 = (inp[7]) ? node7241 : node7212;
										assign node7212 = (inp[15]) ? node7230 : node7213;
											assign node7213 = (inp[5]) ? node7223 : node7214;
												assign node7214 = (inp[0]) ? node7220 : node7215;
													assign node7215 = (inp[14]) ? 4'b0010 : node7216;
														assign node7216 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node7220 = (inp[3]) ? 4'b0001 : 4'b0000;
												assign node7223 = (inp[14]) ? node7227 : node7224;
													assign node7224 = (inp[0]) ? 4'b0010 : 4'b0001;
													assign node7227 = (inp[2]) ? 4'b0011 : 4'b0001;
											assign node7230 = (inp[8]) ? node7234 : node7231;
												assign node7231 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node7234 = (inp[0]) ? 4'b0011 : node7235;
													assign node7235 = (inp[3]) ? node7237 : 4'b0001;
														assign node7237 = (inp[5]) ? 4'b0011 : 4'b0001;
										assign node7241 = (inp[8]) ? node7265 : node7242;
											assign node7242 = (inp[2]) ? node7254 : node7243;
												assign node7243 = (inp[14]) ? node7251 : node7244;
													assign node7244 = (inp[3]) ? node7246 : 4'b0010;
														assign node7246 = (inp[15]) ? node7248 : 4'b0000;
															assign node7248 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node7251 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node7254 = (inp[5]) ? node7260 : node7255;
													assign node7255 = (inp[14]) ? node7257 : 4'b0011;
														assign node7257 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node7260 = (inp[14]) ? node7262 : 4'b0001;
														assign node7262 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node7265 = (inp[2]) ? node7275 : node7266;
												assign node7266 = (inp[14]) ? 4'b0010 : node7267;
													assign node7267 = (inp[15]) ? 4'b0011 : node7268;
														assign node7268 = (inp[0]) ? 4'b0001 : node7269;
															assign node7269 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node7275 = (inp[3]) ? node7283 : node7276;
													assign node7276 = (inp[14]) ? 4'b0010 : node7277;
														assign node7277 = (inp[0]) ? 4'b0000 : node7278;
															assign node7278 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node7283 = (inp[15]) ? 4'b0010 : node7284;
														assign node7284 = (inp[14]) ? node7288 : node7285;
															assign node7285 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node7288 = (inp[0]) ? 4'b0000 : 4'b0010;
									assign node7292 = (inp[7]) ? node7330 : node7293;
										assign node7293 = (inp[8]) ? node7309 : node7294;
											assign node7294 = (inp[15]) ? node7302 : node7295;
												assign node7295 = (inp[0]) ? 4'b0000 : node7296;
													assign node7296 = (inp[2]) ? 4'b0010 : node7297;
														assign node7297 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node7302 = (inp[0]) ? 4'b0011 : node7303;
													assign node7303 = (inp[14]) ? 4'b0000 : node7304;
														assign node7304 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node7309 = (inp[0]) ? node7317 : node7310;
												assign node7310 = (inp[15]) ? 4'b1111 : node7311;
													assign node7311 = (inp[5]) ? 4'b1101 : node7312;
														assign node7312 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node7317 = (inp[14]) ? node7323 : node7318;
													assign node7318 = (inp[3]) ? 4'b0000 : node7319;
														assign node7319 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node7323 = (inp[2]) ? 4'b1101 : node7324;
														assign node7324 = (inp[15]) ? 4'b1111 : node7325;
															assign node7325 = (inp[3]) ? 4'b1111 : 4'b1101;
										assign node7330 = (inp[8]) ? node7352 : node7331;
											assign node7331 = (inp[14]) ? node7341 : node7332;
												assign node7332 = (inp[2]) ? node7334 : 4'b0010;
													assign node7334 = (inp[5]) ? 4'b1111 : node7335;
														assign node7335 = (inp[3]) ? 4'b1101 : node7336;
															assign node7336 = (inp[15]) ? 4'b1101 : 4'b1101;
												assign node7341 = (inp[15]) ? node7345 : node7342;
													assign node7342 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node7345 = (inp[0]) ? node7347 : 4'b1111;
														assign node7347 = (inp[3]) ? 4'b1101 : node7348;
															assign node7348 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node7352 = (inp[2]) ? node7364 : node7353;
												assign node7353 = (inp[14]) ? node7359 : node7354;
													assign node7354 = (inp[5]) ? 4'b1101 : node7355;
														assign node7355 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node7359 = (inp[0]) ? node7361 : 4'b1100;
														assign node7361 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node7364 = (inp[3]) ? 4'b1100 : node7365;
													assign node7365 = (inp[0]) ? node7367 : 4'b1110;
														assign node7367 = (inp[14]) ? node7371 : node7368;
															assign node7368 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node7371 = (inp[5]) ? 4'b1110 : 4'b1100;
							assign node7375 = (inp[6]) ? node7529 : node7376;
								assign node7376 = (inp[1]) ? node7446 : node7377;
									assign node7377 = (inp[7]) ? node7419 : node7378;
										assign node7378 = (inp[8]) ? node7392 : node7379;
											assign node7379 = (inp[2]) ? node7389 : node7380;
												assign node7380 = (inp[14]) ? 4'b0000 : node7381;
													assign node7381 = (inp[15]) ? node7383 : 4'b0001;
														assign node7383 = (inp[3]) ? node7385 : 4'b0011;
															assign node7385 = (inp[0]) ? 4'b0001 : 4'b0001;
												assign node7389 = (inp[14]) ? 4'b0000 : 4'b0010;
											assign node7392 = (inp[2]) ? node7406 : node7393;
												assign node7393 = (inp[14]) ? node7399 : node7394;
													assign node7394 = (inp[3]) ? node7396 : 4'b0010;
														assign node7396 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node7399 = (inp[0]) ? 4'b0001 : node7400;
														assign node7400 = (inp[5]) ? 4'b0011 : node7401;
															assign node7401 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node7406 = (inp[0]) ? node7412 : node7407;
													assign node7407 = (inp[15]) ? node7409 : 4'b0011;
														assign node7409 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node7412 = (inp[14]) ? node7414 : 4'b0011;
														assign node7414 = (inp[5]) ? 4'b0001 : node7415;
															assign node7415 = (inp[3]) ? 4'b0011 : 4'b0001;
										assign node7419 = (inp[8]) ? node7431 : node7420;
											assign node7420 = (inp[14]) ? node7428 : node7421;
												assign node7421 = (inp[2]) ? node7425 : node7422;
													assign node7422 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node7425 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node7428 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node7431 = (inp[2]) ? node7441 : node7432;
												assign node7432 = (inp[14]) ? node7436 : node7433;
													assign node7433 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node7436 = (inp[3]) ? node7438 : 4'b0010;
														assign node7438 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node7441 = (inp[5]) ? 4'b0000 : node7442;
													assign node7442 = (inp[15]) ? 4'b0010 : 4'b0000;
									assign node7446 = (inp[8]) ? node7484 : node7447;
										assign node7447 = (inp[7]) ? node7465 : node7448;
											assign node7448 = (inp[2]) ? node7456 : node7449;
												assign node7449 = (inp[15]) ? node7453 : node7450;
													assign node7450 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node7453 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node7456 = (inp[3]) ? node7458 : 4'b0010;
													assign node7458 = (inp[0]) ? node7460 : 4'b0000;
														assign node7460 = (inp[5]) ? 4'b0010 : node7461;
															assign node7461 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node7465 = (inp[14]) ? node7477 : node7466;
												assign node7466 = (inp[0]) ? node7468 : 4'b1111;
													assign node7468 = (inp[5]) ? node7472 : node7469;
														assign node7469 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node7472 = (inp[15]) ? node7474 : 4'b0010;
															assign node7474 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node7477 = (inp[3]) ? node7479 : 4'b1111;
													assign node7479 = (inp[15]) ? node7481 : 4'b1101;
														assign node7481 = (inp[0]) ? 4'b1101 : 4'b1111;
										assign node7484 = (inp[7]) ? node7502 : node7485;
											assign node7485 = (inp[14]) ? node7493 : node7486;
												assign node7486 = (inp[2]) ? node7490 : node7487;
													assign node7487 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node7490 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node7493 = (inp[0]) ? node7497 : node7494;
													assign node7494 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node7497 = (inp[15]) ? 4'b1101 : node7498;
														assign node7498 = (inp[2]) ? 4'b1101 : 4'b1111;
											assign node7502 = (inp[14]) ? node7516 : node7503;
												assign node7503 = (inp[2]) ? node7509 : node7504;
													assign node7504 = (inp[15]) ? 4'b1101 : node7505;
														assign node7505 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node7509 = (inp[15]) ? node7511 : 4'b1100;
														assign node7511 = (inp[3]) ? 4'b1110 : node7512;
															assign node7512 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node7516 = (inp[2]) ? node7524 : node7517;
													assign node7517 = (inp[0]) ? 4'b1100 : node7518;
														assign node7518 = (inp[15]) ? 4'b1110 : node7519;
															assign node7519 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node7524 = (inp[15]) ? 4'b1110 : node7525;
														assign node7525 = (inp[0]) ? 4'b1110 : 4'b1100;
								assign node7529 = (inp[1]) ? node7611 : node7530;
									assign node7530 = (inp[15]) ? node7574 : node7531;
										assign node7531 = (inp[0]) ? node7555 : node7532;
											assign node7532 = (inp[5]) ? node7542 : node7533;
												assign node7533 = (inp[3]) ? node7539 : node7534;
													assign node7534 = (inp[7]) ? node7536 : 4'b1110;
														assign node7536 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node7539 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node7542 = (inp[8]) ? node7548 : node7543;
													assign node7543 = (inp[3]) ? 4'b1101 : node7544;
														assign node7544 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node7548 = (inp[14]) ? 4'b1100 : node7549;
														assign node7549 = (inp[3]) ? 4'b1100 : node7550;
															assign node7550 = (inp[7]) ? 4'b1101 : 4'b1100;
											assign node7555 = (inp[3]) ? node7565 : node7556;
												assign node7556 = (inp[5]) ? 4'b1111 : node7557;
													assign node7557 = (inp[14]) ? 4'b1101 : node7558;
														assign node7558 = (inp[2]) ? node7560 : 4'b1100;
															assign node7560 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node7565 = (inp[14]) ? 4'b1111 : node7566;
													assign node7566 = (inp[8]) ? node7568 : 4'b1110;
														assign node7568 = (inp[2]) ? node7570 : 4'b1111;
															assign node7570 = (inp[7]) ? 4'b1110 : 4'b1111;
										assign node7574 = (inp[2]) ? node7596 : node7575;
											assign node7575 = (inp[8]) ? node7587 : node7576;
												assign node7576 = (inp[0]) ? node7578 : 4'b1111;
													assign node7578 = (inp[3]) ? node7584 : node7579;
														assign node7579 = (inp[7]) ? 4'b1110 : node7580;
															assign node7580 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node7584 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node7587 = (inp[5]) ? 4'b1101 : node7588;
													assign node7588 = (inp[3]) ? 4'b1100 : node7589;
														assign node7589 = (inp[0]) ? 4'b1111 : node7590;
															assign node7590 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node7596 = (inp[7]) ? node7598 : 4'b1100;
												assign node7598 = (inp[8]) ? node7602 : node7599;
													assign node7599 = (inp[14]) ? 4'b1111 : 4'b1101;
													assign node7602 = (inp[3]) ? 4'b1100 : node7603;
														assign node7603 = (inp[14]) ? node7607 : node7604;
															assign node7604 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node7607 = (inp[5]) ? 4'b1100 : 4'b1110;
									assign node7611 = (inp[7]) ? node7653 : node7612;
										assign node7612 = (inp[8]) ? node7632 : node7613;
											assign node7613 = (inp[14]) ? node7623 : node7614;
												assign node7614 = (inp[2]) ? node7618 : node7615;
													assign node7615 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node7618 = (inp[0]) ? 4'b1110 : node7619;
														assign node7619 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node7623 = (inp[5]) ? 4'b1100 : node7624;
													assign node7624 = (inp[2]) ? 4'b1110 : node7625;
														assign node7625 = (inp[0]) ? node7627 : 4'b1100;
															assign node7627 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node7632 = (inp[14]) ? node7640 : node7633;
												assign node7633 = (inp[2]) ? 4'b0101 : node7634;
													assign node7634 = (inp[3]) ? node7636 : 4'b1100;
														assign node7636 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node7640 = (inp[5]) ? node7646 : node7641;
													assign node7641 = (inp[15]) ? node7643 : 4'b0111;
														assign node7643 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node7646 = (inp[3]) ? 4'b0101 : node7647;
														assign node7647 = (inp[0]) ? 4'b0111 : node7648;
															assign node7648 = (inp[15]) ? 4'b0111 : 4'b0101;
										assign node7653 = (inp[8]) ? node7675 : node7654;
											assign node7654 = (inp[14]) ? node7662 : node7655;
												assign node7655 = (inp[2]) ? node7659 : node7656;
													assign node7656 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node7659 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node7662 = (inp[5]) ? node7668 : node7663;
													assign node7663 = (inp[15]) ? 4'b0101 : node7664;
														assign node7664 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node7668 = (inp[3]) ? 4'b0111 : node7669;
														assign node7669 = (inp[15]) ? node7671 : 4'b0101;
															assign node7671 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node7675 = (inp[14]) ? node7689 : node7676;
												assign node7676 = (inp[2]) ? node7678 : 4'b0101;
													assign node7678 = (inp[15]) ? node7684 : node7679;
														assign node7679 = (inp[0]) ? 4'b0110 : node7680;
															assign node7680 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node7684 = (inp[5]) ? node7686 : 4'b0100;
															assign node7686 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node7689 = (inp[3]) ? node7691 : 4'b0110;
													assign node7691 = (inp[2]) ? 4'b0100 : 4'b0110;
						assign node7694 = (inp[7]) ? node8020 : node7695;
							assign node7695 = (inp[8]) ? node7847 : node7696;
								assign node7696 = (inp[14]) ? node7780 : node7697;
									assign node7697 = (inp[2]) ? node7733 : node7698;
										assign node7698 = (inp[15]) ? node7714 : node7699;
											assign node7699 = (inp[5]) ? node7709 : node7700;
												assign node7700 = (inp[0]) ? node7704 : node7701;
													assign node7701 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node7704 = (inp[6]) ? 4'b0111 : node7705;
														assign node7705 = (inp[1]) ? 4'b1101 : 4'b0101;
												assign node7709 = (inp[11]) ? node7711 : 4'b0101;
													assign node7711 = (inp[6]) ? 4'b1101 : 4'b0101;
											assign node7714 = (inp[0]) ? node7726 : node7715;
												assign node7715 = (inp[1]) ? node7721 : node7716;
													assign node7716 = (inp[11]) ? node7718 : 4'b0111;
														assign node7718 = (inp[6]) ? 4'b1111 : 4'b0111;
													assign node7721 = (inp[3]) ? 4'b1111 : node7722;
														assign node7722 = (inp[6]) ? 4'b1111 : 4'b0111;
												assign node7726 = (inp[3]) ? node7730 : node7727;
													assign node7727 = (inp[6]) ? 4'b1111 : 4'b0111;
													assign node7730 = (inp[1]) ? 4'b1101 : 4'b0101;
										assign node7733 = (inp[15]) ? node7753 : node7734;
											assign node7734 = (inp[0]) ? node7742 : node7735;
												assign node7735 = (inp[5]) ? 4'b1100 : node7736;
													assign node7736 = (inp[11]) ? 4'b0100 : node7737;
														assign node7737 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node7742 = (inp[1]) ? node7746 : node7743;
													assign node7743 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node7746 = (inp[11]) ? node7750 : node7747;
														assign node7747 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node7750 = (inp[6]) ? 4'b1110 : 4'b0110;
											assign node7753 = (inp[0]) ? node7761 : node7754;
												assign node7754 = (inp[3]) ? 4'b1110 : node7755;
													assign node7755 = (inp[11]) ? node7757 : 4'b0110;
														assign node7757 = (inp[6]) ? 4'b1110 : 4'b0110;
												assign node7761 = (inp[3]) ? node7767 : node7762;
													assign node7762 = (inp[5]) ? node7764 : 4'b0110;
														assign node7764 = (inp[6]) ? 4'b1100 : 4'b0100;
													assign node7767 = (inp[1]) ? node7773 : node7768;
														assign node7768 = (inp[6]) ? node7770 : 4'b1100;
															assign node7770 = (inp[5]) ? 4'b1100 : 4'b0100;
														assign node7773 = (inp[6]) ? node7777 : node7774;
															assign node7774 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node7777 = (inp[11]) ? 4'b1100 : 4'b0100;
									assign node7780 = (inp[6]) ? node7812 : node7781;
										assign node7781 = (inp[11]) ? node7793 : node7782;
											assign node7782 = (inp[0]) ? node7788 : node7783;
												assign node7783 = (inp[15]) ? node7785 : 4'b1100;
													assign node7785 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node7788 = (inp[15]) ? node7790 : 4'b1110;
													assign node7790 = (inp[1]) ? 4'b1110 : 4'b1100;
											assign node7793 = (inp[5]) ? node7807 : node7794;
												assign node7794 = (inp[15]) ? node7800 : node7795;
													assign node7795 = (inp[3]) ? node7797 : 4'b0110;
														assign node7797 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node7800 = (inp[1]) ? node7802 : 4'b0100;
														assign node7802 = (inp[0]) ? 4'b0110 : node7803;
															assign node7803 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node7807 = (inp[15]) ? 4'b0100 : node7808;
													assign node7808 = (inp[0]) ? 4'b0110 : 4'b0100;
										assign node7812 = (inp[11]) ? node7834 : node7813;
											assign node7813 = (inp[1]) ? node7829 : node7814;
												assign node7814 = (inp[3]) ? node7822 : node7815;
													assign node7815 = (inp[5]) ? 4'b0110 : node7816;
														assign node7816 = (inp[2]) ? node7818 : 4'b0110;
															assign node7818 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node7822 = (inp[0]) ? node7826 : node7823;
														assign node7823 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node7826 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node7829 = (inp[0]) ? 4'b0110 : node7830;
													assign node7830 = (inp[15]) ? 4'b0110 : 4'b0100;
											assign node7834 = (inp[5]) ? node7842 : node7835;
												assign node7835 = (inp[0]) ? node7837 : 4'b1100;
													assign node7837 = (inp[2]) ? node7839 : 4'b1100;
														assign node7839 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node7842 = (inp[3]) ? node7844 : 4'b1110;
													assign node7844 = (inp[0]) ? 4'b1110 : 4'b1100;
								assign node7847 = (inp[2]) ? node7921 : node7848;
									assign node7848 = (inp[14]) ? node7882 : node7849;
										assign node7849 = (inp[11]) ? node7867 : node7850;
											assign node7850 = (inp[6]) ? node7860 : node7851;
												assign node7851 = (inp[0]) ? 4'b1110 : node7852;
													assign node7852 = (inp[1]) ? 4'b1100 : node7853;
														assign node7853 = (inp[5]) ? 4'b1100 : node7854;
															assign node7854 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node7860 = (inp[0]) ? node7862 : 4'b0100;
													assign node7862 = (inp[3]) ? 4'b0110 : node7863;
														assign node7863 = (inp[1]) ? 4'b0110 : 4'b0100;
											assign node7867 = (inp[6]) ? node7869 : 4'b0110;
												assign node7869 = (inp[0]) ? node7875 : node7870;
													assign node7870 = (inp[15]) ? 4'b1110 : node7871;
														assign node7871 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node7875 = (inp[15]) ? node7879 : node7876;
														assign node7876 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node7879 = (inp[5]) ? 4'b1100 : 4'b1110;
										assign node7882 = (inp[5]) ? node7906 : node7883;
											assign node7883 = (inp[3]) ? node7895 : node7884;
												assign node7884 = (inp[15]) ? node7890 : node7885;
													assign node7885 = (inp[11]) ? node7887 : 4'b0111;
														assign node7887 = (inp[6]) ? 4'b1111 : 4'b0111;
													assign node7890 = (inp[0]) ? 4'b1111 : node7891;
														assign node7891 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node7895 = (inp[6]) ? node7903 : node7896;
													assign node7896 = (inp[0]) ? node7900 : node7897;
														assign node7897 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node7900 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node7903 = (inp[0]) ? 4'b0101 : 4'b1101;
											assign node7906 = (inp[6]) ? node7910 : node7907;
												assign node7907 = (inp[11]) ? 4'b1101 : 4'b0101;
												assign node7910 = (inp[3]) ? node7918 : node7911;
													assign node7911 = (inp[15]) ? 4'b0111 : node7912;
														assign node7912 = (inp[1]) ? 4'b0101 : node7913;
															assign node7913 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node7918 = (inp[1]) ? 4'b1101 : 4'b0111;
									assign node7921 = (inp[1]) ? node7967 : node7922;
										assign node7922 = (inp[0]) ? node7942 : node7923;
											assign node7923 = (inp[15]) ? node7935 : node7924;
												assign node7924 = (inp[5]) ? node7932 : node7925;
													assign node7925 = (inp[3]) ? 4'b1101 : node7926;
														assign node7926 = (inp[11]) ? node7928 : 4'b0111;
															assign node7928 = (inp[6]) ? 4'b1111 : 4'b0111;
													assign node7932 = (inp[3]) ? 4'b0101 : 4'b1101;
												assign node7935 = (inp[3]) ? node7937 : 4'b0111;
													assign node7937 = (inp[6]) ? node7939 : 4'b1111;
														assign node7939 = (inp[11]) ? 4'b1111 : 4'b0111;
											assign node7942 = (inp[15]) ? node7958 : node7943;
												assign node7943 = (inp[3]) ? node7953 : node7944;
													assign node7944 = (inp[5]) ? node7948 : node7945;
														assign node7945 = (inp[6]) ? 4'b1101 : 4'b0101;
														assign node7948 = (inp[6]) ? 4'b1111 : node7949;
															assign node7949 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node7953 = (inp[6]) ? 4'b0111 : node7954;
														assign node7954 = (inp[14]) ? 4'b0111 : 4'b1111;
												assign node7958 = (inp[3]) ? node7962 : node7959;
													assign node7959 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node7962 = (inp[6]) ? node7964 : 4'b1101;
														assign node7964 = (inp[11]) ? 4'b1101 : 4'b0101;
										assign node7967 = (inp[0]) ? node7999 : node7968;
											assign node7968 = (inp[15]) ? node7988 : node7969;
												assign node7969 = (inp[3]) ? node7977 : node7970;
													assign node7970 = (inp[14]) ? node7972 : 4'b0111;
														assign node7972 = (inp[6]) ? node7974 : 4'b1101;
															assign node7974 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node7977 = (inp[5]) ? node7983 : node7978;
														assign node7978 = (inp[6]) ? 4'b1101 : node7979;
															assign node7979 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node7983 = (inp[11]) ? node7985 : 4'b0101;
															assign node7985 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node7988 = (inp[14]) ? node7990 : 4'b0111;
													assign node7990 = (inp[11]) ? node7996 : node7991;
														assign node7991 = (inp[6]) ? node7993 : 4'b0111;
															assign node7993 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node7996 = (inp[6]) ? 4'b0111 : 4'b1111;
											assign node7999 = (inp[15]) ? node8009 : node8000;
												assign node8000 = (inp[3]) ? node8004 : node8001;
													assign node8001 = (inp[5]) ? 4'b0111 : 4'b1101;
													assign node8004 = (inp[5]) ? 4'b1111 : node8005;
														assign node8005 = (inp[11]) ? 4'b1111 : 4'b0111;
												assign node8009 = (inp[3]) ? node8013 : node8010;
													assign node8010 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node8013 = (inp[6]) ? node8017 : node8014;
														assign node8014 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node8017 = (inp[11]) ? 4'b0101 : 4'b1101;
							assign node8020 = (inp[8]) ? node8202 : node8021;
								assign node8021 = (inp[2]) ? node8099 : node8022;
									assign node8022 = (inp[14]) ? node8062 : node8023;
										assign node8023 = (inp[15]) ? node8041 : node8024;
											assign node8024 = (inp[0]) ? node8032 : node8025;
												assign node8025 = (inp[3]) ? node8027 : 4'b0110;
													assign node8027 = (inp[11]) ? node8029 : 4'b0100;
														assign node8029 = (inp[6]) ? 4'b1100 : 4'b0100;
												assign node8032 = (inp[5]) ? node8036 : node8033;
													assign node8033 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node8036 = (inp[1]) ? 4'b0110 : node8037;
														assign node8037 = (inp[11]) ? 4'b1110 : 4'b0110;
											assign node8041 = (inp[0]) ? node8055 : node8042;
												assign node8042 = (inp[3]) ? node8052 : node8043;
													assign node8043 = (inp[5]) ? node8049 : node8044;
														assign node8044 = (inp[1]) ? 4'b1100 : node8045;
															assign node8045 = (inp[11]) ? 4'b0100 : 4'b1100;
														assign node8049 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node8052 = (inp[1]) ? 4'b0110 : 4'b1110;
												assign node8055 = (inp[5]) ? 4'b0100 : node8056;
													assign node8056 = (inp[6]) ? 4'b1110 : node8057;
														assign node8057 = (inp[11]) ? 4'b0110 : 4'b1110;
										assign node8062 = (inp[1]) ? node8084 : node8063;
											assign node8063 = (inp[0]) ? node8079 : node8064;
												assign node8064 = (inp[5]) ? 4'b0101 : node8065;
													assign node8065 = (inp[15]) ? node8071 : node8066;
														assign node8066 = (inp[3]) ? 4'b0101 : node8067;
															assign node8067 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node8071 = (inp[3]) ? node8075 : node8072;
															assign node8072 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node8075 = (inp[11]) ? 4'b1111 : 4'b0111;
												assign node8079 = (inp[15]) ? 4'b1101 : node8080;
													assign node8080 = (inp[6]) ? 4'b0101 : 4'b1111;
											assign node8084 = (inp[0]) ? 4'b1111 : node8085;
												assign node8085 = (inp[15]) ? node8093 : node8086;
													assign node8086 = (inp[6]) ? node8090 : node8087;
														assign node8087 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node8090 = (inp[5]) ? 4'b0101 : 4'b1101;
													assign node8093 = (inp[11]) ? 4'b0111 : node8094;
														assign node8094 = (inp[3]) ? 4'b1111 : 4'b1101;
									assign node8099 = (inp[3]) ? node8149 : node8100;
										assign node8100 = (inp[11]) ? node8134 : node8101;
											assign node8101 = (inp[15]) ? node8117 : node8102;
												assign node8102 = (inp[1]) ? node8110 : node8103;
													assign node8103 = (inp[6]) ? 4'b0101 : node8104;
														assign node8104 = (inp[14]) ? 4'b1101 : node8105;
															assign node8105 = (inp[0]) ? 4'b1101 : 4'b1101;
													assign node8110 = (inp[6]) ? 4'b1101 : node8111;
														assign node8111 = (inp[0]) ? node8113 : 4'b0101;
															assign node8113 = (inp[14]) ? 4'b0101 : 4'b0111;
												assign node8117 = (inp[14]) ? node8127 : node8118;
													assign node8118 = (inp[1]) ? node8122 : node8119;
														assign node8119 = (inp[0]) ? 4'b1101 : 4'b0101;
														assign node8122 = (inp[6]) ? 4'b1101 : node8123;
															assign node8123 = (inp[0]) ? 4'b0101 : 4'b0101;
													assign node8127 = (inp[6]) ? node8131 : node8128;
														assign node8128 = (inp[1]) ? 4'b0101 : 4'b1101;
														assign node8131 = (inp[1]) ? 4'b1111 : 4'b0111;
											assign node8134 = (inp[5]) ? node8136 : 4'b0111;
												assign node8136 = (inp[15]) ? node8140 : node8137;
													assign node8137 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node8140 = (inp[0]) ? node8144 : node8141;
														assign node8141 = (inp[6]) ? 4'b0111 : 4'b1111;
														assign node8144 = (inp[1]) ? 4'b0101 : node8145;
															assign node8145 = (inp[6]) ? 4'b1101 : 4'b0101;
										assign node8149 = (inp[14]) ? node8171 : node8150;
											assign node8150 = (inp[6]) ? node8162 : node8151;
												assign node8151 = (inp[5]) ? node8157 : node8152;
													assign node8152 = (inp[0]) ? node8154 : 4'b1111;
														assign node8154 = (inp[15]) ? 4'b0101 : 4'b1111;
													assign node8157 = (inp[1]) ? 4'b1111 : node8158;
														assign node8158 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node8162 = (inp[11]) ? node8166 : node8163;
													assign node8163 = (inp[1]) ? 4'b1111 : 4'b0111;
													assign node8166 = (inp[1]) ? node8168 : 4'b1101;
														assign node8168 = (inp[5]) ? 4'b0111 : 4'b0101;
											assign node8171 = (inp[5]) ? node8187 : node8172;
												assign node8172 = (inp[11]) ? node8180 : node8173;
													assign node8173 = (inp[0]) ? node8175 : 4'b0111;
														assign node8175 = (inp[15]) ? 4'b1101 : node8176;
															assign node8176 = (inp[1]) ? 4'b0111 : 4'b1111;
													assign node8180 = (inp[1]) ? node8184 : node8181;
														assign node8181 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node8184 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node8187 = (inp[15]) ? node8195 : node8188;
													assign node8188 = (inp[0]) ? 4'b0111 : node8189;
														assign node8189 = (inp[1]) ? node8191 : 4'b0101;
															assign node8191 = (inp[11]) ? 4'b0101 : 4'b0101;
													assign node8195 = (inp[0]) ? node8197 : 4'b1111;
														assign node8197 = (inp[11]) ? node8199 : 4'b1101;
															assign node8199 = (inp[1]) ? 4'b0101 : 4'b1101;
								assign node8202 = (inp[2]) ? node8296 : node8203;
									assign node8203 = (inp[14]) ? node8259 : node8204;
										assign node8204 = (inp[0]) ? node8236 : node8205;
											assign node8205 = (inp[15]) ? node8221 : node8206;
												assign node8206 = (inp[3]) ? node8214 : node8207;
													assign node8207 = (inp[5]) ? 4'b0101 : node8208;
														assign node8208 = (inp[6]) ? 4'b1111 : node8209;
															assign node8209 = (inp[11]) ? 4'b1111 : 4'b0111;
													assign node8214 = (inp[11]) ? node8216 : 4'b0101;
														assign node8216 = (inp[6]) ? node8218 : 4'b1101;
															assign node8218 = (inp[5]) ? 4'b0101 : 4'b1101;
												assign node8221 = (inp[6]) ? 4'b0111 : node8222;
													assign node8222 = (inp[5]) ? node8228 : node8223;
														assign node8223 = (inp[11]) ? 4'b0101 : node8224;
															assign node8224 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node8228 = (inp[11]) ? node8232 : node8229;
															assign node8229 = (inp[1]) ? 4'b0111 : 4'b1111;
															assign node8232 = (inp[1]) ? 4'b1111 : 4'b0111;
											assign node8236 = (inp[15]) ? node8252 : node8237;
												assign node8237 = (inp[3]) ? node8247 : node8238;
													assign node8238 = (inp[5]) ? 4'b1111 : node8239;
														assign node8239 = (inp[6]) ? node8243 : node8240;
															assign node8240 = (inp[1]) ? 4'b1101 : 4'b0101;
															assign node8243 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node8247 = (inp[11]) ? 4'b0111 : node8248;
														assign node8248 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node8252 = (inp[1]) ? 4'b0101 : node8253;
													assign node8253 = (inp[11]) ? node8255 : 4'b1101;
														assign node8255 = (inp[6]) ? 4'b1101 : 4'b0101;
										assign node8259 = (inp[15]) ? node8279 : node8260;
											assign node8260 = (inp[6]) ? node8270 : node8261;
												assign node8261 = (inp[1]) ? node8265 : node8262;
													assign node8262 = (inp[11]) ? 4'b0110 : 4'b1100;
													assign node8265 = (inp[0]) ? node8267 : 4'b1100;
														assign node8267 = (inp[11]) ? 4'b1110 : 4'b0110;
												assign node8270 = (inp[11]) ? node8272 : 4'b1100;
													assign node8272 = (inp[1]) ? node8274 : 4'b1100;
														assign node8274 = (inp[5]) ? 4'b0100 : node8275;
															assign node8275 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node8279 = (inp[6]) ? node8291 : node8280;
												assign node8280 = (inp[5]) ? node8286 : node8281;
													assign node8281 = (inp[0]) ? 4'b0110 : node8282;
														assign node8282 = (inp[1]) ? 4'b1100 : 4'b0100;
													assign node8286 = (inp[11]) ? 4'b0100 : node8287;
														assign node8287 = (inp[1]) ? 4'b0100 : 4'b1100;
												assign node8291 = (inp[0]) ? 4'b0100 : node8292;
													assign node8292 = (inp[5]) ? 4'b0110 : 4'b0100;
									assign node8296 = (inp[5]) ? node8336 : node8297;
										assign node8297 = (inp[11]) ? node8319 : node8298;
											assign node8298 = (inp[1]) ? node8302 : node8299;
												assign node8299 = (inp[6]) ? 4'b0100 : 4'b1100;
												assign node8302 = (inp[6]) ? node8312 : node8303;
													assign node8303 = (inp[14]) ? 4'b0110 : node8304;
														assign node8304 = (inp[15]) ? node8308 : node8305;
															assign node8305 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node8308 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node8312 = (inp[0]) ? node8314 : 4'b1100;
														assign node8314 = (inp[3]) ? 4'b1100 : node8315;
															assign node8315 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node8319 = (inp[0]) ? node8331 : node8320;
												assign node8320 = (inp[14]) ? 4'b1100 : node8321;
													assign node8321 = (inp[3]) ? 4'b1100 : node8322;
														assign node8322 = (inp[1]) ? node8326 : node8323;
															assign node8323 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node8326 = (inp[6]) ? 4'b0100 : 4'b1100;
												assign node8331 = (inp[3]) ? 4'b1110 : node8332;
													assign node8332 = (inp[15]) ? 4'b1110 : 4'b1100;
										assign node8336 = (inp[15]) ? node8354 : node8337;
											assign node8337 = (inp[0]) ? node8343 : node8338;
												assign node8338 = (inp[6]) ? node8340 : 4'b0100;
													assign node8340 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node8343 = (inp[3]) ? 4'b0110 : node8344;
													assign node8344 = (inp[6]) ? node8346 : 4'b0110;
														assign node8346 = (inp[14]) ? node8350 : node8347;
															assign node8347 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node8350 = (inp[1]) ? 4'b0110 : 4'b0110;
											assign node8354 = (inp[0]) ? node8368 : node8355;
												assign node8355 = (inp[6]) ? node8361 : node8356;
													assign node8356 = (inp[14]) ? 4'b1110 : node8357;
														assign node8357 = (inp[11]) ? 4'b1110 : 4'b0110;
													assign node8361 = (inp[1]) ? node8365 : node8362;
														assign node8362 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node8365 = (inp[11]) ? 4'b0110 : 4'b1110;
												assign node8368 = (inp[14]) ? node8378 : node8369;
													assign node8369 = (inp[6]) ? node8375 : node8370;
														assign node8370 = (inp[3]) ? node8372 : 4'b1100;
															assign node8372 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node8375 = (inp[3]) ? 4'b1100 : 4'b0100;
													assign node8378 = (inp[1]) ? 4'b1100 : 4'b0100;
				assign node8381 = (inp[12]) ? node9837 : node8382;
					assign node8382 = (inp[10]) ? node9138 : node8383;
						assign node8383 = (inp[5]) ? node8775 : node8384;
							assign node8384 = (inp[11]) ? node8584 : node8385;
								assign node8385 = (inp[6]) ? node8489 : node8386;
									assign node8386 = (inp[1]) ? node8440 : node8387;
										assign node8387 = (inp[2]) ? node8413 : node8388;
											assign node8388 = (inp[3]) ? node8404 : node8389;
												assign node8389 = (inp[7]) ? node8393 : node8390;
													assign node8390 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node8393 = (inp[15]) ? node8401 : node8394;
														assign node8394 = (inp[0]) ? node8398 : node8395;
															assign node8395 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node8398 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node8401 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node8404 = (inp[0]) ? node8410 : node8405;
													assign node8405 = (inp[14]) ? 4'b1110 : node8406;
														assign node8406 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node8410 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node8413 = (inp[0]) ? node8427 : node8414;
												assign node8414 = (inp[7]) ? node8424 : node8415;
													assign node8415 = (inp[8]) ? node8419 : node8416;
														assign node8416 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node8419 = (inp[15]) ? node8421 : 4'b1101;
															assign node8421 = (inp[14]) ? 4'b1101 : 4'b1111;
													assign node8424 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node8427 = (inp[15]) ? node8435 : node8428;
													assign node8428 = (inp[3]) ? node8430 : 4'b1100;
														assign node8430 = (inp[7]) ? 4'b1110 : node8431;
															assign node8431 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node8435 = (inp[14]) ? node8437 : 4'b1110;
														assign node8437 = (inp[7]) ? 4'b1101 : 4'b1100;
										assign node8440 = (inp[7]) ? node8468 : node8441;
											assign node8441 = (inp[8]) ? node8459 : node8442;
												assign node8442 = (inp[2]) ? node8452 : node8443;
													assign node8443 = (inp[14]) ? node8445 : 4'b1101;
														assign node8445 = (inp[3]) ? node8449 : node8446;
															assign node8446 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node8449 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node8452 = (inp[14]) ? node8454 : 4'b1110;
														assign node8454 = (inp[3]) ? node8456 : 4'b1110;
															assign node8456 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node8459 = (inp[14]) ? node8463 : node8460;
													assign node8460 = (inp[2]) ? 4'b0111 : 4'b1110;
													assign node8463 = (inp[2]) ? 4'b0111 : node8464;
														assign node8464 = (inp[0]) ? 4'b0111 : 4'b0101;
											assign node8468 = (inp[8]) ? node8480 : node8469;
												assign node8469 = (inp[2]) ? node8473 : node8470;
													assign node8470 = (inp[0]) ? 4'b0111 : 4'b1110;
													assign node8473 = (inp[0]) ? 4'b0111 : node8474;
														assign node8474 = (inp[3]) ? node8476 : 4'b0101;
															assign node8476 = (inp[14]) ? 4'b0111 : 4'b0101;
												assign node8480 = (inp[14]) ? node8482 : 4'b0101;
													assign node8482 = (inp[0]) ? node8484 : 4'b0100;
														assign node8484 = (inp[3]) ? node8486 : 4'b0100;
															assign node8486 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node8489 = (inp[1]) ? node8533 : node8490;
										assign node8490 = (inp[3]) ? node8510 : node8491;
											assign node8491 = (inp[14]) ? node8505 : node8492;
												assign node8492 = (inp[7]) ? 4'b0100 : node8493;
													assign node8493 = (inp[15]) ? node8499 : node8494;
														assign node8494 = (inp[0]) ? node8496 : 4'b0111;
															assign node8496 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node8499 = (inp[0]) ? 4'b0111 : node8500;
															assign node8500 = (inp[8]) ? 4'b0101 : 4'b0100;
												assign node8505 = (inp[15]) ? node8507 : 4'b0101;
													assign node8507 = (inp[0]) ? 4'b0111 : 4'b0101;
											assign node8510 = (inp[7]) ? node8528 : node8511;
												assign node8511 = (inp[8]) ? node8521 : node8512;
													assign node8512 = (inp[2]) ? node8518 : node8513;
														assign node8513 = (inp[14]) ? 4'b0110 : node8514;
															assign node8514 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node8518 = (inp[14]) ? 4'b0100 : 4'b0110;
													assign node8521 = (inp[2]) ? node8523 : 4'b0110;
														assign node8523 = (inp[15]) ? 4'b0101 : node8524;
															assign node8524 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node8528 = (inp[15]) ? node8530 : 4'b0101;
													assign node8530 = (inp[8]) ? 4'b0110 : 4'b0100;
										assign node8533 = (inp[14]) ? node8561 : node8534;
											assign node8534 = (inp[3]) ? node8548 : node8535;
												assign node8535 = (inp[8]) ? node8543 : node8536;
													assign node8536 = (inp[7]) ? node8538 : 4'b0111;
														assign node8538 = (inp[0]) ? node8540 : 4'b1111;
															assign node8540 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node8543 = (inp[2]) ? node8545 : 4'b1101;
														assign node8545 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node8548 = (inp[2]) ? node8558 : node8549;
													assign node8549 = (inp[8]) ? node8555 : node8550;
														assign node8550 = (inp[7]) ? 4'b0110 : node8551;
															assign node8551 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node8555 = (inp[15]) ? 4'b0110 : 4'b1111;
													assign node8558 = (inp[8]) ? 4'b1101 : 4'b0100;
											assign node8561 = (inp[8]) ? node8569 : node8562;
												assign node8562 = (inp[15]) ? 4'b1111 : node8563;
													assign node8563 = (inp[0]) ? node8565 : 4'b1111;
														assign node8565 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node8569 = (inp[7]) ? node8577 : node8570;
													assign node8570 = (inp[15]) ? node8572 : 4'b1111;
														assign node8572 = (inp[2]) ? 4'b1101 : node8573;
															assign node8573 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node8577 = (inp[2]) ? node8579 : 4'b1110;
														assign node8579 = (inp[3]) ? 4'b1100 : node8580;
															assign node8580 = (inp[15]) ? 4'b1110 : 4'b1100;
								assign node8584 = (inp[6]) ? node8664 : node8585;
									assign node8585 = (inp[1]) ? node8633 : node8586;
										assign node8586 = (inp[0]) ? node8612 : node8587;
											assign node8587 = (inp[14]) ? node8597 : node8588;
												assign node8588 = (inp[3]) ? node8594 : node8589;
													assign node8589 = (inp[15]) ? 4'b0101 : node8590;
														assign node8590 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node8594 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node8597 = (inp[2]) ? node8607 : node8598;
													assign node8598 = (inp[7]) ? node8602 : node8599;
														assign node8599 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node8602 = (inp[8]) ? node8604 : 4'b0111;
															assign node8604 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node8607 = (inp[15]) ? node8609 : 4'b0111;
														assign node8609 = (inp[8]) ? 4'b0101 : 4'b0100;
											assign node8612 = (inp[15]) ? node8624 : node8613;
												assign node8613 = (inp[3]) ? node8621 : node8614;
													assign node8614 = (inp[2]) ? 4'b0101 : node8615;
														assign node8615 = (inp[7]) ? node8617 : 4'b0101;
															assign node8617 = (inp[8]) ? 4'b0100 : 4'b0100;
													assign node8621 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node8624 = (inp[3]) ? node8626 : 4'b0110;
													assign node8626 = (inp[14]) ? node8628 : 4'b0100;
														assign node8628 = (inp[7]) ? 4'b0100 : node8629;
															assign node8629 = (inp[8]) ? 4'b0101 : 4'b0100;
										assign node8633 = (inp[8]) ? node8645 : node8634;
											assign node8634 = (inp[7]) ? node8638 : node8635;
												assign node8635 = (inp[14]) ? 4'b0100 : 4'b0110;
												assign node8638 = (inp[3]) ? 4'b1101 : node8639;
													assign node8639 = (inp[0]) ? 4'b1111 : node8640;
														assign node8640 = (inp[2]) ? 4'b1101 : 4'b1111;
											assign node8645 = (inp[7]) ? node8659 : node8646;
												assign node8646 = (inp[3]) ? node8650 : node8647;
													assign node8647 = (inp[2]) ? 4'b1111 : 4'b1101;
													assign node8650 = (inp[14]) ? node8652 : 4'b1101;
														assign node8652 = (inp[2]) ? node8656 : node8653;
															assign node8653 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node8656 = (inp[0]) ? 4'b1101 : 4'b1101;
												assign node8659 = (inp[2]) ? 4'b1100 : node8660;
													assign node8660 = (inp[15]) ? 4'b1111 : 4'b1100;
									assign node8664 = (inp[1]) ? node8716 : node8665;
										assign node8665 = (inp[2]) ? node8695 : node8666;
											assign node8666 = (inp[8]) ? node8680 : node8667;
												assign node8667 = (inp[7]) ? node8675 : node8668;
													assign node8668 = (inp[14]) ? 4'b1110 : node8669;
														assign node8669 = (inp[3]) ? 4'b1111 : node8670;
															assign node8670 = (inp[0]) ? 4'b1101 : 4'b1101;
													assign node8675 = (inp[15]) ? node8677 : 4'b1101;
														assign node8677 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node8680 = (inp[15]) ? node8688 : node8681;
													assign node8681 = (inp[7]) ? node8685 : node8682;
														assign node8682 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node8685 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node8688 = (inp[0]) ? node8692 : node8689;
														assign node8689 = (inp[14]) ? 4'b1100 : 4'b1110;
														assign node8692 = (inp[14]) ? 4'b1110 : 4'b1111;
											assign node8695 = (inp[8]) ? node8701 : node8696;
												assign node8696 = (inp[7]) ? node8698 : 4'b1100;
													assign node8698 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node8701 = (inp[14]) ? node8709 : node8702;
													assign node8702 = (inp[3]) ? 4'b1101 : node8703;
														assign node8703 = (inp[0]) ? 4'b1101 : node8704;
															assign node8704 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node8709 = (inp[7]) ? 4'b1110 : node8710;
														assign node8710 = (inp[15]) ? node8712 : 4'b1111;
															assign node8712 = (inp[3]) ? 4'b1111 : 4'b1101;
										assign node8716 = (inp[7]) ? node8746 : node8717;
											assign node8717 = (inp[8]) ? node8731 : node8718;
												assign node8718 = (inp[0]) ? node8728 : node8719;
													assign node8719 = (inp[14]) ? node8723 : node8720;
														assign node8720 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node8723 = (inp[15]) ? node8725 : 4'b1100;
															assign node8725 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node8728 = (inp[14]) ? 4'b1110 : 4'b1101;
												assign node8731 = (inp[2]) ? node8741 : node8732;
													assign node8732 = (inp[14]) ? node8738 : node8733;
														assign node8733 = (inp[3]) ? node8735 : 4'b1100;
															assign node8735 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node8738 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node8741 = (inp[14]) ? node8743 : 4'b0101;
														assign node8743 = (inp[3]) ? 4'b0111 : 4'b0101;
											assign node8746 = (inp[8]) ? node8758 : node8747;
												assign node8747 = (inp[14]) ? node8751 : node8748;
													assign node8748 = (inp[2]) ? 4'b0101 : 4'b1100;
													assign node8751 = (inp[15]) ? node8753 : 4'b0111;
														assign node8753 = (inp[0]) ? node8755 : 4'b0111;
															assign node8755 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node8758 = (inp[14]) ? node8762 : node8759;
													assign node8759 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node8762 = (inp[15]) ? node8770 : node8763;
														assign node8763 = (inp[3]) ? node8767 : node8764;
															assign node8764 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node8767 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node8770 = (inp[3]) ? node8772 : 4'b0100;
															assign node8772 = (inp[0]) ? 4'b0100 : 4'b0110;
							assign node8775 = (inp[7]) ? node8957 : node8776;
								assign node8776 = (inp[8]) ? node8856 : node8777;
									assign node8777 = (inp[2]) ? node8813 : node8778;
										assign node8778 = (inp[14]) ? node8800 : node8779;
											assign node8779 = (inp[11]) ? node8787 : node8780;
												assign node8780 = (inp[6]) ? 4'b0111 : node8781;
													assign node8781 = (inp[0]) ? 4'b1111 : node8782;
														assign node8782 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node8787 = (inp[6]) ? node8793 : node8788;
													assign node8788 = (inp[15]) ? node8790 : 4'b0101;
														assign node8790 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node8793 = (inp[0]) ? node8797 : node8794;
														assign node8794 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node8797 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node8800 = (inp[3]) ? node8808 : node8801;
												assign node8801 = (inp[15]) ? 4'b1100 : node8802;
													assign node8802 = (inp[1]) ? node8804 : 4'b1110;
														assign node8804 = (inp[6]) ? 4'b1110 : 4'b0110;
												assign node8808 = (inp[15]) ? node8810 : 4'b0110;
													assign node8810 = (inp[0]) ? 4'b0100 : 4'b0110;
										assign node8813 = (inp[1]) ? node8837 : node8814;
											assign node8814 = (inp[3]) ? node8830 : node8815;
												assign node8815 = (inp[15]) ? node8823 : node8816;
													assign node8816 = (inp[0]) ? node8818 : 4'b1100;
														assign node8818 = (inp[11]) ? 4'b1110 : node8819;
															assign node8819 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node8823 = (inp[6]) ? node8827 : node8824;
														assign node8824 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node8827 = (inp[11]) ? 4'b1110 : 4'b0110;
												assign node8830 = (inp[0]) ? node8834 : node8831;
													assign node8831 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node8834 = (inp[11]) ? 4'b1110 : 4'b0110;
											assign node8837 = (inp[11]) ? node8847 : node8838;
												assign node8838 = (inp[6]) ? node8844 : node8839;
													assign node8839 = (inp[0]) ? 4'b1100 : node8840;
														assign node8840 = (inp[14]) ? 4'b1110 : 4'b1100;
													assign node8844 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node8847 = (inp[6]) ? node8853 : node8848;
													assign node8848 = (inp[0]) ? 4'b0100 : node8849;
														assign node8849 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node8853 = (inp[14]) ? 4'b1100 : 4'b1110;
									assign node8856 = (inp[2]) ? node8908 : node8857;
										assign node8857 = (inp[14]) ? node8883 : node8858;
											assign node8858 = (inp[6]) ? node8872 : node8859;
												assign node8859 = (inp[11]) ? node8867 : node8860;
													assign node8860 = (inp[1]) ? 4'b1100 : node8861;
														assign node8861 = (inp[0]) ? 4'b1110 : node8862;
															assign node8862 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node8867 = (inp[1]) ? 4'b0100 : node8868;
														assign node8868 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node8872 = (inp[11]) ? node8874 : 4'b0100;
													assign node8874 = (inp[1]) ? node8878 : node8875;
														assign node8875 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node8878 = (inp[3]) ? 4'b1110 : node8879;
															assign node8879 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node8883 = (inp[11]) ? node8893 : node8884;
												assign node8884 = (inp[6]) ? 4'b1101 : node8885;
													assign node8885 = (inp[1]) ? 4'b0111 : node8886;
														assign node8886 = (inp[0]) ? 4'b1111 : node8887;
															assign node8887 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node8893 = (inp[15]) ? node8901 : node8894;
													assign node8894 = (inp[1]) ? node8898 : node8895;
														assign node8895 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node8898 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node8901 = (inp[0]) ? 4'b0101 : node8902;
														assign node8902 = (inp[1]) ? 4'b0111 : node8903;
															assign node8903 = (inp[6]) ? 4'b1111 : 4'b0111;
										assign node8908 = (inp[0]) ? node8926 : node8909;
											assign node8909 = (inp[15]) ? node8921 : node8910;
												assign node8910 = (inp[1]) ? node8916 : node8911;
													assign node8911 = (inp[6]) ? node8913 : 4'b1101;
														assign node8913 = (inp[14]) ? 4'b1101 : 4'b0101;
													assign node8916 = (inp[11]) ? node8918 : 4'b0101;
														assign node8918 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node8921 = (inp[3]) ? node8923 : 4'b0111;
													assign node8923 = (inp[14]) ? 4'b1111 : 4'b0111;
											assign node8926 = (inp[15]) ? node8948 : node8927;
												assign node8927 = (inp[14]) ? node8939 : node8928;
													assign node8928 = (inp[11]) ? node8934 : node8929;
														assign node8929 = (inp[6]) ? 4'b0111 : node8930;
															assign node8930 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node8934 = (inp[1]) ? 4'b1111 : node8935;
															assign node8935 = (inp[6]) ? 4'b1111 : 4'b0111;
													assign node8939 = (inp[1]) ? 4'b0111 : node8940;
														assign node8940 = (inp[11]) ? node8944 : node8941;
															assign node8941 = (inp[3]) ? 4'b1111 : 4'b0111;
															assign node8944 = (inp[6]) ? 4'b1111 : 4'b0111;
												assign node8948 = (inp[14]) ? node8950 : 4'b1101;
													assign node8950 = (inp[6]) ? node8952 : 4'b0101;
														assign node8952 = (inp[3]) ? 4'b1101 : node8953;
															assign node8953 = (inp[11]) ? 4'b0101 : 4'b1101;
								assign node8957 = (inp[8]) ? node9039 : node8958;
									assign node8958 = (inp[14]) ? node8996 : node8959;
										assign node8959 = (inp[2]) ? node8979 : node8960;
											assign node8960 = (inp[1]) ? node8970 : node8961;
												assign node8961 = (inp[3]) ? 4'b0110 : node8962;
													assign node8962 = (inp[6]) ? 4'b1110 : node8963;
														assign node8963 = (inp[0]) ? 4'b1100 : node8964;
															assign node8964 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node8970 = (inp[11]) ? node8976 : node8971;
													assign node8971 = (inp[3]) ? node8973 : 4'b0110;
														assign node8973 = (inp[0]) ? 4'b1100 : 4'b0100;
													assign node8976 = (inp[6]) ? 4'b1100 : 4'b0110;
											assign node8979 = (inp[15]) ? node8987 : node8980;
												assign node8980 = (inp[0]) ? node8984 : node8981;
													assign node8981 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node8984 = (inp[11]) ? 4'b0111 : 4'b1111;
												assign node8987 = (inp[0]) ? node8989 : 4'b0111;
													assign node8989 = (inp[11]) ? node8991 : 4'b0101;
														assign node8991 = (inp[6]) ? 4'b1101 : node8992;
															assign node8992 = (inp[1]) ? 4'b1101 : 4'b0101;
										assign node8996 = (inp[0]) ? node9022 : node8997;
											assign node8997 = (inp[15]) ? node9007 : node8998;
												assign node8998 = (inp[11]) ? node9004 : node8999;
													assign node8999 = (inp[1]) ? node9001 : 4'b1101;
														assign node9001 = (inp[2]) ? 4'b0101 : 4'b1101;
													assign node9004 = (inp[2]) ? 4'b1101 : 4'b0101;
												assign node9007 = (inp[6]) ? node9015 : node9008;
													assign node9008 = (inp[3]) ? node9010 : 4'b0111;
														assign node9010 = (inp[2]) ? 4'b1111 : node9011;
															assign node9011 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node9015 = (inp[3]) ? node9017 : 4'b1111;
														assign node9017 = (inp[11]) ? 4'b1111 : node9018;
															assign node9018 = (inp[2]) ? 4'b0111 : 4'b1111;
											assign node9022 = (inp[15]) ? node9036 : node9023;
												assign node9023 = (inp[1]) ? node9031 : node9024;
													assign node9024 = (inp[6]) ? node9028 : node9025;
														assign node9025 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node9028 = (inp[11]) ? 4'b1111 : 4'b0111;
													assign node9031 = (inp[3]) ? 4'b0111 : node9032;
														assign node9032 = (inp[11]) ? 4'b0111 : 4'b1111;
												assign node9036 = (inp[3]) ? 4'b0101 : 4'b1101;
									assign node9039 = (inp[14]) ? node9093 : node9040;
										assign node9040 = (inp[2]) ? node9074 : node9041;
											assign node9041 = (inp[3]) ? node9059 : node9042;
												assign node9042 = (inp[1]) ? node9054 : node9043;
													assign node9043 = (inp[0]) ? node9051 : node9044;
														assign node9044 = (inp[15]) ? node9048 : node9045;
															assign node9045 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node9048 = (inp[6]) ? 4'b0111 : 4'b0111;
														assign node9051 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node9054 = (inp[15]) ? 4'b1101 : node9055;
														assign node9055 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node9059 = (inp[15]) ? node9067 : node9060;
													assign node9060 = (inp[0]) ? node9062 : 4'b1101;
														assign node9062 = (inp[6]) ? node9064 : 4'b1111;
															assign node9064 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node9067 = (inp[0]) ? node9069 : 4'b0111;
														assign node9069 = (inp[6]) ? node9071 : 4'b0101;
															assign node9071 = (inp[1]) ? 4'b0101 : 4'b1101;
											assign node9074 = (inp[6]) ? node9084 : node9075;
												assign node9075 = (inp[1]) ? node9077 : 4'b0100;
													assign node9077 = (inp[11]) ? node9079 : 4'b0100;
														assign node9079 = (inp[3]) ? node9081 : 4'b1100;
															assign node9081 = (inp[15]) ? 4'b1100 : 4'b1100;
												assign node9084 = (inp[15]) ? node9086 : 4'b0110;
													assign node9086 = (inp[0]) ? node9088 : 4'b0110;
														assign node9088 = (inp[11]) ? node9090 : 4'b1100;
															assign node9090 = (inp[1]) ? 4'b0100 : 4'b1100;
										assign node9093 = (inp[11]) ? node9121 : node9094;
											assign node9094 = (inp[1]) ? node9102 : node9095;
												assign node9095 = (inp[6]) ? 4'b0100 : node9096;
													assign node9096 = (inp[0]) ? node9098 : 4'b1100;
														assign node9098 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node9102 = (inp[6]) ? node9110 : node9103;
													assign node9103 = (inp[2]) ? node9105 : 4'b0100;
														assign node9105 = (inp[3]) ? 4'b0110 : node9106;
															assign node9106 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node9110 = (inp[3]) ? node9116 : node9111;
														assign node9111 = (inp[0]) ? node9113 : 4'b1110;
															assign node9113 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node9116 = (inp[0]) ? 4'b1100 : node9117;
															assign node9117 = (inp[2]) ? 4'b1110 : 4'b1100;
											assign node9121 = (inp[15]) ? node9129 : node9122;
												assign node9122 = (inp[0]) ? node9124 : 4'b0100;
													assign node9124 = (inp[1]) ? node9126 : 4'b0110;
														assign node9126 = (inp[3]) ? 4'b0110 : 4'b1110;
												assign node9129 = (inp[0]) ? 4'b0100 : node9130;
													assign node9130 = (inp[3]) ? node9132 : 4'b1110;
														assign node9132 = (inp[2]) ? 4'b0110 : node9133;
															assign node9133 = (inp[6]) ? 4'b0110 : 4'b1110;
						assign node9138 = (inp[11]) ? node9480 : node9139;
							assign node9139 = (inp[6]) ? node9307 : node9140;
								assign node9140 = (inp[1]) ? node9216 : node9141;
									assign node9141 = (inp[7]) ? node9171 : node9142;
										assign node9142 = (inp[8]) ? node9160 : node9143;
											assign node9143 = (inp[2]) ? node9151 : node9144;
												assign node9144 = (inp[14]) ? 4'b1110 : node9145;
													assign node9145 = (inp[15]) ? node9147 : 4'b1111;
														assign node9147 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node9151 = (inp[3]) ? node9153 : 4'b1110;
													assign node9153 = (inp[15]) ? node9157 : node9154;
														assign node9154 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node9157 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node9160 = (inp[14]) ? node9164 : node9161;
												assign node9161 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node9164 = (inp[3]) ? 4'b1111 : node9165;
													assign node9165 = (inp[2]) ? node9167 : 4'b1101;
														assign node9167 = (inp[5]) ? 4'b1101 : 4'b1111;
										assign node9171 = (inp[8]) ? node9201 : node9172;
											assign node9172 = (inp[14]) ? node9180 : node9173;
												assign node9173 = (inp[2]) ? node9177 : node9174;
													assign node9174 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node9177 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node9180 = (inp[5]) ? node9194 : node9181;
													assign node9181 = (inp[2]) ? node9189 : node9182;
														assign node9182 = (inp[0]) ? node9186 : node9183;
															assign node9183 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node9186 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node9189 = (inp[0]) ? 4'b1111 : node9190;
															assign node9190 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node9194 = (inp[3]) ? node9196 : 4'b1101;
														assign node9196 = (inp[2]) ? node9198 : 4'b1111;
															assign node9198 = (inp[15]) ? 4'b1101 : 4'b1101;
											assign node9201 = (inp[14]) ? node9211 : node9202;
												assign node9202 = (inp[2]) ? 4'b1110 : node9203;
													assign node9203 = (inp[5]) ? node9205 : 4'b1111;
														assign node9205 = (inp[15]) ? 4'b1101 : node9206;
															assign node9206 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node9211 = (inp[2]) ? node9213 : 4'b1100;
													assign node9213 = (inp[5]) ? 4'b1110 : 4'b1100;
									assign node9216 = (inp[7]) ? node9266 : node9217;
										assign node9217 = (inp[8]) ? node9239 : node9218;
											assign node9218 = (inp[14]) ? node9228 : node9219;
												assign node9219 = (inp[2]) ? node9223 : node9220;
													assign node9220 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node9223 = (inp[0]) ? 4'b1110 : node9224;
														assign node9224 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node9228 = (inp[15]) ? node9234 : node9229;
													assign node9229 = (inp[0]) ? 4'b1110 : node9230;
														assign node9230 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node9234 = (inp[0]) ? 4'b1100 : node9235;
														assign node9235 = (inp[3]) ? 4'b1110 : 4'b1100;
											assign node9239 = (inp[14]) ? node9251 : node9240;
												assign node9240 = (inp[2]) ? node9248 : node9241;
													assign node9241 = (inp[5]) ? node9243 : 4'b1100;
														assign node9243 = (inp[15]) ? node9245 : 4'b1100;
															assign node9245 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node9248 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node9251 = (inp[15]) ? node9257 : node9252;
													assign node9252 = (inp[3]) ? 4'b0111 : node9253;
														assign node9253 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node9257 = (inp[0]) ? node9261 : node9258;
														assign node9258 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node9261 = (inp[3]) ? 4'b0101 : node9262;
															assign node9262 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node9266 = (inp[8]) ? node9282 : node9267;
											assign node9267 = (inp[2]) ? node9273 : node9268;
												assign node9268 = (inp[14]) ? node9270 : 4'b1110;
													assign node9270 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node9273 = (inp[14]) ? node9275 : 4'b0101;
													assign node9275 = (inp[15]) ? 4'b0111 : node9276;
														assign node9276 = (inp[0]) ? 4'b0101 : node9277;
															assign node9277 = (inp[5]) ? 4'b0101 : 4'b0111;
											assign node9282 = (inp[14]) ? node9296 : node9283;
												assign node9283 = (inp[2]) ? node9289 : node9284;
													assign node9284 = (inp[15]) ? 4'b0101 : node9285;
														assign node9285 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node9289 = (inp[3]) ? node9291 : 4'b0110;
														assign node9291 = (inp[0]) ? node9293 : 4'b0100;
															assign node9293 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node9296 = (inp[2]) ? 4'b0100 : node9297;
													assign node9297 = (inp[5]) ? 4'b0100 : node9298;
														assign node9298 = (inp[3]) ? node9302 : node9299;
															assign node9299 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node9302 = (inp[0]) ? 4'b0100 : 4'b0110;
								assign node9307 = (inp[1]) ? node9387 : node9308;
									assign node9308 = (inp[0]) ? node9346 : node9309;
										assign node9309 = (inp[15]) ? node9327 : node9310;
											assign node9310 = (inp[3]) ? node9322 : node9311;
												assign node9311 = (inp[5]) ? node9319 : node9312;
													assign node9312 = (inp[14]) ? node9314 : 4'b0110;
														assign node9314 = (inp[7]) ? node9316 : 4'b0110;
															assign node9316 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node9319 = (inp[8]) ? 4'b0101 : 4'b0100;
												assign node9322 = (inp[8]) ? node9324 : 4'b0100;
													assign node9324 = (inp[14]) ? 4'b0101 : 4'b0100;
											assign node9327 = (inp[3]) ? node9339 : node9328;
												assign node9328 = (inp[5]) ? node9330 : 4'b0100;
													assign node9330 = (inp[7]) ? 4'b0110 : node9331;
														assign node9331 = (inp[8]) ? node9335 : node9332;
															assign node9332 = (inp[2]) ? 4'b0110 : 4'b0110;
															assign node9335 = (inp[14]) ? 4'b0111 : 4'b0110;
												assign node9339 = (inp[5]) ? node9341 : 4'b0111;
													assign node9341 = (inp[14]) ? node9343 : 4'b0111;
														assign node9343 = (inp[8]) ? 4'b0111 : 4'b0110;
										assign node9346 = (inp[15]) ? node9364 : node9347;
											assign node9347 = (inp[3]) ? node9357 : node9348;
												assign node9348 = (inp[5]) ? 4'b0111 : node9349;
													assign node9349 = (inp[2]) ? 4'b0101 : node9350;
														assign node9350 = (inp[8]) ? 4'b0100 : node9351;
															assign node9351 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node9357 = (inp[8]) ? node9359 : 4'b0111;
													assign node9359 = (inp[2]) ? 4'b0110 : node9360;
														assign node9360 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node9364 = (inp[3]) ? node9380 : node9365;
												assign node9365 = (inp[5]) ? node9377 : node9366;
													assign node9366 = (inp[14]) ? node9372 : node9367;
														assign node9367 = (inp[8]) ? 4'b0111 : node9368;
															assign node9368 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node9372 = (inp[2]) ? 4'b0110 : node9373;
															assign node9373 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node9377 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node9380 = (inp[7]) ? 4'b0100 : node9381;
													assign node9381 = (inp[8]) ? 4'b0101 : node9382;
														assign node9382 = (inp[2]) ? 4'b0100 : 4'b0101;
									assign node9387 = (inp[7]) ? node9431 : node9388;
										assign node9388 = (inp[8]) ? node9416 : node9389;
											assign node9389 = (inp[14]) ? node9401 : node9390;
												assign node9390 = (inp[2]) ? node9398 : node9391;
													assign node9391 = (inp[0]) ? 4'b0101 : node9392;
														assign node9392 = (inp[5]) ? 4'b0101 : node9393;
															assign node9393 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node9398 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node9401 = (inp[15]) ? node9411 : node9402;
													assign node9402 = (inp[3]) ? node9408 : node9403;
														assign node9403 = (inp[0]) ? node9405 : 4'b0110;
															assign node9405 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node9408 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node9411 = (inp[3]) ? node9413 : 4'b0100;
														assign node9413 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node9416 = (inp[14]) ? node9422 : node9417;
												assign node9417 = (inp[2]) ? 4'b1011 : node9418;
													assign node9418 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node9422 = (inp[2]) ? 4'b1011 : node9423;
													assign node9423 = (inp[3]) ? 4'b1001 : node9424;
														assign node9424 = (inp[15]) ? node9426 : 4'b1011;
															assign node9426 = (inp[0]) ? 4'b1001 : 4'b1001;
										assign node9431 = (inp[8]) ? node9459 : node9432;
											assign node9432 = (inp[14]) ? node9444 : node9433;
												assign node9433 = (inp[2]) ? node9437 : node9434;
													assign node9434 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node9437 = (inp[3]) ? 4'b1001 : node9438;
														assign node9438 = (inp[15]) ? node9440 : 4'b1011;
															assign node9440 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node9444 = (inp[2]) ? node9450 : node9445;
													assign node9445 = (inp[0]) ? 4'b1011 : node9446;
														assign node9446 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node9450 = (inp[0]) ? 4'b1001 : node9451;
														assign node9451 = (inp[3]) ? node9455 : node9452;
															assign node9452 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node9455 = (inp[15]) ? 4'b1011 : 4'b1001;
											assign node9459 = (inp[2]) ? node9475 : node9460;
												assign node9460 = (inp[14]) ? node9472 : node9461;
													assign node9461 = (inp[5]) ? node9467 : node9462;
														assign node9462 = (inp[15]) ? 4'b1011 : node9463;
															assign node9463 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node9467 = (inp[15]) ? 4'b1001 : node9468;
															assign node9468 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node9472 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node9475 = (inp[5]) ? 4'b1010 : node9476;
													assign node9476 = (inp[14]) ? 4'b1010 : 4'b1000;
							assign node9480 = (inp[6]) ? node9668 : node9481;
								assign node9481 = (inp[1]) ? node9575 : node9482;
									assign node9482 = (inp[0]) ? node9528 : node9483;
										assign node9483 = (inp[8]) ? node9501 : node9484;
											assign node9484 = (inp[7]) ? node9494 : node9485;
												assign node9485 = (inp[5]) ? node9491 : node9486;
													assign node9486 = (inp[14]) ? 4'b0100 : node9487;
														assign node9487 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node9491 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node9494 = (inp[3]) ? 4'b0101 : node9495;
													assign node9495 = (inp[2]) ? node9497 : 4'b0101;
														assign node9497 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node9501 = (inp[7]) ? node9513 : node9502;
												assign node9502 = (inp[3]) ? 4'b0111 : node9503;
													assign node9503 = (inp[5]) ? node9507 : node9504;
														assign node9504 = (inp[14]) ? 4'b0101 : 4'b0111;
														assign node9507 = (inp[14]) ? 4'b0101 : node9508;
															assign node9508 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node9513 = (inp[15]) ? node9521 : node9514;
													assign node9514 = (inp[2]) ? node9518 : node9515;
														assign node9515 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node9518 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node9521 = (inp[3]) ? node9525 : node9522;
														assign node9522 = (inp[14]) ? 4'b0100 : 4'b0110;
														assign node9525 = (inp[14]) ? 4'b0110 : 4'b0111;
										assign node9528 = (inp[15]) ? node9548 : node9529;
											assign node9529 = (inp[2]) ? node9539 : node9530;
												assign node9530 = (inp[8]) ? node9534 : node9531;
													assign node9531 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node9534 = (inp[7]) ? node9536 : 4'b0110;
														assign node9536 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node9539 = (inp[5]) ? 4'b0111 : node9540;
													assign node9540 = (inp[14]) ? node9542 : 4'b0110;
														assign node9542 = (inp[7]) ? node9544 : 4'b0111;
															assign node9544 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node9548 = (inp[5]) ? node9562 : node9549;
												assign node9549 = (inp[3]) ? node9555 : node9550;
													assign node9550 = (inp[7]) ? node9552 : 4'b0110;
														assign node9552 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node9555 = (inp[8]) ? node9557 : 4'b0100;
														assign node9557 = (inp[2]) ? node9559 : 4'b0100;
															assign node9559 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node9562 = (inp[2]) ? node9570 : node9563;
													assign node9563 = (inp[3]) ? 4'b0100 : node9564;
														assign node9564 = (inp[7]) ? 4'b0101 : node9565;
															assign node9565 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node9570 = (inp[8]) ? 4'b0100 : node9571;
														assign node9571 = (inp[7]) ? 4'b0101 : 4'b0100;
									assign node9575 = (inp[7]) ? node9625 : node9576;
										assign node9576 = (inp[8]) ? node9608 : node9577;
											assign node9577 = (inp[14]) ? node9593 : node9578;
												assign node9578 = (inp[2]) ? node9586 : node9579;
													assign node9579 = (inp[3]) ? node9581 : 4'b0101;
														assign node9581 = (inp[0]) ? 4'b0111 : node9582;
															assign node9582 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node9586 = (inp[15]) ? node9590 : node9587;
														assign node9587 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node9590 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node9593 = (inp[3]) ? node9601 : node9594;
													assign node9594 = (inp[15]) ? node9596 : 4'b0100;
														assign node9596 = (inp[5]) ? node9598 : 4'b0110;
															assign node9598 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node9601 = (inp[15]) ? node9605 : node9602;
														assign node9602 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node9605 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node9608 = (inp[2]) ? node9616 : node9609;
												assign node9609 = (inp[14]) ? node9613 : node9610;
													assign node9610 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node9613 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node9616 = (inp[15]) ? node9618 : 4'b1001;
													assign node9618 = (inp[3]) ? 4'b1001 : node9619;
														assign node9619 = (inp[0]) ? 4'b1011 : node9620;
															assign node9620 = (inp[5]) ? 4'b1011 : 4'b1001;
										assign node9625 = (inp[8]) ? node9645 : node9626;
											assign node9626 = (inp[14]) ? node9634 : node9627;
												assign node9627 = (inp[2]) ? node9631 : node9628;
													assign node9628 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node9631 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node9634 = (inp[0]) ? node9640 : node9635;
													assign node9635 = (inp[15]) ? node9637 : 4'b1001;
														assign node9637 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node9640 = (inp[5]) ? node9642 : 4'b1001;
														assign node9642 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node9645 = (inp[14]) ? node9655 : node9646;
												assign node9646 = (inp[2]) ? node9652 : node9647;
													assign node9647 = (inp[5]) ? node9649 : 4'b1011;
														assign node9649 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node9652 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node9655 = (inp[2]) ? node9661 : node9656;
													assign node9656 = (inp[0]) ? node9658 : 4'b1000;
														assign node9658 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node9661 = (inp[15]) ? 4'b1010 : node9662;
														assign node9662 = (inp[5]) ? 4'b1010 : node9663;
															assign node9663 = (inp[3]) ? 4'b1010 : 4'b1000;
								assign node9668 = (inp[1]) ? node9746 : node9669;
									assign node9669 = (inp[15]) ? node9725 : node9670;
										assign node9670 = (inp[0]) ? node9698 : node9671;
											assign node9671 = (inp[3]) ? node9689 : node9672;
												assign node9672 = (inp[5]) ? node9684 : node9673;
													assign node9673 = (inp[8]) ? node9679 : node9674;
														assign node9674 = (inp[14]) ? 4'b1010 : node9675;
															assign node9675 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node9679 = (inp[14]) ? 4'b1011 : node9680;
															assign node9680 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node9684 = (inp[7]) ? node9686 : 4'b1001;
														assign node9686 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node9689 = (inp[14]) ? node9691 : 4'b1000;
													assign node9691 = (inp[5]) ? 4'b1001 : node9692;
														assign node9692 = (inp[7]) ? 4'b1000 : node9693;
															assign node9693 = (inp[8]) ? 4'b1001 : 4'b1000;
											assign node9698 = (inp[3]) ? node9712 : node9699;
												assign node9699 = (inp[5]) ? node9707 : node9700;
													assign node9700 = (inp[8]) ? 4'b1001 : node9701;
														assign node9701 = (inp[7]) ? node9703 : 4'b1000;
															assign node9703 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node9707 = (inp[2]) ? node9709 : 4'b1011;
														assign node9709 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node9712 = (inp[14]) ? 4'b1011 : node9713;
													assign node9713 = (inp[7]) ? node9719 : node9714;
														assign node9714 = (inp[8]) ? 4'b1011 : node9715;
															assign node9715 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node9719 = (inp[8]) ? node9721 : 4'b1010;
															assign node9721 = (inp[2]) ? 4'b1010 : 4'b1011;
										assign node9725 = (inp[0]) ? node9735 : node9726;
											assign node9726 = (inp[7]) ? node9732 : node9727;
												assign node9727 = (inp[2]) ? node9729 : 4'b1011;
													assign node9729 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node9732 = (inp[14]) ? 4'b1010 : 4'b1000;
											assign node9735 = (inp[7]) ? node9741 : node9736;
												assign node9736 = (inp[3]) ? 4'b1000 : node9737;
													assign node9737 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node9741 = (inp[2]) ? 4'b1001 : node9742;
													assign node9742 = (inp[3]) ? 4'b1000 : 4'b1001;
									assign node9746 = (inp[8]) ? node9782 : node9747;
										assign node9747 = (inp[7]) ? node9767 : node9748;
											assign node9748 = (inp[14]) ? node9760 : node9749;
												assign node9749 = (inp[2]) ? node9757 : node9750;
													assign node9750 = (inp[15]) ? 4'b1001 : node9751;
														assign node9751 = (inp[5]) ? node9753 : 4'b1011;
															assign node9753 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node9757 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node9760 = (inp[5]) ? node9762 : 4'b1010;
													assign node9762 = (inp[15]) ? 4'b1000 : node9763;
														assign node9763 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node9767 = (inp[2]) ? node9773 : node9768;
												assign node9768 = (inp[14]) ? 4'b0001 : node9769;
													assign node9769 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node9773 = (inp[0]) ? node9777 : node9774;
													assign node9774 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node9777 = (inp[3]) ? node9779 : 4'b0011;
														assign node9779 = (inp[5]) ? 4'b0011 : 4'b0001;
										assign node9782 = (inp[7]) ? node9806 : node9783;
											assign node9783 = (inp[14]) ? node9793 : node9784;
												assign node9784 = (inp[2]) ? node9786 : 4'b1000;
													assign node9786 = (inp[0]) ? 4'b0011 : node9787;
														assign node9787 = (inp[5]) ? 4'b0011 : node9788;
															assign node9788 = (inp[3]) ? 4'b0001 : 4'b0001;
												assign node9793 = (inp[5]) ? node9801 : node9794;
													assign node9794 = (inp[3]) ? node9796 : 4'b0001;
														assign node9796 = (inp[2]) ? 4'b0001 : node9797;
															assign node9797 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node9801 = (inp[15]) ? node9803 : 4'b0011;
														assign node9803 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node9806 = (inp[2]) ? node9822 : node9807;
												assign node9807 = (inp[14]) ? node9817 : node9808;
													assign node9808 = (inp[0]) ? 4'b0001 : node9809;
														assign node9809 = (inp[15]) ? node9813 : node9810;
															assign node9810 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node9813 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node9817 = (inp[5]) ? node9819 : 4'b0010;
														assign node9819 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node9822 = (inp[14]) ? node9830 : node9823;
													assign node9823 = (inp[5]) ? node9825 : 4'b0000;
														assign node9825 = (inp[15]) ? node9827 : 4'b0010;
															assign node9827 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node9830 = (inp[15]) ? 4'b0010 : node9831;
														assign node9831 = (inp[5]) ? 4'b0000 : node9832;
															assign node9832 = (inp[0]) ? 4'b0000 : 4'b0010;
					assign node9837 = (inp[10]) ? node10493 : node9838;
						assign node9838 = (inp[6]) ? node10154 : node9839;
							assign node9839 = (inp[11]) ? node10003 : node9840;
								assign node9840 = (inp[1]) ? node9932 : node9841;
									assign node9841 = (inp[5]) ? node9891 : node9842;
										assign node9842 = (inp[7]) ? node9860 : node9843;
											assign node9843 = (inp[8]) ? node9849 : node9844;
												assign node9844 = (inp[14]) ? 4'b1100 : node9845;
													assign node9845 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node9849 = (inp[3]) ? 4'b1111 : node9850;
													assign node9850 = (inp[2]) ? node9854 : node9851;
														assign node9851 = (inp[0]) ? 4'b1110 : 4'b1101;
														assign node9854 = (inp[0]) ? 4'b1101 : node9855;
															assign node9855 = (inp[14]) ? 4'b1111 : 4'b1101;
											assign node9860 = (inp[8]) ? node9878 : node9861;
												assign node9861 = (inp[2]) ? node9869 : node9862;
													assign node9862 = (inp[3]) ? node9866 : node9863;
														assign node9863 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node9866 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node9869 = (inp[14]) ? node9875 : node9870;
														assign node9870 = (inp[3]) ? 4'b1111 : node9871;
															assign node9871 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node9875 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node9878 = (inp[0]) ? node9884 : node9879;
													assign node9879 = (inp[15]) ? 4'b1110 : node9880;
														assign node9880 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node9884 = (inp[3]) ? node9888 : node9885;
														assign node9885 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node9888 = (inp[14]) ? 4'b1100 : 4'b1101;
										assign node9891 = (inp[8]) ? node9915 : node9892;
											assign node9892 = (inp[7]) ? node9908 : node9893;
												assign node9893 = (inp[2]) ? node9903 : node9894;
													assign node9894 = (inp[3]) ? node9898 : node9895;
														assign node9895 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node9898 = (inp[15]) ? 4'b1100 : node9899;
															assign node9899 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node9903 = (inp[0]) ? 4'b1110 : node9904;
														assign node9904 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node9908 = (inp[0]) ? node9910 : 4'b1111;
													assign node9910 = (inp[2]) ? 4'b1101 : node9911;
														assign node9911 = (inp[3]) ? 4'b1110 : 4'b1100;
											assign node9915 = (inp[7]) ? node9925 : node9916;
												assign node9916 = (inp[2]) ? node9920 : node9917;
													assign node9917 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node9920 = (inp[15]) ? 4'b1111 : node9921;
														assign node9921 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node9925 = (inp[2]) ? node9927 : 4'b1101;
													assign node9927 = (inp[0]) ? node9929 : 4'b1100;
														assign node9929 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node9932 = (inp[7]) ? node9966 : node9933;
										assign node9933 = (inp[8]) ? node9953 : node9934;
											assign node9934 = (inp[2]) ? node9944 : node9935;
												assign node9935 = (inp[14]) ? 4'b1100 : node9936;
													assign node9936 = (inp[3]) ? 4'b1101 : node9937;
														assign node9937 = (inp[0]) ? 4'b1111 : node9938;
															assign node9938 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node9944 = (inp[3]) ? node9946 : 4'b1100;
													assign node9946 = (inp[0]) ? node9950 : node9947;
														assign node9947 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node9950 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node9953 = (inp[14]) ? node9959 : node9954;
												assign node9954 = (inp[2]) ? 4'b0111 : node9955;
													assign node9955 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node9959 = (inp[3]) ? 4'b0111 : node9960;
													assign node9960 = (inp[15]) ? 4'b0101 : node9961;
														assign node9961 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node9966 = (inp[8]) ? node9986 : node9967;
											assign node9967 = (inp[2]) ? node9979 : node9968;
												assign node9968 = (inp[14]) ? node9974 : node9969;
													assign node9969 = (inp[0]) ? 4'b1100 : node9970;
														assign node9970 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node9974 = (inp[3]) ? node9976 : 4'b0101;
														assign node9976 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node9979 = (inp[5]) ? 4'b0101 : node9980;
													assign node9980 = (inp[0]) ? node9982 : 4'b0111;
														assign node9982 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node9986 = (inp[5]) ? node9998 : node9987;
												assign node9987 = (inp[14]) ? node9993 : node9988;
													assign node9988 = (inp[2]) ? 4'b0110 : node9989;
														assign node9989 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node9993 = (inp[15]) ? node9995 : 4'b0110;
														assign node9995 = (inp[2]) ? 4'b0110 : 4'b0100;
												assign node9998 = (inp[2]) ? 4'b0100 : node9999;
													assign node9999 = (inp[14]) ? 4'b0100 : 4'b0101;
								assign node10003 = (inp[1]) ? node10071 : node10004;
									assign node10004 = (inp[0]) ? node10036 : node10005;
										assign node10005 = (inp[15]) ? node10015 : node10006;
											assign node10006 = (inp[5]) ? 4'b0101 : node10007;
												assign node10007 = (inp[7]) ? 4'b0100 : node10008;
													assign node10008 = (inp[8]) ? 4'b0101 : node10009;
														assign node10009 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node10015 = (inp[3]) ? node10027 : node10016;
												assign node10016 = (inp[5]) ? node10022 : node10017;
													assign node10017 = (inp[8]) ? node10019 : 4'b0100;
														assign node10019 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node10022 = (inp[2]) ? 4'b0111 : node10023;
														assign node10023 = (inp[14]) ? 4'b0111 : 4'b0110;
												assign node10027 = (inp[8]) ? node10029 : 4'b0111;
													assign node10029 = (inp[7]) ? 4'b0110 : node10030;
														assign node10030 = (inp[2]) ? 4'b0111 : node10031;
															assign node10031 = (inp[14]) ? 4'b0111 : 4'b0110;
										assign node10036 = (inp[15]) ? node10052 : node10037;
											assign node10037 = (inp[5]) ? node10047 : node10038;
												assign node10038 = (inp[3]) ? 4'b0110 : node10039;
													assign node10039 = (inp[2]) ? node10041 : 4'b0101;
														assign node10041 = (inp[8]) ? node10043 : 4'b0100;
															assign node10043 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node10047 = (inp[7]) ? 4'b0111 : node10048;
													assign node10048 = (inp[3]) ? 4'b0110 : 4'b0111;
											assign node10052 = (inp[5]) ? node10060 : node10053;
												assign node10053 = (inp[3]) ? node10057 : node10054;
													assign node10054 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node10057 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node10060 = (inp[2]) ? node10066 : node10061;
													assign node10061 = (inp[8]) ? 4'b0100 : node10062;
														assign node10062 = (inp[3]) ? 4'b0100 : 4'b0101;
													assign node10066 = (inp[7]) ? 4'b0101 : node10067;
														assign node10067 = (inp[8]) ? 4'b0101 : 4'b0100;
									assign node10071 = (inp[7]) ? node10117 : node10072;
										assign node10072 = (inp[8]) ? node10096 : node10073;
											assign node10073 = (inp[2]) ? node10087 : node10074;
												assign node10074 = (inp[14]) ? node10080 : node10075;
													assign node10075 = (inp[5]) ? 4'b0101 : node10076;
														assign node10076 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node10080 = (inp[5]) ? node10082 : 4'b0110;
														assign node10082 = (inp[15]) ? 4'b0100 : node10083;
															assign node10083 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node10087 = (inp[14]) ? node10089 : 4'b0110;
													assign node10089 = (inp[5]) ? node10091 : 4'b0100;
														assign node10091 = (inp[15]) ? 4'b0110 : node10092;
															assign node10092 = (inp[0]) ? 4'b0110 : 4'b0100;
											assign node10096 = (inp[14]) ? node10104 : node10097;
												assign node10097 = (inp[2]) ? node10101 : node10098;
													assign node10098 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node10101 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node10104 = (inp[0]) ? node10112 : node10105;
													assign node10105 = (inp[3]) ? 4'b1011 : node10106;
														assign node10106 = (inp[2]) ? node10108 : 4'b1011;
															assign node10108 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node10112 = (inp[3]) ? node10114 : 4'b1001;
														assign node10114 = (inp[15]) ? 4'b1001 : 4'b1011;
										assign node10117 = (inp[8]) ? node10133 : node10118;
											assign node10118 = (inp[14]) ? node10126 : node10119;
												assign node10119 = (inp[2]) ? node10123 : node10120;
													assign node10120 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node10123 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node10126 = (inp[15]) ? node10130 : node10127;
													assign node10127 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node10130 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node10133 = (inp[2]) ? node10139 : node10134;
												assign node10134 = (inp[5]) ? node10136 : 4'b1011;
													assign node10136 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node10139 = (inp[5]) ? node10147 : node10140;
													assign node10140 = (inp[14]) ? 4'b1010 : node10141;
														assign node10141 = (inp[15]) ? node10143 : 4'b1010;
															assign node10143 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node10147 = (inp[3]) ? node10149 : 4'b1010;
														assign node10149 = (inp[14]) ? 4'b1000 : node10150;
															assign node10150 = (inp[15]) ? 4'b1000 : 4'b1010;
							assign node10154 = (inp[11]) ? node10316 : node10155;
								assign node10155 = (inp[1]) ? node10231 : node10156;
									assign node10156 = (inp[0]) ? node10192 : node10157;
										assign node10157 = (inp[15]) ? node10173 : node10158;
											assign node10158 = (inp[3]) ? node10166 : node10159;
												assign node10159 = (inp[5]) ? node10163 : node10160;
													assign node10160 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node10163 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node10166 = (inp[7]) ? 4'b0100 : node10167;
													assign node10167 = (inp[8]) ? 4'b0101 : node10168;
														assign node10168 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node10173 = (inp[8]) ? node10183 : node10174;
												assign node10174 = (inp[3]) ? node10178 : node10175;
													assign node10175 = (inp[2]) ? 4'b0100 : 4'b0110;
													assign node10178 = (inp[7]) ? node10180 : 4'b0110;
														assign node10180 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node10183 = (inp[5]) ? node10187 : node10184;
													assign node10184 = (inp[14]) ? 4'b0101 : 4'b0111;
													assign node10187 = (inp[14]) ? 4'b0110 : node10188;
														assign node10188 = (inp[2]) ? 4'b0110 : 4'b0111;
										assign node10192 = (inp[15]) ? node10210 : node10193;
											assign node10193 = (inp[3]) ? node10201 : node10194;
												assign node10194 = (inp[5]) ? 4'b0110 : node10195;
													assign node10195 = (inp[14]) ? 4'b0101 : node10196;
														assign node10196 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node10201 = (inp[5]) ? node10203 : 4'b0111;
													assign node10203 = (inp[8]) ? node10205 : 4'b0110;
														assign node10205 = (inp[7]) ? node10207 : 4'b0111;
															assign node10207 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node10210 = (inp[3]) ? node10220 : node10211;
												assign node10211 = (inp[5]) ? node10213 : 4'b0111;
													assign node10213 = (inp[2]) ? 4'b0101 : node10214;
														assign node10214 = (inp[14]) ? 4'b0100 : node10215;
															assign node10215 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node10220 = (inp[8]) ? node10224 : node10221;
													assign node10221 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node10224 = (inp[7]) ? 4'b0100 : node10225;
														assign node10225 = (inp[2]) ? 4'b0101 : node10226;
															assign node10226 = (inp[14]) ? 4'b0101 : 4'b0100;
									assign node10231 = (inp[2]) ? node10281 : node10232;
										assign node10232 = (inp[14]) ? node10262 : node10233;
											assign node10233 = (inp[7]) ? node10247 : node10234;
												assign node10234 = (inp[8]) ? node10242 : node10235;
													assign node10235 = (inp[15]) ? node10237 : 4'b0111;
														assign node10237 = (inp[0]) ? 4'b0101 : node10238;
															assign node10238 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node10242 = (inp[5]) ? node10244 : 4'b0110;
														assign node10244 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node10247 = (inp[8]) ? node10259 : node10248;
													assign node10248 = (inp[15]) ? node10254 : node10249;
														assign node10249 = (inp[0]) ? node10251 : 4'b0100;
															assign node10251 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node10254 = (inp[0]) ? node10256 : 4'b0110;
															assign node10256 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node10259 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node10262 = (inp[7]) ? node10270 : node10263;
												assign node10263 = (inp[8]) ? node10265 : 4'b0110;
													assign node10265 = (inp[15]) ? 4'b1011 : node10266;
														assign node10266 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node10270 = (inp[8]) ? node10276 : node10271;
													assign node10271 = (inp[15]) ? 4'b1001 : node10272;
														assign node10272 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node10276 = (inp[15]) ? 4'b1000 : node10277;
														assign node10277 = (inp[5]) ? 4'b1010 : 4'b1000;
										assign node10281 = (inp[7]) ? node10299 : node10282;
											assign node10282 = (inp[8]) ? node10286 : node10283;
												assign node10283 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node10286 = (inp[15]) ? node10294 : node10287;
													assign node10287 = (inp[0]) ? node10291 : node10288;
														assign node10288 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node10291 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node10294 = (inp[0]) ? 4'b1001 : node10295;
														assign node10295 = (inp[5]) ? 4'b1011 : 4'b1001;
											assign node10299 = (inp[8]) ? node10309 : node10300;
												assign node10300 = (inp[15]) ? node10302 : 4'b1011;
													assign node10302 = (inp[0]) ? node10306 : node10303;
														assign node10303 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node10306 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node10309 = (inp[0]) ? 4'b1000 : node10310;
													assign node10310 = (inp[3]) ? 4'b1010 : node10311;
														assign node10311 = (inp[14]) ? 4'b1010 : 4'b1000;
								assign node10316 = (inp[1]) ? node10396 : node10317;
									assign node10317 = (inp[15]) ? node10359 : node10318;
										assign node10318 = (inp[0]) ? node10340 : node10319;
											assign node10319 = (inp[5]) ? node10325 : node10320;
												assign node10320 = (inp[3]) ? node10322 : 4'b1011;
													assign node10322 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node10325 = (inp[2]) ? node10335 : node10326;
													assign node10326 = (inp[7]) ? 4'b1001 : node10327;
														assign node10327 = (inp[8]) ? node10331 : node10328;
															assign node10328 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node10331 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node10335 = (inp[7]) ? node10337 : 4'b1001;
														assign node10337 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node10340 = (inp[5]) ? node10348 : node10341;
												assign node10341 = (inp[3]) ? 4'b1010 : node10342;
													assign node10342 = (inp[8]) ? node10344 : 4'b1001;
														assign node10344 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node10348 = (inp[8]) ? node10354 : node10349;
													assign node10349 = (inp[3]) ? node10351 : 4'b1010;
														assign node10351 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node10354 = (inp[7]) ? node10356 : 4'b1011;
														assign node10356 = (inp[3]) ? 4'b1010 : 4'b1011;
										assign node10359 = (inp[0]) ? node10383 : node10360;
											assign node10360 = (inp[3]) ? node10368 : node10361;
												assign node10361 = (inp[5]) ? 4'b1011 : node10362;
													assign node10362 = (inp[14]) ? node10364 : 4'b1000;
														assign node10364 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node10368 = (inp[2]) ? node10376 : node10369;
													assign node10369 = (inp[7]) ? node10371 : 4'b1011;
														assign node10371 = (inp[8]) ? node10373 : 4'b1010;
															assign node10373 = (inp[5]) ? 4'b1010 : 4'b1011;
													assign node10376 = (inp[5]) ? 4'b1010 : node10377;
														assign node10377 = (inp[14]) ? 4'b1010 : node10378;
															assign node10378 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node10383 = (inp[5]) ? node10391 : node10384;
												assign node10384 = (inp[3]) ? node10388 : node10385;
													assign node10385 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node10388 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node10391 = (inp[14]) ? node10393 : 4'b1000;
													assign node10393 = (inp[3]) ? 4'b1000 : 4'b1001;
									assign node10396 = (inp[7]) ? node10450 : node10397;
										assign node10397 = (inp[8]) ? node10425 : node10398;
											assign node10398 = (inp[14]) ? node10412 : node10399;
												assign node10399 = (inp[2]) ? node10405 : node10400;
													assign node10400 = (inp[0]) ? node10402 : 4'b1011;
														assign node10402 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node10405 = (inp[3]) ? node10407 : 4'b1010;
														assign node10407 = (inp[15]) ? 4'b1010 : node10408;
															assign node10408 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node10412 = (inp[2]) ? node10420 : node10413;
													assign node10413 = (inp[0]) ? node10415 : 4'b1000;
														assign node10415 = (inp[15]) ? node10417 : 4'b1010;
															assign node10417 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node10420 = (inp[5]) ? 4'b1010 : node10421;
														assign node10421 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node10425 = (inp[14]) ? node10441 : node10426;
												assign node10426 = (inp[2]) ? node10436 : node10427;
													assign node10427 = (inp[15]) ? 4'b1010 : node10428;
														assign node10428 = (inp[5]) ? node10432 : node10429;
															assign node10429 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node10432 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node10436 = (inp[0]) ? node10438 : 4'b0001;
														assign node10438 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node10441 = (inp[2]) ? 4'b0001 : node10442;
													assign node10442 = (inp[5]) ? 4'b0011 : node10443;
														assign node10443 = (inp[0]) ? 4'b0001 : node10444;
															assign node10444 = (inp[3]) ? 4'b0001 : 4'b0001;
										assign node10450 = (inp[8]) ? node10472 : node10451;
											assign node10451 = (inp[2]) ? node10461 : node10452;
												assign node10452 = (inp[14]) ? 4'b0001 : node10453;
													assign node10453 = (inp[0]) ? 4'b1000 : node10454;
														assign node10454 = (inp[15]) ? 4'b1010 : node10455;
															assign node10455 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node10461 = (inp[15]) ? node10463 : 4'b0011;
													assign node10463 = (inp[3]) ? node10469 : node10464;
														assign node10464 = (inp[0]) ? node10466 : 4'b0001;
															assign node10466 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node10469 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node10472 = (inp[2]) ? node10484 : node10473;
												assign node10473 = (inp[14]) ? node10481 : node10474;
													assign node10474 = (inp[0]) ? 4'b0011 : node10475;
														assign node10475 = (inp[15]) ? 4'b0001 : node10476;
															assign node10476 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node10481 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node10484 = (inp[5]) ? node10486 : 4'b0010;
													assign node10486 = (inp[3]) ? node10488 : 4'b0010;
														assign node10488 = (inp[15]) ? node10490 : 4'b0000;
															assign node10490 = (inp[0]) ? 4'b0000 : 4'b0010;
						assign node10493 = (inp[0]) ? node10859 : node10494;
							assign node10494 = (inp[15]) ? node10678 : node10495;
								assign node10495 = (inp[5]) ? node10591 : node10496;
									assign node10496 = (inp[3]) ? node10536 : node10497;
										assign node10497 = (inp[2]) ? node10519 : node10498;
											assign node10498 = (inp[8]) ? node10512 : node10499;
												assign node10499 = (inp[11]) ? node10507 : node10500;
													assign node10500 = (inp[6]) ? 4'b0011 : node10501;
														assign node10501 = (inp[1]) ? node10503 : 4'b1010;
															assign node10503 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node10507 = (inp[6]) ? node10509 : 4'b0011;
														assign node10509 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node10512 = (inp[6]) ? node10516 : node10513;
													assign node10513 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node10516 = (inp[14]) ? 4'b0011 : 4'b0010;
											assign node10519 = (inp[6]) ? node10531 : node10520;
												assign node10520 = (inp[11]) ? node10522 : 4'b1011;
													assign node10522 = (inp[7]) ? node10526 : node10523;
														assign node10523 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node10526 = (inp[1]) ? node10528 : 4'b0011;
															assign node10528 = (inp[14]) ? 4'b1011 : 4'b1010;
												assign node10531 = (inp[14]) ? 4'b0010 : node10532;
													assign node10532 = (inp[11]) ? 4'b1010 : 4'b0010;
										assign node10536 = (inp[14]) ? node10564 : node10537;
											assign node10537 = (inp[1]) ? node10549 : node10538;
												assign node10538 = (inp[7]) ? node10542 : node10539;
													assign node10539 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node10542 = (inp[2]) ? node10546 : node10543;
														assign node10543 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node10546 = (inp[6]) ? 4'b1001 : 4'b0001;
												assign node10549 = (inp[7]) ? node10557 : node10550;
													assign node10550 = (inp[2]) ? 4'b1000 : node10551;
														assign node10551 = (inp[8]) ? node10553 : 4'b0001;
															assign node10553 = (inp[6]) ? 4'b0000 : 4'b0000;
													assign node10557 = (inp[11]) ? node10559 : 4'b1001;
														assign node10559 = (inp[8]) ? 4'b1000 : node10560;
															assign node10560 = (inp[6]) ? 4'b1000 : 4'b1001;
											assign node10564 = (inp[2]) ? node10580 : node10565;
												assign node10565 = (inp[11]) ? node10577 : node10566;
													assign node10566 = (inp[7]) ? node10574 : node10567;
														assign node10567 = (inp[1]) ? node10571 : node10568;
															assign node10568 = (inp[6]) ? 4'b0001 : 4'b1001;
															assign node10571 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node10574 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node10577 = (inp[1]) ? 4'b0001 : 4'b1000;
												assign node10580 = (inp[11]) ? node10584 : node10581;
													assign node10581 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node10584 = (inp[1]) ? 4'b0001 : node10585;
														assign node10585 = (inp[8]) ? node10587 : 4'b0000;
															assign node10587 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node10591 = (inp[2]) ? node10631 : node10592;
										assign node10592 = (inp[11]) ? node10612 : node10593;
											assign node10593 = (inp[7]) ? node10603 : node10594;
												assign node10594 = (inp[6]) ? node10600 : node10595;
													assign node10595 = (inp[8]) ? 4'b1000 : node10596;
														assign node10596 = (inp[3]) ? 4'b1000 : 4'b1001;
													assign node10600 = (inp[3]) ? 4'b0001 : 4'b1001;
												assign node10603 = (inp[3]) ? node10605 : 4'b0001;
													assign node10605 = (inp[6]) ? node10607 : 4'b1001;
														assign node10607 = (inp[8]) ? node10609 : 4'b0000;
															assign node10609 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node10612 = (inp[6]) ? node10626 : node10613;
												assign node10613 = (inp[7]) ? node10615 : 4'b0000;
													assign node10615 = (inp[3]) ? node10621 : node10616;
														assign node10616 = (inp[1]) ? 4'b1001 : node10617;
															assign node10617 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node10621 = (inp[14]) ? node10623 : 4'b0000;
															assign node10623 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node10626 = (inp[8]) ? node10628 : 4'b1000;
													assign node10628 = (inp[1]) ? 4'b0000 : 4'b1001;
										assign node10631 = (inp[1]) ? node10651 : node10632;
											assign node10632 = (inp[6]) ? node10642 : node10633;
												assign node10633 = (inp[11]) ? 4'b0000 : node10634;
													assign node10634 = (inp[14]) ? node10636 : 4'b1000;
														assign node10636 = (inp[3]) ? 4'b1000 : node10637;
															assign node10637 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node10642 = (inp[11]) ? node10644 : 4'b0000;
													assign node10644 = (inp[14]) ? node10646 : 4'b1001;
														assign node10646 = (inp[7]) ? node10648 : 4'b1000;
															assign node10648 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node10651 = (inp[3]) ? node10667 : node10652;
												assign node10652 = (inp[6]) ? node10656 : node10653;
													assign node10653 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node10656 = (inp[8]) ? node10660 : node10657;
														assign node10657 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node10660 = (inp[7]) ? node10664 : node10661;
															assign node10661 = (inp[14]) ? 4'b1001 : 4'b0001;
															assign node10664 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node10667 = (inp[8]) ? node10671 : node10668;
													assign node10668 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node10671 = (inp[7]) ? node10673 : 4'b0001;
														assign node10673 = (inp[6]) ? node10675 : 4'b0000;
															assign node10675 = (inp[11]) ? 4'b0000 : 4'b1000;
								assign node10678 = (inp[3]) ? node10766 : node10679;
									assign node10679 = (inp[5]) ? node10723 : node10680;
										assign node10680 = (inp[7]) ? node10696 : node10681;
											assign node10681 = (inp[8]) ? node10687 : node10682;
												assign node10682 = (inp[11]) ? 4'b0000 : node10683;
													assign node10683 = (inp[6]) ? 4'b0000 : 4'b1000;
												assign node10687 = (inp[1]) ? node10689 : 4'b0001;
													assign node10689 = (inp[6]) ? node10691 : 4'b0000;
														assign node10691 = (inp[14]) ? 4'b1001 : node10692;
															assign node10692 = (inp[2]) ? 4'b1001 : 4'b0000;
											assign node10696 = (inp[11]) ? node10710 : node10697;
												assign node10697 = (inp[6]) ? node10705 : node10698;
													assign node10698 = (inp[14]) ? 4'b0000 : node10699;
														assign node10699 = (inp[8]) ? node10701 : 4'b0001;
															assign node10701 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node10705 = (inp[2]) ? 4'b0001 : node10706;
														assign node10706 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node10710 = (inp[1]) ? node10716 : node10711;
													assign node10711 = (inp[6]) ? 4'b1000 : node10712;
														assign node10712 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node10716 = (inp[6]) ? node10718 : 4'b1001;
														assign node10718 = (inp[2]) ? 4'b0001 : node10719;
															assign node10719 = (inp[8]) ? 4'b0001 : 4'b0000;
										assign node10723 = (inp[7]) ? node10747 : node10724;
											assign node10724 = (inp[8]) ? node10736 : node10725;
												assign node10725 = (inp[14]) ? 4'b0010 : node10726;
													assign node10726 = (inp[2]) ? node10732 : node10727;
														assign node10727 = (inp[11]) ? 4'b0011 : node10728;
															assign node10728 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node10732 = (inp[1]) ? 4'b0010 : 4'b1010;
												assign node10736 = (inp[1]) ? node10742 : node10737;
													assign node10737 = (inp[11]) ? 4'b0011 : node10738;
														assign node10738 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node10742 = (inp[6]) ? 4'b0010 : node10743;
														assign node10743 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node10747 = (inp[8]) ? node10759 : node10748;
												assign node10748 = (inp[14]) ? node10752 : node10749;
													assign node10749 = (inp[11]) ? 4'b1010 : 4'b0011;
													assign node10752 = (inp[6]) ? node10754 : 4'b1011;
														assign node10754 = (inp[11]) ? 4'b0011 : node10755;
															assign node10755 = (inp[1]) ? 4'b1011 : 4'b0011;
												assign node10759 = (inp[6]) ? node10761 : 4'b1010;
													assign node10761 = (inp[11]) ? 4'b0010 : node10762;
														assign node10762 = (inp[1]) ? 4'b1010 : 4'b0010;
									assign node10766 = (inp[8]) ? node10814 : node10767;
										assign node10767 = (inp[7]) ? node10787 : node10768;
											assign node10768 = (inp[2]) ? node10780 : node10769;
												assign node10769 = (inp[14]) ? node10777 : node10770;
													assign node10770 = (inp[1]) ? node10772 : 4'b1011;
														assign node10772 = (inp[11]) ? 4'b0011 : node10773;
															assign node10773 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node10777 = (inp[11]) ? 4'b1010 : 4'b0010;
												assign node10780 = (inp[1]) ? 4'b0010 : node10781;
													assign node10781 = (inp[6]) ? node10783 : 4'b1010;
														assign node10783 = (inp[11]) ? 4'b1010 : 4'b0010;
											assign node10787 = (inp[14]) ? node10797 : node10788;
												assign node10788 = (inp[2]) ? node10794 : node10789;
													assign node10789 = (inp[1]) ? node10791 : 4'b0010;
														assign node10791 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node10794 = (inp[5]) ? 4'b0011 : 4'b1011;
												assign node10797 = (inp[1]) ? node10807 : node10798;
													assign node10798 = (inp[2]) ? 4'b1011 : node10799;
														assign node10799 = (inp[5]) ? node10803 : node10800;
															assign node10800 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node10803 = (inp[11]) ? 4'b1011 : 4'b0011;
													assign node10807 = (inp[6]) ? node10811 : node10808;
														assign node10808 = (inp[5]) ? 4'b1011 : 4'b0011;
														assign node10811 = (inp[11]) ? 4'b0011 : 4'b1011;
										assign node10814 = (inp[7]) ? node10832 : node10815;
											assign node10815 = (inp[14]) ? node10825 : node10816;
												assign node10816 = (inp[2]) ? 4'b1011 : node10817;
													assign node10817 = (inp[1]) ? node10819 : 4'b1010;
														assign node10819 = (inp[11]) ? 4'b1010 : node10820;
															assign node10820 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node10825 = (inp[2]) ? node10829 : node10826;
													assign node10826 = (inp[6]) ? 4'b1011 : 4'b0011;
													assign node10829 = (inp[6]) ? 4'b0011 : 4'b1011;
											assign node10832 = (inp[2]) ? node10844 : node10833;
												assign node10833 = (inp[14]) ? node10839 : node10834;
													assign node10834 = (inp[1]) ? node10836 : 4'b1011;
														assign node10836 = (inp[5]) ? 4'b1011 : 4'b0011;
													assign node10839 = (inp[5]) ? 4'b1010 : node10840;
														assign node10840 = (inp[11]) ? 4'b1010 : 4'b0010;
												assign node10844 = (inp[11]) ? node10852 : node10845;
													assign node10845 = (inp[14]) ? 4'b1010 : node10846;
														assign node10846 = (inp[1]) ? 4'b0010 : node10847;
															assign node10847 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node10852 = (inp[14]) ? 4'b0010 : node10853;
														assign node10853 = (inp[5]) ? node10855 : 4'b1010;
															assign node10855 = (inp[1]) ? 4'b0010 : 4'b0010;
							assign node10859 = (inp[15]) ? node11037 : node10860;
								assign node10860 = (inp[5]) ? node10940 : node10861;
									assign node10861 = (inp[3]) ? node10901 : node10862;
										assign node10862 = (inp[2]) ? node10886 : node10863;
											assign node10863 = (inp[14]) ? node10879 : node10864;
												assign node10864 = (inp[8]) ? node10870 : node10865;
													assign node10865 = (inp[6]) ? node10867 : 4'b0001;
														assign node10867 = (inp[11]) ? 4'b1001 : 4'b0001;
													assign node10870 = (inp[7]) ? node10876 : node10871;
														assign node10871 = (inp[11]) ? node10873 : 4'b1000;
															assign node10873 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node10876 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node10879 = (inp[8]) ? node10883 : node10880;
													assign node10880 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node10883 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node10886 = (inp[11]) ? node10892 : node10887;
												assign node10887 = (inp[14]) ? node10889 : 4'b0000;
													assign node10889 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node10892 = (inp[6]) ? node10896 : node10893;
													assign node10893 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node10896 = (inp[8]) ? node10898 : 4'b1000;
														assign node10898 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node10901 = (inp[8]) ? node10913 : node10902;
											assign node10902 = (inp[14]) ? node10910 : node10903;
												assign node10903 = (inp[1]) ? 4'b1011 : node10904;
													assign node10904 = (inp[11]) ? 4'b0010 : node10905;
														assign node10905 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node10910 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node10913 = (inp[7]) ? node10925 : node10914;
												assign node10914 = (inp[11]) ? node10916 : 4'b1011;
													assign node10916 = (inp[14]) ? node10920 : node10917;
														assign node10917 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node10920 = (inp[6]) ? 4'b1011 : node10921;
															assign node10921 = (inp[1]) ? 4'b1011 : 4'b0011;
												assign node10925 = (inp[2]) ? node10929 : node10926;
													assign node10926 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node10929 = (inp[14]) ? node10935 : node10930;
														assign node10930 = (inp[1]) ? 4'b0010 : node10931;
															assign node10931 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node10935 = (inp[11]) ? node10937 : 4'b1010;
															assign node10937 = (inp[6]) ? 4'b1010 : 4'b0010;
									assign node10940 = (inp[3]) ? node10992 : node10941;
										assign node10941 = (inp[7]) ? node10963 : node10942;
											assign node10942 = (inp[8]) ? node10958 : node10943;
												assign node10943 = (inp[1]) ? node10955 : node10944;
													assign node10944 = (inp[2]) ? node10950 : node10945;
														assign node10945 = (inp[14]) ? node10947 : 4'b1011;
															assign node10947 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node10950 = (inp[6]) ? node10952 : 4'b1010;
															assign node10952 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node10955 = (inp[11]) ? 4'b0010 : 4'b1010;
												assign node10958 = (inp[14]) ? 4'b1011 : node10959;
													assign node10959 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node10963 = (inp[8]) ? node10979 : node10964;
												assign node10964 = (inp[2]) ? node10972 : node10965;
													assign node10965 = (inp[1]) ? node10967 : 4'b1010;
														assign node10967 = (inp[11]) ? 4'b1011 : node10968;
															assign node10968 = (inp[6]) ? 4'b1011 : 4'b0011;
													assign node10972 = (inp[14]) ? 4'b1011 : node10973;
														assign node10973 = (inp[11]) ? node10975 : 4'b1011;
															assign node10975 = (inp[6]) ? 4'b0011 : 4'b0011;
												assign node10979 = (inp[2]) ? node10987 : node10980;
													assign node10980 = (inp[6]) ? node10984 : node10981;
														assign node10981 = (inp[1]) ? 4'b0011 : 4'b1011;
														assign node10984 = (inp[1]) ? 4'b1011 : 4'b0011;
													assign node10987 = (inp[14]) ? 4'b0010 : node10988;
														assign node10988 = (inp[1]) ? 4'b1010 : 4'b0010;
										assign node10992 = (inp[1]) ? node11018 : node10993;
											assign node10993 = (inp[7]) ? node11005 : node10994;
												assign node10994 = (inp[14]) ? node11000 : node10995;
													assign node10995 = (inp[6]) ? 4'b1011 : node10996;
														assign node10996 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node11000 = (inp[8]) ? node11002 : 4'b1010;
														assign node11002 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node11005 = (inp[11]) ? node11013 : node11006;
													assign node11006 = (inp[6]) ? node11008 : 4'b1010;
														assign node11008 = (inp[2]) ? 4'b0010 : node11009;
															assign node11009 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node11013 = (inp[6]) ? node11015 : 4'b0011;
														assign node11015 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node11018 = (inp[2]) ? node11028 : node11019;
												assign node11019 = (inp[11]) ? node11025 : node11020;
													assign node11020 = (inp[8]) ? 4'b0010 : node11021;
														assign node11021 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node11025 = (inp[6]) ? 4'b0011 : 4'b0010;
												assign node11028 = (inp[7]) ? node11034 : node11029;
													assign node11029 = (inp[8]) ? 4'b0011 : node11030;
														assign node11030 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node11034 = (inp[6]) ? 4'b1011 : 4'b0011;
								assign node11037 = (inp[3]) ? node11143 : node11038;
									assign node11038 = (inp[5]) ? node11096 : node11039;
										assign node11039 = (inp[7]) ? node11069 : node11040;
											assign node11040 = (inp[6]) ? node11054 : node11041;
												assign node11041 = (inp[14]) ? node11049 : node11042;
													assign node11042 = (inp[11]) ? 4'b0011 : node11043;
														assign node11043 = (inp[2]) ? node11045 : 4'b1010;
															assign node11045 = (inp[1]) ? 4'b0011 : 4'b1010;
													assign node11049 = (inp[1]) ? node11051 : 4'b1011;
														assign node11051 = (inp[2]) ? 4'b1011 : 4'b0011;
												assign node11054 = (inp[8]) ? node11060 : node11055;
													assign node11055 = (inp[11]) ? 4'b1010 : node11056;
														assign node11056 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node11060 = (inp[14]) ? node11064 : node11061;
														assign node11061 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node11064 = (inp[1]) ? node11066 : 4'b0011;
															assign node11066 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node11069 = (inp[8]) ? node11085 : node11070;
												assign node11070 = (inp[2]) ? node11078 : node11071;
													assign node11071 = (inp[11]) ? node11075 : node11072;
														assign node11072 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node11075 = (inp[6]) ? 4'b1010 : 4'b0010;
													assign node11078 = (inp[6]) ? 4'b0011 : node11079;
														assign node11079 = (inp[11]) ? node11081 : 4'b1011;
															assign node11081 = (inp[1]) ? 4'b1011 : 4'b0011;
												assign node11085 = (inp[2]) ? node11089 : node11086;
													assign node11086 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node11089 = (inp[14]) ? 4'b0010 : node11090;
														assign node11090 = (inp[1]) ? 4'b1010 : node11091;
															assign node11091 = (inp[6]) ? 4'b0010 : 4'b0010;
										assign node11096 = (inp[8]) ? node11128 : node11097;
											assign node11097 = (inp[7]) ? node11109 : node11098;
												assign node11098 = (inp[6]) ? node11106 : node11099;
													assign node11099 = (inp[11]) ? 4'b0000 : node11100;
														assign node11100 = (inp[14]) ? 4'b1000 : node11101;
															assign node11101 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node11106 = (inp[11]) ? 4'b1000 : 4'b0000;
												assign node11109 = (inp[6]) ? node11117 : node11110;
													assign node11110 = (inp[11]) ? node11114 : node11111;
														assign node11111 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node11114 = (inp[14]) ? 4'b1001 : 4'b0001;
													assign node11117 = (inp[2]) ? node11123 : node11118;
														assign node11118 = (inp[14]) ? node11120 : 4'b1000;
															assign node11120 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node11123 = (inp[1]) ? node11125 : 4'b1001;
															assign node11125 = (inp[11]) ? 4'b0001 : 4'b1001;
											assign node11128 = (inp[7]) ? node11138 : node11129;
												assign node11129 = (inp[14]) ? 4'b1001 : node11130;
													assign node11130 = (inp[2]) ? 4'b0001 : node11131;
														assign node11131 = (inp[6]) ? 4'b0000 : node11132;
															assign node11132 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node11138 = (inp[11]) ? 4'b0000 : node11139;
													assign node11139 = (inp[14]) ? 4'b1000 : 4'b0000;
									assign node11143 = (inp[1]) ? node11199 : node11144;
										assign node11144 = (inp[11]) ? node11172 : node11145;
											assign node11145 = (inp[6]) ? node11163 : node11146;
												assign node11146 = (inp[5]) ? node11158 : node11147;
													assign node11147 = (inp[7]) ? node11151 : node11148;
														assign node11148 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node11151 = (inp[14]) ? node11155 : node11152;
															assign node11152 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node11155 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node11158 = (inp[14]) ? node11160 : 4'b1001;
														assign node11160 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node11163 = (inp[2]) ? node11165 : 4'b0000;
													assign node11165 = (inp[8]) ? node11169 : node11166;
														assign node11166 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node11169 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node11172 = (inp[6]) ? node11190 : node11173;
												assign node11173 = (inp[2]) ? node11185 : node11174;
													assign node11174 = (inp[5]) ? node11180 : node11175;
														assign node11175 = (inp[8]) ? node11177 : 4'b0000;
															assign node11177 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node11180 = (inp[8]) ? node11182 : 4'b0001;
															assign node11182 = (inp[14]) ? 4'b0000 : 4'b0000;
													assign node11185 = (inp[5]) ? node11187 : 4'b0001;
														assign node11187 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node11190 = (inp[7]) ? node11196 : node11191;
													assign node11191 = (inp[8]) ? 4'b1001 : node11192;
														assign node11192 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node11196 = (inp[8]) ? 4'b1000 : 4'b1001;
										assign node11199 = (inp[2]) ? node11233 : node11200;
											assign node11200 = (inp[11]) ? node11218 : node11201;
												assign node11201 = (inp[8]) ? node11209 : node11202;
													assign node11202 = (inp[6]) ? node11204 : 4'b1000;
														assign node11204 = (inp[14]) ? 4'b0000 : node11205;
															assign node11205 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node11209 = (inp[6]) ? node11213 : node11210;
														assign node11210 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node11213 = (inp[5]) ? 4'b1001 : node11214;
															assign node11214 = (inp[7]) ? 4'b1000 : 4'b0000;
												assign node11218 = (inp[7]) ? node11228 : node11219;
													assign node11219 = (inp[5]) ? 4'b1001 : node11220;
														assign node11220 = (inp[6]) ? node11224 : node11221;
															assign node11221 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node11224 = (inp[14]) ? 4'b1000 : 4'b1000;
													assign node11228 = (inp[6]) ? 4'b0001 : node11229;
														assign node11229 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node11233 = (inp[5]) ? node11243 : node11234;
												assign node11234 = (inp[8]) ? node11238 : node11235;
													assign node11235 = (inp[7]) ? 4'b0001 : 4'b1000;
													assign node11238 = (inp[7]) ? node11240 : 4'b0001;
														assign node11240 = (inp[6]) ? 4'b0000 : 4'b1000;
												assign node11243 = (inp[11]) ? 4'b0001 : node11244;
													assign node11244 = (inp[6]) ? node11250 : node11245;
														assign node11245 = (inp[7]) ? node11247 : 4'b0001;
															assign node11247 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node11250 = (inp[14]) ? 4'b1001 : 4'b0000;
		assign node11254 = (inp[10]) ? node16684 : node11255;
			assign node11255 = (inp[4]) ? node13893 : node11256;
				assign node11256 = (inp[9]) ? node12562 : node11257;
					assign node11257 = (inp[12]) ? node11885 : node11258;
						assign node11258 = (inp[7]) ? node11578 : node11259;
							assign node11259 = (inp[8]) ? node11433 : node11260;
								assign node11260 = (inp[2]) ? node11350 : node11261;
									assign node11261 = (inp[14]) ? node11315 : node11262;
										assign node11262 = (inp[6]) ? node11296 : node11263;
											assign node11263 = (inp[15]) ? node11275 : node11264;
												assign node11264 = (inp[3]) ? node11270 : node11265;
													assign node11265 = (inp[11]) ? node11267 : 4'b1101;
														assign node11267 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node11270 = (inp[11]) ? 4'b0101 : node11271;
														assign node11271 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node11275 = (inp[0]) ? node11285 : node11276;
													assign node11276 = (inp[5]) ? node11282 : node11277;
														assign node11277 = (inp[11]) ? 4'b1101 : node11278;
															assign node11278 = (inp[1]) ? 4'b0101 : 4'b1101;
														assign node11282 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node11285 = (inp[5]) ? node11293 : node11286;
														assign node11286 = (inp[11]) ? node11290 : node11287;
															assign node11287 = (inp[1]) ? 4'b0111 : 4'b1111;
															assign node11290 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node11293 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node11296 = (inp[3]) ? node11304 : node11297;
												assign node11297 = (inp[1]) ? node11301 : node11298;
													assign node11298 = (inp[11]) ? 4'b1111 : 4'b0111;
													assign node11301 = (inp[0]) ? 4'b1111 : 4'b0101;
												assign node11304 = (inp[15]) ? node11306 : 4'b1111;
													assign node11306 = (inp[0]) ? node11310 : node11307;
														assign node11307 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node11310 = (inp[5]) ? 4'b1101 : node11311;
															assign node11311 = (inp[11]) ? 4'b1111 : 4'b0111;
										assign node11315 = (inp[0]) ? node11331 : node11316;
											assign node11316 = (inp[1]) ? node11324 : node11317;
												assign node11317 = (inp[5]) ? node11319 : 4'b0100;
													assign node11319 = (inp[3]) ? 4'b1110 : node11320;
														assign node11320 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node11324 = (inp[3]) ? 4'b1100 : node11325;
													assign node11325 = (inp[11]) ? 4'b0100 : node11326;
														assign node11326 = (inp[6]) ? 4'b1100 : 4'b0100;
											assign node11331 = (inp[11]) ? node11339 : node11332;
												assign node11332 = (inp[3]) ? 4'b0110 : node11333;
													assign node11333 = (inp[6]) ? node11335 : 4'b0110;
														assign node11335 = (inp[1]) ? 4'b1110 : 4'b0110;
												assign node11339 = (inp[1]) ? node11347 : node11340;
													assign node11340 = (inp[6]) ? node11344 : node11341;
														assign node11341 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node11344 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node11347 = (inp[6]) ? 4'b0110 : 4'b1110;
									assign node11350 = (inp[1]) ? node11396 : node11351;
										assign node11351 = (inp[0]) ? node11377 : node11352;
											assign node11352 = (inp[15]) ? node11362 : node11353;
												assign node11353 = (inp[14]) ? node11355 : 4'b1110;
													assign node11355 = (inp[6]) ? node11359 : node11356;
														assign node11356 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node11359 = (inp[11]) ? 4'b1100 : 4'b0100;
												assign node11362 = (inp[5]) ? node11368 : node11363;
													assign node11363 = (inp[6]) ? 4'b1100 : node11364;
														assign node11364 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node11368 = (inp[3]) ? node11372 : node11369;
														assign node11369 = (inp[6]) ? 4'b0100 : 4'b1100;
														assign node11372 = (inp[6]) ? node11374 : 4'b0110;
															assign node11374 = (inp[11]) ? 4'b1110 : 4'b0110;
											assign node11377 = (inp[15]) ? node11387 : node11378;
												assign node11378 = (inp[6]) ? node11384 : node11379;
													assign node11379 = (inp[5]) ? node11381 : 4'b0100;
														assign node11381 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node11384 = (inp[11]) ? 4'b1100 : 4'b0100;
												assign node11387 = (inp[6]) ? node11393 : node11388;
													assign node11388 = (inp[11]) ? 4'b0110 : node11389;
														assign node11389 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node11393 = (inp[3]) ? 4'b0100 : 4'b0110;
										assign node11396 = (inp[0]) ? node11414 : node11397;
											assign node11397 = (inp[6]) ? node11405 : node11398;
												assign node11398 = (inp[11]) ? 4'b1110 : node11399;
													assign node11399 = (inp[5]) ? node11401 : 4'b0110;
														assign node11401 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node11405 = (inp[11]) ? node11411 : node11406;
													assign node11406 = (inp[5]) ? 4'b1100 : node11407;
														assign node11407 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node11411 = (inp[5]) ? 4'b0110 : 4'b0100;
											assign node11414 = (inp[15]) ? node11426 : node11415;
												assign node11415 = (inp[5]) ? node11423 : node11416;
													assign node11416 = (inp[11]) ? node11420 : node11417;
														assign node11417 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node11420 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node11423 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node11426 = (inp[5]) ? node11428 : 4'b1110;
													assign node11428 = (inp[14]) ? 4'b0100 : node11429;
														assign node11429 = (inp[11]) ? 4'b1100 : 4'b0100;
								assign node11433 = (inp[14]) ? node11519 : node11434;
									assign node11434 = (inp[2]) ? node11476 : node11435;
										assign node11435 = (inp[15]) ? node11453 : node11436;
											assign node11436 = (inp[0]) ? node11446 : node11437;
												assign node11437 = (inp[3]) ? node11443 : node11438;
													assign node11438 = (inp[11]) ? node11440 : 4'b1110;
														assign node11440 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node11443 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node11446 = (inp[6]) ? node11448 : 4'b1100;
													assign node11448 = (inp[11]) ? 4'b0100 : node11449;
														assign node11449 = (inp[1]) ? 4'b1100 : 4'b0100;
											assign node11453 = (inp[3]) ? node11459 : node11454;
												assign node11454 = (inp[6]) ? node11456 : 4'b0100;
													assign node11456 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node11459 = (inp[6]) ? node11465 : node11460;
													assign node11460 = (inp[0]) ? node11462 : 4'b1110;
														assign node11462 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node11465 = (inp[11]) ? node11471 : node11466;
														assign node11466 = (inp[1]) ? 4'b1110 : node11467;
															assign node11467 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node11471 = (inp[1]) ? 4'b0100 : node11472;
															assign node11472 = (inp[5]) ? 4'b1110 : 4'b1100;
										assign node11476 = (inp[15]) ? node11504 : node11477;
											assign node11477 = (inp[3]) ? node11495 : node11478;
												assign node11478 = (inp[0]) ? node11482 : node11479;
													assign node11479 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node11482 = (inp[5]) ? node11490 : node11483;
														assign node11483 = (inp[1]) ? node11487 : node11484;
															assign node11484 = (inp[6]) ? 4'b0101 : 4'b1101;
															assign node11487 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node11490 = (inp[11]) ? 4'b0101 : node11491;
															assign node11491 = (inp[6]) ? 4'b1101 : 4'b0101;
												assign node11495 = (inp[11]) ? node11497 : 4'b1111;
													assign node11497 = (inp[1]) ? node11499 : 4'b1101;
														assign node11499 = (inp[5]) ? node11501 : 4'b1101;
															assign node11501 = (inp[0]) ? 4'b1111 : 4'b1101;
											assign node11504 = (inp[0]) ? node11512 : node11505;
												assign node11505 = (inp[3]) ? node11509 : node11506;
													assign node11506 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node11509 = (inp[6]) ? 4'b1111 : 4'b0111;
												assign node11512 = (inp[3]) ? 4'b0101 : node11513;
													assign node11513 = (inp[1]) ? node11515 : 4'b0111;
														assign node11515 = (inp[11]) ? 4'b1111 : 4'b0111;
									assign node11519 = (inp[6]) ? node11553 : node11520;
										assign node11520 = (inp[11]) ? node11534 : node11521;
											assign node11521 = (inp[0]) ? node11527 : node11522;
												assign node11522 = (inp[15]) ? node11524 : 4'b0111;
													assign node11524 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node11527 = (inp[5]) ? node11531 : node11528;
													assign node11528 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node11531 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node11534 = (inp[2]) ? node11548 : node11535;
												assign node11535 = (inp[5]) ? node11541 : node11536;
													assign node11536 = (inp[3]) ? 4'b1101 : node11537;
														assign node11537 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node11541 = (inp[1]) ? 4'b1111 : node11542;
														assign node11542 = (inp[3]) ? node11544 : 4'b1101;
															assign node11544 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node11548 = (inp[0]) ? node11550 : 4'b1111;
													assign node11550 = (inp[15]) ? 4'b1111 : 4'b1101;
										assign node11553 = (inp[11]) ? node11563 : node11554;
											assign node11554 = (inp[2]) ? node11556 : 4'b1111;
												assign node11556 = (inp[1]) ? 4'b1101 : node11557;
													assign node11557 = (inp[5]) ? 4'b1111 : node11558;
														assign node11558 = (inp[0]) ? 4'b1111 : 4'b1101;
											assign node11563 = (inp[15]) ? node11571 : node11564;
												assign node11564 = (inp[2]) ? node11566 : 4'b0111;
													assign node11566 = (inp[3]) ? node11568 : 4'b0111;
														assign node11568 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node11571 = (inp[3]) ? node11575 : node11572;
													assign node11572 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node11575 = (inp[0]) ? 4'b0101 : 4'b0111;
							assign node11578 = (inp[8]) ? node11736 : node11579;
								assign node11579 = (inp[2]) ? node11669 : node11580;
									assign node11580 = (inp[14]) ? node11636 : node11581;
										assign node11581 = (inp[5]) ? node11601 : node11582;
											assign node11582 = (inp[1]) ? node11588 : node11583;
												assign node11583 = (inp[0]) ? 4'b0100 : node11584;
													assign node11584 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node11588 = (inp[3]) ? node11592 : node11589;
													assign node11589 = (inp[6]) ? 4'b1100 : 4'b0100;
													assign node11592 = (inp[0]) ? node11596 : node11593;
														assign node11593 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node11596 = (inp[11]) ? 4'b1110 : node11597;
															assign node11597 = (inp[6]) ? 4'b1110 : 4'b0110;
											assign node11601 = (inp[1]) ? node11621 : node11602;
												assign node11602 = (inp[0]) ? node11612 : node11603;
													assign node11603 = (inp[11]) ? node11609 : node11604;
														assign node11604 = (inp[6]) ? 4'b0110 : node11605;
															assign node11605 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node11609 = (inp[6]) ? 4'b1110 : 4'b0100;
													assign node11612 = (inp[11]) ? node11616 : node11613;
														assign node11613 = (inp[6]) ? 4'b0100 : 4'b1100;
														assign node11616 = (inp[6]) ? 4'b1110 : node11617;
															assign node11617 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node11621 = (inp[0]) ? node11627 : node11622;
													assign node11622 = (inp[15]) ? 4'b1110 : node11623;
														assign node11623 = (inp[11]) ? 4'b0100 : 4'b1110;
													assign node11627 = (inp[3]) ? node11633 : node11628;
														assign node11628 = (inp[11]) ? 4'b1100 : node11629;
															assign node11629 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node11633 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node11636 = (inp[3]) ? node11648 : node11637;
											assign node11637 = (inp[5]) ? 4'b1101 : node11638;
												assign node11638 = (inp[15]) ? node11640 : 4'b0101;
													assign node11640 = (inp[0]) ? 4'b1111 : node11641;
														assign node11641 = (inp[11]) ? 4'b1101 : node11642;
															assign node11642 = (inp[6]) ? 4'b1101 : 4'b0101;
											assign node11648 = (inp[0]) ? node11664 : node11649;
												assign node11649 = (inp[1]) ? node11659 : node11650;
													assign node11650 = (inp[5]) ? node11654 : node11651;
														assign node11651 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node11654 = (inp[15]) ? 4'b1111 : node11655;
															assign node11655 = (inp[6]) ? 4'b0101 : 4'b0101;
													assign node11659 = (inp[6]) ? 4'b0101 : node11660;
														assign node11660 = (inp[11]) ? 4'b1101 : 4'b0101;
												assign node11664 = (inp[11]) ? node11666 : 4'b1111;
													assign node11666 = (inp[1]) ? 4'b1101 : 4'b1111;
									assign node11669 = (inp[14]) ? node11709 : node11670;
										assign node11670 = (inp[1]) ? node11684 : node11671;
											assign node11671 = (inp[5]) ? node11681 : node11672;
												assign node11672 = (inp[15]) ? node11676 : node11673;
													assign node11673 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node11676 = (inp[0]) ? 4'b1111 : node11677;
														assign node11677 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node11681 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node11684 = (inp[6]) ? node11690 : node11685;
												assign node11685 = (inp[11]) ? 4'b1101 : node11686;
													assign node11686 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node11690 = (inp[11]) ? node11696 : node11691;
													assign node11691 = (inp[3]) ? node11693 : 4'b1111;
														assign node11693 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node11696 = (inp[15]) ? node11702 : node11697;
														assign node11697 = (inp[5]) ? 4'b0111 : node11698;
															assign node11698 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node11702 = (inp[0]) ? node11706 : node11703;
															assign node11703 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node11706 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node11709 = (inp[11]) ? node11723 : node11710;
											assign node11710 = (inp[6]) ? node11714 : node11711;
												assign node11711 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node11714 = (inp[0]) ? node11716 : 4'b1101;
													assign node11716 = (inp[15]) ? 4'b1111 : node11717;
														assign node11717 = (inp[3]) ? node11719 : 4'b1101;
															assign node11719 = (inp[5]) ? 4'b1111 : 4'b1101;
											assign node11723 = (inp[6]) ? node11731 : node11724;
												assign node11724 = (inp[15]) ? 4'b1101 : node11725;
													assign node11725 = (inp[0]) ? node11727 : 4'b1111;
														assign node11727 = (inp[1]) ? 4'b1111 : 4'b1101;
												assign node11731 = (inp[3]) ? 4'b0101 : node11732;
													assign node11732 = (inp[0]) ? 4'b0101 : 4'b0111;
								assign node11736 = (inp[2]) ? node11814 : node11737;
									assign node11737 = (inp[14]) ? node11773 : node11738;
										assign node11738 = (inp[6]) ? node11754 : node11739;
											assign node11739 = (inp[11]) ? 4'b1101 : node11740;
												assign node11740 = (inp[1]) ? node11748 : node11741;
													assign node11741 = (inp[0]) ? 4'b0101 : node11742;
														assign node11742 = (inp[3]) ? node11744 : 4'b0111;
															assign node11744 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node11748 = (inp[0]) ? 4'b0111 : node11749;
														assign node11749 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node11754 = (inp[11]) ? node11768 : node11755;
												assign node11755 = (inp[0]) ? node11765 : node11756;
													assign node11756 = (inp[3]) ? node11758 : 4'b1101;
														assign node11758 = (inp[5]) ? node11762 : node11759;
															assign node11759 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node11762 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node11765 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node11768 = (inp[3]) ? 4'b0101 : node11769;
													assign node11769 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node11773 = (inp[6]) ? node11795 : node11774;
											assign node11774 = (inp[11]) ? node11788 : node11775;
												assign node11775 = (inp[1]) ? 4'b0100 : node11776;
													assign node11776 = (inp[0]) ? node11782 : node11777;
														assign node11777 = (inp[3]) ? 4'b0100 : node11778;
															assign node11778 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node11782 = (inp[5]) ? node11784 : 4'b0110;
															assign node11784 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node11788 = (inp[0]) ? 4'b1100 : node11789;
													assign node11789 = (inp[3]) ? node11791 : 4'b1110;
														assign node11791 = (inp[1]) ? 4'b1110 : 4'b1100;
											assign node11795 = (inp[11]) ? node11807 : node11796;
												assign node11796 = (inp[3]) ? node11798 : 4'b1100;
													assign node11798 = (inp[0]) ? 4'b1100 : node11799;
														assign node11799 = (inp[1]) ? node11803 : node11800;
															assign node11800 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node11803 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node11807 = (inp[15]) ? node11809 : 4'b0100;
													assign node11809 = (inp[5]) ? 4'b0100 : node11810;
														assign node11810 = (inp[3]) ? 4'b0110 : 4'b0100;
									assign node11814 = (inp[0]) ? node11856 : node11815;
										assign node11815 = (inp[15]) ? node11833 : node11816;
											assign node11816 = (inp[5]) ? node11824 : node11817;
												assign node11817 = (inp[6]) ? node11821 : node11818;
													assign node11818 = (inp[11]) ? 4'b1110 : 4'b0110;
													assign node11821 = (inp[11]) ? 4'b0110 : 4'b1110;
												assign node11824 = (inp[3]) ? node11830 : node11825;
													assign node11825 = (inp[1]) ? 4'b1110 : node11826;
														assign node11826 = (inp[14]) ? 4'b1110 : 4'b0110;
													assign node11830 = (inp[1]) ? 4'b1100 : 4'b0100;
											assign node11833 = (inp[5]) ? node11841 : node11834;
												assign node11834 = (inp[11]) ? node11838 : node11835;
													assign node11835 = (inp[6]) ? 4'b1100 : 4'b0100;
													assign node11838 = (inp[6]) ? 4'b0100 : 4'b1100;
												assign node11841 = (inp[3]) ? node11847 : node11842;
													assign node11842 = (inp[6]) ? node11844 : 4'b1100;
														assign node11844 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node11847 = (inp[1]) ? node11849 : 4'b1110;
														assign node11849 = (inp[11]) ? node11853 : node11850;
															assign node11850 = (inp[14]) ? 4'b1110 : 4'b0110;
															assign node11853 = (inp[6]) ? 4'b0110 : 4'b1110;
										assign node11856 = (inp[15]) ? node11868 : node11857;
											assign node11857 = (inp[11]) ? node11865 : node11858;
												assign node11858 = (inp[6]) ? 4'b1100 : node11859;
													assign node11859 = (inp[5]) ? node11861 : 4'b0100;
														assign node11861 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node11865 = (inp[6]) ? 4'b0100 : 4'b1100;
											assign node11868 = (inp[5]) ? node11880 : node11869;
												assign node11869 = (inp[3]) ? node11875 : node11870;
													assign node11870 = (inp[1]) ? node11872 : 4'b0110;
														assign node11872 = (inp[14]) ? 4'b0110 : 4'b1110;
													assign node11875 = (inp[11]) ? 4'b1110 : node11876;
														assign node11876 = (inp[14]) ? 4'b0110 : 4'b1110;
												assign node11880 = (inp[3]) ? node11882 : 4'b1110;
													assign node11882 = (inp[6]) ? 4'b1100 : 4'b0100;
						assign node11885 = (inp[11]) ? node12233 : node11886;
							assign node11886 = (inp[6]) ? node12056 : node11887;
								assign node11887 = (inp[1]) ? node11967 : node11888;
									assign node11888 = (inp[8]) ? node11932 : node11889;
										assign node11889 = (inp[7]) ? node11907 : node11890;
											assign node11890 = (inp[15]) ? node11902 : node11891;
												assign node11891 = (inp[2]) ? node11899 : node11892;
													assign node11892 = (inp[14]) ? node11896 : node11893;
														assign node11893 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node11896 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node11899 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node11902 = (inp[14]) ? 4'b1110 : node11903;
													assign node11903 = (inp[5]) ? 4'b1111 : 4'b1110;
											assign node11907 = (inp[14]) ? node11921 : node11908;
												assign node11908 = (inp[2]) ? node11918 : node11909;
													assign node11909 = (inp[5]) ? 4'b1100 : node11910;
														assign node11910 = (inp[0]) ? node11914 : node11911;
															assign node11911 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node11914 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node11918 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node11921 = (inp[15]) ? node11929 : node11922;
													assign node11922 = (inp[3]) ? node11924 : 4'b0111;
														assign node11924 = (inp[2]) ? node11926 : 4'b0111;
															assign node11926 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node11929 = (inp[0]) ? 4'b0111 : 4'b0101;
										assign node11932 = (inp[7]) ? node11952 : node11933;
											assign node11933 = (inp[2]) ? node11943 : node11934;
												assign node11934 = (inp[14]) ? node11940 : node11935;
													assign node11935 = (inp[5]) ? node11937 : 4'b1110;
														assign node11937 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node11940 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node11943 = (inp[14]) ? 4'b0111 : node11944;
													assign node11944 = (inp[0]) ? node11946 : 4'b0111;
														assign node11946 = (inp[5]) ? node11948 : 4'b0101;
															assign node11948 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node11952 = (inp[14]) ? node11962 : node11953;
												assign node11953 = (inp[2]) ? 4'b0100 : node11954;
													assign node11954 = (inp[5]) ? 4'b0101 : node11955;
														assign node11955 = (inp[0]) ? 4'b0111 : node11956;
															assign node11956 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node11962 = (inp[3]) ? node11964 : 4'b0110;
													assign node11964 = (inp[2]) ? 4'b0110 : 4'b0100;
									assign node11967 = (inp[14]) ? node12015 : node11968;
										assign node11968 = (inp[15]) ? node11996 : node11969;
											assign node11969 = (inp[7]) ? node11987 : node11970;
												assign node11970 = (inp[2]) ? node11980 : node11971;
													assign node11971 = (inp[8]) ? node11975 : node11972;
														assign node11972 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node11975 = (inp[5]) ? node11977 : 4'b0110;
															assign node11977 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node11980 = (inp[8]) ? node11982 : 4'b0110;
														assign node11982 = (inp[0]) ? 4'b0101 : node11983;
															assign node11983 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node11987 = (inp[8]) ? node11991 : node11988;
													assign node11988 = (inp[2]) ? 4'b0101 : 4'b0110;
													assign node11991 = (inp[2]) ? 4'b0110 : node11992;
														assign node11992 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node11996 = (inp[0]) ? node12008 : node11997;
												assign node11997 = (inp[3]) ? node12003 : node11998;
													assign node11998 = (inp[8]) ? node12000 : 4'b0100;
														assign node12000 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node12003 = (inp[7]) ? node12005 : 4'b0101;
														assign node12005 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node12008 = (inp[5]) ? node12012 : node12009;
													assign node12009 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node12012 = (inp[3]) ? 4'b0100 : 4'b0110;
										assign node12015 = (inp[8]) ? node12039 : node12016;
											assign node12016 = (inp[7]) ? node12030 : node12017;
												assign node12017 = (inp[3]) ? node12019 : 4'b0100;
													assign node12019 = (inp[5]) ? node12025 : node12020;
														assign node12020 = (inp[0]) ? 4'b0100 : node12021;
															assign node12021 = (inp[2]) ? 4'b0100 : 4'b0110;
														assign node12025 = (inp[0]) ? 4'b0110 : node12026;
															assign node12026 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node12030 = (inp[15]) ? node12032 : 4'b0101;
													assign node12032 = (inp[2]) ? node12036 : node12033;
														assign node12033 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node12036 = (inp[0]) ? 4'b0111 : 4'b0101;
											assign node12039 = (inp[7]) ? node12049 : node12040;
												assign node12040 = (inp[5]) ? 4'b0111 : node12041;
													assign node12041 = (inp[15]) ? node12045 : node12042;
														assign node12042 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node12045 = (inp[2]) ? 4'b0101 : 4'b0111;
												assign node12049 = (inp[5]) ? node12051 : 4'b0100;
													assign node12051 = (inp[2]) ? node12053 : 4'b0110;
														assign node12053 = (inp[15]) ? 4'b0110 : 4'b0100;
								assign node12056 = (inp[1]) ? node12136 : node12057;
									assign node12057 = (inp[8]) ? node12099 : node12058;
										assign node12058 = (inp[7]) ? node12082 : node12059;
											assign node12059 = (inp[0]) ? node12071 : node12060;
												assign node12060 = (inp[14]) ? 4'b0100 : node12061;
													assign node12061 = (inp[2]) ? node12067 : node12062;
														assign node12062 = (inp[3]) ? 4'b0101 : node12063;
															assign node12063 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node12067 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node12071 = (inp[15]) ? node12077 : node12072;
													assign node12072 = (inp[14]) ? node12074 : 4'b0100;
														assign node12074 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node12077 = (inp[14]) ? 4'b0110 : node12078;
														assign node12078 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node12082 = (inp[14]) ? node12092 : node12083;
												assign node12083 = (inp[2]) ? 4'b1001 : node12084;
													assign node12084 = (inp[5]) ? 4'b0110 : node12085;
														assign node12085 = (inp[3]) ? 4'b0100 : node12086;
															assign node12086 = (inp[0]) ? 4'b0100 : 4'b0100;
												assign node12092 = (inp[2]) ? node12094 : 4'b1011;
													assign node12094 = (inp[3]) ? node12096 : 4'b1001;
														assign node12096 = (inp[15]) ? 4'b1011 : 4'b1001;
										assign node12099 = (inp[7]) ? node12117 : node12100;
											assign node12100 = (inp[14]) ? node12108 : node12101;
												assign node12101 = (inp[2]) ? node12103 : 4'b0100;
													assign node12103 = (inp[0]) ? 4'b1001 : node12104;
														assign node12104 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node12108 = (inp[15]) ? node12110 : 4'b1011;
													assign node12110 = (inp[2]) ? node12112 : 4'b1001;
														assign node12112 = (inp[5]) ? node12114 : 4'b1011;
															assign node12114 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node12117 = (inp[2]) ? node12125 : node12118;
												assign node12118 = (inp[14]) ? 4'b1010 : node12119;
													assign node12119 = (inp[3]) ? node12121 : 4'b1011;
														assign node12121 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node12125 = (inp[0]) ? 4'b1000 : node12126;
													assign node12126 = (inp[14]) ? node12132 : node12127;
														assign node12127 = (inp[3]) ? node12129 : 4'b1010;
															assign node12129 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node12132 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node12136 = (inp[14]) ? node12196 : node12137;
										assign node12137 = (inp[3]) ? node12165 : node12138;
											assign node12138 = (inp[7]) ? node12154 : node12139;
												assign node12139 = (inp[5]) ? node12149 : node12140;
													assign node12140 = (inp[8]) ? node12144 : node12141;
														assign node12141 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node12144 = (inp[2]) ? 4'b1011 : node12145;
															assign node12145 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node12149 = (inp[15]) ? node12151 : 4'b1000;
														assign node12151 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node12154 = (inp[5]) ? node12158 : node12155;
													assign node12155 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node12158 = (inp[0]) ? node12162 : node12159;
														assign node12159 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node12162 = (inp[15]) ? 4'b1011 : 4'b1001;
											assign node12165 = (inp[5]) ? node12185 : node12166;
												assign node12166 = (inp[0]) ? node12176 : node12167;
													assign node12167 = (inp[15]) ? node12171 : node12168;
														assign node12168 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node12171 = (inp[2]) ? 4'b1000 : node12172;
															assign node12172 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node12176 = (inp[15]) ? node12180 : node12177;
														assign node12177 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node12180 = (inp[8]) ? 4'b1010 : node12181;
															assign node12181 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node12185 = (inp[0]) ? node12193 : node12186;
													assign node12186 = (inp[15]) ? node12188 : 4'b1000;
														assign node12188 = (inp[8]) ? 4'b1011 : node12189;
															assign node12189 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node12193 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node12196 = (inp[0]) ? node12216 : node12197;
											assign node12197 = (inp[15]) ? node12209 : node12198;
												assign node12198 = (inp[3]) ? node12200 : 4'b1011;
													assign node12200 = (inp[5]) ? node12206 : node12201;
														assign node12201 = (inp[8]) ? node12203 : 4'b1010;
															assign node12203 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node12206 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node12209 = (inp[3]) ? 4'b1011 : node12210;
													assign node12210 = (inp[7]) ? node12212 : 4'b1001;
														assign node12212 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node12216 = (inp[3]) ? node12224 : node12217;
												assign node12217 = (inp[15]) ? node12219 : 4'b1000;
													assign node12219 = (inp[7]) ? 4'b1010 : node12220;
														assign node12220 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node12224 = (inp[5]) ? node12228 : node12225;
													assign node12225 = (inp[2]) ? 4'b1000 : 4'b1010;
													assign node12228 = (inp[8]) ? 4'b1000 : node12229;
														assign node12229 = (inp[2]) ? 4'b1000 : 4'b1001;
							assign node12233 = (inp[6]) ? node12403 : node12234;
								assign node12234 = (inp[1]) ? node12320 : node12235;
									assign node12235 = (inp[2]) ? node12281 : node12236;
										assign node12236 = (inp[7]) ? node12262 : node12237;
											assign node12237 = (inp[8]) ? node12251 : node12238;
												assign node12238 = (inp[14]) ? node12244 : node12239;
													assign node12239 = (inp[5]) ? 4'b0111 : node12240;
														assign node12240 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node12244 = (inp[3]) ? 4'b0110 : node12245;
														assign node12245 = (inp[15]) ? node12247 : 4'b0100;
															assign node12247 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node12251 = (inp[15]) ? node12253 : 4'b0110;
													assign node12253 = (inp[3]) ? node12257 : node12254;
														assign node12254 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node12257 = (inp[5]) ? node12259 : 4'b0100;
															assign node12259 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node12262 = (inp[8]) ? node12270 : node12263;
												assign node12263 = (inp[14]) ? 4'b1011 : node12264;
													assign node12264 = (inp[5]) ? 4'b0110 : node12265;
														assign node12265 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node12270 = (inp[14]) ? node12278 : node12271;
													assign node12271 = (inp[3]) ? node12273 : 4'b1011;
														assign node12273 = (inp[5]) ? 4'b1001 : node12274;
															assign node12274 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node12278 = (inp[5]) ? 4'b1010 : 4'b1000;
										assign node12281 = (inp[8]) ? node12299 : node12282;
											assign node12282 = (inp[7]) ? node12290 : node12283;
												assign node12283 = (inp[5]) ? 4'b0110 : node12284;
													assign node12284 = (inp[0]) ? node12286 : 4'b0110;
														assign node12286 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node12290 = (inp[15]) ? node12296 : node12291;
													assign node12291 = (inp[0]) ? 4'b1001 : node12292;
														assign node12292 = (inp[14]) ? 4'b1001 : 4'b1011;
													assign node12296 = (inp[14]) ? 4'b1011 : 4'b1001;
											assign node12299 = (inp[7]) ? node12311 : node12300;
												assign node12300 = (inp[0]) ? node12302 : 4'b1001;
													assign node12302 = (inp[14]) ? node12304 : 4'b1001;
														assign node12304 = (inp[3]) ? node12308 : node12305;
															assign node12305 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node12308 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node12311 = (inp[5]) ? 4'b1000 : node12312;
													assign node12312 = (inp[0]) ? node12316 : node12313;
														assign node12313 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node12316 = (inp[15]) ? 4'b1010 : 4'b1000;
									assign node12320 = (inp[3]) ? node12350 : node12321;
										assign node12321 = (inp[7]) ? node12335 : node12322;
											assign node12322 = (inp[0]) ? node12326 : node12323;
												assign node12323 = (inp[5]) ? 4'b1000 : 4'b1001;
												assign node12326 = (inp[15]) ? node12330 : node12327;
													assign node12327 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node12330 = (inp[8]) ? 4'b1011 : node12331;
														assign node12331 = (inp[5]) ? 4'b1010 : 4'b1011;
											assign node12335 = (inp[8]) ? node12341 : node12336;
												assign node12336 = (inp[0]) ? 4'b1010 : node12337;
													assign node12337 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node12341 = (inp[0]) ? node12347 : node12342;
													assign node12342 = (inp[2]) ? node12344 : 4'b1011;
														assign node12344 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node12347 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node12350 = (inp[2]) ? node12378 : node12351;
											assign node12351 = (inp[7]) ? node12367 : node12352;
												assign node12352 = (inp[0]) ? node12358 : node12353;
													assign node12353 = (inp[8]) ? node12355 : 4'b1011;
														assign node12355 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node12358 = (inp[8]) ? node12362 : node12359;
														assign node12359 = (inp[14]) ? 4'b1010 : 4'b1001;
														assign node12362 = (inp[14]) ? node12364 : 4'b1000;
															assign node12364 = (inp[5]) ? 4'b1001 : 4'b1001;
												assign node12367 = (inp[8]) ? 4'b1000 : node12368;
													assign node12368 = (inp[14]) ? node12374 : node12369;
														assign node12369 = (inp[5]) ? 4'b1010 : node12370;
															assign node12370 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node12374 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node12378 = (inp[0]) ? node12392 : node12379;
												assign node12379 = (inp[5]) ? node12387 : node12380;
													assign node12380 = (inp[15]) ? node12382 : 4'b1011;
														assign node12382 = (inp[14]) ? node12384 : 4'b1001;
															assign node12384 = (inp[8]) ? 4'b1000 : 4'b1000;
													assign node12387 = (inp[15]) ? 4'b1011 : node12388;
														assign node12388 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node12392 = (inp[8]) ? node12398 : node12393;
													assign node12393 = (inp[7]) ? node12395 : 4'b1000;
														assign node12395 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node12398 = (inp[14]) ? node12400 : 4'b1000;
														assign node12400 = (inp[7]) ? 4'b1010 : 4'b1011;
								assign node12403 = (inp[1]) ? node12489 : node12404;
									assign node12404 = (inp[8]) ? node12448 : node12405;
										assign node12405 = (inp[7]) ? node12425 : node12406;
											assign node12406 = (inp[2]) ? node12414 : node12407;
												assign node12407 = (inp[14]) ? node12409 : 4'b1011;
													assign node12409 = (inp[15]) ? 4'b1010 : node12410;
														assign node12410 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node12414 = (inp[0]) ? node12418 : node12415;
													assign node12415 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node12418 = (inp[5]) ? node12420 : 4'b1000;
														assign node12420 = (inp[3]) ? node12422 : 4'b1000;
															assign node12422 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node12425 = (inp[2]) ? node12439 : node12426;
												assign node12426 = (inp[14]) ? 4'b0001 : node12427;
													assign node12427 = (inp[5]) ? node12433 : node12428;
														assign node12428 = (inp[15]) ? node12430 : 4'b1000;
															assign node12430 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node12433 = (inp[15]) ? node12435 : 4'b1010;
															assign node12435 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node12439 = (inp[3]) ? node12441 : 4'b0011;
													assign node12441 = (inp[14]) ? 4'b0001 : node12442;
														assign node12442 = (inp[15]) ? 4'b0011 : node12443;
															assign node12443 = (inp[0]) ? 4'b0001 : 4'b0001;
										assign node12448 = (inp[7]) ? node12474 : node12449;
											assign node12449 = (inp[14]) ? node12463 : node12450;
												assign node12450 = (inp[2]) ? node12458 : node12451;
													assign node12451 = (inp[3]) ? 4'b1010 : node12452;
														assign node12452 = (inp[5]) ? node12454 : 4'b1000;
															assign node12454 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node12458 = (inp[0]) ? node12460 : 4'b0001;
														assign node12460 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node12463 = (inp[15]) ? node12469 : node12464;
													assign node12464 = (inp[5]) ? node12466 : 4'b0011;
														assign node12466 = (inp[2]) ? 4'b0001 : 4'b0011;
													assign node12469 = (inp[0]) ? node12471 : 4'b0001;
														assign node12471 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node12474 = (inp[14]) ? node12484 : node12475;
												assign node12475 = (inp[2]) ? node12477 : 4'b0001;
													assign node12477 = (inp[15]) ? 4'b0010 : node12478;
														assign node12478 = (inp[5]) ? node12480 : 4'b0000;
															assign node12480 = (inp[3]) ? 4'b0000 : 4'b0000;
												assign node12484 = (inp[3]) ? node12486 : 4'b0000;
													assign node12486 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node12489 = (inp[7]) ? node12537 : node12490;
										assign node12490 = (inp[8]) ? node12516 : node12491;
											assign node12491 = (inp[14]) ? node12499 : node12492;
												assign node12492 = (inp[2]) ? node12494 : 4'b0001;
													assign node12494 = (inp[3]) ? node12496 : 4'b0000;
														assign node12496 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node12499 = (inp[2]) ? node12511 : node12500;
													assign node12500 = (inp[3]) ? node12506 : node12501;
														assign node12501 = (inp[5]) ? 4'b0010 : node12502;
															assign node12502 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node12506 = (inp[5]) ? 4'b0000 : node12507;
															assign node12507 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node12511 = (inp[5]) ? node12513 : 4'b0000;
														assign node12513 = (inp[3]) ? 4'b0010 : 4'b0000;
											assign node12516 = (inp[3]) ? 4'b0010 : node12517;
												assign node12517 = (inp[14]) ? node12527 : node12518;
													assign node12518 = (inp[2]) ? node12522 : node12519;
														assign node12519 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node12522 = (inp[5]) ? 4'b0001 : node12523;
															assign node12523 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node12527 = (inp[2]) ? 4'b0011 : node12528;
														assign node12528 = (inp[0]) ? node12532 : node12529;
															assign node12529 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node12532 = (inp[15]) ? 4'b0011 : 4'b0001;
										assign node12537 = (inp[8]) ? node12549 : node12538;
											assign node12538 = (inp[2]) ? node12544 : node12539;
												assign node12539 = (inp[5]) ? 4'b0010 : node12540;
													assign node12540 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node12544 = (inp[5]) ? node12546 : 4'b0011;
													assign node12546 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node12549 = (inp[2]) ? node12557 : node12550;
												assign node12550 = (inp[14]) ? 4'b0010 : node12551;
													assign node12551 = (inp[0]) ? 4'b0001 : node12552;
														assign node12552 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node12557 = (inp[15]) ? node12559 : 4'b0000;
													assign node12559 = (inp[0]) ? 4'b0010 : 4'b0000;
					assign node12562 = (inp[12]) ? node13240 : node12563;
						assign node12563 = (inp[14]) ? node12987 : node12564;
							assign node12564 = (inp[0]) ? node12772 : node12565;
								assign node12565 = (inp[15]) ? node12673 : node12566;
									assign node12566 = (inp[3]) ? node12616 : node12567;
										assign node12567 = (inp[11]) ? node12591 : node12568;
											assign node12568 = (inp[5]) ? node12578 : node12569;
												assign node12569 = (inp[2]) ? node12571 : 4'b1010;
													assign node12571 = (inp[1]) ? 4'b1010 : node12572;
														assign node12572 = (inp[7]) ? 4'b0010 : node12573;
															assign node12573 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node12578 = (inp[7]) ? node12582 : node12579;
													assign node12579 = (inp[8]) ? 4'b0011 : 4'b1011;
													assign node12582 = (inp[2]) ? node12588 : node12583;
														assign node12583 = (inp[6]) ? node12585 : 4'b0010;
															assign node12585 = (inp[1]) ? 4'b1010 : 4'b0010;
														assign node12588 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node12591 = (inp[6]) ? node12609 : node12592;
												assign node12592 = (inp[1]) ? node12598 : node12593;
													assign node12593 = (inp[7]) ? node12595 : 4'b0010;
														assign node12595 = (inp[8]) ? 4'b1011 : 4'b0010;
													assign node12598 = (inp[2]) ? node12604 : node12599;
														assign node12599 = (inp[8]) ? node12601 : 4'b1010;
															assign node12601 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node12604 = (inp[7]) ? 4'b1011 : node12605;
															assign node12605 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node12609 = (inp[7]) ? 4'b0011 : node12610;
													assign node12610 = (inp[1]) ? 4'b0010 : node12611;
														assign node12611 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node12616 = (inp[5]) ? node12642 : node12617;
											assign node12617 = (inp[2]) ? node12627 : node12618;
												assign node12618 = (inp[1]) ? node12624 : node12619;
													assign node12619 = (inp[7]) ? 4'b1010 : node12620;
														assign node12620 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node12624 = (inp[11]) ? 4'b0010 : 4'b1010;
												assign node12627 = (inp[6]) ? node12637 : node12628;
													assign node12628 = (inp[11]) ? node12634 : node12629;
														assign node12629 = (inp[1]) ? node12631 : 4'b0010;
															assign node12631 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node12634 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node12637 = (inp[7]) ? 4'b1011 : node12638;
														assign node12638 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node12642 = (inp[7]) ? node12658 : node12643;
												assign node12643 = (inp[2]) ? node12653 : node12644;
													assign node12644 = (inp[8]) ? node12648 : node12645;
														assign node12645 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node12648 = (inp[6]) ? node12650 : 4'b0000;
															assign node12650 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node12653 = (inp[8]) ? node12655 : 4'b0000;
														assign node12655 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node12658 = (inp[6]) ? node12666 : node12659;
													assign node12659 = (inp[11]) ? node12661 : 4'b0001;
														assign node12661 = (inp[8]) ? 4'b1001 : node12662;
															assign node12662 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node12666 = (inp[2]) ? node12670 : node12667;
														assign node12667 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node12670 = (inp[8]) ? 4'b1000 : 4'b1001;
									assign node12673 = (inp[3]) ? node12725 : node12674;
										assign node12674 = (inp[8]) ? node12698 : node12675;
											assign node12675 = (inp[11]) ? node12687 : node12676;
												assign node12676 = (inp[6]) ? node12682 : node12677;
													assign node12677 = (inp[2]) ? node12679 : 4'b0001;
														assign node12679 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node12682 = (inp[2]) ? 4'b0000 : node12683;
														assign node12683 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node12687 = (inp[6]) ? node12691 : node12688;
													assign node12688 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node12691 = (inp[1]) ? node12693 : 4'b1001;
														assign node12693 = (inp[2]) ? node12695 : 4'b0000;
															assign node12695 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node12698 = (inp[11]) ? node12708 : node12699;
												assign node12699 = (inp[2]) ? node12705 : node12700;
													assign node12700 = (inp[1]) ? node12702 : 4'b0000;
														assign node12702 = (inp[6]) ? 4'b1001 : 4'b0001;
													assign node12705 = (inp[6]) ? 4'b1000 : 4'b0000;
												assign node12708 = (inp[6]) ? node12720 : node12709;
													assign node12709 = (inp[5]) ? node12715 : node12710;
														assign node12710 = (inp[2]) ? node12712 : 4'b1000;
															assign node12712 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node12715 = (inp[7]) ? node12717 : 4'b1001;
															assign node12717 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node12720 = (inp[7]) ? 4'b0001 : node12721;
														assign node12721 = (inp[2]) ? 4'b0001 : 4'b0000;
										assign node12725 = (inp[5]) ? node12749 : node12726;
											assign node12726 = (inp[2]) ? node12734 : node12727;
												assign node12727 = (inp[1]) ? node12731 : node12728;
													assign node12728 = (inp[7]) ? 4'b0001 : 4'b1001;
													assign node12731 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node12734 = (inp[1]) ? node12742 : node12735;
													assign node12735 = (inp[11]) ? 4'b0000 : node12736;
														assign node12736 = (inp[7]) ? node12738 : 4'b0001;
															assign node12738 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node12742 = (inp[8]) ? node12746 : node12743;
														assign node12743 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node12746 = (inp[6]) ? 4'b1000 : 4'b1001;
											assign node12749 = (inp[8]) ? node12765 : node12750;
												assign node12750 = (inp[2]) ? node12758 : node12751;
													assign node12751 = (inp[11]) ? 4'b1011 : node12752;
														assign node12752 = (inp[6]) ? 4'b0010 : node12753;
															assign node12753 = (inp[1]) ? 4'b0010 : 4'b1010;
													assign node12758 = (inp[7]) ? node12760 : 4'b1010;
														assign node12760 = (inp[1]) ? 4'b1011 : node12761;
															assign node12761 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node12765 = (inp[11]) ? node12767 : 4'b0011;
													assign node12767 = (inp[6]) ? node12769 : 4'b0010;
														assign node12769 = (inp[2]) ? 4'b0010 : 4'b0011;
								assign node12772 = (inp[15]) ? node12906 : node12773;
									assign node12773 = (inp[5]) ? node12841 : node12774;
										assign node12774 = (inp[7]) ? node12806 : node12775;
											assign node12775 = (inp[3]) ? node12789 : node12776;
												assign node12776 = (inp[6]) ? node12784 : node12777;
													assign node12777 = (inp[8]) ? 4'b1001 : node12778;
														assign node12778 = (inp[1]) ? 4'b1001 : node12779;
															assign node12779 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node12784 = (inp[2]) ? node12786 : 4'b0000;
														assign node12786 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node12789 = (inp[2]) ? node12797 : node12790;
													assign node12790 = (inp[8]) ? node12792 : 4'b1001;
														assign node12792 = (inp[1]) ? 4'b1000 : node12793;
															assign node12793 = (inp[6]) ? 4'b0000 : 4'b0000;
													assign node12797 = (inp[8]) ? node12801 : node12798;
														assign node12798 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node12801 = (inp[6]) ? node12803 : 4'b1001;
															assign node12803 = (inp[1]) ? 4'b0001 : 4'b1001;
											assign node12806 = (inp[1]) ? node12822 : node12807;
												assign node12807 = (inp[6]) ? node12815 : node12808;
													assign node12808 = (inp[11]) ? node12812 : node12809;
														assign node12809 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node12812 = (inp[8]) ? 4'b1000 : 4'b0000;
													assign node12815 = (inp[2]) ? 4'b1000 : node12816;
														assign node12816 = (inp[8]) ? node12818 : 4'b1000;
															assign node12818 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node12822 = (inp[8]) ? node12834 : node12823;
													assign node12823 = (inp[2]) ? node12829 : node12824;
														assign node12824 = (inp[3]) ? 4'b0000 : node12825;
															assign node12825 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node12829 = (inp[6]) ? node12831 : 4'b1001;
															assign node12831 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node12834 = (inp[2]) ? node12836 : 4'b0001;
														assign node12836 = (inp[3]) ? 4'b0000 : node12837;
															assign node12837 = (inp[6]) ? 4'b1000 : 4'b0000;
										assign node12841 = (inp[3]) ? node12879 : node12842;
											assign node12842 = (inp[8]) ? node12860 : node12843;
												assign node12843 = (inp[11]) ? node12853 : node12844;
													assign node12844 = (inp[1]) ? node12850 : node12845;
														assign node12845 = (inp[2]) ? 4'b1000 : node12846;
															assign node12846 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node12850 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node12853 = (inp[7]) ? node12855 : 4'b1000;
														assign node12855 = (inp[2]) ? node12857 : 4'b1000;
															assign node12857 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node12860 = (inp[2]) ? node12872 : node12861;
													assign node12861 = (inp[7]) ? node12869 : node12862;
														assign node12862 = (inp[11]) ? node12866 : node12863;
															assign node12863 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node12866 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node12869 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node12872 = (inp[11]) ? node12876 : node12873;
														assign node12873 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node12876 = (inp[6]) ? 4'b0001 : 4'b1001;
											assign node12879 = (inp[8]) ? node12889 : node12880;
												assign node12880 = (inp[1]) ? 4'b1011 : node12881;
													assign node12881 = (inp[11]) ? node12883 : 4'b0010;
														assign node12883 = (inp[2]) ? node12885 : 4'b0011;
															assign node12885 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node12889 = (inp[6]) ? node12897 : node12890;
													assign node12890 = (inp[7]) ? 4'b0010 : node12891;
														assign node12891 = (inp[2]) ? node12893 : 4'b0010;
															assign node12893 = (inp[11]) ? 4'b1011 : 4'b0011;
													assign node12897 = (inp[2]) ? node12903 : node12898;
														assign node12898 = (inp[7]) ? node12900 : 4'b1010;
															assign node12900 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node12903 = (inp[11]) ? 4'b0010 : 4'b1010;
									assign node12906 = (inp[5]) ? node12950 : node12907;
										assign node12907 = (inp[2]) ? node12933 : node12908;
											assign node12908 = (inp[3]) ? node12916 : node12909;
												assign node12909 = (inp[1]) ? node12911 : 4'b0010;
													assign node12911 = (inp[6]) ? 4'b1010 : node12912;
														assign node12912 = (inp[11]) ? 4'b1010 : 4'b0011;
												assign node12916 = (inp[8]) ? node12924 : node12917;
													assign node12917 = (inp[6]) ? 4'b1011 : node12918;
														assign node12918 = (inp[11]) ? node12920 : 4'b0011;
															assign node12920 = (inp[1]) ? 4'b1011 : 4'b0011;
													assign node12924 = (inp[7]) ? node12928 : node12925;
														assign node12925 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node12928 = (inp[6]) ? node12930 : 4'b1011;
															assign node12930 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node12933 = (inp[11]) ? node12939 : node12934;
												assign node12934 = (inp[6]) ? node12936 : 4'b0010;
													assign node12936 = (inp[7]) ? 4'b1010 : 4'b0010;
												assign node12939 = (inp[6]) ? node12947 : node12940;
													assign node12940 = (inp[1]) ? 4'b1010 : node12941;
														assign node12941 = (inp[3]) ? node12943 : 4'b1011;
															assign node12943 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node12947 = (inp[8]) ? 4'b0010 : 4'b1010;
										assign node12950 = (inp[3]) ? node12964 : node12951;
											assign node12951 = (inp[1]) ? node12953 : 4'b1010;
												assign node12953 = (inp[6]) ? node12959 : node12954;
													assign node12954 = (inp[8]) ? 4'b1010 : node12955;
														assign node12955 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node12959 = (inp[7]) ? 4'b1010 : node12960;
														assign node12960 = (inp[8]) ? 4'b0011 : 4'b0010;
											assign node12964 = (inp[2]) ? node12978 : node12965;
												assign node12965 = (inp[7]) ? node12967 : 4'b1001;
													assign node12967 = (inp[8]) ? node12971 : node12968;
														assign node12968 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node12971 = (inp[11]) ? node12975 : node12972;
															assign node12972 = (inp[1]) ? 4'b0001 : 4'b1001;
															assign node12975 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node12978 = (inp[11]) ? node12982 : node12979;
													assign node12979 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node12982 = (inp[1]) ? 4'b0000 : node12983;
														assign node12983 = (inp[7]) ? 4'b1000 : 4'b0000;
							assign node12987 = (inp[11]) ? node13121 : node12988;
								assign node12988 = (inp[6]) ? node13060 : node12989;
									assign node12989 = (inp[1]) ? node13011 : node12990;
										assign node12990 = (inp[7]) ? node13000 : node12991;
											assign node12991 = (inp[8]) ? node12997 : node12992;
												assign node12992 = (inp[2]) ? 4'b1000 : node12993;
													assign node12993 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node12997 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node13000 = (inp[8]) ? node13008 : node13001;
												assign node13001 = (inp[2]) ? 4'b0011 : node13002;
													assign node13002 = (inp[0]) ? 4'b0001 : node13003;
														assign node13003 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node13008 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node13011 = (inp[0]) ? node13039 : node13012;
											assign node13012 = (inp[15]) ? node13026 : node13013;
												assign node13013 = (inp[3]) ? node13021 : node13014;
													assign node13014 = (inp[5]) ? 4'b0011 : node13015;
														assign node13015 = (inp[8]) ? 4'b0010 : node13016;
															assign node13016 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node13021 = (inp[7]) ? node13023 : 4'b0000;
														assign node13023 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node13026 = (inp[5]) ? node13034 : node13027;
													assign node13027 = (inp[7]) ? node13031 : node13028;
														assign node13028 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node13031 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node13034 = (inp[3]) ? node13036 : 4'b0000;
														assign node13036 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node13039 = (inp[15]) ? node13051 : node13040;
												assign node13040 = (inp[3]) ? node13046 : node13041;
													assign node13041 = (inp[7]) ? node13043 : 4'b0001;
														assign node13043 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node13046 = (inp[8]) ? 4'b0010 : node13047;
														assign node13047 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node13051 = (inp[5]) ? node13057 : node13052;
													assign node13052 = (inp[3]) ? node13054 : 4'b0010;
														assign node13054 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node13057 = (inp[3]) ? 4'b0001 : 4'b0011;
									assign node13060 = (inp[8]) ? node13092 : node13061;
										assign node13061 = (inp[7]) ? node13069 : node13062;
											assign node13062 = (inp[1]) ? node13064 : 4'b0010;
												assign node13064 = (inp[15]) ? 4'b1000 : node13065;
													assign node13065 = (inp[3]) ? 4'b1010 : 4'b1000;
											assign node13069 = (inp[0]) ? node13079 : node13070;
												assign node13070 = (inp[2]) ? node13074 : node13071;
													assign node13071 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node13074 = (inp[15]) ? node13076 : 4'b1001;
														assign node13076 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node13079 = (inp[2]) ? node13087 : node13080;
													assign node13080 = (inp[3]) ? node13082 : 4'b1011;
														assign node13082 = (inp[15]) ? 4'b1001 : node13083;
															assign node13083 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node13087 = (inp[15]) ? 4'b1011 : node13088;
														assign node13088 = (inp[5]) ? 4'b1011 : 4'b1001;
										assign node13092 = (inp[7]) ? node13114 : node13093;
											assign node13093 = (inp[5]) ? node13101 : node13094;
												assign node13094 = (inp[0]) ? node13098 : node13095;
													assign node13095 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node13098 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node13101 = (inp[1]) ? 4'b1001 : node13102;
													assign node13102 = (inp[15]) ? node13108 : node13103;
														assign node13103 = (inp[2]) ? 4'b1001 : node13104;
															assign node13104 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node13108 = (inp[2]) ? node13110 : 4'b1001;
															assign node13110 = (inp[0]) ? 4'b1001 : 4'b1001;
											assign node13114 = (inp[2]) ? node13116 : 4'b1010;
												assign node13116 = (inp[0]) ? node13118 : 4'b1000;
													assign node13118 = (inp[15]) ? 4'b1010 : 4'b1000;
								assign node13121 = (inp[6]) ? node13183 : node13122;
									assign node13122 = (inp[7]) ? node13148 : node13123;
										assign node13123 = (inp[8]) ? node13139 : node13124;
											assign node13124 = (inp[1]) ? node13132 : node13125;
												assign node13125 = (inp[0]) ? node13127 : 4'b0000;
													assign node13127 = (inp[2]) ? node13129 : 4'b0010;
														assign node13129 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node13132 = (inp[0]) ? node13134 : 4'b1000;
													assign node13134 = (inp[3]) ? 4'b1010 : node13135;
														assign node13135 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node13139 = (inp[0]) ? 4'b1011 : node13140;
												assign node13140 = (inp[15]) ? 4'b1001 : node13141;
													assign node13141 = (inp[5]) ? node13143 : 4'b1011;
														assign node13143 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node13148 = (inp[8]) ? node13170 : node13149;
											assign node13149 = (inp[1]) ? node13163 : node13150;
												assign node13150 = (inp[3]) ? node13152 : 4'b1011;
													assign node13152 = (inp[2]) ? node13158 : node13153;
														assign node13153 = (inp[0]) ? 4'b1001 : node13154;
															assign node13154 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node13158 = (inp[5]) ? node13160 : 4'b1001;
															assign node13160 = (inp[15]) ? 4'b1001 : 4'b1001;
												assign node13163 = (inp[15]) ? node13165 : 4'b1001;
													assign node13165 = (inp[0]) ? 4'b1011 : node13166;
														assign node13166 = (inp[3]) ? 4'b1011 : 4'b1001;
											assign node13170 = (inp[15]) ? node13176 : node13171;
												assign node13171 = (inp[5]) ? 4'b1000 : node13172;
													assign node13172 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node13176 = (inp[0]) ? 4'b1010 : node13177;
													assign node13177 = (inp[5]) ? node13179 : 4'b1000;
														assign node13179 = (inp[3]) ? 4'b1010 : 4'b1000;
									assign node13183 = (inp[7]) ? node13207 : node13184;
										assign node13184 = (inp[8]) ? node13200 : node13185;
											assign node13185 = (inp[1]) ? node13195 : node13186;
												assign node13186 = (inp[15]) ? 4'b1000 : node13187;
													assign node13187 = (inp[5]) ? node13189 : 4'b1010;
														assign node13189 = (inp[2]) ? 4'b1000 : node13190;
															assign node13190 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node13195 = (inp[0]) ? node13197 : 4'b0000;
													assign node13197 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node13200 = (inp[3]) ? node13202 : 4'b0011;
												assign node13202 = (inp[15]) ? 4'b0001 : node13203;
													assign node13203 = (inp[0]) ? 4'b0011 : 4'b0001;
										assign node13207 = (inp[8]) ? node13227 : node13208;
											assign node13208 = (inp[2]) ? node13222 : node13209;
												assign node13209 = (inp[5]) ? node13215 : node13210;
													assign node13210 = (inp[15]) ? 4'b0011 : node13211;
														assign node13211 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node13215 = (inp[1]) ? node13217 : 4'b0001;
														assign node13217 = (inp[15]) ? 4'b0001 : node13218;
															assign node13218 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node13222 = (inp[3]) ? node13224 : 4'b0011;
													assign node13224 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node13227 = (inp[15]) ? node13235 : node13228;
												assign node13228 = (inp[0]) ? node13230 : 4'b0010;
													assign node13230 = (inp[2]) ? node13232 : 4'b0000;
														assign node13232 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node13235 = (inp[0]) ? node13237 : 4'b0000;
													assign node13237 = (inp[5]) ? 4'b0000 : 4'b0010;
						assign node13240 = (inp[11]) ? node13572 : node13241;
							assign node13241 = (inp[6]) ? node13403 : node13242;
								assign node13242 = (inp[1]) ? node13334 : node13243;
									assign node13243 = (inp[7]) ? node13285 : node13244;
										assign node13244 = (inp[8]) ? node13270 : node13245;
											assign node13245 = (inp[14]) ? node13255 : node13246;
												assign node13246 = (inp[2]) ? node13250 : node13247;
													assign node13247 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node13250 = (inp[3]) ? 4'b1000 : node13251;
														assign node13251 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node13255 = (inp[0]) ? node13261 : node13256;
													assign node13256 = (inp[15]) ? node13258 : 4'b1010;
														assign node13258 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node13261 = (inp[15]) ? node13267 : node13262;
														assign node13262 = (inp[3]) ? node13264 : 4'b1000;
															assign node13264 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node13267 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node13270 = (inp[2]) ? node13276 : node13271;
												assign node13271 = (inp[14]) ? 4'b0011 : node13272;
													assign node13272 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node13276 = (inp[0]) ? node13282 : node13277;
													assign node13277 = (inp[3]) ? 4'b0001 : node13278;
														assign node13278 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node13282 = (inp[15]) ? 4'b0011 : 4'b0001;
										assign node13285 = (inp[8]) ? node13309 : node13286;
											assign node13286 = (inp[14]) ? node13298 : node13287;
												assign node13287 = (inp[2]) ? node13293 : node13288;
													assign node13288 = (inp[0]) ? 4'b1000 : node13289;
														assign node13289 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node13293 = (inp[15]) ? 4'b0001 : node13294;
														assign node13294 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node13298 = (inp[5]) ? node13304 : node13299;
													assign node13299 = (inp[3]) ? node13301 : 4'b0011;
														assign node13301 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node13304 = (inp[15]) ? 4'b0001 : node13305;
														assign node13305 = (inp[3]) ? 4'b0011 : 4'b0001;
											assign node13309 = (inp[2]) ? node13317 : node13310;
												assign node13310 = (inp[14]) ? node13314 : node13311;
													assign node13311 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node13314 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node13317 = (inp[14]) ? node13329 : node13318;
													assign node13318 = (inp[0]) ? node13324 : node13319;
														assign node13319 = (inp[15]) ? 4'b0000 : node13320;
															assign node13320 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node13324 = (inp[5]) ? 4'b0010 : node13325;
															assign node13325 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node13329 = (inp[3]) ? node13331 : 4'b0010;
														assign node13331 = (inp[15]) ? 4'b0010 : 4'b0000;
									assign node13334 = (inp[3]) ? node13354 : node13335;
										assign node13335 = (inp[0]) ? node13345 : node13336;
											assign node13336 = (inp[15]) ? node13342 : node13337;
												assign node13337 = (inp[8]) ? 4'b0010 : node13338;
													assign node13338 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node13342 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node13345 = (inp[15]) ? 4'b0010 : node13346;
												assign node13346 = (inp[14]) ? node13348 : 4'b0001;
													assign node13348 = (inp[7]) ? 4'b0000 : node13349;
														assign node13349 = (inp[8]) ? 4'b0001 : 4'b0000;
										assign node13354 = (inp[7]) ? node13378 : node13355;
											assign node13355 = (inp[14]) ? node13367 : node13356;
												assign node13356 = (inp[8]) ? node13360 : node13357;
													assign node13357 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node13360 = (inp[2]) ? 4'b0011 : node13361;
														assign node13361 = (inp[0]) ? 4'b0010 : node13362;
															assign node13362 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node13367 = (inp[8]) ? node13371 : node13368;
													assign node13368 = (inp[2]) ? 4'b0010 : 4'b0000;
													assign node13371 = (inp[15]) ? 4'b0011 : node13372;
														assign node13372 = (inp[5]) ? node13374 : 4'b0001;
															assign node13374 = (inp[2]) ? 4'b0001 : 4'b0011;
											assign node13378 = (inp[14]) ? node13396 : node13379;
												assign node13379 = (inp[15]) ? node13387 : node13380;
													assign node13380 = (inp[8]) ? 4'b0011 : node13381;
														assign node13381 = (inp[5]) ? 4'b0001 : node13382;
															assign node13382 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node13387 = (inp[8]) ? node13389 : 4'b0011;
														assign node13389 = (inp[0]) ? node13393 : node13390;
															assign node13390 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node13393 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node13396 = (inp[8]) ? node13398 : 4'b0011;
													assign node13398 = (inp[15]) ? node13400 : 4'b0000;
														assign node13400 = (inp[5]) ? 4'b0010 : 4'b0000;
								assign node13403 = (inp[1]) ? node13499 : node13404;
									assign node13404 = (inp[7]) ? node13446 : node13405;
										assign node13405 = (inp[8]) ? node13423 : node13406;
											assign node13406 = (inp[0]) ? node13410 : node13407;
												assign node13407 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node13410 = (inp[15]) ? 4'b0010 : node13411;
													assign node13411 = (inp[2]) ? node13417 : node13412;
														assign node13412 = (inp[3]) ? node13414 : 4'b0001;
															assign node13414 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node13417 = (inp[3]) ? node13419 : 4'b0000;
															assign node13419 = (inp[14]) ? 4'b0000 : 4'b0010;
											assign node13423 = (inp[14]) ? node13437 : node13424;
												assign node13424 = (inp[2]) ? node13428 : node13425;
													assign node13425 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node13428 = (inp[0]) ? node13432 : node13429;
														assign node13429 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node13432 = (inp[15]) ? node13434 : 4'b1111;
															assign node13434 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node13437 = (inp[0]) ? node13439 : 4'b1101;
													assign node13439 = (inp[15]) ? 4'b1101 : node13440;
														assign node13440 = (inp[5]) ? 4'b1111 : node13441;
															assign node13441 = (inp[3]) ? 4'b1111 : 4'b1101;
										assign node13446 = (inp[8]) ? node13478 : node13447;
											assign node13447 = (inp[14]) ? node13465 : node13448;
												assign node13448 = (inp[2]) ? node13454 : node13449;
													assign node13449 = (inp[15]) ? node13451 : 4'b0010;
														assign node13451 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node13454 = (inp[0]) ? node13460 : node13455;
														assign node13455 = (inp[5]) ? 4'b1101 : node13456;
															assign node13456 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node13460 = (inp[15]) ? 4'b1111 : node13461;
															assign node13461 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node13465 = (inp[15]) ? node13471 : node13466;
													assign node13466 = (inp[0]) ? node13468 : 4'b1101;
														assign node13468 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node13471 = (inp[0]) ? node13473 : 4'b1111;
														assign node13473 = (inp[3]) ? 4'b1101 : node13474;
															assign node13474 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node13478 = (inp[2]) ? node13494 : node13479;
												assign node13479 = (inp[14]) ? node13487 : node13480;
													assign node13480 = (inp[3]) ? node13484 : node13481;
														assign node13481 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node13484 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node13487 = (inp[0]) ? 4'b1100 : node13488;
														assign node13488 = (inp[15]) ? 4'b1110 : node13489;
															assign node13489 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node13494 = (inp[5]) ? node13496 : 4'b1100;
													assign node13496 = (inp[0]) ? 4'b1110 : 4'b1100;
									assign node13499 = (inp[5]) ? node13539 : node13500;
										assign node13500 = (inp[14]) ? node13522 : node13501;
											assign node13501 = (inp[15]) ? node13513 : node13502;
												assign node13502 = (inp[8]) ? 4'b1100 : node13503;
													assign node13503 = (inp[3]) ? node13507 : node13504;
														assign node13504 = (inp[2]) ? 4'b1100 : 4'b1110;
														assign node13507 = (inp[7]) ? node13509 : 4'b1110;
															assign node13509 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node13513 = (inp[2]) ? 4'b1101 : node13514;
													assign node13514 = (inp[3]) ? 4'b1111 : node13515;
														assign node13515 = (inp[0]) ? node13517 : 4'b1100;
															assign node13517 = (inp[7]) ? 4'b1110 : 4'b1110;
											assign node13522 = (inp[3]) ? node13532 : node13523;
												assign node13523 = (inp[2]) ? node13525 : 4'b1101;
													assign node13525 = (inp[0]) ? 4'b1100 : node13526;
														assign node13526 = (inp[15]) ? node13528 : 4'b1111;
															assign node13528 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node13532 = (inp[2]) ? 4'b1101 : node13533;
													assign node13533 = (inp[8]) ? 4'b1100 : node13534;
														assign node13534 = (inp[7]) ? 4'b1101 : 4'b1100;
										assign node13539 = (inp[8]) ? node13559 : node13540;
											assign node13540 = (inp[7]) ? node13544 : node13541;
												assign node13541 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node13544 = (inp[2]) ? node13548 : node13545;
													assign node13545 = (inp[14]) ? 4'b1111 : 4'b1100;
													assign node13548 = (inp[3]) ? node13554 : node13549;
														assign node13549 = (inp[0]) ? 4'b1111 : node13550;
															assign node13550 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node13554 = (inp[0]) ? node13556 : 4'b1101;
															assign node13556 = (inp[14]) ? 4'b1111 : 4'b1101;
											assign node13559 = (inp[3]) ? node13569 : node13560;
												assign node13560 = (inp[0]) ? 4'b1111 : node13561;
													assign node13561 = (inp[15]) ? 4'b1111 : node13562;
														assign node13562 = (inp[14]) ? 4'b1101 : node13563;
															assign node13563 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node13569 = (inp[7]) ? 4'b1110 : 4'b1111;
							assign node13572 = (inp[6]) ? node13732 : node13573;
								assign node13573 = (inp[1]) ? node13661 : node13574;
									assign node13574 = (inp[7]) ? node13614 : node13575;
										assign node13575 = (inp[8]) ? node13597 : node13576;
											assign node13576 = (inp[3]) ? node13584 : node13577;
												assign node13577 = (inp[5]) ? 4'b0010 : node13578;
													assign node13578 = (inp[0]) ? 4'b0010 : node13579;
														assign node13579 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node13584 = (inp[14]) ? node13592 : node13585;
													assign node13585 = (inp[2]) ? node13589 : node13586;
														assign node13586 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node13589 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node13592 = (inp[15]) ? 4'b0000 : node13593;
														assign node13593 = (inp[5]) ? 4'b0010 : 4'b0000;
											assign node13597 = (inp[2]) ? node13607 : node13598;
												assign node13598 = (inp[14]) ? 4'b1101 : node13599;
													assign node13599 = (inp[5]) ? node13601 : 4'b0010;
														assign node13601 = (inp[0]) ? node13603 : 4'b0010;
															assign node13603 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node13607 = (inp[14]) ? 4'b1111 : node13608;
													assign node13608 = (inp[5]) ? 4'b1101 : node13609;
														assign node13609 = (inp[0]) ? 4'b1111 : 4'b1101;
										assign node13614 = (inp[8]) ? node13636 : node13615;
											assign node13615 = (inp[14]) ? node13627 : node13616;
												assign node13616 = (inp[2]) ? node13624 : node13617;
													assign node13617 = (inp[15]) ? node13619 : 4'b0000;
														assign node13619 = (inp[5]) ? node13621 : 4'b0010;
															assign node13621 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node13624 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node13627 = (inp[0]) ? node13629 : 4'b1111;
													assign node13629 = (inp[5]) ? 4'b1101 : node13630;
														assign node13630 = (inp[15]) ? 4'b1111 : node13631;
															assign node13631 = (inp[3]) ? 4'b1111 : 4'b1101;
											assign node13636 = (inp[2]) ? node13650 : node13637;
												assign node13637 = (inp[14]) ? node13645 : node13638;
													assign node13638 = (inp[15]) ? node13642 : node13639;
														assign node13639 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node13642 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node13645 = (inp[3]) ? 4'b1110 : node13646;
														assign node13646 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node13650 = (inp[15]) ? 4'b1100 : node13651;
													assign node13651 = (inp[0]) ? node13655 : node13652;
														assign node13652 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node13655 = (inp[14]) ? 4'b1110 : node13656;
															assign node13656 = (inp[5]) ? 4'b1110 : 4'b1100;
									assign node13661 = (inp[14]) ? node13697 : node13662;
										assign node13662 = (inp[3]) ? node13684 : node13663;
											assign node13663 = (inp[5]) ? node13673 : node13664;
												assign node13664 = (inp[7]) ? 4'b1111 : node13665;
													assign node13665 = (inp[0]) ? node13667 : 4'b1110;
														assign node13667 = (inp[8]) ? 4'b1101 : node13668;
															assign node13668 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node13673 = (inp[8]) ? node13679 : node13674;
													assign node13674 = (inp[7]) ? node13676 : 4'b1110;
														assign node13676 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node13679 = (inp[0]) ? node13681 : 4'b1100;
														assign node13681 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node13684 = (inp[15]) ? node13694 : node13685;
												assign node13685 = (inp[0]) ? node13689 : node13686;
													assign node13686 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node13689 = (inp[7]) ? 4'b1111 : node13690;
														assign node13690 = (inp[5]) ? 4'b1111 : 4'b1110;
												assign node13694 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node13697 = (inp[8]) ? node13717 : node13698;
											assign node13698 = (inp[7]) ? node13710 : node13699;
												assign node13699 = (inp[15]) ? node13707 : node13700;
													assign node13700 = (inp[2]) ? node13702 : 4'b1100;
														assign node13702 = (inp[3]) ? 4'b1100 : node13703;
															assign node13703 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node13707 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node13710 = (inp[5]) ? 4'b1101 : node13711;
													assign node13711 = (inp[2]) ? 4'b1101 : node13712;
														assign node13712 = (inp[15]) ? 4'b1111 : 4'b1101;
											assign node13717 = (inp[7]) ? node13727 : node13718;
												assign node13718 = (inp[0]) ? 4'b1111 : node13719;
													assign node13719 = (inp[3]) ? 4'b1101 : node13720;
														assign node13720 = (inp[15]) ? 4'b1101 : node13721;
															assign node13721 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node13727 = (inp[0]) ? node13729 : 4'b1110;
													assign node13729 = (inp[15]) ? 4'b1100 : 4'b1110;
								assign node13732 = (inp[1]) ? node13818 : node13733;
									assign node13733 = (inp[7]) ? node13775 : node13734;
										assign node13734 = (inp[8]) ? node13752 : node13735;
											assign node13735 = (inp[14]) ? node13743 : node13736;
												assign node13736 = (inp[2]) ? node13738 : 4'b1101;
													assign node13738 = (inp[0]) ? 4'b1100 : node13739;
														assign node13739 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node13743 = (inp[15]) ? node13749 : node13744;
													assign node13744 = (inp[3]) ? 4'b1110 : node13745;
														assign node13745 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node13749 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node13752 = (inp[14]) ? node13764 : node13753;
												assign node13753 = (inp[2]) ? node13761 : node13754;
													assign node13754 = (inp[3]) ? 4'b1110 : node13755;
														assign node13755 = (inp[15]) ? 4'b1110 : node13756;
															assign node13756 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node13761 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node13764 = (inp[0]) ? node13768 : node13765;
													assign node13765 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node13768 = (inp[15]) ? node13770 : 4'b0111;
														assign node13770 = (inp[5]) ? 4'b0101 : node13771;
															assign node13771 = (inp[3]) ? 4'b0101 : 4'b0111;
										assign node13775 = (inp[8]) ? node13799 : node13776;
											assign node13776 = (inp[2]) ? node13784 : node13777;
												assign node13777 = (inp[14]) ? 4'b0101 : node13778;
													assign node13778 = (inp[3]) ? node13780 : 4'b1100;
														assign node13780 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node13784 = (inp[14]) ? node13794 : node13785;
													assign node13785 = (inp[5]) ? node13787 : 4'b0101;
														assign node13787 = (inp[0]) ? node13791 : node13788;
															assign node13788 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node13791 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node13794 = (inp[3]) ? 4'b0111 : node13795;
														assign node13795 = (inp[15]) ? 4'b0111 : 4'b0101;
											assign node13799 = (inp[14]) ? node13809 : node13800;
												assign node13800 = (inp[2]) ? node13804 : node13801;
													assign node13801 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node13804 = (inp[15]) ? node13806 : 4'b0100;
														assign node13806 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node13809 = (inp[0]) ? node13815 : node13810;
													assign node13810 = (inp[15]) ? 4'b0110 : node13811;
														assign node13811 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node13815 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node13818 = (inp[2]) ? node13850 : node13819;
										assign node13819 = (inp[0]) ? node13835 : node13820;
											assign node13820 = (inp[5]) ? node13830 : node13821;
												assign node13821 = (inp[15]) ? 4'b0101 : node13822;
													assign node13822 = (inp[7]) ? 4'b0111 : node13823;
														assign node13823 = (inp[14]) ? 4'b0110 : node13824;
															assign node13824 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node13830 = (inp[15]) ? 4'b0110 : node13831;
													assign node13831 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node13835 = (inp[8]) ? node13847 : node13836;
												assign node13836 = (inp[3]) ? node13840 : node13837;
													assign node13837 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node13840 = (inp[14]) ? node13844 : node13841;
														assign node13841 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node13844 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node13847 = (inp[7]) ? 4'b0111 : 4'b0110;
										assign node13850 = (inp[14]) ? node13876 : node13851;
											assign node13851 = (inp[15]) ? node13867 : node13852;
												assign node13852 = (inp[0]) ? node13862 : node13853;
													assign node13853 = (inp[5]) ? node13857 : node13854;
														assign node13854 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node13857 = (inp[7]) ? 4'b0100 : node13858;
															assign node13858 = (inp[3]) ? 4'b0101 : 4'b0100;
													assign node13862 = (inp[8]) ? node13864 : 4'b0101;
														assign node13864 = (inp[3]) ? 4'b0110 : 4'b0111;
												assign node13867 = (inp[5]) ? node13869 : 4'b0100;
													assign node13869 = (inp[0]) ? node13871 : 4'b0111;
														assign node13871 = (inp[7]) ? 4'b0100 : node13872;
															assign node13872 = (inp[8]) ? 4'b0101 : 4'b0100;
											assign node13876 = (inp[7]) ? node13886 : node13877;
												assign node13877 = (inp[15]) ? node13879 : 4'b0110;
													assign node13879 = (inp[0]) ? 4'b0100 : node13880;
														assign node13880 = (inp[3]) ? 4'b0110 : node13881;
															assign node13881 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node13886 = (inp[8]) ? node13890 : node13887;
													assign node13887 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node13890 = (inp[0]) ? 4'b0100 : 4'b0110;
				assign node13893 = (inp[9]) ? node15287 : node13894;
					assign node13894 = (inp[12]) ? node14584 : node13895;
						assign node13895 = (inp[7]) ? node14243 : node13896;
							assign node13896 = (inp[8]) ? node14068 : node13897;
								assign node13897 = (inp[2]) ? node13977 : node13898;
									assign node13898 = (inp[14]) ? node13952 : node13899;
										assign node13899 = (inp[3]) ? node13931 : node13900;
											assign node13900 = (inp[11]) ? node13912 : node13901;
												assign node13901 = (inp[5]) ? node13907 : node13902;
													assign node13902 = (inp[0]) ? 4'b0011 : node13903;
														assign node13903 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node13907 = (inp[6]) ? node13909 : 4'b0001;
														assign node13909 = (inp[1]) ? 4'b1001 : 4'b0001;
												assign node13912 = (inp[6]) ? node13922 : node13913;
													assign node13913 = (inp[1]) ? node13917 : node13914;
														assign node13914 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node13917 = (inp[15]) ? 4'b1001 : node13918;
															assign node13918 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node13922 = (inp[1]) ? node13926 : node13923;
														assign node13923 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node13926 = (inp[15]) ? 4'b0011 : node13927;
															assign node13927 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node13931 = (inp[5]) ? node13947 : node13932;
												assign node13932 = (inp[1]) ? node13938 : node13933;
													assign node13933 = (inp[11]) ? 4'b1001 : node13934;
														assign node13934 = (inp[6]) ? 4'b0011 : 4'b1001;
													assign node13938 = (inp[0]) ? node13942 : node13939;
														assign node13939 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node13942 = (inp[6]) ? node13944 : 4'b0001;
															assign node13944 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node13947 = (inp[6]) ? node13949 : 4'b1011;
													assign node13949 = (inp[1]) ? 4'b0011 : 4'b1011;
										assign node13952 = (inp[0]) ? node13970 : node13953;
											assign node13953 = (inp[15]) ? node13961 : node13954;
												assign node13954 = (inp[5]) ? node13958 : node13955;
													assign node13955 = (inp[1]) ? 4'b1010 : 4'b0010;
													assign node13958 = (inp[1]) ? 4'b0000 : 4'b1010;
												assign node13961 = (inp[6]) ? node13963 : 4'b1000;
													assign node13963 = (inp[5]) ? 4'b0000 : node13964;
														assign node13964 = (inp[11]) ? node13966 : 4'b0000;
															assign node13966 = (inp[1]) ? 4'b0000 : 4'b1000;
											assign node13970 = (inp[15]) ? node13972 : 4'b0000;
												assign node13972 = (inp[1]) ? 4'b0010 : node13973;
													assign node13973 = (inp[11]) ? 4'b1000 : 4'b0000;
									assign node13977 = (inp[5]) ? node14019 : node13978;
										assign node13978 = (inp[15]) ? node13996 : node13979;
											assign node13979 = (inp[0]) ? node13991 : node13980;
												assign node13980 = (inp[14]) ? node13982 : 4'b0010;
													assign node13982 = (inp[11]) ? 4'b0010 : node13983;
														assign node13983 = (inp[6]) ? node13987 : node13984;
															assign node13984 = (inp[1]) ? 4'b0010 : 4'b1010;
															assign node13987 = (inp[1]) ? 4'b1010 : 4'b0010;
												assign node13991 = (inp[11]) ? node13993 : 4'b0000;
													assign node13993 = (inp[14]) ? 4'b1000 : 4'b0000;
											assign node13996 = (inp[0]) ? node14006 : node13997;
												assign node13997 = (inp[6]) ? node14001 : node13998;
													assign node13998 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node14001 = (inp[14]) ? node14003 : 4'b1000;
														assign node14003 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node14006 = (inp[6]) ? 4'b0010 : node14007;
													assign node14007 = (inp[3]) ? node14011 : node14008;
														assign node14008 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node14011 = (inp[14]) ? node14015 : node14012;
															assign node14012 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node14015 = (inp[1]) ? 4'b0010 : 4'b0010;
										assign node14019 = (inp[15]) ? node14039 : node14020;
											assign node14020 = (inp[3]) ? node14028 : node14021;
												assign node14021 = (inp[0]) ? node14023 : 4'b1010;
													assign node14023 = (inp[14]) ? node14025 : 4'b1000;
														assign node14025 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node14028 = (inp[0]) ? node14034 : node14029;
													assign node14029 = (inp[6]) ? 4'b1000 : node14030;
														assign node14030 = (inp[14]) ? 4'b1000 : 4'b0000;
													assign node14034 = (inp[11]) ? node14036 : 4'b1010;
														assign node14036 = (inp[1]) ? 4'b0010 : 4'b1010;
											assign node14039 = (inp[1]) ? node14053 : node14040;
												assign node14040 = (inp[11]) ? node14048 : node14041;
													assign node14041 = (inp[6]) ? 4'b0000 : node14042;
														assign node14042 = (inp[3]) ? 4'b1000 : node14043;
															assign node14043 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node14048 = (inp[6]) ? node14050 : 4'b0010;
														assign node14050 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node14053 = (inp[11]) ? node14061 : node14054;
													assign node14054 = (inp[6]) ? 4'b1010 : node14055;
														assign node14055 = (inp[0]) ? 4'b0010 : node14056;
															assign node14056 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node14061 = (inp[6]) ? node14063 : 4'b1000;
														assign node14063 = (inp[14]) ? 4'b0000 : node14064;
															assign node14064 = (inp[3]) ? 4'b0000 : 4'b0010;
								assign node14068 = (inp[2]) ? node14146 : node14069;
									assign node14069 = (inp[14]) ? node14109 : node14070;
										assign node14070 = (inp[15]) ? node14086 : node14071;
											assign node14071 = (inp[0]) ? node14083 : node14072;
												assign node14072 = (inp[1]) ? node14078 : node14073;
													assign node14073 = (inp[11]) ? 4'b1010 : node14074;
														assign node14074 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node14078 = (inp[3]) ? 4'b0010 : node14079;
														assign node14079 = (inp[6]) ? 4'b1010 : 4'b0010;
												assign node14083 = (inp[3]) ? 4'b1010 : 4'b1000;
											assign node14086 = (inp[0]) ? node14104 : node14087;
												assign node14087 = (inp[6]) ? node14093 : node14088;
													assign node14088 = (inp[1]) ? 4'b1000 : node14089;
														assign node14089 = (inp[3]) ? 4'b1000 : 4'b0000;
													assign node14093 = (inp[5]) ? node14101 : node14094;
														assign node14094 = (inp[3]) ? node14098 : node14095;
															assign node14095 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node14098 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node14101 = (inp[3]) ? 4'b0010 : 4'b1000;
												assign node14104 = (inp[3]) ? node14106 : 4'b1010;
													assign node14106 = (inp[11]) ? 4'b1000 : 4'b0010;
										assign node14109 = (inp[15]) ? node14121 : node14110;
											assign node14110 = (inp[0]) ? node14116 : node14111;
												assign node14111 = (inp[3]) ? node14113 : 4'b0011;
													assign node14113 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node14116 = (inp[6]) ? 4'b0001 : node14117;
													assign node14117 = (inp[11]) ? 4'b1001 : 4'b0001;
											assign node14121 = (inp[6]) ? node14133 : node14122;
												assign node14122 = (inp[11]) ? node14128 : node14123;
													assign node14123 = (inp[3]) ? 4'b0001 : node14124;
														assign node14124 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node14128 = (inp[1]) ? node14130 : 4'b1001;
														assign node14130 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node14133 = (inp[11]) ? node14143 : node14134;
													assign node14134 = (inp[3]) ? node14138 : node14135;
														assign node14135 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node14138 = (inp[0]) ? 4'b1001 : node14139;
															assign node14139 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node14143 = (inp[0]) ? 4'b0011 : 4'b0001;
									assign node14146 = (inp[14]) ? node14194 : node14147;
										assign node14147 = (inp[5]) ? node14173 : node14148;
											assign node14148 = (inp[11]) ? node14164 : node14149;
												assign node14149 = (inp[6]) ? node14159 : node14150;
													assign node14150 = (inp[1]) ? node14152 : 4'b0011;
														assign node14152 = (inp[15]) ? node14156 : node14153;
															assign node14153 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node14156 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node14159 = (inp[1]) ? 4'b1011 : node14160;
														assign node14160 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node14164 = (inp[6]) ? node14170 : node14165;
													assign node14165 = (inp[1]) ? node14167 : 4'b1001;
														assign node14167 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node14170 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node14173 = (inp[3]) ? node14185 : node14174;
												assign node14174 = (inp[15]) ? node14180 : node14175;
													assign node14175 = (inp[6]) ? node14177 : 4'b0011;
														assign node14177 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node14180 = (inp[0]) ? 4'b0011 : node14181;
														assign node14181 = (inp[6]) ? 4'b1001 : 4'b0001;
												assign node14185 = (inp[6]) ? node14189 : node14186;
													assign node14186 = (inp[11]) ? 4'b1001 : 4'b0001;
													assign node14189 = (inp[15]) ? 4'b0011 : node14190;
														assign node14190 = (inp[11]) ? 4'b0001 : 4'b1001;
										assign node14194 = (inp[1]) ? node14220 : node14195;
											assign node14195 = (inp[15]) ? node14207 : node14196;
												assign node14196 = (inp[0]) ? node14202 : node14197;
													assign node14197 = (inp[3]) ? node14199 : 4'b0011;
														assign node14199 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node14202 = (inp[3]) ? 4'b1011 : node14203;
														assign node14203 = (inp[5]) ? 4'b0001 : 4'b1001;
												assign node14207 = (inp[0]) ? node14213 : node14208;
													assign node14208 = (inp[3]) ? node14210 : 4'b1001;
														assign node14210 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node14213 = (inp[6]) ? node14217 : node14214;
														assign node14214 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node14217 = (inp[5]) ? 4'b1001 : 4'b0011;
											assign node14220 = (inp[5]) ? node14234 : node14221;
												assign node14221 = (inp[3]) ? node14227 : node14222;
													assign node14222 = (inp[0]) ? node14224 : 4'b1001;
														assign node14224 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node14227 = (inp[6]) ? node14231 : node14228;
														assign node14228 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node14231 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node14234 = (inp[0]) ? node14236 : 4'b1011;
													assign node14236 = (inp[11]) ? node14238 : 4'b1001;
														assign node14238 = (inp[6]) ? 4'b0011 : node14239;
															assign node14239 = (inp[15]) ? 4'b1001 : 4'b1011;
							assign node14243 = (inp[8]) ? node14393 : node14244;
								assign node14244 = (inp[14]) ? node14318 : node14245;
									assign node14245 = (inp[2]) ? node14289 : node14246;
										assign node14246 = (inp[3]) ? node14274 : node14247;
											assign node14247 = (inp[6]) ? node14265 : node14248;
												assign node14248 = (inp[15]) ? node14256 : node14249;
													assign node14249 = (inp[0]) ? 4'b1000 : node14250;
														assign node14250 = (inp[11]) ? node14252 : 4'b1010;
															assign node14252 = (inp[1]) ? 4'b1010 : 4'b0010;
													assign node14256 = (inp[0]) ? 4'b0010 : node14257;
														assign node14257 = (inp[5]) ? node14261 : node14258;
															assign node14258 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node14261 = (inp[11]) ? 4'b1000 : 4'b0000;
												assign node14265 = (inp[15]) ? node14271 : node14266;
													assign node14266 = (inp[1]) ? node14268 : 4'b1000;
														assign node14268 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node14271 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node14274 = (inp[1]) ? node14282 : node14275;
												assign node14275 = (inp[15]) ? 4'b0010 : node14276;
													assign node14276 = (inp[0]) ? node14278 : 4'b0010;
														assign node14278 = (inp[11]) ? 4'b0010 : 4'b1010;
												assign node14282 = (inp[5]) ? node14286 : node14283;
													assign node14283 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node14286 = (inp[15]) ? 4'b1010 : 4'b0010;
										assign node14289 = (inp[15]) ? node14305 : node14290;
											assign node14290 = (inp[0]) ? node14298 : node14291;
												assign node14291 = (inp[5]) ? node14295 : node14292;
													assign node14292 = (inp[3]) ? 4'b1011 : 4'b0011;
													assign node14295 = (inp[3]) ? 4'b0001 : 4'b1011;
												assign node14298 = (inp[11]) ? node14300 : 4'b1001;
													assign node14300 = (inp[6]) ? node14302 : 4'b1001;
														assign node14302 = (inp[3]) ? 4'b0011 : 4'b0001;
											assign node14305 = (inp[11]) ? node14309 : node14306;
												assign node14306 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node14309 = (inp[6]) ? 4'b0011 : node14310;
													assign node14310 = (inp[5]) ? node14312 : 4'b1011;
														assign node14312 = (inp[3]) ? node14314 : 4'b1001;
															assign node14314 = (inp[0]) ? 4'b1001 : 4'b1011;
									assign node14318 = (inp[1]) ? node14354 : node14319;
										assign node14319 = (inp[6]) ? node14341 : node14320;
											assign node14320 = (inp[11]) ? node14334 : node14321;
												assign node14321 = (inp[2]) ? node14331 : node14322;
													assign node14322 = (inp[15]) ? node14324 : 4'b0011;
														assign node14324 = (inp[3]) ? node14328 : node14325;
															assign node14325 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node14328 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node14331 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node14334 = (inp[3]) ? 4'b1011 : node14335;
													assign node14335 = (inp[15]) ? node14337 : 4'b1001;
														assign node14337 = (inp[0]) ? 4'b1011 : 4'b1001;
											assign node14341 = (inp[11]) ? node14351 : node14342;
												assign node14342 = (inp[5]) ? node14344 : 4'b1011;
													assign node14344 = (inp[2]) ? 4'b1001 : node14345;
														assign node14345 = (inp[0]) ? 4'b1011 : node14346;
															assign node14346 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node14351 = (inp[0]) ? 4'b0011 : 4'b0001;
										assign node14354 = (inp[0]) ? node14370 : node14355;
											assign node14355 = (inp[5]) ? node14361 : node14356;
												assign node14356 = (inp[6]) ? node14358 : 4'b1011;
													assign node14358 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node14361 = (inp[11]) ? node14363 : 4'b0011;
													assign node14363 = (inp[6]) ? node14365 : 4'b1001;
														assign node14365 = (inp[15]) ? 4'b0011 : node14366;
															assign node14366 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node14370 = (inp[15]) ? node14388 : node14371;
												assign node14371 = (inp[2]) ? node14385 : node14372;
													assign node14372 = (inp[5]) ? node14380 : node14373;
														assign node14373 = (inp[6]) ? node14377 : node14374;
															assign node14374 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node14377 = (inp[3]) ? 4'b1001 : 4'b0001;
														assign node14380 = (inp[6]) ? 4'b0001 : node14381;
															assign node14381 = (inp[11]) ? 4'b1001 : 4'b0001;
													assign node14385 = (inp[11]) ? 4'b0011 : 4'b0001;
												assign node14388 = (inp[6]) ? node14390 : 4'b1011;
													assign node14390 = (inp[5]) ? 4'b0001 : 4'b0011;
								assign node14393 = (inp[2]) ? node14473 : node14394;
									assign node14394 = (inp[14]) ? node14432 : node14395;
										assign node14395 = (inp[5]) ? node14415 : node14396;
											assign node14396 = (inp[0]) ? node14408 : node14397;
												assign node14397 = (inp[15]) ? node14403 : node14398;
													assign node14398 = (inp[1]) ? node14400 : 4'b0011;
														assign node14400 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node14403 = (inp[11]) ? node14405 : 4'b0001;
														assign node14405 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node14408 = (inp[15]) ? node14410 : 4'b0001;
													assign node14410 = (inp[6]) ? node14412 : 4'b0011;
														assign node14412 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node14415 = (inp[6]) ? node14421 : node14416;
												assign node14416 = (inp[11]) ? 4'b1001 : node14417;
													assign node14417 = (inp[1]) ? 4'b0011 : 4'b0001;
												assign node14421 = (inp[11]) ? node14423 : 4'b1011;
													assign node14423 = (inp[1]) ? 4'b0001 : node14424;
														assign node14424 = (inp[3]) ? node14428 : node14425;
															assign node14425 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node14428 = (inp[0]) ? 4'b0001 : 4'b0011;
										assign node14432 = (inp[5]) ? node14452 : node14433;
											assign node14433 = (inp[15]) ? node14441 : node14434;
												assign node14434 = (inp[6]) ? node14438 : node14435;
													assign node14435 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node14438 = (inp[11]) ? 4'b0010 : 4'b1010;
												assign node14441 = (inp[0]) ? node14447 : node14442;
													assign node14442 = (inp[11]) ? node14444 : 4'b1000;
														assign node14444 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node14447 = (inp[3]) ? 4'b1010 : node14448;
														assign node14448 = (inp[6]) ? 4'b0010 : 4'b1010;
											assign node14452 = (inp[15]) ? node14464 : node14453;
												assign node14453 = (inp[1]) ? node14455 : 4'b0000;
													assign node14455 = (inp[0]) ? node14459 : node14456;
														assign node14456 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node14459 = (inp[3]) ? node14461 : 4'b1000;
															assign node14461 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node14464 = (inp[1]) ? 4'b0010 : node14465;
													assign node14465 = (inp[6]) ? 4'b1010 : node14466;
														assign node14466 = (inp[0]) ? 4'b0000 : node14467;
															assign node14467 = (inp[11]) ? 4'b1010 : 4'b0010;
									assign node14473 = (inp[1]) ? node14533 : node14474;
										assign node14474 = (inp[5]) ? node14502 : node14475;
											assign node14475 = (inp[6]) ? node14487 : node14476;
												assign node14476 = (inp[11]) ? 4'b1010 : node14477;
													assign node14477 = (inp[14]) ? node14479 : 4'b0010;
														assign node14479 = (inp[15]) ? node14483 : node14480;
															assign node14480 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node14483 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node14487 = (inp[11]) ? node14495 : node14488;
													assign node14488 = (inp[0]) ? node14492 : node14489;
														assign node14489 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node14492 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node14495 = (inp[15]) ? node14499 : node14496;
														assign node14496 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node14499 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node14502 = (inp[0]) ? node14520 : node14503;
												assign node14503 = (inp[6]) ? node14509 : node14504;
													assign node14504 = (inp[11]) ? node14506 : 4'b0000;
														assign node14506 = (inp[14]) ? 4'b1000 : 4'b1010;
													assign node14509 = (inp[14]) ? node14515 : node14510;
														assign node14510 = (inp[3]) ? node14512 : 4'b1010;
															assign node14512 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node14515 = (inp[3]) ? node14517 : 4'b1000;
															assign node14517 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node14520 = (inp[6]) ? node14526 : node14521;
													assign node14521 = (inp[15]) ? node14523 : 4'b0010;
														assign node14523 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node14526 = (inp[11]) ? node14528 : 4'b1000;
														assign node14528 = (inp[15]) ? 4'b0000 : node14529;
															assign node14529 = (inp[3]) ? 4'b0010 : 4'b0000;
										assign node14533 = (inp[11]) ? node14559 : node14534;
											assign node14534 = (inp[6]) ? node14552 : node14535;
												assign node14535 = (inp[14]) ? node14543 : node14536;
													assign node14536 = (inp[3]) ? node14538 : 4'b0010;
														assign node14538 = (inp[5]) ? node14540 : 4'b0000;
															assign node14540 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node14543 = (inp[3]) ? node14549 : node14544;
														assign node14544 = (inp[5]) ? 4'b0000 : node14545;
															assign node14545 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node14549 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node14552 = (inp[3]) ? 4'b1010 : node14553;
													assign node14553 = (inp[15]) ? node14555 : 4'b1010;
														assign node14555 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node14559 = (inp[6]) ? node14573 : node14560;
												assign node14560 = (inp[3]) ? node14566 : node14561;
													assign node14561 = (inp[5]) ? 4'b1000 : node14562;
														assign node14562 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node14566 = (inp[14]) ? 4'b1010 : node14567;
														assign node14567 = (inp[15]) ? 4'b1010 : node14568;
															assign node14568 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node14573 = (inp[5]) ? node14575 : 4'b0000;
													assign node14575 = (inp[14]) ? node14579 : node14576;
														assign node14576 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node14579 = (inp[15]) ? node14581 : 4'b0000;
															assign node14581 = (inp[0]) ? 4'b0000 : 4'b0000;
						assign node14584 = (inp[6]) ? node14946 : node14585;
							assign node14585 = (inp[11]) ? node14765 : node14586;
								assign node14586 = (inp[1]) ? node14680 : node14587;
									assign node14587 = (inp[7]) ? node14633 : node14588;
										assign node14588 = (inp[8]) ? node14608 : node14589;
											assign node14589 = (inp[14]) ? node14599 : node14590;
												assign node14590 = (inp[2]) ? node14594 : node14591;
													assign node14591 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node14594 = (inp[0]) ? node14596 : 4'b1000;
														assign node14596 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node14599 = (inp[3]) ? 4'b1010 : node14600;
													assign node14600 = (inp[0]) ? node14604 : node14601;
														assign node14601 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node14604 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node14608 = (inp[2]) ? node14618 : node14609;
												assign node14609 = (inp[14]) ? 4'b0011 : node14610;
													assign node14610 = (inp[0]) ? 4'b1010 : node14611;
														assign node14611 = (inp[5]) ? node14613 : 4'b1000;
															assign node14613 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node14618 = (inp[3]) ? node14624 : node14619;
													assign node14619 = (inp[15]) ? 4'b0001 : node14620;
														assign node14620 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node14624 = (inp[15]) ? 4'b0011 : node14625;
														assign node14625 = (inp[14]) ? node14629 : node14626;
															assign node14626 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node14629 = (inp[0]) ? 4'b0001 : 4'b0001;
										assign node14633 = (inp[8]) ? node14661 : node14634;
											assign node14634 = (inp[2]) ? node14648 : node14635;
												assign node14635 = (inp[14]) ? node14643 : node14636;
													assign node14636 = (inp[15]) ? node14638 : 4'b1010;
														assign node14638 = (inp[5]) ? 4'b1000 : node14639;
															assign node14639 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node14643 = (inp[15]) ? node14645 : 4'b0001;
														assign node14645 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node14648 = (inp[5]) ? node14656 : node14649;
													assign node14649 = (inp[14]) ? 4'b0011 : node14650;
														assign node14650 = (inp[15]) ? node14652 : 4'b0001;
															assign node14652 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node14656 = (inp[0]) ? node14658 : 4'b0001;
														assign node14658 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node14661 = (inp[2]) ? node14671 : node14662;
												assign node14662 = (inp[14]) ? 4'b0010 : node14663;
													assign node14663 = (inp[3]) ? node14667 : node14664;
														assign node14664 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node14667 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node14671 = (inp[5]) ? 4'b0010 : node14672;
													assign node14672 = (inp[14]) ? 4'b0000 : node14673;
														assign node14673 = (inp[0]) ? 4'b0000 : node14674;
															assign node14674 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node14680 = (inp[3]) ? node14722 : node14681;
										assign node14681 = (inp[0]) ? node14705 : node14682;
											assign node14682 = (inp[15]) ? node14692 : node14683;
												assign node14683 = (inp[5]) ? node14685 : 4'b0011;
													assign node14685 = (inp[8]) ? node14687 : 4'b0010;
														assign node14687 = (inp[2]) ? 4'b0011 : node14688;
															assign node14688 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node14692 = (inp[2]) ? node14702 : node14693;
													assign node14693 = (inp[7]) ? node14695 : 4'b0000;
														assign node14695 = (inp[14]) ? node14699 : node14696;
															assign node14696 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node14699 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node14702 = (inp[5]) ? 4'b0001 : 4'b0000;
											assign node14705 = (inp[15]) ? node14713 : node14706;
												assign node14706 = (inp[8]) ? node14708 : 4'b0001;
													assign node14708 = (inp[2]) ? 4'b0001 : node14709;
														assign node14709 = (inp[14]) ? 4'b0001 : 4'b0000;
												assign node14713 = (inp[2]) ? 4'b0011 : node14714;
													assign node14714 = (inp[5]) ? node14716 : 4'b0010;
														assign node14716 = (inp[8]) ? 4'b0011 : node14717;
															assign node14717 = (inp[14]) ? 4'b0011 : 4'b0010;
										assign node14722 = (inp[14]) ? node14750 : node14723;
											assign node14723 = (inp[7]) ? node14739 : node14724;
												assign node14724 = (inp[2]) ? node14732 : node14725;
													assign node14725 = (inp[8]) ? node14727 : 4'b0011;
														assign node14727 = (inp[15]) ? 4'b0010 : node14728;
															assign node14728 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node14732 = (inp[8]) ? 4'b0011 : node14733;
														assign node14733 = (inp[0]) ? 4'b0000 : node14734;
															assign node14734 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node14739 = (inp[0]) ? 4'b0000 : node14740;
													assign node14740 = (inp[8]) ? node14746 : node14741;
														assign node14741 = (inp[2]) ? 4'b0001 : node14742;
															assign node14742 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node14746 = (inp[15]) ? 4'b0010 : 4'b0001;
											assign node14750 = (inp[2]) ? node14758 : node14751;
												assign node14751 = (inp[0]) ? 4'b0000 : node14752;
													assign node14752 = (inp[5]) ? 4'b0011 : node14753;
														assign node14753 = (inp[7]) ? 4'b0000 : 4'b0010;
												assign node14758 = (inp[7]) ? node14762 : node14759;
													assign node14759 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node14762 = (inp[8]) ? 4'b0010 : 4'b0011;
								assign node14765 = (inp[1]) ? node14857 : node14766;
									assign node14766 = (inp[7]) ? node14802 : node14767;
										assign node14767 = (inp[8]) ? node14785 : node14768;
											assign node14768 = (inp[14]) ? node14778 : node14769;
												assign node14769 = (inp[2]) ? 4'b0000 : node14770;
													assign node14770 = (inp[15]) ? 4'b0001 : node14771;
														assign node14771 = (inp[3]) ? node14773 : 4'b0011;
															assign node14773 = (inp[5]) ? 4'b0001 : 4'b0001;
												assign node14778 = (inp[3]) ? 4'b0010 : node14779;
													assign node14779 = (inp[5]) ? node14781 : 4'b0000;
														assign node14781 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node14785 = (inp[14]) ? node14795 : node14786;
												assign node14786 = (inp[2]) ? 4'b1111 : node14787;
													assign node14787 = (inp[15]) ? 4'b0000 : node14788;
														assign node14788 = (inp[0]) ? node14790 : 4'b0010;
															assign node14790 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node14795 = (inp[0]) ? 4'b1111 : node14796;
													assign node14796 = (inp[5]) ? 4'b1101 : node14797;
														assign node14797 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node14802 = (inp[8]) ? node14830 : node14803;
											assign node14803 = (inp[2]) ? node14817 : node14804;
												assign node14804 = (inp[14]) ? node14810 : node14805;
													assign node14805 = (inp[0]) ? 4'b0000 : node14806;
														assign node14806 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node14810 = (inp[3]) ? node14812 : 4'b1101;
														assign node14812 = (inp[15]) ? node14814 : 4'b1111;
															assign node14814 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node14817 = (inp[5]) ? 4'b1101 : node14818;
													assign node14818 = (inp[3]) ? node14824 : node14819;
														assign node14819 = (inp[15]) ? 4'b1101 : node14820;
															assign node14820 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node14824 = (inp[0]) ? node14826 : 4'b1111;
															assign node14826 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node14830 = (inp[14]) ? node14842 : node14831;
												assign node14831 = (inp[2]) ? node14835 : node14832;
													assign node14832 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node14835 = (inp[15]) ? node14837 : 4'b1110;
														assign node14837 = (inp[0]) ? 4'b1100 : node14838;
															assign node14838 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node14842 = (inp[3]) ? node14848 : node14843;
													assign node14843 = (inp[15]) ? 4'b1110 : node14844;
														assign node14844 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node14848 = (inp[5]) ? node14852 : node14849;
														assign node14849 = (inp[2]) ? 4'b1110 : 4'b1100;
														assign node14852 = (inp[15]) ? node14854 : 4'b1100;
															assign node14854 = (inp[0]) ? 4'b1100 : 4'b1110;
									assign node14857 = (inp[7]) ? node14903 : node14858;
										assign node14858 = (inp[8]) ? node14880 : node14859;
											assign node14859 = (inp[14]) ? node14869 : node14860;
												assign node14860 = (inp[2]) ? node14864 : node14861;
													assign node14861 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node14864 = (inp[3]) ? 4'b1110 : node14865;
														assign node14865 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node14869 = (inp[15]) ? 4'b1110 : node14870;
													assign node14870 = (inp[0]) ? node14876 : node14871;
														assign node14871 = (inp[3]) ? 4'b1100 : node14872;
															assign node14872 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node14876 = (inp[3]) ? 4'b1110 : 4'b1100;
											assign node14880 = (inp[2]) ? node14896 : node14881;
												assign node14881 = (inp[14]) ? node14889 : node14882;
													assign node14882 = (inp[15]) ? node14886 : node14883;
														assign node14883 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node14886 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node14889 = (inp[15]) ? node14891 : 4'b1101;
														assign node14891 = (inp[5]) ? 4'b1111 : node14892;
															assign node14892 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node14896 = (inp[15]) ? node14898 : 4'b1111;
													assign node14898 = (inp[0]) ? node14900 : 4'b1111;
														assign node14900 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node14903 = (inp[8]) ? node14927 : node14904;
											assign node14904 = (inp[14]) ? node14918 : node14905;
												assign node14905 = (inp[2]) ? node14913 : node14906;
													assign node14906 = (inp[5]) ? 4'b1110 : node14907;
														assign node14907 = (inp[0]) ? 4'b1100 : node14908;
															assign node14908 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node14913 = (inp[15]) ? 4'b1101 : node14914;
														assign node14914 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node14918 = (inp[0]) ? 4'b1101 : node14919;
													assign node14919 = (inp[15]) ? 4'b1111 : node14920;
														assign node14920 = (inp[3]) ? 4'b1101 : node14921;
															assign node14921 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node14927 = (inp[14]) ? node14935 : node14928;
												assign node14928 = (inp[2]) ? node14932 : node14929;
													assign node14929 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node14932 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node14935 = (inp[0]) ? node14941 : node14936;
													assign node14936 = (inp[15]) ? node14938 : 4'b1100;
														assign node14938 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node14941 = (inp[15]) ? node14943 : 4'b1110;
														assign node14943 = (inp[3]) ? 4'b1100 : 4'b1110;
							assign node14946 = (inp[11]) ? node15136 : node14947;
								assign node14947 = (inp[1]) ? node15029 : node14948;
									assign node14948 = (inp[2]) ? node14996 : node14949;
										assign node14949 = (inp[8]) ? node14967 : node14950;
											assign node14950 = (inp[15]) ? node14962 : node14951;
												assign node14951 = (inp[7]) ? node14957 : node14952;
													assign node14952 = (inp[14]) ? 4'b0010 : node14953;
														assign node14953 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node14957 = (inp[14]) ? 4'b1101 : node14958;
														assign node14958 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node14962 = (inp[14]) ? node14964 : 4'b0000;
													assign node14964 = (inp[7]) ? 4'b1111 : 4'b0000;
											assign node14967 = (inp[7]) ? node14979 : node14968;
												assign node14968 = (inp[14]) ? node14976 : node14969;
													assign node14969 = (inp[5]) ? 4'b0010 : node14970;
														assign node14970 = (inp[15]) ? node14972 : 4'b0000;
															assign node14972 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node14976 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node14979 = (inp[14]) ? node14991 : node14980;
													assign node14980 = (inp[3]) ? node14986 : node14981;
														assign node14981 = (inp[5]) ? node14983 : 4'b1111;
															assign node14983 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node14986 = (inp[15]) ? node14988 : 4'b1101;
															assign node14988 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node14991 = (inp[3]) ? 4'b1110 : node14992;
														assign node14992 = (inp[5]) ? 4'b1110 : 4'b1100;
										assign node14996 = (inp[8]) ? node15010 : node14997;
											assign node14997 = (inp[7]) ? node14999 : 4'b0010;
												assign node14999 = (inp[3]) ? node15005 : node15000;
													assign node15000 = (inp[0]) ? node15002 : 4'b1111;
														assign node15002 = (inp[14]) ? 4'b1111 : 4'b1101;
													assign node15005 = (inp[15]) ? 4'b1101 : node15006;
														assign node15006 = (inp[0]) ? 4'b1111 : 4'b1101;
											assign node15010 = (inp[7]) ? node15022 : node15011;
												assign node15011 = (inp[15]) ? 4'b1111 : node15012;
													assign node15012 = (inp[3]) ? 4'b1101 : node15013;
														assign node15013 = (inp[0]) ? node15017 : node15014;
															assign node15014 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node15017 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node15022 = (inp[14]) ? 4'b1100 : node15023;
													assign node15023 = (inp[15]) ? 4'b1110 : node15024;
														assign node15024 = (inp[3]) ? 4'b1110 : 4'b1100;
									assign node15029 = (inp[3]) ? node15079 : node15030;
										assign node15030 = (inp[15]) ? node15050 : node15031;
											assign node15031 = (inp[0]) ? node15043 : node15032;
												assign node15032 = (inp[5]) ? node15034 : 4'b1110;
													assign node15034 = (inp[7]) ? node15036 : 4'b1100;
														assign node15036 = (inp[2]) ? node15040 : node15037;
															assign node15037 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node15040 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node15043 = (inp[5]) ? node15045 : 4'b1101;
													assign node15045 = (inp[14]) ? node15047 : 4'b1111;
														assign node15047 = (inp[7]) ? 4'b1111 : 4'b1110;
											assign node15050 = (inp[8]) ? node15060 : node15051;
												assign node15051 = (inp[2]) ? 4'b1111 : node15052;
													assign node15052 = (inp[7]) ? node15054 : 4'b1111;
														assign node15054 = (inp[14]) ? node15056 : 4'b1100;
															assign node15056 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node15060 = (inp[7]) ? node15068 : node15061;
													assign node15061 = (inp[2]) ? node15063 : 4'b1110;
														assign node15063 = (inp[0]) ? node15065 : 4'b1111;
															assign node15065 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node15068 = (inp[2]) ? node15074 : node15069;
														assign node15069 = (inp[0]) ? 4'b1111 : node15070;
															assign node15070 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node15074 = (inp[5]) ? node15076 : 4'b1110;
															assign node15076 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node15079 = (inp[14]) ? node15109 : node15080;
											assign node15080 = (inp[7]) ? node15094 : node15081;
												assign node15081 = (inp[8]) ? node15091 : node15082;
													assign node15082 = (inp[2]) ? node15084 : 4'b1101;
														assign node15084 = (inp[0]) ? node15088 : node15085;
															assign node15085 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node15088 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node15091 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node15094 = (inp[8]) ? node15106 : node15095;
													assign node15095 = (inp[2]) ? node15101 : node15096;
														assign node15096 = (inp[0]) ? node15098 : 4'b1100;
															assign node15098 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node15101 = (inp[0]) ? 4'b1101 : node15102;
															assign node15102 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node15106 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node15109 = (inp[15]) ? node15123 : node15110;
												assign node15110 = (inp[0]) ? node15118 : node15111;
													assign node15111 = (inp[5]) ? 4'b1101 : node15112;
														assign node15112 = (inp[8]) ? node15114 : 4'b1100;
															assign node15114 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node15118 = (inp[8]) ? node15120 : 4'b1111;
														assign node15120 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node15123 = (inp[0]) ? node15129 : node15124;
													assign node15124 = (inp[7]) ? node15126 : 4'b1110;
														assign node15126 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node15129 = (inp[7]) ? node15133 : node15130;
														assign node15130 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node15133 = (inp[8]) ? 4'b1100 : 4'b1101;
								assign node15136 = (inp[1]) ? node15214 : node15137;
									assign node15137 = (inp[7]) ? node15173 : node15138;
										assign node15138 = (inp[8]) ? node15160 : node15139;
											assign node15139 = (inp[2]) ? node15153 : node15140;
												assign node15140 = (inp[14]) ? node15148 : node15141;
													assign node15141 = (inp[5]) ? 4'b1111 : node15142;
														assign node15142 = (inp[3]) ? 4'b1101 : node15143;
															assign node15143 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node15148 = (inp[0]) ? node15150 : 4'b1110;
														assign node15150 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node15153 = (inp[3]) ? node15155 : 4'b1110;
													assign node15155 = (inp[0]) ? node15157 : 4'b1100;
														assign node15157 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node15160 = (inp[14]) ? node15166 : node15161;
												assign node15161 = (inp[2]) ? node15163 : 4'b1100;
													assign node15163 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node15166 = (inp[3]) ? node15168 : 4'b0111;
													assign node15168 = (inp[0]) ? 4'b0101 : node15169;
														assign node15169 = (inp[15]) ? 4'b0111 : 4'b0101;
										assign node15173 = (inp[8]) ? node15189 : node15174;
											assign node15174 = (inp[0]) ? node15180 : node15175;
												assign node15175 = (inp[15]) ? 4'b0111 : node15176;
													assign node15176 = (inp[14]) ? 4'b0111 : 4'b0101;
												assign node15180 = (inp[14]) ? node15182 : 4'b1100;
													assign node15182 = (inp[5]) ? 4'b0101 : node15183;
														assign node15183 = (inp[15]) ? 4'b0111 : node15184;
															assign node15184 = (inp[3]) ? 4'b0111 : 4'b0101;
											assign node15189 = (inp[14]) ? node15201 : node15190;
												assign node15190 = (inp[2]) ? node15198 : node15191;
													assign node15191 = (inp[5]) ? node15193 : 4'b0111;
														assign node15193 = (inp[3]) ? node15195 : 4'b0101;
															assign node15195 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node15198 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node15201 = (inp[3]) ? node15207 : node15202;
													assign node15202 = (inp[15]) ? node15204 : 4'b0110;
														assign node15204 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node15207 = (inp[2]) ? 4'b0100 : node15208;
														assign node15208 = (inp[0]) ? 4'b0100 : node15209;
															assign node15209 = (inp[5]) ? 4'b0110 : 4'b0100;
									assign node15214 = (inp[15]) ? node15248 : node15215;
										assign node15215 = (inp[0]) ? node15233 : node15216;
											assign node15216 = (inp[5]) ? node15224 : node15217;
												assign node15217 = (inp[3]) ? node15219 : 4'b0110;
													assign node15219 = (inp[7]) ? node15221 : 4'b0101;
														assign node15221 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node15224 = (inp[7]) ? node15230 : node15225;
													assign node15225 = (inp[8]) ? node15227 : 4'b0100;
														assign node15227 = (inp[3]) ? 4'b0100 : 4'b0101;
													assign node15230 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node15233 = (inp[3]) ? node15241 : node15234;
												assign node15234 = (inp[5]) ? 4'b0110 : node15235;
													assign node15235 = (inp[7]) ? node15237 : 4'b0100;
														assign node15237 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node15241 = (inp[2]) ? node15243 : 4'b0110;
													assign node15243 = (inp[7]) ? node15245 : 4'b0110;
														assign node15245 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node15248 = (inp[0]) ? node15274 : node15249;
											assign node15249 = (inp[5]) ? node15265 : node15250;
												assign node15250 = (inp[3]) ? node15262 : node15251;
													assign node15251 = (inp[7]) ? node15257 : node15252;
														assign node15252 = (inp[2]) ? 4'b0101 : node15253;
															assign node15253 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node15257 = (inp[2]) ? 4'b0100 : node15258;
															assign node15258 = (inp[8]) ? 4'b0100 : 4'b0100;
													assign node15262 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node15265 = (inp[8]) ? node15269 : node15266;
													assign node15266 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node15269 = (inp[2]) ? node15271 : 4'b0110;
														assign node15271 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node15274 = (inp[5]) ? node15280 : node15275;
												assign node15275 = (inp[3]) ? 4'b0101 : node15276;
													assign node15276 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node15280 = (inp[8]) ? node15282 : 4'b0101;
													assign node15282 = (inp[7]) ? node15284 : 4'b0101;
														assign node15284 = (inp[14]) ? 4'b0100 : 4'b0101;
					assign node15287 = (inp[12]) ? node15945 : node15288;
						assign node15288 = (inp[3]) ? node15640 : node15289;
							assign node15289 = (inp[15]) ? node15485 : node15290;
								assign node15290 = (inp[7]) ? node15400 : node15291;
									assign node15291 = (inp[8]) ? node15349 : node15292;
										assign node15292 = (inp[14]) ? node15324 : node15293;
											assign node15293 = (inp[2]) ? node15311 : node15294;
												assign node15294 = (inp[0]) ? node15302 : node15295;
													assign node15295 = (inp[5]) ? node15297 : 4'b1111;
														assign node15297 = (inp[6]) ? node15299 : 4'b1101;
															assign node15299 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node15302 = (inp[5]) ? node15304 : 4'b0101;
														assign node15304 = (inp[1]) ? node15308 : node15305;
															assign node15305 = (inp[6]) ? 4'b1111 : 4'b0111;
															assign node15308 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node15311 = (inp[11]) ? node15319 : node15312;
													assign node15312 = (inp[0]) ? node15316 : node15313;
														assign node15313 = (inp[1]) ? 4'b1110 : 4'b0110;
														assign node15316 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node15319 = (inp[1]) ? node15321 : 4'b0110;
														assign node15321 = (inp[5]) ? 4'b1100 : 4'b0110;
											assign node15324 = (inp[1]) ? node15338 : node15325;
												assign node15325 = (inp[2]) ? 4'b0110 : node15326;
													assign node15326 = (inp[5]) ? node15332 : node15327;
														assign node15327 = (inp[0]) ? 4'b0100 : node15328;
															assign node15328 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node15332 = (inp[6]) ? 4'b1110 : node15333;
															assign node15333 = (inp[11]) ? 4'b0110 : 4'b1110;
												assign node15338 = (inp[5]) ? node15346 : node15339;
													assign node15339 = (inp[0]) ? node15341 : 4'b1110;
														assign node15341 = (inp[11]) ? 4'b0100 : node15342;
															assign node15342 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node15346 = (inp[2]) ? 4'b0110 : 4'b0100;
										assign node15349 = (inp[2]) ? node15377 : node15350;
											assign node15350 = (inp[14]) ? node15366 : node15351;
												assign node15351 = (inp[6]) ? node15357 : node15352;
													assign node15352 = (inp[5]) ? 4'b0100 : node15353;
														assign node15353 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node15357 = (inp[0]) ? node15363 : node15358;
														assign node15358 = (inp[5]) ? 4'b1100 : node15359;
															assign node15359 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node15363 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node15366 = (inp[11]) ? node15372 : node15367;
													assign node15367 = (inp[5]) ? node15369 : 4'b1111;
														assign node15369 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node15372 = (inp[5]) ? 4'b0101 : node15373;
														assign node15373 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node15377 = (inp[14]) ? node15393 : node15378;
												assign node15378 = (inp[0]) ? node15390 : node15379;
													assign node15379 = (inp[5]) ? node15385 : node15380;
														assign node15380 = (inp[1]) ? node15382 : 4'b0111;
															assign node15382 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node15385 = (inp[6]) ? node15387 : 4'b1101;
															assign node15387 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node15390 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node15393 = (inp[6]) ? 4'b1111 : node15394;
													assign node15394 = (inp[0]) ? node15396 : 4'b1111;
														assign node15396 = (inp[5]) ? 4'b0111 : 4'b0101;
									assign node15400 = (inp[8]) ? node15440 : node15401;
										assign node15401 = (inp[2]) ? node15421 : node15402;
											assign node15402 = (inp[14]) ? node15418 : node15403;
												assign node15403 = (inp[6]) ? node15409 : node15404;
													assign node15404 = (inp[11]) ? node15406 : 4'b0110;
														assign node15406 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node15409 = (inp[0]) ? node15413 : node15410;
														assign node15410 = (inp[1]) ? 4'b0110 : 4'b1110;
														assign node15413 = (inp[5]) ? node15415 : 4'b1100;
															assign node15415 = (inp[11]) ? 4'b1110 : 4'b0110;
												assign node15418 = (inp[6]) ? 4'b0101 : 4'b1111;
											assign node15421 = (inp[0]) ? node15429 : node15422;
												assign node15422 = (inp[5]) ? node15424 : 4'b1111;
													assign node15424 = (inp[6]) ? 4'b1101 : node15425;
														assign node15425 = (inp[11]) ? 4'b1101 : 4'b0101;
												assign node15429 = (inp[5]) ? node15433 : node15430;
													assign node15430 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node15433 = (inp[14]) ? node15435 : 4'b0111;
														assign node15435 = (inp[11]) ? node15437 : 4'b1111;
															assign node15437 = (inp[6]) ? 4'b0111 : 4'b1111;
										assign node15440 = (inp[2]) ? node15466 : node15441;
											assign node15441 = (inp[14]) ? node15453 : node15442;
												assign node15442 = (inp[5]) ? node15448 : node15443;
													assign node15443 = (inp[1]) ? 4'b1101 : node15444;
														assign node15444 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node15448 = (inp[0]) ? node15450 : 4'b0101;
														assign node15450 = (inp[1]) ? 4'b1111 : 4'b0111;
												assign node15453 = (inp[1]) ? node15461 : node15454;
													assign node15454 = (inp[5]) ? node15458 : node15455;
														assign node15455 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node15458 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node15461 = (inp[6]) ? node15463 : 4'b1110;
														assign node15463 = (inp[5]) ? 4'b1110 : 4'b1100;
											assign node15466 = (inp[0]) ? node15474 : node15467;
												assign node15467 = (inp[5]) ? node15469 : 4'b0110;
													assign node15469 = (inp[14]) ? 4'b0100 : node15470;
														assign node15470 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node15474 = (inp[5]) ? node15476 : 4'b0100;
													assign node15476 = (inp[1]) ? 4'b1110 : node15477;
														assign node15477 = (inp[6]) ? node15481 : node15478;
															assign node15478 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node15481 = (inp[11]) ? 4'b0110 : 4'b1110;
								assign node15485 = (inp[11]) ? node15553 : node15486;
									assign node15486 = (inp[6]) ? node15522 : node15487;
										assign node15487 = (inp[1]) ? node15509 : node15488;
											assign node15488 = (inp[8]) ? node15502 : node15489;
												assign node15489 = (inp[7]) ? node15497 : node15490;
													assign node15490 = (inp[0]) ? 4'b1110 : node15491;
														assign node15491 = (inp[14]) ? node15493 : 4'b1101;
															assign node15493 = (inp[2]) ? 4'b1100 : 4'b1110;
													assign node15497 = (inp[2]) ? 4'b0111 : node15498;
														assign node15498 = (inp[14]) ? 4'b0111 : 4'b1110;
												assign node15502 = (inp[0]) ? node15506 : node15503;
													assign node15503 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node15506 = (inp[5]) ? 4'b0101 : 4'b0111;
											assign node15509 = (inp[0]) ? node15519 : node15510;
												assign node15510 = (inp[5]) ? node15512 : 4'b0101;
													assign node15512 = (inp[14]) ? node15514 : 4'b0111;
														assign node15514 = (inp[8]) ? 4'b0111 : node15515;
															assign node15515 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node15519 = (inp[5]) ? 4'b0100 : 4'b0110;
										assign node15522 = (inp[7]) ? node15544 : node15523;
											assign node15523 = (inp[8]) ? node15539 : node15524;
												assign node15524 = (inp[1]) ? node15530 : node15525;
													assign node15525 = (inp[0]) ? node15527 : 4'b0110;
														assign node15527 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node15530 = (inp[5]) ? node15534 : node15531;
														assign node15531 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node15534 = (inp[2]) ? 4'b1100 : node15535;
															assign node15535 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node15539 = (inp[0]) ? node15541 : 4'b1101;
													assign node15541 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node15544 = (inp[8]) ? node15550 : node15545;
												assign node15545 = (inp[0]) ? 4'b1101 : node15546;
													assign node15546 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node15550 = (inp[5]) ? 4'b1100 : 4'b1110;
									assign node15553 = (inp[6]) ? node15599 : node15554;
										assign node15554 = (inp[1]) ? node15574 : node15555;
											assign node15555 = (inp[14]) ? node15561 : node15556;
												assign node15556 = (inp[2]) ? 4'b0100 : node15557;
													assign node15557 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node15561 = (inp[7]) ? node15567 : node15562;
													assign node15562 = (inp[2]) ? 4'b1101 : node15563;
														assign node15563 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node15567 = (inp[8]) ? node15569 : 4'b1101;
														assign node15569 = (inp[0]) ? 4'b1100 : node15570;
															assign node15570 = (inp[5]) ? 4'b1110 : 4'b1100;
											assign node15574 = (inp[5]) ? node15582 : node15575;
												assign node15575 = (inp[0]) ? 4'b1111 : node15576;
													assign node15576 = (inp[8]) ? node15578 : 4'b1101;
														assign node15578 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node15582 = (inp[0]) ? node15592 : node15583;
													assign node15583 = (inp[14]) ? node15587 : node15584;
														assign node15584 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node15587 = (inp[2]) ? node15589 : 4'b1111;
															assign node15589 = (inp[8]) ? 4'b1110 : 4'b1110;
													assign node15592 = (inp[7]) ? node15594 : 4'b1100;
														assign node15594 = (inp[2]) ? node15596 : 4'b1100;
															assign node15596 = (inp[8]) ? 4'b1100 : 4'b1101;
										assign node15599 = (inp[1]) ? node15619 : node15600;
											assign node15600 = (inp[8]) ? node15612 : node15601;
												assign node15601 = (inp[7]) ? 4'b0111 : node15602;
													assign node15602 = (inp[5]) ? node15604 : 4'b1100;
														assign node15604 = (inp[0]) ? node15608 : node15605;
															assign node15605 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node15608 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node15612 = (inp[2]) ? 4'b0111 : node15613;
													assign node15613 = (inp[5]) ? 4'b1100 : node15614;
														assign node15614 = (inp[0]) ? 4'b0111 : 4'b0100;
											assign node15619 = (inp[8]) ? node15629 : node15620;
												assign node15620 = (inp[7]) ? node15622 : 4'b0100;
													assign node15622 = (inp[14]) ? node15624 : 4'b0111;
														assign node15624 = (inp[2]) ? 4'b0101 : node15625;
															assign node15625 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node15629 = (inp[5]) ? node15633 : node15630;
													assign node15630 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node15633 = (inp[14]) ? 4'b0111 : node15634;
														assign node15634 = (inp[7]) ? 4'b0111 : node15635;
															assign node15635 = (inp[2]) ? 4'b0111 : 4'b0110;
							assign node15640 = (inp[2]) ? node15806 : node15641;
								assign node15641 = (inp[15]) ? node15725 : node15642;
									assign node15642 = (inp[0]) ? node15698 : node15643;
										assign node15643 = (inp[6]) ? node15667 : node15644;
											assign node15644 = (inp[5]) ? node15660 : node15645;
												assign node15645 = (inp[11]) ? node15653 : node15646;
													assign node15646 = (inp[14]) ? node15648 : 4'b1100;
														assign node15648 = (inp[8]) ? 4'b0101 : node15649;
															assign node15649 = (inp[1]) ? 4'b0100 : 4'b1100;
													assign node15653 = (inp[1]) ? node15655 : 4'b1101;
														assign node15655 = (inp[14]) ? 4'b1101 : node15656;
															assign node15656 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node15660 = (inp[8]) ? 4'b1100 : node15661;
													assign node15661 = (inp[14]) ? node15663 : 4'b1100;
														assign node15663 = (inp[11]) ? 4'b0100 : 4'b1100;
											assign node15667 = (inp[11]) ? node15685 : node15668;
												assign node15668 = (inp[1]) ? node15676 : node15669;
													assign node15669 = (inp[14]) ? node15673 : node15670;
														assign node15670 = (inp[7]) ? 4'b1101 : 4'b0101;
														assign node15673 = (inp[8]) ? 4'b1100 : 4'b0100;
													assign node15676 = (inp[14]) ? node15682 : node15677;
														assign node15677 = (inp[5]) ? 4'b1100 : node15678;
															assign node15678 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node15682 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node15685 = (inp[7]) ? node15693 : node15686;
													assign node15686 = (inp[8]) ? node15690 : node15687;
														assign node15687 = (inp[1]) ? 4'b0101 : 4'b1101;
														assign node15690 = (inp[5]) ? 4'b0100 : 4'b1100;
													assign node15693 = (inp[5]) ? 4'b0101 : node15694;
														assign node15694 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node15698 = (inp[8]) ? node15712 : node15699;
											assign node15699 = (inp[5]) ? node15705 : node15700;
												assign node15700 = (inp[7]) ? node15702 : 4'b1110;
													assign node15702 = (inp[14]) ? 4'b0111 : 4'b1110;
												assign node15705 = (inp[6]) ? node15707 : 4'b0111;
													assign node15707 = (inp[7]) ? node15709 : 4'b1110;
														assign node15709 = (inp[1]) ? 4'b1110 : 4'b0110;
											assign node15712 = (inp[5]) ? node15720 : node15713;
												assign node15713 = (inp[1]) ? node15715 : 4'b1111;
													assign node15715 = (inp[14]) ? node15717 : 4'b0111;
														assign node15717 = (inp[7]) ? 4'b1110 : 4'b0111;
												assign node15720 = (inp[1]) ? 4'b1110 : node15721;
													assign node15721 = (inp[11]) ? 4'b1110 : 4'b1111;
									assign node15725 = (inp[0]) ? node15747 : node15726;
										assign node15726 = (inp[1]) ? node15730 : node15727;
											assign node15727 = (inp[7]) ? 4'b0110 : 4'b1110;
											assign node15730 = (inp[5]) ? node15738 : node15731;
												assign node15731 = (inp[8]) ? node15733 : 4'b1111;
													assign node15733 = (inp[6]) ? 4'b0111 : node15734;
														assign node15734 = (inp[11]) ? 4'b1110 : 4'b0111;
												assign node15738 = (inp[7]) ? node15740 : 4'b0110;
													assign node15740 = (inp[8]) ? node15744 : node15741;
														assign node15741 = (inp[6]) ? 4'b1110 : 4'b0110;
														assign node15744 = (inp[11]) ? 4'b1111 : 4'b0111;
										assign node15747 = (inp[1]) ? node15781 : node15748;
											assign node15748 = (inp[5]) ? node15760 : node15749;
												assign node15749 = (inp[11]) ? node15757 : node15750;
													assign node15750 = (inp[8]) ? node15752 : 4'b1100;
														assign node15752 = (inp[6]) ? 4'b1100 : node15753;
															assign node15753 = (inp[7]) ? 4'b0101 : 4'b1100;
													assign node15757 = (inp[6]) ? 4'b0101 : 4'b0100;
												assign node15760 = (inp[11]) ? node15770 : node15761;
													assign node15761 = (inp[8]) ? 4'b0101 : node15762;
														assign node15762 = (inp[6]) ? node15766 : node15763;
															assign node15763 = (inp[7]) ? 4'b0101 : 4'b1100;
															assign node15766 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node15770 = (inp[7]) ? node15776 : node15771;
														assign node15771 = (inp[8]) ? 4'b1101 : node15772;
															assign node15772 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node15776 = (inp[6]) ? 4'b1100 : node15777;
															assign node15777 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node15781 = (inp[6]) ? node15793 : node15782;
												assign node15782 = (inp[11]) ? node15790 : node15783;
													assign node15783 = (inp[5]) ? 4'b0101 : node15784;
														assign node15784 = (inp[7]) ? node15786 : 4'b0100;
															assign node15786 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node15790 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node15793 = (inp[11]) ? node15801 : node15794;
													assign node15794 = (inp[14]) ? 4'b1101 : node15795;
														assign node15795 = (inp[7]) ? 4'b1100 : node15796;
															assign node15796 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node15801 = (inp[7]) ? node15803 : 4'b0100;
														assign node15803 = (inp[8]) ? 4'b0101 : 4'b0100;
								assign node15806 = (inp[7]) ? node15884 : node15807;
									assign node15807 = (inp[8]) ? node15855 : node15808;
										assign node15808 = (inp[6]) ? node15834 : node15809;
											assign node15809 = (inp[11]) ? node15827 : node15810;
												assign node15810 = (inp[1]) ? node15820 : node15811;
													assign node15811 = (inp[14]) ? 4'b1110 : node15812;
														assign node15812 = (inp[15]) ? node15816 : node15813;
															assign node15813 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node15816 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node15820 = (inp[15]) ? node15824 : node15821;
														assign node15821 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node15824 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node15827 = (inp[1]) ? node15829 : 4'b0100;
													assign node15829 = (inp[15]) ? node15831 : 4'b1100;
														assign node15831 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node15834 = (inp[0]) ? node15844 : node15835;
												assign node15835 = (inp[15]) ? node15841 : node15836;
													assign node15836 = (inp[1]) ? node15838 : 4'b1100;
														assign node15838 = (inp[5]) ? 4'b0100 : 4'b1100;
													assign node15841 = (inp[5]) ? 4'b0110 : 4'b1110;
												assign node15844 = (inp[15]) ? 4'b1100 : node15845;
													assign node15845 = (inp[5]) ? node15847 : 4'b0110;
														assign node15847 = (inp[1]) ? node15851 : node15848;
															assign node15848 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node15851 = (inp[14]) ? 4'b1110 : 4'b0110;
										assign node15855 = (inp[6]) ? node15871 : node15856;
											assign node15856 = (inp[11]) ? node15864 : node15857;
												assign node15857 = (inp[0]) ? node15861 : node15858;
													assign node15858 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node15861 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node15864 = (inp[14]) ? node15868 : node15865;
													assign node15865 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node15868 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node15871 = (inp[11]) ? node15879 : node15872;
												assign node15872 = (inp[0]) ? node15876 : node15873;
													assign node15873 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node15876 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node15879 = (inp[15]) ? node15881 : 4'b0101;
													assign node15881 = (inp[0]) ? 4'b0101 : 4'b0111;
									assign node15884 = (inp[8]) ? node15920 : node15885;
										assign node15885 = (inp[11]) ? node15903 : node15886;
											assign node15886 = (inp[6]) ? node15898 : node15887;
												assign node15887 = (inp[5]) ? node15895 : node15888;
													assign node15888 = (inp[1]) ? node15890 : 4'b0111;
														assign node15890 = (inp[15]) ? node15892 : 4'b0101;
															assign node15892 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node15895 = (inp[1]) ? 4'b0111 : 4'b0101;
												assign node15898 = (inp[5]) ? node15900 : 4'b1101;
													assign node15900 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node15903 = (inp[6]) ? node15905 : 4'b1111;
												assign node15905 = (inp[1]) ? node15911 : node15906;
													assign node15906 = (inp[15]) ? node15908 : 4'b0101;
														assign node15908 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node15911 = (inp[5]) ? node15915 : node15912;
														assign node15912 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node15915 = (inp[15]) ? node15917 : 4'b0111;
															assign node15917 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node15920 = (inp[6]) ? node15932 : node15921;
											assign node15921 = (inp[11]) ? node15927 : node15922;
												assign node15922 = (inp[0]) ? 4'b0110 : node15923;
													assign node15923 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node15927 = (inp[0]) ? 4'b1110 : node15928;
													assign node15928 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node15932 = (inp[11]) ? node15940 : node15933;
												assign node15933 = (inp[0]) ? node15937 : node15934;
													assign node15934 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node15937 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node15940 = (inp[14]) ? node15942 : 4'b0100;
													assign node15942 = (inp[1]) ? 4'b0100 : 4'b0110;
						assign node15945 = (inp[6]) ? node16325 : node15946;
							assign node15946 = (inp[11]) ? node16142 : node15947;
								assign node15947 = (inp[1]) ? node16031 : node15948;
									assign node15948 = (inp[8]) ? node15986 : node15949;
										assign node15949 = (inp[7]) ? node15973 : node15950;
											assign node15950 = (inp[14]) ? node15964 : node15951;
												assign node15951 = (inp[2]) ? node15957 : node15952;
													assign node15952 = (inp[15]) ? node15954 : 4'b1101;
														assign node15954 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node15957 = (inp[5]) ? node15959 : 4'b1100;
														assign node15959 = (inp[0]) ? 4'b1110 : node15960;
															assign node15960 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node15964 = (inp[2]) ? 4'b1100 : node15965;
													assign node15965 = (inp[15]) ? node15969 : node15966;
														assign node15966 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node15969 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node15973 = (inp[2]) ? node15981 : node15974;
												assign node15974 = (inp[14]) ? node15976 : 4'b1110;
													assign node15976 = (inp[15]) ? node15978 : 4'b0111;
														assign node15978 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node15981 = (inp[15]) ? 4'b0101 : node15982;
													assign node15982 = (inp[5]) ? 4'b0111 : 4'b0101;
										assign node15986 = (inp[7]) ? node16010 : node15987;
											assign node15987 = (inp[2]) ? node15999 : node15988;
												assign node15988 = (inp[14]) ? node15996 : node15989;
													assign node15989 = (inp[0]) ? node15991 : 4'b1110;
														assign node15991 = (inp[3]) ? 4'b1110 : node15992;
															assign node15992 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node15996 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node15999 = (inp[3]) ? node16005 : node16000;
													assign node16000 = (inp[0]) ? 4'b0111 : node16001;
														assign node16001 = (inp[14]) ? 4'b0111 : 4'b0101;
													assign node16005 = (inp[15]) ? node16007 : 4'b0101;
														assign node16007 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node16010 = (inp[14]) ? node16020 : node16011;
												assign node16011 = (inp[2]) ? node16013 : 4'b0101;
													assign node16013 = (inp[5]) ? node16015 : 4'b0100;
														assign node16015 = (inp[0]) ? node16017 : 4'b0100;
															assign node16017 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node16020 = (inp[5]) ? node16024 : node16021;
													assign node16021 = (inp[2]) ? 4'b0100 : 4'b0110;
													assign node16024 = (inp[2]) ? 4'b0110 : node16025;
														assign node16025 = (inp[15]) ? node16027 : 4'b0100;
															assign node16027 = (inp[0]) ? 4'b0100 : 4'b0110;
									assign node16031 = (inp[14]) ? node16091 : node16032;
										assign node16032 = (inp[7]) ? node16072 : node16033;
											assign node16033 = (inp[3]) ? node16053 : node16034;
												assign node16034 = (inp[2]) ? node16046 : node16035;
													assign node16035 = (inp[8]) ? node16039 : node16036;
														assign node16036 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node16039 = (inp[15]) ? node16043 : node16040;
															assign node16040 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node16043 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node16046 = (inp[8]) ? 4'b0111 : node16047;
														assign node16047 = (inp[5]) ? 4'b0110 : node16048;
															assign node16048 = (inp[0]) ? 4'b0100 : 4'b0100;
												assign node16053 = (inp[2]) ? node16063 : node16054;
													assign node16054 = (inp[8]) ? node16060 : node16055;
														assign node16055 = (inp[15]) ? node16057 : 4'b0111;
															assign node16057 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node16060 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node16063 = (inp[8]) ? node16069 : node16064;
														assign node16064 = (inp[15]) ? node16066 : 4'b0100;
															assign node16066 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node16069 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node16072 = (inp[15]) ? node16084 : node16073;
												assign node16073 = (inp[0]) ? node16081 : node16074;
													assign node16074 = (inp[2]) ? node16078 : node16075;
														assign node16075 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node16078 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node16081 = (inp[3]) ? 4'b0111 : 4'b0100;
												assign node16084 = (inp[3]) ? 4'b0110 : node16085;
													assign node16085 = (inp[0]) ? 4'b0100 : node16086;
														assign node16086 = (inp[2]) ? 4'b0110 : 4'b0100;
										assign node16091 = (inp[2]) ? node16119 : node16092;
											assign node16092 = (inp[15]) ? node16108 : node16093;
												assign node16093 = (inp[0]) ? node16101 : node16094;
													assign node16094 = (inp[5]) ? node16096 : 4'b0110;
														assign node16096 = (inp[8]) ? node16098 : 4'b0100;
															assign node16098 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node16101 = (inp[5]) ? node16103 : 4'b0101;
														assign node16103 = (inp[3]) ? node16105 : 4'b0110;
															assign node16105 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node16108 = (inp[0]) ? node16114 : node16109;
													assign node16109 = (inp[5]) ? 4'b0111 : node16110;
														assign node16110 = (inp[8]) ? 4'b0101 : 4'b0111;
													assign node16114 = (inp[8]) ? node16116 : 4'b0100;
														assign node16116 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node16119 = (inp[3]) ? node16131 : node16120;
												assign node16120 = (inp[8]) ? node16128 : node16121;
													assign node16121 = (inp[7]) ? node16123 : 4'b0100;
														assign node16123 = (inp[5]) ? node16125 : 4'b0101;
															assign node16125 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node16128 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node16131 = (inp[15]) ? node16135 : node16132;
													assign node16132 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node16135 = (inp[0]) ? node16137 : 4'b0111;
														assign node16137 = (inp[8]) ? node16139 : 4'b0101;
															assign node16139 = (inp[7]) ? 4'b0100 : 4'b0101;
								assign node16142 = (inp[1]) ? node16232 : node16143;
									assign node16143 = (inp[8]) ? node16193 : node16144;
										assign node16144 = (inp[7]) ? node16170 : node16145;
											assign node16145 = (inp[14]) ? node16155 : node16146;
												assign node16146 = (inp[2]) ? 4'b0100 : node16147;
													assign node16147 = (inp[3]) ? 4'b0101 : node16148;
														assign node16148 = (inp[5]) ? 4'b0111 : node16149;
															assign node16149 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node16155 = (inp[0]) ? node16165 : node16156;
													assign node16156 = (inp[5]) ? 4'b0100 : node16157;
														assign node16157 = (inp[2]) ? node16161 : node16158;
															assign node16158 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node16161 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node16165 = (inp[15]) ? node16167 : 4'b0110;
														assign node16167 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node16170 = (inp[2]) ? node16186 : node16171;
												assign node16171 = (inp[14]) ? node16183 : node16172;
													assign node16172 = (inp[3]) ? node16178 : node16173;
														assign node16173 = (inp[0]) ? 4'b0100 : node16174;
															assign node16174 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node16178 = (inp[0]) ? 4'b0110 : node16179;
															assign node16179 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node16183 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node16186 = (inp[15]) ? 4'b1011 : node16187;
													assign node16187 = (inp[0]) ? 4'b1001 : node16188;
														assign node16188 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node16193 = (inp[7]) ? node16211 : node16194;
											assign node16194 = (inp[14]) ? node16206 : node16195;
												assign node16195 = (inp[2]) ? node16203 : node16196;
													assign node16196 = (inp[3]) ? node16198 : 4'b0100;
														assign node16198 = (inp[5]) ? 4'b0110 : node16199;
															assign node16199 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node16203 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node16206 = (inp[2]) ? 4'b1001 : node16207;
													assign node16207 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node16211 = (inp[2]) ? node16223 : node16212;
												assign node16212 = (inp[14]) ? node16216 : node16213;
													assign node16213 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node16216 = (inp[3]) ? 4'b1010 : node16217;
														assign node16217 = (inp[5]) ? node16219 : 4'b1000;
															assign node16219 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node16223 = (inp[5]) ? node16229 : node16224;
													assign node16224 = (inp[3]) ? 4'b1010 : node16225;
														assign node16225 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node16229 = (inp[3]) ? 4'b1000 : 4'b1010;
									assign node16232 = (inp[8]) ? node16278 : node16233;
										assign node16233 = (inp[7]) ? node16255 : node16234;
											assign node16234 = (inp[5]) ? node16246 : node16235;
												assign node16235 = (inp[2]) ? node16239 : node16236;
													assign node16236 = (inp[15]) ? 4'b1000 : 4'b1001;
													assign node16239 = (inp[15]) ? 4'b1000 : node16240;
														assign node16240 = (inp[0]) ? 4'b1010 : node16241;
															assign node16241 = (inp[14]) ? 4'b1000 : 4'b1010;
												assign node16246 = (inp[3]) ? 4'b1010 : node16247;
													assign node16247 = (inp[0]) ? node16251 : node16248;
														assign node16248 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node16251 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node16255 = (inp[2]) ? node16275 : node16256;
												assign node16256 = (inp[14]) ? node16270 : node16257;
													assign node16257 = (inp[5]) ? node16263 : node16258;
														assign node16258 = (inp[15]) ? node16260 : 4'b1000;
															assign node16260 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node16263 = (inp[15]) ? node16267 : node16264;
															assign node16264 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node16267 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node16270 = (inp[5]) ? node16272 : 4'b1001;
														assign node16272 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node16275 = (inp[0]) ? 4'b1011 : 4'b1001;
										assign node16278 = (inp[7]) ? node16304 : node16279;
											assign node16279 = (inp[14]) ? node16289 : node16280;
												assign node16280 = (inp[2]) ? node16282 : 4'b1010;
													assign node16282 = (inp[0]) ? node16284 : 4'b1011;
														assign node16284 = (inp[3]) ? 4'b1001 : node16285;
															assign node16285 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node16289 = (inp[2]) ? node16295 : node16290;
													assign node16290 = (inp[15]) ? 4'b1001 : node16291;
														assign node16291 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node16295 = (inp[5]) ? node16301 : node16296;
														assign node16296 = (inp[0]) ? node16298 : 4'b1001;
															assign node16298 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node16301 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node16304 = (inp[2]) ? node16316 : node16305;
												assign node16305 = (inp[14]) ? node16313 : node16306;
													assign node16306 = (inp[5]) ? 4'b1001 : node16307;
														assign node16307 = (inp[0]) ? node16309 : 4'b1011;
															assign node16309 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node16313 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node16316 = (inp[15]) ? 4'b1000 : node16317;
													assign node16317 = (inp[5]) ? 4'b1010 : node16318;
														assign node16318 = (inp[14]) ? 4'b1010 : node16319;
															assign node16319 = (inp[3]) ? 4'b1000 : 4'b1000;
							assign node16325 = (inp[11]) ? node16513 : node16326;
								assign node16326 = (inp[1]) ? node16420 : node16327;
									assign node16327 = (inp[8]) ? node16359 : node16328;
										assign node16328 = (inp[7]) ? node16344 : node16329;
											assign node16329 = (inp[2]) ? node16339 : node16330;
												assign node16330 = (inp[3]) ? node16336 : node16331;
													assign node16331 = (inp[0]) ? 4'b0101 : node16332;
														assign node16332 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node16336 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node16339 = (inp[15]) ? node16341 : 4'b0110;
													assign node16341 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node16344 = (inp[14]) ? node16350 : node16345;
												assign node16345 = (inp[2]) ? 4'b1001 : node16346;
													assign node16346 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node16350 = (inp[5]) ? 4'b1011 : node16351;
													assign node16351 = (inp[3]) ? 4'b1001 : node16352;
														assign node16352 = (inp[0]) ? node16354 : 4'b1011;
															assign node16354 = (inp[15]) ? 4'b1011 : 4'b1001;
										assign node16359 = (inp[7]) ? node16389 : node16360;
											assign node16360 = (inp[14]) ? node16378 : node16361;
												assign node16361 = (inp[2]) ? node16371 : node16362;
													assign node16362 = (inp[3]) ? 4'b0100 : node16363;
														assign node16363 = (inp[0]) ? node16367 : node16364;
															assign node16364 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node16367 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node16371 = (inp[15]) ? node16373 : 4'b1001;
														assign node16373 = (inp[5]) ? 4'b1001 : node16374;
															assign node16374 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node16378 = (inp[3]) ? node16384 : node16379;
													assign node16379 = (inp[5]) ? 4'b1001 : node16380;
														assign node16380 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node16384 = (inp[2]) ? 4'b1011 : node16385;
														assign node16385 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node16389 = (inp[14]) ? node16405 : node16390;
												assign node16390 = (inp[2]) ? node16400 : node16391;
													assign node16391 = (inp[15]) ? node16397 : node16392;
														assign node16392 = (inp[5]) ? 4'b1011 : node16393;
															assign node16393 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node16397 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node16400 = (inp[3]) ? 4'b1010 : node16401;
														assign node16401 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node16405 = (inp[3]) ? node16413 : node16406;
													assign node16406 = (inp[0]) ? node16408 : 4'b1000;
														assign node16408 = (inp[2]) ? node16410 : 4'b1010;
															assign node16410 = (inp[5]) ? 4'b1000 : 4'b1000;
													assign node16413 = (inp[0]) ? node16417 : node16414;
														assign node16414 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node16417 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node16420 = (inp[5]) ? node16476 : node16421;
										assign node16421 = (inp[2]) ? node16443 : node16422;
											assign node16422 = (inp[3]) ? node16432 : node16423;
												assign node16423 = (inp[0]) ? 4'b1001 : node16424;
													assign node16424 = (inp[14]) ? node16426 : 4'b1010;
														assign node16426 = (inp[8]) ? 4'b1001 : node16427;
															assign node16427 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node16432 = (inp[14]) ? node16436 : node16433;
													assign node16433 = (inp[15]) ? 4'b1001 : 4'b1000;
													assign node16436 = (inp[7]) ? node16440 : node16437;
														assign node16437 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node16440 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node16443 = (inp[14]) ? node16457 : node16444;
												assign node16444 = (inp[7]) ? node16452 : node16445;
													assign node16445 = (inp[8]) ? 4'b1001 : node16446;
														assign node16446 = (inp[3]) ? 4'b1010 : node16447;
															assign node16447 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node16452 = (inp[8]) ? 4'b1010 : node16453;
														assign node16453 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node16457 = (inp[3]) ? node16467 : node16458;
													assign node16458 = (inp[7]) ? node16462 : node16459;
														assign node16459 = (inp[15]) ? 4'b1010 : 4'b1011;
														assign node16462 = (inp[8]) ? node16464 : 4'b1001;
															assign node16464 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node16467 = (inp[7]) ? node16471 : node16468;
														assign node16468 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node16471 = (inp[15]) ? node16473 : 4'b1000;
															assign node16473 = (inp[0]) ? 4'b1000 : 4'b1010;
										assign node16476 = (inp[2]) ? node16496 : node16477;
											assign node16477 = (inp[3]) ? node16487 : node16478;
												assign node16478 = (inp[8]) ? node16480 : 4'b1010;
													assign node16480 = (inp[7]) ? node16482 : 4'b1010;
														assign node16482 = (inp[15]) ? 4'b1001 : node16483;
															assign node16483 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node16487 = (inp[14]) ? node16489 : 4'b1000;
													assign node16489 = (inp[15]) ? node16491 : 4'b1000;
														assign node16491 = (inp[0]) ? node16493 : 4'b1011;
															assign node16493 = (inp[8]) ? 4'b1001 : 4'b1000;
											assign node16496 = (inp[3]) ? node16506 : node16497;
												assign node16497 = (inp[15]) ? node16503 : node16498;
													assign node16498 = (inp[8]) ? 4'b1000 : node16499;
														assign node16499 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node16503 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node16506 = (inp[0]) ? node16510 : node16507;
													assign node16507 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node16510 = (inp[15]) ? 4'b1001 : 4'b1011;
								assign node16513 = (inp[1]) ? node16593 : node16514;
									assign node16514 = (inp[8]) ? node16548 : node16515;
										assign node16515 = (inp[7]) ? node16531 : node16516;
											assign node16516 = (inp[2]) ? node16526 : node16517;
												assign node16517 = (inp[14]) ? node16521 : node16518;
													assign node16518 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node16521 = (inp[5]) ? 4'b1000 : node16522;
														assign node16522 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node16526 = (inp[14]) ? 4'b1010 : node16527;
													assign node16527 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node16531 = (inp[2]) ? node16539 : node16532;
												assign node16532 = (inp[14]) ? 4'b0001 : node16533;
													assign node16533 = (inp[0]) ? node16535 : 4'b1010;
														assign node16535 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node16539 = (inp[15]) ? 4'b0001 : node16540;
													assign node16540 = (inp[5]) ? 4'b0011 : node16541;
														assign node16541 = (inp[0]) ? node16543 : 4'b0001;
															assign node16543 = (inp[14]) ? 4'b0001 : 4'b0011;
										assign node16548 = (inp[7]) ? node16572 : node16549;
											assign node16549 = (inp[2]) ? node16563 : node16550;
												assign node16550 = (inp[14]) ? node16558 : node16551;
													assign node16551 = (inp[0]) ? node16553 : 4'b1000;
														assign node16553 = (inp[5]) ? 4'b1010 : node16554;
															assign node16554 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node16558 = (inp[0]) ? 4'b0011 : node16559;
														assign node16559 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node16563 = (inp[0]) ? node16565 : 4'b0011;
													assign node16565 = (inp[15]) ? 4'b0001 : node16566;
														assign node16566 = (inp[3]) ? 4'b0011 : node16567;
															assign node16567 = (inp[5]) ? 4'b0011 : 4'b0001;
											assign node16572 = (inp[2]) ? node16584 : node16573;
												assign node16573 = (inp[14]) ? 4'b0000 : node16574;
													assign node16574 = (inp[0]) ? node16578 : node16575;
														assign node16575 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node16578 = (inp[5]) ? 4'b0011 : node16579;
															assign node16579 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node16584 = (inp[14]) ? node16586 : 4'b0000;
													assign node16586 = (inp[3]) ? 4'b0010 : node16587;
														assign node16587 = (inp[0]) ? 4'b0010 : node16588;
															assign node16588 = (inp[15]) ? 4'b0000 : 4'b0000;
									assign node16593 = (inp[0]) ? node16647 : node16594;
										assign node16594 = (inp[15]) ? node16618 : node16595;
											assign node16595 = (inp[3]) ? node16607 : node16596;
												assign node16596 = (inp[5]) ? node16604 : node16597;
													assign node16597 = (inp[14]) ? 4'b0011 : node16598;
														assign node16598 = (inp[8]) ? node16600 : 4'b0010;
															assign node16600 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node16604 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node16607 = (inp[2]) ? node16613 : node16608;
													assign node16608 = (inp[5]) ? node16610 : 4'b0001;
														assign node16610 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node16613 = (inp[5]) ? node16615 : 4'b0000;
														assign node16615 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node16618 = (inp[3]) ? node16632 : node16619;
												assign node16619 = (inp[5]) ? node16625 : node16620;
													assign node16620 = (inp[8]) ? 4'b0001 : node16621;
														assign node16621 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node16625 = (inp[7]) ? node16627 : 4'b0011;
														assign node16627 = (inp[8]) ? node16629 : 4'b0011;
															assign node16629 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node16632 = (inp[7]) ? node16640 : node16633;
													assign node16633 = (inp[8]) ? 4'b0011 : node16634;
														assign node16634 = (inp[5]) ? node16636 : 4'b0010;
															assign node16636 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node16640 = (inp[14]) ? 4'b0011 : node16641;
														assign node16641 = (inp[2]) ? node16643 : 4'b0010;
															assign node16643 = (inp[8]) ? 4'b0010 : 4'b0011;
										assign node16647 = (inp[15]) ? node16671 : node16648;
											assign node16648 = (inp[5]) ? node16658 : node16649;
												assign node16649 = (inp[3]) ? node16653 : node16650;
													assign node16650 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node16653 = (inp[7]) ? node16655 : 4'b0010;
														assign node16655 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node16658 = (inp[8]) ? node16664 : node16659;
													assign node16659 = (inp[14]) ? node16661 : 4'b0010;
														assign node16661 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node16664 = (inp[7]) ? 4'b0010 : node16665;
														assign node16665 = (inp[2]) ? 4'b0011 : node16666;
															assign node16666 = (inp[14]) ? 4'b0011 : 4'b0010;
											assign node16671 = (inp[3]) ? node16675 : node16672;
												assign node16672 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node16675 = (inp[8]) ? node16679 : node16676;
													assign node16676 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node16679 = (inp[7]) ? 4'b0000 : node16680;
														assign node16680 = (inp[2]) ? 4'b0001 : 4'b0000;
			assign node16684 = (inp[15]) ? node19608 : node16685;
				assign node16685 = (inp[0]) ? node18149 : node16686;
					assign node16686 = (inp[5]) ? node17360 : node16687;
						assign node16687 = (inp[3]) ? node17033 : node16688;
							assign node16688 = (inp[9]) ? node16852 : node16689;
								assign node16689 = (inp[4]) ? node16785 : node16690;
									assign node16690 = (inp[12]) ? node16732 : node16691;
										assign node16691 = (inp[11]) ? node16713 : node16692;
											assign node16692 = (inp[6]) ? node16700 : node16693;
												assign node16693 = (inp[1]) ? node16695 : 4'b1111;
													assign node16695 = (inp[8]) ? node16697 : 4'b0110;
														assign node16697 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node16700 = (inp[1]) ? node16710 : node16701;
													assign node16701 = (inp[14]) ? node16707 : node16702;
														assign node16702 = (inp[2]) ? node16704 : 4'b0110;
															assign node16704 = (inp[8]) ? 4'b1011 : 4'b0110;
														assign node16707 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node16710 = (inp[7]) ? 4'b1011 : 4'b1010;
											assign node16713 = (inp[6]) ? node16721 : node16714;
												assign node16714 = (inp[8]) ? node16718 : node16715;
													assign node16715 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node16718 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node16721 = (inp[1]) ? 4'b0011 : node16722;
													assign node16722 = (inp[8]) ? 4'b0010 : node16723;
														assign node16723 = (inp[2]) ? node16727 : node16724;
															assign node16724 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node16727 = (inp[7]) ? 4'b0011 : 4'b1010;
										assign node16732 = (inp[7]) ? node16762 : node16733;
											assign node16733 = (inp[8]) ? node16749 : node16734;
												assign node16734 = (inp[2]) ? node16742 : node16735;
													assign node16735 = (inp[14]) ? node16739 : node16736;
														assign node16736 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node16739 = (inp[1]) ? 4'b0010 : 4'b1010;
													assign node16742 = (inp[1]) ? 4'b0010 : node16743;
														assign node16743 = (inp[11]) ? node16745 : 4'b0010;
															assign node16745 = (inp[6]) ? 4'b1010 : 4'b0010;
												assign node16749 = (inp[14]) ? node16757 : node16750;
													assign node16750 = (inp[2]) ? 4'b0011 : node16751;
														assign node16751 = (inp[6]) ? 4'b0010 : node16752;
															assign node16752 = (inp[1]) ? 4'b0010 : 4'b1010;
													assign node16757 = (inp[11]) ? 4'b0011 : node16758;
														assign node16758 = (inp[6]) ? 4'b1011 : 4'b0011;
											assign node16762 = (inp[8]) ? node16778 : node16763;
												assign node16763 = (inp[2]) ? node16771 : node16764;
													assign node16764 = (inp[14]) ? node16766 : 4'b1010;
														assign node16766 = (inp[11]) ? node16768 : 4'b1011;
															assign node16768 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node16771 = (inp[1]) ? node16773 : 4'b0011;
														assign node16773 = (inp[6]) ? node16775 : 4'b1011;
															assign node16775 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node16778 = (inp[14]) ? node16780 : 4'b1011;
													assign node16780 = (inp[6]) ? 4'b1010 : node16781;
														assign node16781 = (inp[2]) ? 4'b1010 : 4'b0010;
									assign node16785 = (inp[11]) ? node16811 : node16786;
										assign node16786 = (inp[12]) ? node16802 : node16787;
											assign node16787 = (inp[6]) ? 4'b1111 : node16788;
												assign node16788 = (inp[7]) ? node16794 : node16789;
													assign node16789 = (inp[8]) ? 4'b0011 : node16790;
														assign node16790 = (inp[1]) ? 4'b0010 : 4'b1010;
													assign node16794 = (inp[8]) ? node16796 : 4'b0011;
														assign node16796 = (inp[2]) ? 4'b0010 : node16797;
															assign node16797 = (inp[14]) ? 4'b0010 : 4'b0011;
											assign node16802 = (inp[1]) ? node16804 : 4'b1110;
												assign node16804 = (inp[6]) ? 4'b1110 : node16805;
													assign node16805 = (inp[8]) ? node16807 : 4'b0110;
														assign node16807 = (inp[7]) ? 4'b0110 : 4'b0111;
										assign node16811 = (inp[6]) ? node16829 : node16812;
											assign node16812 = (inp[1]) ? node16818 : node16813;
												assign node16813 = (inp[8]) ? node16815 : 4'b0110;
													assign node16815 = (inp[2]) ? 4'b1111 : 4'b0110;
												assign node16818 = (inp[7]) ? 4'b1111 : node16819;
													assign node16819 = (inp[14]) ? 4'b1110 : node16820;
														assign node16820 = (inp[8]) ? node16824 : node16821;
															assign node16821 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node16824 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node16829 = (inp[1]) ? node16843 : node16830;
												assign node16830 = (inp[7]) ? node16838 : node16831;
													assign node16831 = (inp[12]) ? node16833 : 4'b1110;
														assign node16833 = (inp[8]) ? 4'b0111 : node16834;
															assign node16834 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node16838 = (inp[8]) ? node16840 : 4'b0111;
														assign node16840 = (inp[12]) ? 4'b0111 : 4'b0110;
												assign node16843 = (inp[12]) ? node16845 : 4'b0111;
													assign node16845 = (inp[14]) ? node16847 : 4'b0111;
														assign node16847 = (inp[8]) ? node16849 : 4'b0110;
															assign node16849 = (inp[7]) ? 4'b0110 : 4'b0111;
								assign node16852 = (inp[4]) ? node16948 : node16853;
									assign node16853 = (inp[12]) ? node16897 : node16854;
										assign node16854 = (inp[6]) ? node16878 : node16855;
											assign node16855 = (inp[11]) ? node16869 : node16856;
												assign node16856 = (inp[14]) ? node16864 : node16857;
													assign node16857 = (inp[1]) ? node16859 : 4'b1010;
														assign node16859 = (inp[7]) ? node16861 : 4'b0010;
															assign node16861 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node16864 = (inp[1]) ? 4'b0011 : node16865;
														assign node16865 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node16869 = (inp[1]) ? node16871 : 4'b0010;
													assign node16871 = (inp[2]) ? 4'b1111 : node16872;
														assign node16872 = (inp[7]) ? 4'b1110 : node16873;
															assign node16873 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node16878 = (inp[1]) ? node16890 : node16879;
												assign node16879 = (inp[11]) ? node16881 : 4'b0010;
													assign node16881 = (inp[14]) ? node16883 : 4'b1110;
														assign node16883 = (inp[8]) ? node16887 : node16884;
															assign node16884 = (inp[7]) ? 4'b0111 : 4'b1110;
															assign node16887 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node16890 = (inp[11]) ? 4'b0111 : node16891;
													assign node16891 = (inp[2]) ? 4'b1111 : node16892;
														assign node16892 = (inp[14]) ? 4'b1110 : 4'b1111;
										assign node16897 = (inp[8]) ? node16925 : node16898;
											assign node16898 = (inp[6]) ? node16910 : node16899;
												assign node16899 = (inp[14]) ? node16907 : node16900;
													assign node16900 = (inp[1]) ? 4'b1110 : node16901;
														assign node16901 = (inp[2]) ? 4'b0111 : node16902;
															assign node16902 = (inp[11]) ? 4'b0110 : 4'b1110;
													assign node16907 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node16910 = (inp[14]) ? node16920 : node16911;
													assign node16911 = (inp[2]) ? node16917 : node16912;
														assign node16912 = (inp[7]) ? 4'b0110 : node16913;
															assign node16913 = (inp[11]) ? 4'b1111 : 4'b0111;
														assign node16917 = (inp[1]) ? 4'b1111 : 4'b1110;
													assign node16920 = (inp[2]) ? node16922 : 4'b1111;
														assign node16922 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node16925 = (inp[7]) ? node16935 : node16926;
												assign node16926 = (inp[14]) ? 4'b0111 : node16927;
													assign node16927 = (inp[2]) ? node16929 : 4'b0110;
														assign node16929 = (inp[11]) ? node16931 : 4'b0111;
															assign node16931 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node16935 = (inp[2]) ? node16943 : node16936;
													assign node16936 = (inp[14]) ? node16940 : node16937;
														assign node16937 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node16940 = (inp[6]) ? 4'b1110 : 4'b0110;
													assign node16943 = (inp[6]) ? node16945 : 4'b0110;
														assign node16945 = (inp[14]) ? 4'b1110 : 4'b0110;
									assign node16948 = (inp[12]) ? node16986 : node16949;
										assign node16949 = (inp[6]) ? node16965 : node16950;
											assign node16950 = (inp[8]) ? node16960 : node16951;
												assign node16951 = (inp[1]) ? node16955 : node16952;
													assign node16952 = (inp[2]) ? 4'b0111 : 4'b1111;
													assign node16955 = (inp[14]) ? 4'b0111 : node16956;
														assign node16956 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node16960 = (inp[7]) ? node16962 : 4'b1110;
													assign node16962 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node16965 = (inp[11]) ? node16975 : node16966;
												assign node16966 = (inp[1]) ? 4'b1010 : node16967;
													assign node16967 = (inp[7]) ? node16969 : 4'b0110;
														assign node16969 = (inp[14]) ? 4'b1011 : node16970;
															assign node16970 = (inp[2]) ? 4'b1011 : 4'b0010;
												assign node16975 = (inp[7]) ? node16981 : node16976;
													assign node16976 = (inp[8]) ? 4'b0011 : node16977;
														assign node16977 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node16981 = (inp[8]) ? 4'b0010 : node16982;
														assign node16982 = (inp[2]) ? 4'b0011 : 4'b0010;
										assign node16986 = (inp[7]) ? node17012 : node16987;
											assign node16987 = (inp[8]) ? node17003 : node16988;
												assign node16988 = (inp[14]) ? node16998 : node16989;
													assign node16989 = (inp[11]) ? node16993 : node16990;
														assign node16990 = (inp[1]) ? 4'b0010 : 4'b1010;
														assign node16993 = (inp[6]) ? 4'b0011 : node16994;
															assign node16994 = (inp[1]) ? 4'b1011 : 4'b0011;
													assign node16998 = (inp[6]) ? 4'b0010 : node16999;
														assign node16999 = (inp[2]) ? 4'b0010 : 4'b1010;
												assign node17003 = (inp[1]) ? 4'b1011 : node17004;
													assign node17004 = (inp[6]) ? node17008 : node17005;
														assign node17005 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node17008 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node17012 = (inp[1]) ? node17026 : node17013;
												assign node17013 = (inp[11]) ? node17023 : node17014;
													assign node17014 = (inp[6]) ? node17016 : 4'b0010;
														assign node17016 = (inp[2]) ? node17020 : node17017;
															assign node17017 = (inp[14]) ? 4'b1010 : 4'b0010;
															assign node17020 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node17023 = (inp[6]) ? 4'b1010 : 4'b1011;
												assign node17026 = (inp[6]) ? node17030 : node17027;
													assign node17027 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node17030 = (inp[2]) ? 4'b0011 : 4'b0010;
							assign node17033 = (inp[9]) ? node17205 : node17034;
								assign node17034 = (inp[4]) ? node17128 : node17035;
									assign node17035 = (inp[12]) ? node17083 : node17036;
										assign node17036 = (inp[11]) ? node17054 : node17037;
											assign node17037 = (inp[6]) ? node17051 : node17038;
												assign node17038 = (inp[8]) ? node17044 : node17039;
													assign node17039 = (inp[14]) ? 4'b0111 : node17040;
														assign node17040 = (inp[1]) ? 4'b0111 : 4'b1111;
													assign node17044 = (inp[1]) ? node17048 : node17045;
														assign node17045 = (inp[14]) ? 4'b0110 : 4'b1110;
														assign node17048 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node17051 = (inp[1]) ? 4'b1010 : 4'b0110;
											assign node17054 = (inp[6]) ? node17068 : node17055;
												assign node17055 = (inp[14]) ? 4'b1011 : node17056;
													assign node17056 = (inp[8]) ? node17062 : node17057;
														assign node17057 = (inp[1]) ? 4'b1010 : node17058;
															assign node17058 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node17062 = (inp[7]) ? node17064 : 4'b1011;
															assign node17064 = (inp[1]) ? 4'b1011 : 4'b1010;
												assign node17068 = (inp[1]) ? node17076 : node17069;
													assign node17069 = (inp[7]) ? node17073 : node17070;
														assign node17070 = (inp[8]) ? 4'b0011 : 4'b1010;
														assign node17073 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node17076 = (inp[14]) ? 4'b0011 : node17077;
														assign node17077 = (inp[2]) ? node17079 : 4'b0010;
															assign node17079 = (inp[8]) ? 4'b0010 : 4'b0011;
										assign node17083 = (inp[2]) ? node17109 : node17084;
											assign node17084 = (inp[7]) ? node17096 : node17085;
												assign node17085 = (inp[6]) ? node17089 : node17086;
													assign node17086 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node17089 = (inp[11]) ? 4'b0011 : node17090;
														assign node17090 = (inp[8]) ? 4'b1011 : node17091;
															assign node17091 = (inp[1]) ? 4'b1011 : 4'b0011;
												assign node17096 = (inp[1]) ? node17104 : node17097;
													assign node17097 = (inp[14]) ? node17099 : 4'b1010;
														assign node17099 = (inp[8]) ? 4'b1010 : node17100;
															assign node17100 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node17104 = (inp[6]) ? 4'b0010 : node17105;
														assign node17105 = (inp[11]) ? 4'b1011 : 4'b0011;
											assign node17109 = (inp[11]) ? node17115 : node17110;
												assign node17110 = (inp[1]) ? 4'b1010 : node17111;
													assign node17111 = (inp[6]) ? 4'b1011 : 4'b1010;
												assign node17115 = (inp[6]) ? node17123 : node17116;
													assign node17116 = (inp[1]) ? 4'b1011 : node17117;
														assign node17117 = (inp[8]) ? node17119 : 4'b0010;
															assign node17119 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node17123 = (inp[1]) ? 4'b0010 : node17124;
														assign node17124 = (inp[8]) ? 4'b0010 : 4'b1010;
									assign node17128 = (inp[12]) ? node17168 : node17129;
										assign node17129 = (inp[6]) ? node17151 : node17130;
											assign node17130 = (inp[11]) ? node17140 : node17131;
												assign node17131 = (inp[8]) ? 4'b0011 : node17132;
													assign node17132 = (inp[14]) ? 4'b1010 : node17133;
														assign node17133 = (inp[2]) ? 4'b0011 : node17134;
															assign node17134 = (inp[1]) ? 4'b0011 : 4'b1011;
												assign node17140 = (inp[7]) ? node17146 : node17141;
													assign node17141 = (inp[8]) ? 4'b1101 : node17142;
														assign node17142 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node17146 = (inp[14]) ? node17148 : 4'b1101;
														assign node17148 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node17151 = (inp[11]) ? node17159 : node17152;
												assign node17152 = (inp[1]) ? 4'b1100 : node17153;
													assign node17153 = (inp[7]) ? node17155 : 4'b0010;
														assign node17155 = (inp[2]) ? 4'b1100 : 4'b0010;
												assign node17159 = (inp[1]) ? 4'b0100 : node17160;
													assign node17160 = (inp[2]) ? node17162 : 4'b1100;
														assign node17162 = (inp[8]) ? node17164 : 4'b1100;
															assign node17164 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node17168 = (inp[11]) ? node17192 : node17169;
											assign node17169 = (inp[14]) ? node17179 : node17170;
												assign node17170 = (inp[2]) ? 4'b0101 : node17171;
													assign node17171 = (inp[1]) ? node17173 : 4'b1100;
														assign node17173 = (inp[7]) ? node17175 : 4'b0100;
															assign node17175 = (inp[8]) ? 4'b0101 : 4'b0100;
												assign node17179 = (inp[1]) ? node17185 : node17180;
													assign node17180 = (inp[8]) ? 4'b0101 : node17181;
														assign node17181 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node17185 = (inp[2]) ? node17187 : 4'b1101;
														assign node17187 = (inp[7]) ? node17189 : 4'b1100;
															assign node17189 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node17192 = (inp[6]) ? node17200 : node17193;
												assign node17193 = (inp[2]) ? 4'b1101 : node17194;
													assign node17194 = (inp[8]) ? 4'b1101 : node17195;
														assign node17195 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node17200 = (inp[8]) ? 4'b0101 : node17201;
													assign node17201 = (inp[1]) ? 4'b0101 : 4'b1101;
								assign node17205 = (inp[4]) ? node17279 : node17206;
									assign node17206 = (inp[12]) ? node17246 : node17207;
										assign node17207 = (inp[11]) ? node17227 : node17208;
											assign node17208 = (inp[6]) ? node17218 : node17209;
												assign node17209 = (inp[8]) ? node17215 : node17210;
													assign node17210 = (inp[7]) ? 4'b0011 : node17211;
														assign node17211 = (inp[1]) ? 4'b0010 : 4'b1010;
													assign node17215 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node17218 = (inp[1]) ? 4'b1101 : node17219;
													assign node17219 = (inp[14]) ? 4'b1100 : node17220;
														assign node17220 = (inp[8]) ? 4'b0010 : node17221;
															assign node17221 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node17227 = (inp[6]) ? node17241 : node17228;
												assign node17228 = (inp[7]) ? node17234 : node17229;
													assign node17229 = (inp[14]) ? node17231 : 4'b1101;
														assign node17231 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node17234 = (inp[14]) ? 4'b1100 : node17235;
														assign node17235 = (inp[8]) ? node17237 : 4'b1100;
															assign node17237 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node17241 = (inp[7]) ? node17243 : 4'b1100;
													assign node17243 = (inp[8]) ? 4'b0100 : 4'b0101;
										assign node17246 = (inp[11]) ? node17266 : node17247;
											assign node17247 = (inp[6]) ? node17253 : node17248;
												assign node17248 = (inp[7]) ? node17250 : 4'b0101;
													assign node17250 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node17253 = (inp[8]) ? node17261 : node17254;
													assign node17254 = (inp[7]) ? node17258 : node17255;
														assign node17255 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node17258 = (inp[14]) ? 4'b1101 : 4'b0100;
													assign node17261 = (inp[14]) ? node17263 : 4'b1101;
														assign node17263 = (inp[1]) ? 4'b1100 : 4'b1101;
											assign node17266 = (inp[2]) ? node17272 : node17267;
												assign node17267 = (inp[7]) ? node17269 : 4'b0101;
													assign node17269 = (inp[14]) ? 4'b0100 : 4'b1101;
												assign node17272 = (inp[7]) ? node17276 : node17273;
													assign node17273 = (inp[8]) ? 4'b1101 : 4'b0100;
													assign node17276 = (inp[8]) ? 4'b0100 : 4'b0101;
									assign node17279 = (inp[12]) ? node17319 : node17280;
										assign node17280 = (inp[6]) ? node17302 : node17281;
											assign node17281 = (inp[11]) ? node17295 : node17282;
												assign node17282 = (inp[1]) ? node17290 : node17283;
													assign node17283 = (inp[8]) ? 4'b0101 : node17284;
														assign node17284 = (inp[14]) ? node17286 : 4'b1100;
															assign node17286 = (inp[7]) ? 4'b0101 : 4'b1100;
													assign node17290 = (inp[8]) ? 4'b0100 : node17291;
														assign node17291 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node17295 = (inp[14]) ? node17297 : 4'b1001;
													assign node17297 = (inp[7]) ? node17299 : 4'b0100;
														assign node17299 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node17302 = (inp[11]) ? node17312 : node17303;
												assign node17303 = (inp[1]) ? node17309 : node17304;
													assign node17304 = (inp[14]) ? 4'b1001 : node17305;
														assign node17305 = (inp[7]) ? 4'b1001 : 4'b0101;
													assign node17309 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node17312 = (inp[14]) ? node17314 : 4'b0001;
													assign node17314 = (inp[1]) ? 4'b0001 : node17315;
														assign node17315 = (inp[7]) ? 4'b0000 : 4'b1000;
										assign node17319 = (inp[1]) ? node17345 : node17320;
											assign node17320 = (inp[6]) ? node17334 : node17321;
												assign node17321 = (inp[14]) ? node17331 : node17322;
													assign node17322 = (inp[8]) ? node17326 : node17323;
														assign node17323 = (inp[2]) ? 4'b0000 : 4'b1000;
														assign node17326 = (inp[2]) ? node17328 : 4'b0000;
															assign node17328 = (inp[11]) ? 4'b1001 : 4'b0000;
													assign node17331 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node17334 = (inp[2]) ? node17340 : node17335;
													assign node17335 = (inp[8]) ? 4'b1001 : node17336;
														assign node17336 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node17340 = (inp[11]) ? node17342 : 4'b0000;
														assign node17342 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node17345 = (inp[11]) ? node17355 : node17346;
												assign node17346 = (inp[6]) ? node17348 : 4'b0000;
													assign node17348 = (inp[7]) ? node17352 : node17349;
														assign node17349 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node17352 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node17355 = (inp[6]) ? 4'b0000 : node17356;
													assign node17356 = (inp[7]) ? 4'b1001 : 4'b1000;
						assign node17360 = (inp[3]) ? node17710 : node17361;
							assign node17361 = (inp[9]) ? node17543 : node17362;
								assign node17362 = (inp[4]) ? node17460 : node17363;
									assign node17363 = (inp[6]) ? node17413 : node17364;
										assign node17364 = (inp[12]) ? node17386 : node17365;
											assign node17365 = (inp[11]) ? node17381 : node17366;
												assign node17366 = (inp[7]) ? node17374 : node17367;
													assign node17367 = (inp[1]) ? node17369 : 4'b1110;
														assign node17369 = (inp[2]) ? node17371 : 4'b0110;
															assign node17371 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node17374 = (inp[8]) ? node17376 : 4'b0111;
														assign node17376 = (inp[14]) ? 4'b0110 : node17377;
															assign node17377 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node17381 = (inp[8]) ? node17383 : 4'b0110;
													assign node17383 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node17386 = (inp[11]) ? node17404 : node17387;
												assign node17387 = (inp[7]) ? node17399 : node17388;
													assign node17388 = (inp[8]) ? node17394 : node17389;
														assign node17389 = (inp[1]) ? node17391 : 4'b1010;
															assign node17391 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node17394 = (inp[14]) ? 4'b0011 : node17395;
															assign node17395 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node17399 = (inp[8]) ? node17401 : 4'b0011;
														assign node17401 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node17404 = (inp[7]) ? node17410 : node17405;
													assign node17405 = (inp[8]) ? 4'b1011 : node17406;
														assign node17406 = (inp[1]) ? 4'b1010 : 4'b0010;
													assign node17410 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node17413 = (inp[11]) ? node17437 : node17414;
											assign node17414 = (inp[1]) ? node17426 : node17415;
												assign node17415 = (inp[2]) ? node17419 : node17416;
													assign node17416 = (inp[8]) ? 4'b1011 : 4'b0111;
													assign node17419 = (inp[8]) ? node17423 : node17420;
														assign node17420 = (inp[7]) ? 4'b1011 : 4'b0010;
														assign node17423 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node17426 = (inp[8]) ? node17434 : node17427;
													assign node17427 = (inp[7]) ? node17429 : 4'b1010;
														assign node17429 = (inp[14]) ? 4'b1011 : node17430;
															assign node17430 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node17434 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node17437 = (inp[1]) ? node17453 : node17438;
												assign node17438 = (inp[12]) ? node17444 : node17439;
													assign node17439 = (inp[7]) ? 4'b0011 : node17440;
														assign node17440 = (inp[2]) ? 4'b1010 : 4'b0011;
													assign node17444 = (inp[14]) ? node17448 : node17445;
														assign node17445 = (inp[2]) ? 4'b0011 : 4'b1010;
														assign node17448 = (inp[8]) ? node17450 : 4'b1010;
															assign node17450 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node17453 = (inp[14]) ? node17455 : 4'b0010;
													assign node17455 = (inp[8]) ? 4'b0011 : node17456;
														assign node17456 = (inp[7]) ? 4'b0011 : 4'b0010;
									assign node17460 = (inp[12]) ? node17498 : node17461;
										assign node17461 = (inp[11]) ? node17483 : node17462;
											assign node17462 = (inp[6]) ? node17470 : node17463;
												assign node17463 = (inp[7]) ? node17467 : node17464;
													assign node17464 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node17467 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node17470 = (inp[8]) ? node17480 : node17471;
													assign node17471 = (inp[1]) ? node17477 : node17472;
														assign node17472 = (inp[14]) ? 4'b0010 : node17473;
															assign node17473 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node17477 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node17480 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node17483 = (inp[6]) ? node17493 : node17484;
												assign node17484 = (inp[8]) ? node17488 : node17485;
													assign node17485 = (inp[7]) ? 4'b1101 : 4'b0010;
													assign node17488 = (inp[7]) ? node17490 : 4'b1101;
														assign node17490 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node17493 = (inp[14]) ? 4'b0100 : node17494;
													assign node17494 = (inp[8]) ? 4'b0101 : 4'b0100;
										assign node17498 = (inp[7]) ? node17528 : node17499;
											assign node17499 = (inp[8]) ? node17509 : node17500;
												assign node17500 = (inp[2]) ? node17506 : node17501;
													assign node17501 = (inp[14]) ? 4'b0100 : node17502;
														assign node17502 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node17506 = (inp[14]) ? 4'b1100 : 4'b0100;
												assign node17509 = (inp[2]) ? node17517 : node17510;
													assign node17510 = (inp[14]) ? node17512 : 4'b1100;
														assign node17512 = (inp[1]) ? node17514 : 4'b1101;
															assign node17514 = (inp[6]) ? 4'b1101 : 4'b0101;
													assign node17517 = (inp[1]) ? node17523 : node17518;
														assign node17518 = (inp[11]) ? node17520 : 4'b1101;
															assign node17520 = (inp[6]) ? 4'b0101 : 4'b1101;
														assign node17523 = (inp[11]) ? node17525 : 4'b0101;
															assign node17525 = (inp[6]) ? 4'b0101 : 4'b1101;
											assign node17528 = (inp[1]) ? node17532 : node17529;
												assign node17529 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node17532 = (inp[14]) ? 4'b0100 : node17533;
													assign node17533 = (inp[8]) ? node17537 : node17534;
														assign node17534 = (inp[6]) ? 4'b1101 : 4'b0101;
														assign node17537 = (inp[11]) ? node17539 : 4'b0101;
															assign node17539 = (inp[6]) ? 4'b0101 : 4'b1101;
								assign node17543 = (inp[4]) ? node17637 : node17544;
									assign node17544 = (inp[12]) ? node17582 : node17545;
										assign node17545 = (inp[11]) ? node17553 : node17546;
											assign node17546 = (inp[6]) ? node17550 : node17547;
												assign node17547 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node17550 = (inp[7]) ? 4'b1100 : 4'b0010;
											assign node17553 = (inp[6]) ? node17565 : node17554;
												assign node17554 = (inp[1]) ? node17558 : node17555;
													assign node17555 = (inp[2]) ? 4'b1101 : 4'b0010;
													assign node17558 = (inp[7]) ? 4'b1100 : node17559;
														assign node17559 = (inp[2]) ? 4'b1100 : node17560;
															assign node17560 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node17565 = (inp[1]) ? node17573 : node17566;
													assign node17566 = (inp[2]) ? 4'b0101 : node17567;
														assign node17567 = (inp[7]) ? node17569 : 4'b1100;
															assign node17569 = (inp[14]) ? 4'b0100 : 4'b1100;
													assign node17573 = (inp[2]) ? node17579 : node17574;
														assign node17574 = (inp[14]) ? 4'b0101 : node17575;
															assign node17575 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node17579 = (inp[8]) ? 4'b0100 : 4'b0101;
										assign node17582 = (inp[1]) ? node17606 : node17583;
											assign node17583 = (inp[7]) ? node17597 : node17584;
												assign node17584 = (inp[2]) ? node17592 : node17585;
													assign node17585 = (inp[8]) ? node17587 : 4'b0101;
														assign node17587 = (inp[14]) ? 4'b1101 : node17588;
															assign node17588 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node17592 = (inp[8]) ? node17594 : 4'b1100;
														assign node17594 = (inp[14]) ? 4'b0101 : 4'b1101;
												assign node17597 = (inp[8]) ? node17601 : node17598;
													assign node17598 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node17601 = (inp[6]) ? 4'b0100 : node17602;
														assign node17602 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node17606 = (inp[14]) ? node17622 : node17607;
												assign node17607 = (inp[8]) ? node17619 : node17608;
													assign node17608 = (inp[11]) ? node17614 : node17609;
														assign node17609 = (inp[7]) ? 4'b0101 : node17610;
															assign node17610 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node17614 = (inp[7]) ? node17616 : 4'b1101;
															assign node17616 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node17619 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node17622 = (inp[8]) ? node17632 : node17623;
													assign node17623 = (inp[2]) ? node17627 : node17624;
														assign node17624 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node17627 = (inp[11]) ? node17629 : 4'b1100;
															assign node17629 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node17632 = (inp[7]) ? node17634 : 4'b1101;
														assign node17634 = (inp[6]) ? 4'b1100 : 4'b0100;
									assign node17637 = (inp[12]) ? node17675 : node17638;
										assign node17638 = (inp[11]) ? node17656 : node17639;
											assign node17639 = (inp[6]) ? node17649 : node17640;
												assign node17640 = (inp[8]) ? node17642 : 4'b0101;
													assign node17642 = (inp[1]) ? node17644 : 4'b0100;
														assign node17644 = (inp[14]) ? 4'b0101 : node17645;
															assign node17645 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node17649 = (inp[7]) ? node17653 : node17650;
													assign node17650 = (inp[1]) ? 4'b1000 : 4'b0100;
													assign node17653 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node17656 = (inp[6]) ? node17666 : node17657;
												assign node17657 = (inp[14]) ? node17661 : node17658;
													assign node17658 = (inp[7]) ? 4'b1001 : 4'b0100;
													assign node17661 = (inp[7]) ? 4'b1000 : node17662;
														assign node17662 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node17666 = (inp[14]) ? 4'b0001 : node17667;
													assign node17667 = (inp[7]) ? node17671 : node17668;
														assign node17668 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node17671 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node17675 = (inp[11]) ? node17691 : node17676;
											assign node17676 = (inp[6]) ? node17682 : node17677;
												assign node17677 = (inp[7]) ? node17679 : 4'b0001;
													assign node17679 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node17682 = (inp[2]) ? node17688 : node17683;
													assign node17683 = (inp[8]) ? node17685 : 4'b1001;
														assign node17685 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node17688 = (inp[8]) ? 4'b1001 : 4'b0000;
											assign node17691 = (inp[6]) ? node17701 : node17692;
												assign node17692 = (inp[14]) ? 4'b1001 : node17693;
													assign node17693 = (inp[7]) ? 4'b1001 : node17694;
														assign node17694 = (inp[8]) ? 4'b1001 : node17695;
															assign node17695 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node17701 = (inp[8]) ? 4'b0000 : node17702;
													assign node17702 = (inp[14]) ? 4'b0001 : node17703;
														assign node17703 = (inp[1]) ? node17705 : 4'b1000;
															assign node17705 = (inp[7]) ? 4'b0000 : 4'b0001;
							assign node17710 = (inp[14]) ? node17914 : node17711;
								assign node17711 = (inp[1]) ? node17809 : node17712;
									assign node17712 = (inp[2]) ? node17760 : node17713;
										assign node17713 = (inp[7]) ? node17737 : node17714;
											assign node17714 = (inp[8]) ? node17730 : node17715;
												assign node17715 = (inp[12]) ? node17717 : 4'b0001;
													assign node17717 = (inp[6]) ? node17723 : node17718;
														assign node17718 = (inp[11]) ? node17720 : 4'b1001;
															assign node17720 = (inp[9]) ? 4'b0001 : 4'b0001;
														assign node17723 = (inp[9]) ? node17727 : node17724;
															assign node17724 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node17727 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node17730 = (inp[11]) ? node17732 : 4'b1100;
													assign node17732 = (inp[6]) ? 4'b1000 : node17733;
														assign node17733 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node17737 = (inp[8]) ? node17749 : node17738;
												assign node17738 = (inp[4]) ? 4'b1000 : node17739;
													assign node17739 = (inp[11]) ? node17743 : node17740;
														assign node17740 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node17743 = (inp[9]) ? 4'b1100 : node17744;
															assign node17744 = (inp[6]) ? 4'b1000 : 4'b0000;
												assign node17749 = (inp[9]) ? node17753 : node17750;
													assign node17750 = (inp[6]) ? 4'b0001 : 4'b0101;
													assign node17753 = (inp[4]) ? node17755 : 4'b1101;
														assign node17755 = (inp[6]) ? 4'b1001 : node17756;
															assign node17756 = (inp[11]) ? 4'b1001 : 4'b0001;
										assign node17760 = (inp[4]) ? node17786 : node17761;
											assign node17761 = (inp[6]) ? node17775 : node17762;
												assign node17762 = (inp[7]) ? node17770 : node17763;
													assign node17763 = (inp[8]) ? node17765 : 4'b0100;
														assign node17765 = (inp[11]) ? 4'b1001 : node17766;
															assign node17766 = (inp[12]) ? 4'b0001 : 4'b0001;
													assign node17770 = (inp[12]) ? 4'b0001 : node17771;
														assign node17771 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node17775 = (inp[7]) ? node17781 : node17776;
													assign node17776 = (inp[11]) ? node17778 : 4'b0100;
														assign node17778 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node17781 = (inp[11]) ? node17783 : 4'b1101;
														assign node17783 = (inp[9]) ? 4'b0101 : 4'b0001;
											assign node17786 = (inp[9]) ? node17800 : node17787;
												assign node17787 = (inp[6]) ? node17793 : node17788;
													assign node17788 = (inp[7]) ? node17790 : 4'b1100;
														assign node17790 = (inp[12]) ? 4'b1101 : 4'b1100;
													assign node17793 = (inp[12]) ? node17797 : node17794;
														assign node17794 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node17797 = (inp[11]) ? 4'b1100 : 4'b0100;
												assign node17800 = (inp[11]) ? 4'b0001 : node17801;
													assign node17801 = (inp[12]) ? 4'b0000 : node17802;
														assign node17802 = (inp[6]) ? node17804 : 4'b0100;
															assign node17804 = (inp[8]) ? 4'b1001 : 4'b0100;
									assign node17809 = (inp[9]) ? node17865 : node17810;
										assign node17810 = (inp[4]) ? node17836 : node17811;
											assign node17811 = (inp[6]) ? node17823 : node17812;
												assign node17812 = (inp[11]) ? node17818 : node17813;
													assign node17813 = (inp[2]) ? 4'b0100 : node17814;
														assign node17814 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node17818 = (inp[8]) ? 4'b1001 : node17819;
														assign node17819 = (inp[12]) ? 4'b1001 : 4'b1000;
												assign node17823 = (inp[11]) ? node17827 : node17824;
													assign node17824 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node17827 = (inp[2]) ? node17829 : 4'b0000;
														assign node17829 = (inp[7]) ? node17833 : node17830;
															assign node17830 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node17833 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node17836 = (inp[11]) ? node17852 : node17837;
												assign node17837 = (inp[12]) ? node17845 : node17838;
													assign node17838 = (inp[6]) ? 4'b1100 : node17839;
														assign node17839 = (inp[8]) ? 4'b0001 : node17840;
															assign node17840 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node17845 = (inp[2]) ? 4'b0101 : node17846;
														assign node17846 = (inp[8]) ? node17848 : 4'b0100;
															assign node17848 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node17852 = (inp[6]) ? node17858 : node17853;
													assign node17853 = (inp[8]) ? 4'b1100 : node17854;
														assign node17854 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node17858 = (inp[12]) ? 4'b0100 : node17859;
														assign node17859 = (inp[8]) ? 4'b0101 : node17860;
															assign node17860 = (inp[2]) ? 4'b0100 : 4'b0101;
										assign node17865 = (inp[4]) ? node17881 : node17866;
											assign node17866 = (inp[6]) ? node17874 : node17867;
												assign node17867 = (inp[11]) ? 4'b1100 : node17868;
													assign node17868 = (inp[2]) ? node17870 : 4'b0001;
														assign node17870 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node17874 = (inp[11]) ? 4'b0100 : node17875;
													assign node17875 = (inp[7]) ? node17877 : 4'b1101;
														assign node17877 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node17881 = (inp[7]) ? node17895 : node17882;
												assign node17882 = (inp[12]) ? node17890 : node17883;
													assign node17883 = (inp[11]) ? node17887 : node17884;
														assign node17884 = (inp[6]) ? 4'b1001 : 4'b0101;
														assign node17887 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node17890 = (inp[11]) ? node17892 : 4'b1000;
														assign node17892 = (inp[6]) ? 4'b0001 : 4'b1000;
												assign node17895 = (inp[8]) ? node17907 : node17896;
													assign node17896 = (inp[2]) ? node17900 : node17897;
														assign node17897 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node17900 = (inp[12]) ? node17904 : node17901;
															assign node17901 = (inp[11]) ? 4'b0001 : 4'b0101;
															assign node17904 = (inp[6]) ? 4'b0001 : 4'b0001;
													assign node17907 = (inp[2]) ? 4'b1000 : node17908;
														assign node17908 = (inp[12]) ? node17910 : 4'b1001;
															assign node17910 = (inp[6]) ? 4'b0001 : 4'b1001;
								assign node17914 = (inp[2]) ? node18036 : node17915;
									assign node17915 = (inp[12]) ? node17969 : node17916;
										assign node17916 = (inp[1]) ? node17950 : node17917;
											assign node17917 = (inp[6]) ? node17947 : node17918;
												assign node17918 = (inp[11]) ? node17932 : node17919;
													assign node17919 = (inp[7]) ? node17925 : node17920;
														assign node17920 = (inp[8]) ? 4'b0101 : node17921;
															assign node17921 = (inp[9]) ? 4'b1000 : 4'b1000;
														assign node17925 = (inp[8]) ? node17929 : node17926;
															assign node17926 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node17929 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node17932 = (inp[7]) ? node17940 : node17933;
														assign node17933 = (inp[8]) ? node17937 : node17934;
															assign node17934 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node17937 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node17940 = (inp[8]) ? node17944 : node17941;
															assign node17941 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node17944 = (inp[9]) ? 4'b1000 : 4'b1000;
												assign node17947 = (inp[11]) ? 4'b0100 : 4'b1001;
											assign node17950 = (inp[6]) ? node17954 : node17951;
												assign node17951 = (inp[11]) ? 4'b1000 : 4'b0000;
												assign node17954 = (inp[8]) ? node17960 : node17955;
													assign node17955 = (inp[4]) ? 4'b1001 : node17956;
														assign node17956 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node17960 = (inp[7]) ? node17962 : 4'b1101;
														assign node17962 = (inp[9]) ? node17966 : node17963;
															assign node17963 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node17966 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node17969 = (inp[9]) ? node18005 : node17970;
											assign node17970 = (inp[4]) ? node17994 : node17971;
												assign node17971 = (inp[1]) ? node17985 : node17972;
													assign node17972 = (inp[6]) ? node17978 : node17973;
														assign node17973 = (inp[11]) ? 4'b1001 : node17974;
															assign node17974 = (inp[8]) ? 4'b0001 : 4'b1000;
														assign node17978 = (inp[7]) ? node17982 : node17979;
															assign node17979 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node17982 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node17985 = (inp[11]) ? node17989 : node17986;
														assign node17986 = (inp[8]) ? 4'b1001 : 4'b0001;
														assign node17989 = (inp[6]) ? node17991 : 4'b1000;
															assign node17991 = (inp[7]) ? 4'b0000 : 4'b0000;
												assign node17994 = (inp[6]) ? node18002 : node17995;
													assign node17995 = (inp[11]) ? node17997 : 4'b0101;
														assign node17997 = (inp[8]) ? node17999 : 4'b1100;
															assign node17999 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node18002 = (inp[11]) ? 4'b0100 : 4'b1100;
											assign node18005 = (inp[4]) ? node18011 : node18006;
												assign node18006 = (inp[7]) ? 4'b1101 : node18007;
													assign node18007 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node18011 = (inp[1]) ? node18023 : node18012;
													assign node18012 = (inp[6]) ? node18018 : node18013;
														assign node18013 = (inp[11]) ? 4'b1001 : node18014;
															assign node18014 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node18018 = (inp[11]) ? 4'b0000 : node18019;
															assign node18019 = (inp[8]) ? 4'b1001 : 4'b0000;
													assign node18023 = (inp[7]) ? node18029 : node18024;
														assign node18024 = (inp[6]) ? node18026 : 4'b1000;
															assign node18026 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node18029 = (inp[6]) ? node18033 : node18030;
															assign node18030 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node18033 = (inp[11]) ? 4'b0001 : 4'b1001;
									assign node18036 = (inp[12]) ? node18094 : node18037;
										assign node18037 = (inp[7]) ? node18067 : node18038;
											assign node18038 = (inp[8]) ? node18054 : node18039;
												assign node18039 = (inp[4]) ? node18051 : node18040;
													assign node18040 = (inp[1]) ? node18046 : node18041;
														assign node18041 = (inp[6]) ? 4'b1100 : node18042;
															assign node18042 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node18046 = (inp[9]) ? node18048 : 4'b0000;
															assign node18048 = (inp[6]) ? 4'b1100 : 4'b0000;
													assign node18051 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node18054 = (inp[9]) ? node18060 : node18055;
													assign node18055 = (inp[6]) ? 4'b0001 : node18056;
														assign node18056 = (inp[4]) ? 4'b0001 : 4'b1001;
													assign node18060 = (inp[4]) ? node18062 : 4'b1101;
														assign node18062 = (inp[6]) ? 4'b1001 : node18063;
															assign node18063 = (inp[11]) ? 4'b1001 : 4'b0101;
											assign node18067 = (inp[8]) ? node18083 : node18068;
												assign node18068 = (inp[1]) ? node18074 : node18069;
													assign node18069 = (inp[6]) ? node18071 : 4'b0001;
														assign node18071 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node18074 = (inp[6]) ? node18078 : node18075;
														assign node18075 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node18078 = (inp[11]) ? node18080 : 4'b1001;
															assign node18080 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node18083 = (inp[9]) ? node18087 : node18084;
													assign node18084 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node18087 = (inp[6]) ? 4'b0000 : node18088;
														assign node18088 = (inp[11]) ? 4'b1100 : node18089;
															assign node18089 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node18094 = (inp[8]) ? node18118 : node18095;
											assign node18095 = (inp[7]) ? node18109 : node18096;
												assign node18096 = (inp[1]) ? node18102 : node18097;
													assign node18097 = (inp[11]) ? node18099 : 4'b1100;
														assign node18099 = (inp[6]) ? 4'b1100 : 4'b0100;
													assign node18102 = (inp[6]) ? node18104 : 4'b1000;
														assign node18104 = (inp[4]) ? 4'b0000 : node18105;
															assign node18105 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node18109 = (inp[4]) ? node18111 : 4'b0101;
													assign node18111 = (inp[9]) ? node18115 : node18112;
														assign node18112 = (inp[6]) ? 4'b0101 : 4'b1101;
														assign node18115 = (inp[6]) ? 4'b0001 : 4'b1001;
											assign node18118 = (inp[7]) ? node18132 : node18119;
												assign node18119 = (inp[1]) ? node18125 : node18120;
													assign node18120 = (inp[9]) ? 4'b1001 : node18121;
														assign node18121 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node18125 = (inp[11]) ? 4'b0001 : node18126;
														assign node18126 = (inp[9]) ? 4'b1101 : node18127;
															assign node18127 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node18132 = (inp[11]) ? node18140 : node18133;
													assign node18133 = (inp[6]) ? node18135 : 4'b0100;
														assign node18135 = (inp[1]) ? node18137 : 4'b1000;
															assign node18137 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node18140 = (inp[1]) ? node18144 : node18141;
														assign node18141 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node18144 = (inp[4]) ? node18146 : 4'b1000;
															assign node18146 = (inp[9]) ? 4'b1000 : 4'b1100;
					assign node18149 = (inp[3]) ? node18865 : node18150;
						assign node18150 = (inp[5]) ? node18524 : node18151;
							assign node18151 = (inp[1]) ? node18341 : node18152;
								assign node18152 = (inp[4]) ? node18232 : node18153;
									assign node18153 = (inp[9]) ? node18197 : node18154;
										assign node18154 = (inp[8]) ? node18176 : node18155;
											assign node18155 = (inp[7]) ? node18163 : node18156;
												assign node18156 = (inp[14]) ? node18158 : 4'b0101;
													assign node18158 = (inp[11]) ? node18160 : 4'b1100;
														assign node18160 = (inp[6]) ? 4'b1000 : 4'b0000;
												assign node18163 = (inp[6]) ? node18171 : node18164;
													assign node18164 = (inp[11]) ? node18166 : 4'b0101;
														assign node18166 = (inp[2]) ? 4'b1001 : node18167;
															assign node18167 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node18171 = (inp[11]) ? 4'b0001 : node18172;
														assign node18172 = (inp[2]) ? 4'b1001 : 4'b0000;
											assign node18176 = (inp[6]) ? node18190 : node18177;
												assign node18177 = (inp[11]) ? node18183 : node18178;
													assign node18178 = (inp[12]) ? 4'b0001 : node18179;
														assign node18179 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node18183 = (inp[2]) ? 4'b1000 : node18184;
														assign node18184 = (inp[12]) ? node18186 : 4'b1001;
															assign node18186 = (inp[14]) ? 4'b1000 : 4'b0000;
												assign node18190 = (inp[7]) ? node18194 : node18191;
													assign node18191 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node18194 = (inp[11]) ? 4'b0000 : 4'b1000;
										assign node18197 = (inp[7]) ? node18211 : node18198;
											assign node18198 = (inp[8]) ? node18206 : node18199;
												assign node18199 = (inp[12]) ? 4'b1100 : node18200;
													assign node18200 = (inp[6]) ? 4'b1100 : node18201;
														assign node18201 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node18206 = (inp[2]) ? node18208 : 4'b1000;
													assign node18208 = (inp[14]) ? 4'b0101 : 4'b1101;
											assign node18211 = (inp[6]) ? node18219 : node18212;
												assign node18212 = (inp[11]) ? node18214 : 4'b0101;
													assign node18214 = (inp[2]) ? node18216 : 4'b1101;
														assign node18216 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node18219 = (inp[11]) ? node18225 : node18220;
													assign node18220 = (inp[2]) ? node18222 : 4'b0100;
														assign node18222 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node18225 = (inp[14]) ? node18229 : node18226;
														assign node18226 = (inp[8]) ? 4'b0101 : 4'b1100;
														assign node18229 = (inp[8]) ? 4'b0100 : 4'b0101;
									assign node18232 = (inp[9]) ? node18288 : node18233;
										assign node18233 = (inp[11]) ? node18261 : node18234;
											assign node18234 = (inp[12]) ? node18248 : node18235;
												assign node18235 = (inp[14]) ? node18245 : node18236;
													assign node18236 = (inp[8]) ? node18242 : node18237;
														assign node18237 = (inp[6]) ? 4'b1101 : node18238;
															assign node18238 = (inp[7]) ? 4'b0001 : 4'b1001;
														assign node18242 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node18245 = (inp[8]) ? 4'b1101 : 4'b1000;
												assign node18248 = (inp[6]) ? node18252 : node18249;
													assign node18249 = (inp[8]) ? 4'b0100 : 4'b1100;
													assign node18252 = (inp[7]) ? node18258 : node18253;
														assign node18253 = (inp[8]) ? 4'b1101 : node18254;
															assign node18254 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node18258 = (inp[14]) ? 4'b1101 : 4'b1100;
											assign node18261 = (inp[6]) ? node18277 : node18262;
												assign node18262 = (inp[8]) ? node18272 : node18263;
													assign node18263 = (inp[12]) ? node18265 : 4'b0000;
														assign node18265 = (inp[14]) ? node18269 : node18266;
															assign node18266 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node18269 = (inp[7]) ? 4'b1101 : 4'b0100;
													assign node18272 = (inp[12]) ? node18274 : 4'b1100;
														assign node18274 = (inp[2]) ? 4'b1101 : 4'b0100;
												assign node18277 = (inp[12]) ? 4'b0101 : node18278;
													assign node18278 = (inp[7]) ? node18280 : 4'b0101;
														assign node18280 = (inp[8]) ? node18284 : node18281;
															assign node18281 = (inp[2]) ? 4'b0101 : 4'b1100;
															assign node18284 = (inp[14]) ? 4'b0100 : 4'b0100;
										assign node18288 = (inp[12]) ? node18316 : node18289;
											assign node18289 = (inp[11]) ? node18307 : node18290;
												assign node18290 = (inp[14]) ? node18298 : node18291;
													assign node18291 = (inp[6]) ? 4'b1001 : node18292;
														assign node18292 = (inp[2]) ? node18294 : 4'b1100;
															assign node18294 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node18298 = (inp[2]) ? node18302 : node18299;
														assign node18299 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node18302 = (inp[8]) ? 4'b0100 : node18303;
															assign node18303 = (inp[6]) ? 4'b0100 : 4'b1100;
												assign node18307 = (inp[8]) ? node18309 : 4'b1000;
													assign node18309 = (inp[7]) ? node18313 : node18310;
														assign node18310 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node18313 = (inp[6]) ? 4'b0000 : 4'b1000;
											assign node18316 = (inp[2]) ? node18334 : node18317;
												assign node18317 = (inp[7]) ? node18329 : node18318;
													assign node18318 = (inp[8]) ? node18324 : node18319;
														assign node18319 = (inp[14]) ? 4'b1000 : node18320;
															assign node18320 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node18324 = (inp[6]) ? node18326 : 4'b0001;
															assign node18326 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node18329 = (inp[6]) ? node18331 : 4'b0000;
														assign node18331 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node18334 = (inp[8]) ? node18338 : node18335;
													assign node18335 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node18338 = (inp[7]) ? 4'b0000 : 4'b0001;
								assign node18341 = (inp[14]) ? node18435 : node18342;
									assign node18342 = (inp[11]) ? node18380 : node18343;
										assign node18343 = (inp[6]) ? node18369 : node18344;
											assign node18344 = (inp[9]) ? node18358 : node18345;
												assign node18345 = (inp[2]) ? node18355 : node18346;
													assign node18346 = (inp[8]) ? node18352 : node18347;
														assign node18347 = (inp[7]) ? 4'b0100 : node18348;
															assign node18348 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node18352 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node18355 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node18358 = (inp[7]) ? 4'b0100 : node18359;
													assign node18359 = (inp[2]) ? node18363 : node18360;
														assign node18360 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node18363 = (inp[8]) ? 4'b0101 : node18364;
															assign node18364 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node18369 = (inp[2]) ? node18377 : node18370;
												assign node18370 = (inp[8]) ? node18374 : node18371;
													assign node18371 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node18374 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node18377 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node18380 = (inp[6]) ? node18410 : node18381;
											assign node18381 = (inp[8]) ? node18401 : node18382;
												assign node18382 = (inp[12]) ? node18394 : node18383;
													assign node18383 = (inp[2]) ? node18389 : node18384;
														assign node18384 = (inp[7]) ? 4'b1000 : node18385;
															assign node18385 = (inp[4]) ? 4'b1001 : 4'b1001;
														assign node18389 = (inp[7]) ? node18391 : 4'b1100;
															assign node18391 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node18394 = (inp[9]) ? node18396 : 4'b1000;
														assign node18396 = (inp[4]) ? 4'b1000 : node18397;
															assign node18397 = (inp[2]) ? 4'b1100 : 4'b1100;
												assign node18401 = (inp[12]) ? 4'b1101 : node18402;
													assign node18402 = (inp[9]) ? node18404 : 4'b1100;
														assign node18404 = (inp[4]) ? 4'b1001 : node18405;
															assign node18405 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node18410 = (inp[7]) ? node18422 : node18411;
												assign node18411 = (inp[12]) ? node18417 : node18412;
													assign node18412 = (inp[8]) ? node18414 : 4'b0101;
														assign node18414 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node18417 = (inp[9]) ? node18419 : 4'b0100;
														assign node18419 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node18422 = (inp[8]) ? node18428 : node18423;
													assign node18423 = (inp[2]) ? node18425 : 4'b0100;
														assign node18425 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node18428 = (inp[12]) ? 4'b0001 : node18429;
														assign node18429 = (inp[9]) ? node18431 : 4'b0101;
															assign node18431 = (inp[4]) ? 4'b0001 : 4'b0101;
									assign node18435 = (inp[9]) ? node18477 : node18436;
										assign node18436 = (inp[4]) ? node18462 : node18437;
											assign node18437 = (inp[2]) ? node18449 : node18438;
												assign node18438 = (inp[7]) ? node18442 : node18439;
													assign node18439 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node18442 = (inp[12]) ? node18444 : 4'b0001;
														assign node18444 = (inp[6]) ? 4'b1001 : node18445;
															assign node18445 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node18449 = (inp[11]) ? node18453 : node18450;
													assign node18450 = (inp[12]) ? 4'b1000 : 4'b0100;
													assign node18453 = (inp[6]) ? 4'b0001 : node18454;
														assign node18454 = (inp[12]) ? node18458 : node18455;
															assign node18455 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node18458 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node18462 = (inp[7]) ? node18468 : node18463;
												assign node18463 = (inp[8]) ? 4'b1101 : node18464;
													assign node18464 = (inp[12]) ? 4'b0100 : 4'b1100;
												assign node18468 = (inp[8]) ? node18472 : node18469;
													assign node18469 = (inp[2]) ? 4'b1101 : 4'b0101;
													assign node18472 = (inp[2]) ? node18474 : 4'b0100;
														assign node18474 = (inp[11]) ? 4'b1100 : 4'b0100;
										assign node18477 = (inp[4]) ? node18511 : node18478;
											assign node18478 = (inp[12]) ? node18496 : node18479;
												assign node18479 = (inp[6]) ? node18489 : node18480;
													assign node18480 = (inp[11]) ? 4'b1101 : node18481;
														assign node18481 = (inp[8]) ? node18485 : node18482;
															assign node18482 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node18485 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node18489 = (inp[11]) ? node18491 : 4'b1101;
														assign node18491 = (inp[7]) ? node18493 : 4'b0101;
															assign node18493 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node18496 = (inp[7]) ? node18504 : node18497;
													assign node18497 = (inp[8]) ? node18499 : 4'b0100;
														assign node18499 = (inp[6]) ? 4'b0101 : node18500;
															assign node18500 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node18504 = (inp[8]) ? 4'b1100 : node18505;
														assign node18505 = (inp[2]) ? 4'b1101 : node18506;
															assign node18506 = (inp[11]) ? 4'b1101 : 4'b0101;
											assign node18511 = (inp[7]) ? node18515 : node18512;
												assign node18512 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node18515 = (inp[8]) ? 4'b1000 : node18516;
													assign node18516 = (inp[2]) ? 4'b1001 : node18517;
														assign node18517 = (inp[11]) ? 4'b0001 : node18518;
															assign node18518 = (inp[12]) ? 4'b0001 : 4'b0101;
							assign node18524 = (inp[4]) ? node18674 : node18525;
								assign node18525 = (inp[9]) ? node18609 : node18526;
									assign node18526 = (inp[11]) ? node18570 : node18527;
										assign node18527 = (inp[12]) ? node18551 : node18528;
											assign node18528 = (inp[6]) ? node18540 : node18529;
												assign node18529 = (inp[1]) ? node18535 : node18530;
													assign node18530 = (inp[7]) ? node18532 : 4'b0101;
														assign node18532 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node18535 = (inp[7]) ? node18537 : 4'b0100;
														assign node18537 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node18540 = (inp[1]) ? node18548 : node18541;
													assign node18541 = (inp[7]) ? 4'b1001 : node18542;
														assign node18542 = (inp[14]) ? 4'b0100 : node18543;
															assign node18543 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node18548 = (inp[8]) ? 4'b1001 : 4'b1000;
											assign node18551 = (inp[6]) ? node18561 : node18552;
												assign node18552 = (inp[1]) ? node18554 : 4'b0001;
													assign node18554 = (inp[8]) ? node18556 : 4'b0001;
														assign node18556 = (inp[14]) ? node18558 : 4'b0000;
															assign node18558 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node18561 = (inp[8]) ? node18567 : node18562;
													assign node18562 = (inp[14]) ? 4'b1001 : node18563;
														assign node18563 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node18567 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node18570 = (inp[6]) ? node18596 : node18571;
											assign node18571 = (inp[7]) ? node18587 : node18572;
												assign node18572 = (inp[1]) ? node18582 : node18573;
													assign node18573 = (inp[12]) ? node18579 : node18574;
														assign node18574 = (inp[14]) ? 4'b0100 : node18575;
															assign node18575 = (inp[2]) ? 4'b1001 : 4'b0100;
														assign node18579 = (inp[2]) ? 4'b1001 : 4'b0001;
													assign node18582 = (inp[12]) ? 4'b1000 : node18583;
														assign node18583 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node18587 = (inp[8]) ? node18593 : node18588;
													assign node18588 = (inp[14]) ? 4'b1001 : node18589;
														assign node18589 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node18593 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node18596 = (inp[8]) ? node18598 : 4'b0001;
												assign node18598 = (inp[2]) ? node18606 : node18599;
													assign node18599 = (inp[7]) ? 4'b0001 : node18600;
														assign node18600 = (inp[1]) ? node18602 : 4'b1000;
															assign node18602 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node18606 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node18609 = (inp[12]) ? node18645 : node18610;
										assign node18610 = (inp[1]) ? node18630 : node18611;
											assign node18611 = (inp[11]) ? node18619 : node18612;
												assign node18612 = (inp[8]) ? 4'b0000 : node18613;
													assign node18613 = (inp[2]) ? 4'b1111 : node18614;
														assign node18614 = (inp[6]) ? 4'b0000 : 4'b0001;
												assign node18619 = (inp[8]) ? node18623 : node18620;
													assign node18620 = (inp[6]) ? 4'b1110 : 4'b0000;
													assign node18623 = (inp[6]) ? node18627 : node18624;
														assign node18624 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node18627 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node18630 = (inp[11]) ? node18634 : node18631;
												assign node18631 = (inp[6]) ? 4'b1111 : 4'b0001;
												assign node18634 = (inp[6]) ? node18636 : 4'b1111;
													assign node18636 = (inp[14]) ? node18638 : 4'b0110;
														assign node18638 = (inp[7]) ? node18642 : node18639;
															assign node18639 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node18642 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node18645 = (inp[6]) ? node18653 : node18646;
											assign node18646 = (inp[11]) ? 4'b1111 : node18647;
												assign node18647 = (inp[14]) ? 4'b0111 : node18648;
													assign node18648 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node18653 = (inp[11]) ? node18663 : node18654;
												assign node18654 = (inp[1]) ? 4'b1110 : node18655;
													assign node18655 = (inp[7]) ? 4'b1111 : node18656;
														assign node18656 = (inp[14]) ? node18658 : 4'b0110;
															assign node18658 = (inp[8]) ? 4'b1111 : 4'b0110;
												assign node18663 = (inp[8]) ? node18669 : node18664;
													assign node18664 = (inp[14]) ? 4'b1110 : node18665;
														assign node18665 = (inp[7]) ? 4'b0111 : 4'b1111;
													assign node18669 = (inp[7]) ? 4'b0110 : node18670;
														assign node18670 = (inp[14]) ? 4'b0111 : 4'b0110;
								assign node18674 = (inp[9]) ? node18758 : node18675;
									assign node18675 = (inp[12]) ? node18717 : node18676;
										assign node18676 = (inp[6]) ? node18704 : node18677;
											assign node18677 = (inp[11]) ? node18691 : node18678;
												assign node18678 = (inp[2]) ? node18686 : node18679;
													assign node18679 = (inp[1]) ? 4'b0000 : node18680;
														assign node18680 = (inp[8]) ? 4'b1000 : node18681;
															assign node18681 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node18686 = (inp[7]) ? node18688 : 4'b0001;
														assign node18688 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node18691 = (inp[1]) ? node18697 : node18692;
													assign node18692 = (inp[2]) ? 4'b1111 : node18693;
														assign node18693 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node18697 = (inp[8]) ? 4'b1111 : node18698;
														assign node18698 = (inp[7]) ? node18700 : 4'b1110;
															assign node18700 = (inp[14]) ? 4'b1111 : 4'b1110;
											assign node18704 = (inp[11]) ? node18708 : node18705;
												assign node18705 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node18708 = (inp[7]) ? node18712 : node18709;
													assign node18709 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node18712 = (inp[2]) ? node18714 : 4'b0111;
														assign node18714 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node18717 = (inp[7]) ? node18741 : node18718;
											assign node18718 = (inp[8]) ? node18730 : node18719;
												assign node18719 = (inp[6]) ? node18721 : 4'b0110;
													assign node18721 = (inp[1]) ? node18725 : node18722;
														assign node18722 = (inp[2]) ? 4'b0110 : 4'b1110;
														assign node18725 = (inp[11]) ? 4'b0110 : node18726;
															assign node18726 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node18730 = (inp[11]) ? node18732 : 4'b1111;
													assign node18732 = (inp[6]) ? node18738 : node18733;
														assign node18733 = (inp[1]) ? node18735 : 4'b1111;
															assign node18735 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node18738 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node18741 = (inp[14]) ? node18755 : node18742;
												assign node18742 = (inp[6]) ? node18752 : node18743;
													assign node18743 = (inp[11]) ? node18745 : 4'b0111;
														assign node18745 = (inp[1]) ? node18749 : node18746;
															assign node18746 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node18749 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node18752 = (inp[11]) ? 4'b0111 : 4'b1111;
												assign node18755 = (inp[8]) ? 4'b0110 : 4'b0111;
									assign node18758 = (inp[12]) ? node18810 : node18759;
										assign node18759 = (inp[11]) ? node18785 : node18760;
											assign node18760 = (inp[6]) ? node18770 : node18761;
												assign node18761 = (inp[8]) ? node18767 : node18762;
													assign node18762 = (inp[1]) ? 4'b0111 : node18763;
														assign node18763 = (inp[2]) ? 4'b0111 : 4'b1110;
													assign node18767 = (inp[14]) ? 4'b0111 : 4'b0110;
												assign node18770 = (inp[8]) ? node18776 : node18771;
													assign node18771 = (inp[1]) ? 4'b1011 : node18772;
														assign node18772 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node18776 = (inp[14]) ? node18782 : node18777;
														assign node18777 = (inp[1]) ? node18779 : 4'b1011;
															assign node18779 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node18782 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node18785 = (inp[6]) ? node18799 : node18786;
												assign node18786 = (inp[1]) ? node18794 : node18787;
													assign node18787 = (inp[8]) ? 4'b1011 : node18788;
														assign node18788 = (inp[7]) ? 4'b1011 : node18789;
															assign node18789 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node18794 = (inp[7]) ? node18796 : 4'b1011;
														assign node18796 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node18799 = (inp[14]) ? node18807 : node18800;
													assign node18800 = (inp[1]) ? 4'b0011 : node18801;
														assign node18801 = (inp[8]) ? node18803 : 4'b1010;
															assign node18803 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node18807 = (inp[8]) ? 4'b0010 : 4'b1010;
										assign node18810 = (inp[7]) ? node18830 : node18811;
											assign node18811 = (inp[6]) ? node18815 : node18812;
												assign node18812 = (inp[2]) ? 4'b0011 : 4'b1010;
												assign node18815 = (inp[14]) ? node18821 : node18816;
													assign node18816 = (inp[8]) ? 4'b1010 : node18817;
														assign node18817 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node18821 = (inp[8]) ? node18827 : node18822;
														assign node18822 = (inp[11]) ? 4'b0010 : node18823;
															assign node18823 = (inp[1]) ? 4'b1010 : 4'b0010;
														assign node18827 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node18830 = (inp[8]) ? node18850 : node18831;
												assign node18831 = (inp[2]) ? node18839 : node18832;
													assign node18832 = (inp[14]) ? node18834 : 4'b0010;
														assign node18834 = (inp[6]) ? node18836 : 4'b0011;
															assign node18836 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node18839 = (inp[14]) ? node18845 : node18840;
														assign node18840 = (inp[1]) ? 4'b1011 : node18841;
															assign node18841 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node18845 = (inp[11]) ? 4'b0011 : node18846;
															assign node18846 = (inp[6]) ? 4'b1011 : 4'b0011;
												assign node18850 = (inp[2]) ? node18858 : node18851;
													assign node18851 = (inp[14]) ? 4'b1010 : node18852;
														assign node18852 = (inp[6]) ? 4'b0011 : node18853;
															assign node18853 = (inp[11]) ? 4'b1011 : 4'b0011;
													assign node18858 = (inp[1]) ? node18860 : 4'b0010;
														assign node18860 = (inp[14]) ? node18862 : 4'b1010;
															assign node18862 = (inp[6]) ? 4'b0010 : 4'b1010;
						assign node18865 = (inp[5]) ? node19213 : node18866;
							assign node18866 = (inp[4]) ? node19048 : node18867;
								assign node18867 = (inp[9]) ? node18945 : node18868;
									assign node18868 = (inp[12]) ? node18904 : node18869;
										assign node18869 = (inp[11]) ? node18891 : node18870;
											assign node18870 = (inp[6]) ? node18880 : node18871;
												assign node18871 = (inp[1]) ? node18877 : node18872;
													assign node18872 = (inp[7]) ? node18874 : 4'b1100;
														assign node18874 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node18877 = (inp[8]) ? 4'b0101 : 4'b0100;
												assign node18880 = (inp[7]) ? node18888 : node18881;
													assign node18881 = (inp[1]) ? 4'b1001 : node18882;
														assign node18882 = (inp[8]) ? node18884 : 4'b0100;
															assign node18884 = (inp[14]) ? 4'b1001 : 4'b0100;
													assign node18888 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node18891 = (inp[6]) ? node18899 : node18892;
												assign node18892 = (inp[7]) ? node18896 : node18893;
													assign node18893 = (inp[8]) ? 4'b1001 : 4'b0101;
													assign node18896 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node18899 = (inp[8]) ? node18901 : 4'b1000;
													assign node18901 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node18904 = (inp[6]) ? node18922 : node18905;
											assign node18905 = (inp[11]) ? node18915 : node18906;
												assign node18906 = (inp[1]) ? 4'b0001 : node18907;
													assign node18907 = (inp[8]) ? node18909 : 4'b1000;
														assign node18909 = (inp[14]) ? 4'b0001 : node18910;
															assign node18910 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node18915 = (inp[8]) ? node18917 : 4'b1001;
													assign node18917 = (inp[7]) ? node18919 : 4'b0000;
														assign node18919 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node18922 = (inp[11]) ? node18934 : node18923;
												assign node18923 = (inp[8]) ? node18931 : node18924;
													assign node18924 = (inp[1]) ? node18926 : 4'b0000;
														assign node18926 = (inp[7]) ? 4'b1000 : node18927;
															assign node18927 = (inp[14]) ? 4'b1000 : 4'b1000;
													assign node18931 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node18934 = (inp[8]) ? node18936 : 4'b0001;
													assign node18936 = (inp[7]) ? node18940 : node18937;
														assign node18937 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node18940 = (inp[14]) ? 4'b0000 : node18941;
															assign node18941 = (inp[2]) ? 4'b0000 : 4'b0001;
									assign node18945 = (inp[12]) ? node18997 : node18946;
										assign node18946 = (inp[6]) ? node18974 : node18947;
											assign node18947 = (inp[11]) ? node18961 : node18948;
												assign node18948 = (inp[1]) ? node18956 : node18949;
													assign node18949 = (inp[8]) ? node18951 : 4'b1000;
														assign node18951 = (inp[2]) ? node18953 : 4'b1000;
															assign node18953 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node18956 = (inp[7]) ? node18958 : 4'b0001;
														assign node18958 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node18961 = (inp[1]) ? node18967 : node18962;
													assign node18962 = (inp[7]) ? 4'b1110 : node18963;
														assign node18963 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node18967 = (inp[2]) ? 4'b1111 : node18968;
														assign node18968 = (inp[8]) ? 4'b1110 : node18969;
															assign node18969 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node18974 = (inp[11]) ? node18986 : node18975;
												assign node18975 = (inp[1]) ? node18979 : node18976;
													assign node18976 = (inp[14]) ? 4'b1111 : 4'b0001;
													assign node18979 = (inp[14]) ? node18981 : 4'b1110;
														assign node18981 = (inp[7]) ? node18983 : 4'b1111;
															assign node18983 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node18986 = (inp[7]) ? node18988 : 4'b0111;
													assign node18988 = (inp[14]) ? 4'b0110 : node18989;
														assign node18989 = (inp[1]) ? node18993 : node18990;
															assign node18990 = (inp[8]) ? 4'b0111 : 4'b1110;
															assign node18993 = (inp[8]) ? 4'b0110 : 4'b0110;
										assign node18997 = (inp[7]) ? node19021 : node18998;
											assign node18998 = (inp[14]) ? node19010 : node18999;
												assign node18999 = (inp[6]) ? node19005 : node19000;
													assign node19000 = (inp[11]) ? node19002 : 4'b0111;
														assign node19002 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node19005 = (inp[8]) ? node19007 : 4'b0110;
														assign node19007 = (inp[2]) ? 4'b1111 : 4'b0110;
												assign node19010 = (inp[8]) ? node19014 : node19011;
													assign node19011 = (inp[6]) ? 4'b1110 : 4'b0110;
													assign node19014 = (inp[1]) ? node19016 : 4'b1111;
														assign node19016 = (inp[11]) ? 4'b0111 : node19017;
															assign node19017 = (inp[6]) ? 4'b1111 : 4'b0111;
											assign node19021 = (inp[8]) ? node19029 : node19022;
												assign node19022 = (inp[14]) ? 4'b1111 : node19023;
													assign node19023 = (inp[6]) ? 4'b1111 : node19024;
														assign node19024 = (inp[11]) ? 4'b1110 : 4'b0110;
												assign node19029 = (inp[14]) ? node19043 : node19030;
													assign node19030 = (inp[2]) ? node19038 : node19031;
														assign node19031 = (inp[11]) ? node19035 : node19032;
															assign node19032 = (inp[6]) ? 4'b1111 : 4'b0111;
															assign node19035 = (inp[6]) ? 4'b0111 : 4'b1111;
														assign node19038 = (inp[11]) ? node19040 : 4'b1110;
															assign node19040 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node19043 = (inp[11]) ? 4'b0110 : node19044;
														assign node19044 = (inp[6]) ? 4'b1110 : 4'b0110;
								assign node19048 = (inp[9]) ? node19142 : node19049;
									assign node19049 = (inp[12]) ? node19083 : node19050;
										assign node19050 = (inp[11]) ? node19072 : node19051;
											assign node19051 = (inp[6]) ? node19063 : node19052;
												assign node19052 = (inp[2]) ? node19058 : node19053;
													assign node19053 = (inp[1]) ? 4'b0001 : node19054;
														assign node19054 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node19058 = (inp[14]) ? node19060 : 4'b0000;
														assign node19060 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node19063 = (inp[1]) ? node19067 : node19064;
													assign node19064 = (inp[2]) ? 4'b1111 : 4'b0000;
													assign node19067 = (inp[8]) ? 4'b1111 : node19068;
														assign node19068 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node19072 = (inp[6]) ? node19078 : node19073;
												assign node19073 = (inp[2]) ? 4'b1111 : node19074;
													assign node19074 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node19078 = (inp[1]) ? 4'b0111 : node19079;
													assign node19079 = (inp[8]) ? 4'b0111 : 4'b1110;
										assign node19083 = (inp[14]) ? node19117 : node19084;
											assign node19084 = (inp[1]) ? node19104 : node19085;
												assign node19085 = (inp[2]) ? node19095 : node19086;
													assign node19086 = (inp[7]) ? node19088 : 4'b1110;
														assign node19088 = (inp[8]) ? node19092 : node19089;
															assign node19089 = (inp[6]) ? 4'b1110 : 4'b0110;
															assign node19092 = (inp[11]) ? 4'b1111 : 4'b0111;
													assign node19095 = (inp[6]) ? node19097 : 4'b0110;
														assign node19097 = (inp[7]) ? node19101 : node19098;
															assign node19098 = (inp[8]) ? 4'b0111 : 4'b1110;
															assign node19101 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node19104 = (inp[2]) ? node19112 : node19105;
													assign node19105 = (inp[11]) ? node19109 : node19106;
														assign node19106 = (inp[6]) ? 4'b1111 : 4'b0110;
														assign node19109 = (inp[6]) ? 4'b0110 : 4'b1111;
													assign node19112 = (inp[7]) ? node19114 : 4'b1110;
														assign node19114 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node19117 = (inp[2]) ? node19133 : node19118;
												assign node19118 = (inp[6]) ? node19126 : node19119;
													assign node19119 = (inp[11]) ? node19123 : node19120;
														assign node19120 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node19123 = (inp[8]) ? 4'b1110 : 4'b0110;
													assign node19126 = (inp[11]) ? node19128 : 4'b1110;
														assign node19128 = (inp[7]) ? 4'b0110 : node19129;
															assign node19129 = (inp[1]) ? 4'b0110 : 4'b1110;
												assign node19133 = (inp[11]) ? node19135 : 4'b0111;
													assign node19135 = (inp[6]) ? node19139 : node19136;
														assign node19136 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node19139 = (inp[8]) ? 4'b0111 : 4'b0110;
									assign node19142 = (inp[6]) ? node19178 : node19143;
										assign node19143 = (inp[11]) ? node19163 : node19144;
											assign node19144 = (inp[12]) ? node19156 : node19145;
												assign node19145 = (inp[1]) ? node19151 : node19146;
													assign node19146 = (inp[8]) ? 4'b0111 : node19147;
														assign node19147 = (inp[7]) ? 4'b0111 : 4'b1110;
													assign node19151 = (inp[7]) ? 4'b0110 : node19152;
														assign node19152 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node19156 = (inp[7]) ? node19160 : node19157;
													assign node19157 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node19160 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node19163 = (inp[7]) ? node19171 : node19164;
												assign node19164 = (inp[8]) ? 4'b1011 : node19165;
													assign node19165 = (inp[12]) ? node19167 : 4'b0111;
														assign node19167 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node19171 = (inp[8]) ? 4'b1010 : node19172;
													assign node19172 = (inp[14]) ? 4'b1011 : node19173;
														assign node19173 = (inp[2]) ? 4'b1011 : 4'b1010;
										assign node19178 = (inp[11]) ? node19194 : node19179;
											assign node19179 = (inp[14]) ? node19187 : node19180;
												assign node19180 = (inp[12]) ? node19182 : 4'b1011;
													assign node19182 = (inp[8]) ? node19184 : 4'b0010;
														assign node19184 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node19187 = (inp[1]) ? 4'b1010 : node19188;
													assign node19188 = (inp[8]) ? node19190 : 4'b1011;
														assign node19190 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node19194 = (inp[8]) ? node19206 : node19195;
												assign node19195 = (inp[1]) ? node19203 : node19196;
													assign node19196 = (inp[2]) ? 4'b1010 : node19197;
														assign node19197 = (inp[14]) ? 4'b0011 : node19198;
															assign node19198 = (inp[12]) ? 4'b1010 : 4'b1011;
													assign node19203 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node19206 = (inp[7]) ? 4'b0010 : node19207;
													assign node19207 = (inp[2]) ? 4'b0011 : node19208;
														assign node19208 = (inp[14]) ? 4'b0011 : 4'b0010;
							assign node19213 = (inp[2]) ? node19429 : node19214;
								assign node19214 = (inp[8]) ? node19310 : node19215;
									assign node19215 = (inp[9]) ? node19273 : node19216;
										assign node19216 = (inp[4]) ? node19240 : node19217;
											assign node19217 = (inp[7]) ? node19233 : node19218;
												assign node19218 = (inp[14]) ? node19230 : node19219;
													assign node19219 = (inp[12]) ? node19225 : node19220;
														assign node19220 = (inp[11]) ? node19222 : 4'b0111;
															assign node19222 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node19225 = (inp[6]) ? 4'b0011 : node19226;
															assign node19226 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node19230 = (inp[6]) ? 4'b1010 : 4'b0110;
												assign node19233 = (inp[14]) ? node19237 : node19234;
													assign node19234 = (inp[12]) ? 4'b0010 : 4'b1010;
													assign node19237 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node19240 = (inp[6]) ? node19260 : node19241;
												assign node19241 = (inp[12]) ? node19253 : node19242;
													assign node19242 = (inp[7]) ? node19250 : node19243;
														assign node19243 = (inp[14]) ? node19247 : node19244;
															assign node19244 = (inp[11]) ? 4'b1111 : 4'b0011;
															assign node19247 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node19250 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node19253 = (inp[7]) ? 4'b0110 : node19254;
														assign node19254 = (inp[11]) ? node19256 : 4'b0110;
															assign node19256 = (inp[1]) ? 4'b1111 : 4'b0111;
												assign node19260 = (inp[11]) ? node19266 : node19261;
													assign node19261 = (inp[7]) ? node19263 : 4'b0110;
														assign node19263 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node19266 = (inp[14]) ? node19270 : node19267;
														assign node19267 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node19270 = (inp[7]) ? 4'b0111 : 4'b1110;
										assign node19273 = (inp[4]) ? node19297 : node19274;
											assign node19274 = (inp[1]) ? node19286 : node19275;
												assign node19275 = (inp[12]) ? node19283 : node19276;
													assign node19276 = (inp[14]) ? node19280 : node19277;
														assign node19277 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node19280 = (inp[7]) ? 4'b1111 : 4'b0010;
													assign node19283 = (inp[11]) ? 4'b0111 : 4'b1111;
												assign node19286 = (inp[14]) ? node19290 : node19287;
													assign node19287 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node19290 = (inp[6]) ? node19294 : node19291;
														assign node19291 = (inp[12]) ? 4'b0111 : 4'b1111;
														assign node19294 = (inp[11]) ? 4'b0110 : 4'b1110;
											assign node19297 = (inp[14]) ? node19303 : node19298;
												assign node19298 = (inp[7]) ? node19300 : 4'b1011;
													assign node19300 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node19303 = (inp[7]) ? node19305 : 4'b1010;
													assign node19305 = (inp[12]) ? 4'b1011 : node19306;
														assign node19306 = (inp[6]) ? 4'b1011 : 4'b0111;
									assign node19310 = (inp[7]) ? node19374 : node19311;
										assign node19311 = (inp[14]) ? node19349 : node19312;
											assign node19312 = (inp[12]) ? node19332 : node19313;
												assign node19313 = (inp[9]) ? node19323 : node19314;
													assign node19314 = (inp[6]) ? node19318 : node19315;
														assign node19315 = (inp[1]) ? 4'b1010 : 4'b0110;
														assign node19318 = (inp[11]) ? node19320 : 4'b0010;
															assign node19320 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node19323 = (inp[4]) ? node19329 : node19324;
														assign node19324 = (inp[11]) ? 4'b1110 : node19325;
															assign node19325 = (inp[1]) ? 4'b1110 : 4'b0010;
														assign node19329 = (inp[1]) ? 4'b0010 : 4'b1010;
												assign node19332 = (inp[11]) ? node19340 : node19333;
													assign node19333 = (inp[4]) ? node19337 : node19334;
														assign node19334 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node19337 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node19340 = (inp[1]) ? node19346 : node19341;
														assign node19341 = (inp[9]) ? 4'b0010 : node19342;
															assign node19342 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node19346 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node19349 = (inp[6]) ? node19363 : node19350;
												assign node19350 = (inp[11]) ? node19356 : node19351;
													assign node19351 = (inp[9]) ? 4'b0111 : node19352;
														assign node19352 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node19356 = (inp[12]) ? node19358 : 4'b1111;
														assign node19358 = (inp[1]) ? 4'b1011 : node19359;
															assign node19359 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node19363 = (inp[1]) ? node19369 : node19364;
													assign node19364 = (inp[9]) ? node19366 : 4'b1111;
														assign node19366 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node19369 = (inp[12]) ? node19371 : 4'b1011;
														assign node19371 = (inp[4]) ? 4'b1111 : 4'b1011;
										assign node19374 = (inp[14]) ? node19394 : node19375;
											assign node19375 = (inp[4]) ? node19383 : node19376;
												assign node19376 = (inp[12]) ? 4'b0111 : node19377;
													assign node19377 = (inp[9]) ? 4'b1111 : node19378;
														assign node19378 = (inp[1]) ? 4'b1011 : 4'b0111;
												assign node19383 = (inp[12]) ? node19391 : node19384;
													assign node19384 = (inp[9]) ? node19386 : 4'b0011;
														assign node19386 = (inp[6]) ? node19388 : 4'b1011;
															assign node19388 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node19391 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node19394 = (inp[9]) ? node19408 : node19395;
												assign node19395 = (inp[4]) ? node19399 : node19396;
													assign node19396 = (inp[12]) ? 4'b0010 : 4'b1010;
													assign node19399 = (inp[12]) ? 4'b1110 : node19400;
														assign node19400 = (inp[1]) ? node19404 : node19401;
															assign node19401 = (inp[6]) ? 4'b1110 : 4'b0010;
															assign node19404 = (inp[6]) ? 4'b0110 : 4'b1110;
												assign node19408 = (inp[4]) ? node19418 : node19409;
													assign node19409 = (inp[1]) ? node19415 : node19410;
														assign node19410 = (inp[11]) ? node19412 : 4'b1110;
															assign node19412 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node19415 = (inp[11]) ? 4'b1110 : 4'b0010;
													assign node19418 = (inp[1]) ? node19424 : node19419;
														assign node19419 = (inp[6]) ? 4'b0010 : node19420;
															assign node19420 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node19424 = (inp[11]) ? node19426 : 4'b1010;
															assign node19426 = (inp[12]) ? 4'b1010 : 4'b0010;
								assign node19429 = (inp[9]) ? node19515 : node19430;
									assign node19430 = (inp[4]) ? node19476 : node19431;
										assign node19431 = (inp[6]) ? node19461 : node19432;
											assign node19432 = (inp[11]) ? node19448 : node19433;
												assign node19433 = (inp[12]) ? node19441 : node19434;
													assign node19434 = (inp[1]) ? node19436 : 4'b0111;
														assign node19436 = (inp[14]) ? node19438 : 4'b0110;
															assign node19438 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node19441 = (inp[14]) ? node19445 : node19442;
														assign node19442 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node19445 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node19448 = (inp[1]) ? node19454 : node19449;
													assign node19449 = (inp[8]) ? node19451 : 4'b0110;
														assign node19451 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node19454 = (inp[14]) ? node19456 : 4'b1010;
														assign node19456 = (inp[8]) ? 4'b1011 : node19457;
															assign node19457 = (inp[7]) ? 4'b1011 : 4'b1010;
											assign node19461 = (inp[11]) ? node19471 : node19462;
												assign node19462 = (inp[14]) ? 4'b1011 : node19463;
													assign node19463 = (inp[7]) ? node19467 : node19464;
														assign node19464 = (inp[8]) ? 4'b1011 : 4'b0010;
														assign node19467 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node19471 = (inp[12]) ? 4'b0010 : node19472;
													assign node19472 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node19476 = (inp[6]) ? node19494 : node19477;
											assign node19477 = (inp[11]) ? node19487 : node19478;
												assign node19478 = (inp[12]) ? 4'b0110 : node19479;
													assign node19479 = (inp[8]) ? node19483 : node19480;
														assign node19480 = (inp[7]) ? 4'b0011 : 4'b1010;
														assign node19483 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node19487 = (inp[14]) ? node19489 : 4'b1110;
													assign node19489 = (inp[7]) ? node19491 : 4'b1111;
														assign node19491 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node19494 = (inp[11]) ? node19502 : node19495;
												assign node19495 = (inp[8]) ? node19499 : node19496;
													assign node19496 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node19499 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node19502 = (inp[1]) ? node19508 : node19503;
													assign node19503 = (inp[14]) ? node19505 : 4'b0111;
														assign node19505 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node19508 = (inp[8]) ? node19512 : node19509;
														assign node19509 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node19512 = (inp[7]) ? 4'b0110 : 4'b0111;
									assign node19515 = (inp[4]) ? node19565 : node19516;
										assign node19516 = (inp[14]) ? node19548 : node19517;
											assign node19517 = (inp[1]) ? node19533 : node19518;
												assign node19518 = (inp[6]) ? node19522 : node19519;
													assign node19519 = (inp[11]) ? 4'b1111 : 4'b0111;
													assign node19522 = (inp[11]) ? node19528 : node19523;
														assign node19523 = (inp[8]) ? node19525 : 4'b0110;
															assign node19525 = (inp[12]) ? 4'b1110 : 4'b1111;
														assign node19528 = (inp[8]) ? node19530 : 4'b0111;
															assign node19530 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node19533 = (inp[11]) ? node19541 : node19534;
													assign node19534 = (inp[6]) ? 4'b1111 : node19535;
														assign node19535 = (inp[12]) ? 4'b0110 : node19536;
															assign node19536 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node19541 = (inp[6]) ? node19543 : 4'b1110;
														assign node19543 = (inp[8]) ? 4'b0110 : node19544;
															assign node19544 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node19548 = (inp[11]) ? node19562 : node19549;
												assign node19549 = (inp[6]) ? node19557 : node19550;
													assign node19550 = (inp[12]) ? node19552 : 4'b0011;
														assign node19552 = (inp[7]) ? node19554 : 4'b0111;
															assign node19554 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node19557 = (inp[1]) ? 4'b1111 : node19558;
														assign node19558 = (inp[12]) ? 4'b0110 : 4'b1111;
												assign node19562 = (inp[6]) ? 4'b0111 : 4'b1111;
										assign node19565 = (inp[12]) ? node19585 : node19566;
											assign node19566 = (inp[6]) ? node19574 : node19567;
												assign node19567 = (inp[11]) ? 4'b1010 : node19568;
													assign node19568 = (inp[8]) ? node19570 : 4'b0111;
														assign node19570 = (inp[14]) ? 4'b0111 : 4'b0110;
												assign node19574 = (inp[1]) ? node19580 : node19575;
													assign node19575 = (inp[11]) ? node19577 : 4'b0110;
														assign node19577 = (inp[7]) ? 4'b0010 : 4'b1010;
													assign node19580 = (inp[11]) ? 4'b0011 : node19581;
														assign node19581 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node19585 = (inp[7]) ? node19599 : node19586;
												assign node19586 = (inp[8]) ? node19588 : 4'b1010;
													assign node19588 = (inp[1]) ? node19594 : node19589;
														assign node19589 = (inp[11]) ? 4'b0011 : node19590;
															assign node19590 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node19594 = (inp[11]) ? node19596 : 4'b0011;
															assign node19596 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node19599 = (inp[8]) ? node19603 : node19600;
													assign node19600 = (inp[11]) ? 4'b1011 : 4'b0011;
													assign node19603 = (inp[11]) ? 4'b0010 : node19604;
														assign node19604 = (inp[14]) ? 4'b1010 : 4'b0010;
				assign node19608 = (inp[0]) ? node21030 : node19609;
					assign node19609 = (inp[5]) ? node20283 : node19610;
						assign node19610 = (inp[3]) ? node19912 : node19611;
							assign node19611 = (inp[6]) ? node19765 : node19612;
								assign node19612 = (inp[11]) ? node19686 : node19613;
									assign node19613 = (inp[1]) ? node19649 : node19614;
										assign node19614 = (inp[8]) ? node19634 : node19615;
											assign node19615 = (inp[7]) ? node19629 : node19616;
												assign node19616 = (inp[12]) ? node19624 : node19617;
													assign node19617 = (inp[2]) ? 4'b1000 : node19618;
														assign node19618 = (inp[4]) ? node19620 : 4'b1001;
															assign node19620 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node19624 = (inp[4]) ? 4'b1000 : node19625;
														assign node19625 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node19629 = (inp[14]) ? node19631 : 4'b1100;
													assign node19631 = (inp[2]) ? 4'b0101 : 4'b0001;
											assign node19634 = (inp[12]) ? 4'b0101 : node19635;
												assign node19635 = (inp[4]) ? node19643 : node19636;
													assign node19636 = (inp[9]) ? node19640 : node19637;
														assign node19637 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node19640 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node19643 = (inp[2]) ? 4'b0100 : node19644;
														assign node19644 = (inp[9]) ? 4'b1100 : 4'b1000;
										assign node19649 = (inp[14]) ? node19667 : node19650;
											assign node19650 = (inp[2]) ? node19662 : node19651;
												assign node19651 = (inp[9]) ? node19659 : node19652;
													assign node19652 = (inp[12]) ? 4'b0100 : node19653;
														assign node19653 = (inp[4]) ? 4'b0001 : node19654;
															assign node19654 = (inp[7]) ? 4'b0100 : 4'b0100;
													assign node19659 = (inp[7]) ? 4'b0100 : 4'b0001;
												assign node19662 = (inp[9]) ? node19664 : 4'b0000;
													assign node19664 = (inp[8]) ? 4'b0100 : 4'b0000;
											assign node19667 = (inp[7]) ? node19677 : node19668;
												assign node19668 = (inp[8]) ? 4'b0101 : node19669;
													assign node19669 = (inp[9]) ? node19671 : 4'b0000;
														assign node19671 = (inp[2]) ? node19673 : 4'b0100;
															assign node19673 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node19677 = (inp[8]) ? 4'b0000 : node19678;
													assign node19678 = (inp[9]) ? node19680 : 4'b0101;
														assign node19680 = (inp[2]) ? 4'b0101 : node19681;
															assign node19681 = (inp[12]) ? 4'b0001 : 4'b0001;
									assign node19686 = (inp[7]) ? node19720 : node19687;
										assign node19687 = (inp[8]) ? node19705 : node19688;
											assign node19688 = (inp[1]) ? node19694 : node19689;
												assign node19689 = (inp[2]) ? 4'b0100 : node19690;
													assign node19690 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node19694 = (inp[14]) ? node19700 : node19695;
													assign node19695 = (inp[4]) ? 4'b1101 : node19696;
														assign node19696 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node19700 = (inp[12]) ? 4'b1100 : node19701;
														assign node19701 = (inp[9]) ? 4'b1100 : 4'b1000;
											assign node19705 = (inp[2]) ? node19713 : node19706;
												assign node19706 = (inp[14]) ? node19708 : 4'b0000;
													assign node19708 = (inp[9]) ? node19710 : 4'b1001;
														assign node19710 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node19713 = (inp[4]) ? node19717 : node19714;
													assign node19714 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node19717 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node19720 = (inp[8]) ? node19742 : node19721;
											assign node19721 = (inp[12]) ? node19735 : node19722;
												assign node19722 = (inp[1]) ? node19730 : node19723;
													assign node19723 = (inp[14]) ? node19725 : 4'b1101;
														assign node19725 = (inp[4]) ? node19727 : 4'b1001;
															assign node19727 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node19730 = (inp[9]) ? 4'b1001 : node19731;
														assign node19731 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node19735 = (inp[9]) ? node19739 : node19736;
													assign node19736 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node19739 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node19742 = (inp[2]) ? node19752 : node19743;
												assign node19743 = (inp[14]) ? node19745 : 4'b1101;
													assign node19745 = (inp[1]) ? node19747 : 4'b1000;
														assign node19747 = (inp[12]) ? 4'b1100 : node19748;
															assign node19748 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node19752 = (inp[14]) ? node19758 : node19753;
													assign node19753 = (inp[4]) ? node19755 : 4'b1000;
														assign node19755 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node19758 = (inp[1]) ? node19760 : 4'b1000;
														assign node19760 = (inp[4]) ? 4'b1100 : node19761;
															assign node19761 = (inp[9]) ? 4'b1100 : 4'b1000;
								assign node19765 = (inp[11]) ? node19829 : node19766;
									assign node19766 = (inp[1]) ? node19796 : node19767;
										assign node19767 = (inp[8]) ? node19785 : node19768;
											assign node19768 = (inp[7]) ? node19776 : node19769;
												assign node19769 = (inp[14]) ? 4'b0000 : node19770;
													assign node19770 = (inp[2]) ? 4'b0100 : node19771;
														assign node19771 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node19776 = (inp[2]) ? node19782 : node19777;
													assign node19777 = (inp[14]) ? 4'b1101 : node19778;
														assign node19778 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node19782 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node19785 = (inp[7]) ? node19791 : node19786;
												assign node19786 = (inp[9]) ? 4'b1101 : node19787;
													assign node19787 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node19791 = (inp[4]) ? 4'b1000 : node19792;
													assign node19792 = (inp[9]) ? 4'b1101 : 4'b1000;
										assign node19796 = (inp[4]) ? node19812 : node19797;
											assign node19797 = (inp[9]) ? node19807 : node19798;
												assign node19798 = (inp[2]) ? node19800 : 4'b1000;
													assign node19800 = (inp[14]) ? node19802 : 4'b1000;
														assign node19802 = (inp[12]) ? 4'b1001 : node19803;
															assign node19803 = (inp[7]) ? 4'b1000 : 4'b1000;
												assign node19807 = (inp[2]) ? 4'b1100 : node19808;
													assign node19808 = (inp[8]) ? 4'b1101 : 4'b1100;
											assign node19812 = (inp[9]) ? node19818 : node19813;
												assign node19813 = (inp[8]) ? 4'b1101 : node19814;
													assign node19814 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node19818 = (inp[14]) ? node19824 : node19819;
													assign node19819 = (inp[12]) ? node19821 : 4'b1001;
														assign node19821 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node19824 = (inp[2]) ? 4'b1000 : node19825;
														assign node19825 = (inp[12]) ? 4'b1000 : 4'b1001;
									assign node19829 = (inp[1]) ? node19873 : node19830;
										assign node19830 = (inp[8]) ? node19856 : node19831;
											assign node19831 = (inp[7]) ? node19843 : node19832;
												assign node19832 = (inp[2]) ? node19838 : node19833;
													assign node19833 = (inp[14]) ? 4'b1100 : node19834;
														assign node19834 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node19838 = (inp[9]) ? node19840 : 4'b1000;
														assign node19840 = (inp[14]) ? 4'b1000 : 4'b1100;
												assign node19843 = (inp[2]) ? node19849 : node19844;
													assign node19844 = (inp[14]) ? 4'b0101 : node19845;
														assign node19845 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node19849 = (inp[12]) ? node19851 : 4'b0001;
														assign node19851 = (inp[4]) ? node19853 : 4'b0101;
															assign node19853 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node19856 = (inp[7]) ? node19870 : node19857;
												assign node19857 = (inp[2]) ? node19863 : node19858;
													assign node19858 = (inp[14]) ? 4'b0101 : node19859;
														assign node19859 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node19863 = (inp[4]) ? node19867 : node19864;
														assign node19864 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node19867 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node19870 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node19873 = (inp[9]) ? node19895 : node19874;
											assign node19874 = (inp[4]) ? node19884 : node19875;
												assign node19875 = (inp[12]) ? node19877 : 4'b0001;
													assign node19877 = (inp[7]) ? 4'b0000 : node19878;
														assign node19878 = (inp[8]) ? 4'b0000 : node19879;
															assign node19879 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node19884 = (inp[14]) ? node19886 : 4'b0100;
													assign node19886 = (inp[2]) ? 4'b0100 : node19887;
														assign node19887 = (inp[7]) ? node19891 : node19888;
															assign node19888 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node19891 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node19895 = (inp[4]) ? node19907 : node19896;
												assign node19896 = (inp[8]) ? 4'b0101 : node19897;
													assign node19897 = (inp[2]) ? 4'b0101 : node19898;
														assign node19898 = (inp[14]) ? node19902 : node19899;
															assign node19899 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node19902 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node19907 = (inp[14]) ? node19909 : 4'b0001;
													assign node19909 = (inp[2]) ? 4'b0000 : 4'b0001;
							assign node19912 = (inp[9]) ? node20078 : node19913;
								assign node19913 = (inp[4]) ? node19997 : node19914;
									assign node19914 = (inp[12]) ? node19944 : node19915;
										assign node19915 = (inp[1]) ? node19931 : node19916;
											assign node19916 = (inp[2]) ? node19922 : node19917;
												assign node19917 = (inp[11]) ? node19919 : 4'b0101;
													assign node19919 = (inp[6]) ? 4'b0001 : 4'b0100;
												assign node19922 = (inp[8]) ? node19928 : node19923;
													assign node19923 = (inp[6]) ? 4'b0100 : node19924;
														assign node19924 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node19928 = (inp[7]) ? 4'b1000 : 4'b0001;
											assign node19931 = (inp[11]) ? node19935 : node19932;
												assign node19932 = (inp[6]) ? 4'b1001 : 4'b0101;
												assign node19935 = (inp[6]) ? node19941 : node19936;
													assign node19936 = (inp[7]) ? node19938 : 4'b1000;
														assign node19938 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node19941 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node19944 = (inp[1]) ? node19968 : node19945;
											assign node19945 = (inp[8]) ? node19961 : node19946;
												assign node19946 = (inp[7]) ? node19956 : node19947;
													assign node19947 = (inp[2]) ? node19951 : node19948;
														assign node19948 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node19951 = (inp[14]) ? 4'b1000 : node19952;
															assign node19952 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node19956 = (inp[6]) ? node19958 : 4'b0001;
														assign node19958 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node19961 = (inp[11]) ? node19965 : node19962;
													assign node19962 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node19965 = (inp[6]) ? 4'b0001 : 4'b1001;
											assign node19968 = (inp[11]) ? node19980 : node19969;
												assign node19969 = (inp[6]) ? node19973 : node19970;
													assign node19970 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node19973 = (inp[2]) ? 4'b1000 : node19974;
														assign node19974 = (inp[14]) ? 4'b1001 : node19975;
															assign node19975 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node19980 = (inp[6]) ? node19984 : node19981;
													assign node19981 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node19984 = (inp[8]) ? node19990 : node19985;
														assign node19985 = (inp[7]) ? node19987 : 4'b0000;
															assign node19987 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node19990 = (inp[14]) ? node19994 : node19991;
															assign node19991 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node19994 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node19997 = (inp[12]) ? node20045 : node19998;
										assign node19998 = (inp[6]) ? node20028 : node19999;
											assign node19999 = (inp[11]) ? node20017 : node20000;
												assign node20000 = (inp[1]) ? node20008 : node20001;
													assign node20001 = (inp[8]) ? node20003 : 4'b1000;
														assign node20003 = (inp[2]) ? 4'b0001 : node20004;
															assign node20004 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node20008 = (inp[7]) ? node20010 : 4'b0000;
														assign node20010 = (inp[8]) ? node20014 : node20011;
															assign node20011 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node20014 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node20017 = (inp[8]) ? node20019 : 4'b0000;
													assign node20019 = (inp[14]) ? node20025 : node20020;
														assign node20020 = (inp[7]) ? 4'b1111 : node20021;
															assign node20021 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node20025 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node20028 = (inp[14]) ? 4'b1110 : node20029;
												assign node20029 = (inp[11]) ? node20037 : node20030;
													assign node20030 = (inp[1]) ? node20032 : 4'b0000;
														assign node20032 = (inp[8]) ? node20034 : 4'b1111;
															assign node20034 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node20037 = (inp[1]) ? node20039 : 4'b1111;
														assign node20039 = (inp[8]) ? 4'b0110 : node20040;
															assign node20040 = (inp[2]) ? 4'b0111 : 4'b0110;
										assign node20045 = (inp[2]) ? node20065 : node20046;
											assign node20046 = (inp[11]) ? node20054 : node20047;
												assign node20047 = (inp[6]) ? 4'b1111 : node20048;
													assign node20048 = (inp[8]) ? node20050 : 4'b1110;
														assign node20050 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node20054 = (inp[14]) ? 4'b0111 : node20055;
													assign node20055 = (inp[6]) ? node20059 : node20056;
														assign node20056 = (inp[1]) ? 4'b1110 : 4'b0110;
														assign node20059 = (inp[8]) ? 4'b0110 : node20060;
															assign node20060 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node20065 = (inp[11]) ? node20071 : node20066;
												assign node20066 = (inp[7]) ? node20068 : 4'b0110;
													assign node20068 = (inp[6]) ? 4'b1111 : 4'b0111;
												assign node20071 = (inp[7]) ? node20075 : node20072;
													assign node20072 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node20075 = (inp[8]) ? 4'b1110 : 4'b1111;
								assign node20078 = (inp[4]) ? node20180 : node20079;
									assign node20079 = (inp[12]) ? node20123 : node20080;
										assign node20080 = (inp[14]) ? node20104 : node20081;
											assign node20081 = (inp[11]) ? node20091 : node20082;
												assign node20082 = (inp[7]) ? node20088 : node20083;
													assign node20083 = (inp[6]) ? 4'b0000 : node20084;
														assign node20084 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node20088 = (inp[6]) ? 4'b0000 : 4'b0001;
												assign node20091 = (inp[6]) ? node20095 : node20092;
													assign node20092 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node20095 = (inp[2]) ? 4'b0110 : node20096;
														assign node20096 = (inp[7]) ? node20100 : node20097;
															assign node20097 = (inp[8]) ? 4'b1110 : 4'b0111;
															assign node20100 = (inp[8]) ? 4'b0111 : 4'b0110;
											assign node20104 = (inp[11]) ? node20108 : node20105;
												assign node20105 = (inp[6]) ? 4'b1111 : 4'b0001;
												assign node20108 = (inp[6]) ? node20114 : node20109;
													assign node20109 = (inp[2]) ? node20111 : 4'b1111;
														assign node20111 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node20114 = (inp[2]) ? node20118 : node20115;
														assign node20115 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node20118 = (inp[7]) ? 4'b0110 : node20119;
															assign node20119 = (inp[8]) ? 4'b0111 : 4'b0110;
										assign node20123 = (inp[11]) ? node20151 : node20124;
											assign node20124 = (inp[8]) ? node20136 : node20125;
												assign node20125 = (inp[1]) ? 4'b1111 : node20126;
													assign node20126 = (inp[6]) ? node20132 : node20127;
														assign node20127 = (inp[14]) ? 4'b0111 : node20128;
															assign node20128 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node20132 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node20136 = (inp[6]) ? node20146 : node20137;
													assign node20137 = (inp[1]) ? node20141 : node20138;
														assign node20138 = (inp[7]) ? 4'b0111 : 4'b1110;
														assign node20141 = (inp[7]) ? 4'b0110 : node20142;
															assign node20142 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node20146 = (inp[2]) ? 4'b1110 : node20147;
														assign node20147 = (inp[14]) ? 4'b1111 : 4'b0110;
											assign node20151 = (inp[2]) ? node20167 : node20152;
												assign node20152 = (inp[6]) ? node20160 : node20153;
													assign node20153 = (inp[1]) ? 4'b1110 : node20154;
														assign node20154 = (inp[14]) ? 4'b0110 : node20155;
															assign node20155 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node20160 = (inp[1]) ? 4'b0110 : node20161;
														assign node20161 = (inp[8]) ? node20163 : 4'b1110;
															assign node20163 = (inp[14]) ? 4'b0110 : 4'b1110;
												assign node20167 = (inp[14]) ? node20171 : node20168;
													assign node20168 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node20171 = (inp[1]) ? 4'b1110 : node20172;
														assign node20172 = (inp[8]) ? node20176 : node20173;
															assign node20173 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node20176 = (inp[7]) ? 4'b1110 : 4'b1111;
									assign node20180 = (inp[12]) ? node20232 : node20181;
										assign node20181 = (inp[6]) ? node20209 : node20182;
											assign node20182 = (inp[11]) ? node20194 : node20183;
												assign node20183 = (inp[8]) ? node20189 : node20184;
													assign node20184 = (inp[14]) ? 4'b0111 : node20185;
														assign node20185 = (inp[2]) ? 4'b1110 : 4'b0110;
													assign node20189 = (inp[14]) ? node20191 : 4'b0111;
														assign node20191 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node20194 = (inp[1]) ? node20204 : node20195;
													assign node20195 = (inp[7]) ? node20201 : node20196;
														assign node20196 = (inp[8]) ? node20198 : 4'b0110;
															assign node20198 = (inp[14]) ? 4'b1011 : 4'b0110;
														assign node20201 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node20204 = (inp[14]) ? node20206 : 4'b1011;
														assign node20206 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node20209 = (inp[11]) ? node20221 : node20210;
												assign node20210 = (inp[7]) ? node20214 : node20211;
													assign node20211 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node20214 = (inp[2]) ? 4'b1010 : node20215;
														assign node20215 = (inp[8]) ? node20217 : 4'b1010;
															assign node20217 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node20221 = (inp[8]) ? node20227 : node20222;
													assign node20222 = (inp[2]) ? 4'b0010 : node20223;
														assign node20223 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node20227 = (inp[7]) ? node20229 : 4'b0011;
														assign node20229 = (inp[1]) ? 4'b0011 : 4'b0010;
										assign node20232 = (inp[2]) ? node20250 : node20233;
											assign node20233 = (inp[14]) ? node20243 : node20234;
												assign node20234 = (inp[6]) ? node20240 : node20235;
													assign node20235 = (inp[1]) ? node20237 : 4'b0011;
														assign node20237 = (inp[11]) ? 4'b1011 : 4'b0011;
													assign node20240 = (inp[1]) ? 4'b0010 : 4'b1010;
												assign node20243 = (inp[1]) ? 4'b1010 : node20244;
													assign node20244 = (inp[6]) ? node20246 : 4'b0010;
														assign node20246 = (inp[11]) ? 4'b1010 : 4'b0010;
											assign node20250 = (inp[14]) ? node20266 : node20251;
												assign node20251 = (inp[8]) ? node20259 : node20252;
													assign node20252 = (inp[7]) ? node20256 : node20253;
														assign node20253 = (inp[6]) ? 4'b0010 : 4'b1010;
														assign node20256 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node20259 = (inp[7]) ? node20261 : 4'b1011;
														assign node20261 = (inp[6]) ? 4'b1010 : node20262;
															assign node20262 = (inp[11]) ? 4'b1010 : 4'b0010;
												assign node20266 = (inp[6]) ? node20278 : node20267;
													assign node20267 = (inp[11]) ? node20273 : node20268;
														assign node20268 = (inp[7]) ? node20270 : 4'b0011;
															assign node20270 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node20273 = (inp[7]) ? 4'b1011 : node20274;
															assign node20274 = (inp[8]) ? 4'b1011 : 4'b0010;
													assign node20278 = (inp[7]) ? node20280 : 4'b0011;
														assign node20280 = (inp[8]) ? 4'b0010 : 4'b0011;
						assign node20283 = (inp[3]) ? node20647 : node20284;
							assign node20284 = (inp[9]) ? node20468 : node20285;
								assign node20285 = (inp[4]) ? node20377 : node20286;
									assign node20286 = (inp[12]) ? node20326 : node20287;
										assign node20287 = (inp[6]) ? node20303 : node20288;
											assign node20288 = (inp[11]) ? node20296 : node20289;
												assign node20289 = (inp[7]) ? node20293 : node20290;
													assign node20290 = (inp[8]) ? 4'b0101 : 4'b1100;
													assign node20293 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node20296 = (inp[1]) ? node20300 : node20297;
													assign node20297 = (inp[7]) ? 4'b1000 : 4'b0100;
													assign node20300 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node20303 = (inp[11]) ? node20317 : node20304;
												assign node20304 = (inp[1]) ? 4'b1000 : node20305;
													assign node20305 = (inp[2]) ? node20311 : node20306;
														assign node20306 = (inp[7]) ? node20308 : 4'b0100;
															assign node20308 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node20311 = (inp[7]) ? node20313 : 4'b1001;
															assign node20313 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node20317 = (inp[14]) ? node20321 : node20318;
													assign node20318 = (inp[8]) ? 4'b0001 : 4'b1000;
													assign node20321 = (inp[8]) ? 4'b0000 : node20322;
														assign node20322 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node20326 = (inp[8]) ? node20356 : node20327;
											assign node20327 = (inp[6]) ? node20343 : node20328;
												assign node20328 = (inp[11]) ? node20334 : node20329;
													assign node20329 = (inp[7]) ? node20331 : 4'b0000;
														assign node20331 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node20334 = (inp[14]) ? node20340 : node20335;
														assign node20335 = (inp[7]) ? node20337 : 4'b1001;
															assign node20337 = (inp[2]) ? 4'b1001 : 4'b0000;
														assign node20340 = (inp[2]) ? 4'b0000 : 4'b1000;
												assign node20343 = (inp[11]) ? node20351 : node20344;
													assign node20344 = (inp[14]) ? node20348 : node20345;
														assign node20345 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node20348 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node20351 = (inp[1]) ? 4'b0001 : node20352;
														assign node20352 = (inp[14]) ? 4'b0001 : 4'b1000;
											assign node20356 = (inp[2]) ? node20370 : node20357;
												assign node20357 = (inp[1]) ? node20365 : node20358;
													assign node20358 = (inp[6]) ? node20360 : 4'b0001;
														assign node20360 = (inp[11]) ? node20362 : 4'b1000;
															assign node20362 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node20365 = (inp[14]) ? 4'b0001 : node20366;
														assign node20366 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node20370 = (inp[7]) ? node20372 : 4'b1001;
													assign node20372 = (inp[1]) ? node20374 : 4'b1000;
														assign node20374 = (inp[6]) ? 4'b0000 : 4'b1000;
									assign node20377 = (inp[12]) ? node20421 : node20378;
										assign node20378 = (inp[6]) ? node20396 : node20379;
											assign node20379 = (inp[11]) ? node20389 : node20380;
												assign node20380 = (inp[8]) ? node20384 : node20381;
													assign node20381 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node20384 = (inp[2]) ? node20386 : 4'b0001;
														assign node20386 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node20389 = (inp[7]) ? node20393 : node20390;
													assign node20390 = (inp[8]) ? 4'b1111 : 4'b0000;
													assign node20393 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node20396 = (inp[11]) ? node20410 : node20397;
												assign node20397 = (inp[8]) ? node20403 : node20398;
													assign node20398 = (inp[2]) ? node20400 : 4'b0000;
														assign node20400 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node20403 = (inp[7]) ? node20405 : 4'b1111;
														assign node20405 = (inp[2]) ? 4'b1110 : node20406;
															assign node20406 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node20410 = (inp[1]) ? node20414 : node20411;
													assign node20411 = (inp[7]) ? 4'b0111 : 4'b1110;
													assign node20414 = (inp[7]) ? node20416 : 4'b0111;
														assign node20416 = (inp[14]) ? 4'b0111 : node20417;
															assign node20417 = (inp[2]) ? 4'b0110 : 4'b0111;
										assign node20421 = (inp[7]) ? node20445 : node20422;
											assign node20422 = (inp[8]) ? node20436 : node20423;
												assign node20423 = (inp[14]) ? node20429 : node20424;
													assign node20424 = (inp[2]) ? node20426 : 4'b0111;
														assign node20426 = (inp[11]) ? 4'b0110 : 4'b1110;
													assign node20429 = (inp[2]) ? 4'b1110 : node20430;
														assign node20430 = (inp[1]) ? node20432 : 4'b1110;
															assign node20432 = (inp[6]) ? 4'b0110 : 4'b1110;
												assign node20436 = (inp[2]) ? node20442 : node20437;
													assign node20437 = (inp[14]) ? 4'b1111 : node20438;
														assign node20438 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node20442 = (inp[6]) ? 4'b1111 : 4'b0111;
											assign node20445 = (inp[11]) ? node20461 : node20446;
												assign node20446 = (inp[6]) ? node20450 : node20447;
													assign node20447 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node20450 = (inp[1]) ? node20454 : node20451;
														assign node20451 = (inp[2]) ? 4'b1110 : 4'b0110;
														assign node20454 = (inp[8]) ? node20458 : node20455;
															assign node20455 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node20458 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node20461 = (inp[6]) ? node20463 : 4'b1111;
													assign node20463 = (inp[14]) ? node20465 : 4'b0111;
														assign node20465 = (inp[8]) ? 4'b0110 : 4'b0111;
								assign node20468 = (inp[4]) ? node20568 : node20469;
									assign node20469 = (inp[12]) ? node20513 : node20470;
										assign node20470 = (inp[6]) ? node20498 : node20471;
											assign node20471 = (inp[11]) ? node20489 : node20472;
												assign node20472 = (inp[14]) ? node20478 : node20473;
													assign node20473 = (inp[7]) ? node20475 : 4'b1000;
														assign node20475 = (inp[2]) ? 4'b0001 : 4'b1000;
													assign node20478 = (inp[1]) ? node20484 : node20479;
														assign node20479 = (inp[2]) ? 4'b0001 : node20480;
															assign node20480 = (inp[8]) ? 4'b0001 : 4'b1000;
														assign node20484 = (inp[8]) ? node20486 : 4'b0001;
															assign node20486 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node20489 = (inp[14]) ? node20493 : node20490;
													assign node20490 = (inp[1]) ? 4'b1111 : 4'b0000;
													assign node20493 = (inp[8]) ? node20495 : 4'b1111;
														assign node20495 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node20498 = (inp[11]) ? node20510 : node20499;
												assign node20499 = (inp[1]) ? node20503 : node20500;
													assign node20500 = (inp[14]) ? 4'b1111 : 4'b0001;
													assign node20503 = (inp[7]) ? node20507 : node20504;
														assign node20504 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node20507 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node20510 = (inp[1]) ? 4'b0110 : 4'b1110;
										assign node20513 = (inp[14]) ? node20547 : node20514;
											assign node20514 = (inp[8]) ? node20526 : node20515;
												assign node20515 = (inp[2]) ? node20523 : node20516;
													assign node20516 = (inp[7]) ? node20520 : node20517;
														assign node20517 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node20520 = (inp[11]) ? 4'b1110 : 4'b0110;
													assign node20523 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node20526 = (inp[11]) ? node20538 : node20527;
													assign node20527 = (inp[1]) ? node20533 : node20528;
														assign node20528 = (inp[6]) ? node20530 : 4'b1110;
															assign node20530 = (inp[7]) ? 4'b1110 : 4'b0110;
														assign node20533 = (inp[2]) ? node20535 : 4'b1111;
															assign node20535 = (inp[6]) ? 4'b1110 : 4'b0110;
													assign node20538 = (inp[1]) ? 4'b0110 : node20539;
														assign node20539 = (inp[2]) ? node20543 : node20540;
															assign node20540 = (inp[7]) ? 4'b1111 : 4'b0110;
															assign node20543 = (inp[6]) ? 4'b0111 : 4'b1111;
											assign node20547 = (inp[8]) ? node20559 : node20548;
												assign node20548 = (inp[7]) ? node20552 : node20549;
													assign node20549 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node20552 = (inp[1]) ? 4'b1111 : node20553;
														assign node20553 = (inp[6]) ? 4'b0111 : node20554;
															assign node20554 = (inp[11]) ? 4'b1111 : 4'b0111;
												assign node20559 = (inp[7]) ? 4'b1110 : node20560;
													assign node20560 = (inp[11]) ? node20564 : node20561;
														assign node20561 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node20564 = (inp[6]) ? 4'b0111 : 4'b1111;
									assign node20568 = (inp[11]) ? node20610 : node20569;
										assign node20569 = (inp[12]) ? node20595 : node20570;
											assign node20570 = (inp[6]) ? node20588 : node20571;
												assign node20571 = (inp[1]) ? node20579 : node20572;
													assign node20572 = (inp[8]) ? 4'b0111 : node20573;
														assign node20573 = (inp[7]) ? node20575 : 4'b1110;
															assign node20575 = (inp[2]) ? 4'b0111 : 4'b1110;
													assign node20579 = (inp[8]) ? 4'b0110 : node20580;
														assign node20580 = (inp[2]) ? node20584 : node20581;
															assign node20581 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node20584 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node20588 = (inp[8]) ? node20592 : node20589;
													assign node20589 = (inp[1]) ? 4'b1011 : 4'b0110;
													assign node20592 = (inp[14]) ? 4'b1011 : 4'b1010;
											assign node20595 = (inp[8]) ? node20603 : node20596;
												assign node20596 = (inp[2]) ? node20598 : 4'b0010;
													assign node20598 = (inp[1]) ? 4'b1010 : node20599;
														assign node20599 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node20603 = (inp[7]) ? node20607 : node20604;
													assign node20604 = (inp[6]) ? 4'b1011 : 4'b0011;
													assign node20607 = (inp[6]) ? 4'b1010 : 4'b0010;
										assign node20610 = (inp[6]) ? node20626 : node20611;
											assign node20611 = (inp[1]) ? 4'b1010 : node20612;
												assign node20612 = (inp[8]) ? node20618 : node20613;
													assign node20613 = (inp[14]) ? node20615 : 4'b0010;
														assign node20615 = (inp[7]) ? 4'b1011 : 4'b0010;
													assign node20618 = (inp[7]) ? node20620 : 4'b1011;
														assign node20620 = (inp[2]) ? 4'b1010 : node20621;
															assign node20621 = (inp[14]) ? 4'b1010 : 4'b1011;
											assign node20626 = (inp[1]) ? node20642 : node20627;
												assign node20627 = (inp[7]) ? node20631 : node20628;
													assign node20628 = (inp[2]) ? 4'b0011 : 4'b1010;
													assign node20631 = (inp[12]) ? node20637 : node20632;
														assign node20632 = (inp[8]) ? node20634 : 4'b0011;
															assign node20634 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node20637 = (inp[14]) ? 4'b0011 : node20638;
															assign node20638 = (inp[2]) ? 4'b0010 : 4'b1010;
												assign node20642 = (inp[8]) ? node20644 : 4'b0011;
													assign node20644 = (inp[7]) ? 4'b0010 : 4'b0011;
							assign node20647 = (inp[12]) ? node20841 : node20648;
								assign node20648 = (inp[6]) ? node20728 : node20649;
									assign node20649 = (inp[11]) ? node20681 : node20650;
										assign node20650 = (inp[7]) ? node20668 : node20651;
											assign node20651 = (inp[1]) ? node20663 : node20652;
												assign node20652 = (inp[8]) ? node20660 : node20653;
													assign node20653 = (inp[2]) ? 4'b1010 : node20654;
														assign node20654 = (inp[4]) ? 4'b1111 : node20655;
															assign node20655 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node20660 = (inp[14]) ? 4'b0111 : 4'b1010;
												assign node20663 = (inp[4]) ? 4'b0011 : node20664;
													assign node20664 = (inp[2]) ? 4'b0110 : 4'b0010;
											assign node20668 = (inp[14]) ? node20672 : node20669;
												assign node20669 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node20672 = (inp[8]) ? node20676 : node20673;
													assign node20673 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node20676 = (inp[1]) ? 4'b0010 : node20677;
														assign node20677 = (inp[4]) ? 4'b0110 : 4'b0010;
										assign node20681 = (inp[1]) ? node20701 : node20682;
											assign node20682 = (inp[2]) ? node20690 : node20683;
												assign node20683 = (inp[7]) ? 4'b0010 : node20684;
													assign node20684 = (inp[8]) ? 4'b1111 : node20685;
														assign node20685 = (inp[4]) ? 4'b0110 : 4'b0111;
												assign node20690 = (inp[4]) ? node20698 : node20691;
													assign node20691 = (inp[7]) ? node20695 : node20692;
														assign node20692 = (inp[14]) ? 4'b1011 : 4'b0010;
														assign node20695 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node20698 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node20701 = (inp[4]) ? node20723 : node20702;
												assign node20702 = (inp[9]) ? node20714 : node20703;
													assign node20703 = (inp[2]) ? node20709 : node20704;
														assign node20704 = (inp[8]) ? 4'b1010 : node20705;
															assign node20705 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node20709 = (inp[14]) ? 4'b1011 : node20710;
															assign node20710 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node20714 = (inp[14]) ? node20718 : node20715;
														assign node20715 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node20718 = (inp[7]) ? 4'b1110 : node20719;
															assign node20719 = (inp[8]) ? 4'b1111 : 4'b1110;
												assign node20723 = (inp[9]) ? node20725 : 4'b1110;
													assign node20725 = (inp[7]) ? 4'b1011 : 4'b1010;
									assign node20728 = (inp[11]) ? node20782 : node20729;
										assign node20729 = (inp[8]) ? node20753 : node20730;
											assign node20730 = (inp[7]) ? node20742 : node20731;
												assign node20731 = (inp[1]) ? node20737 : node20732;
													assign node20732 = (inp[2]) ? 4'b0010 : node20733;
														assign node20733 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node20737 = (inp[4]) ? 4'b1011 : node20738;
														assign node20738 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node20742 = (inp[1]) ? node20748 : node20743;
													assign node20743 = (inp[2]) ? node20745 : 4'b1111;
														assign node20745 = (inp[14]) ? 4'b1011 : 4'b1111;
													assign node20748 = (inp[2]) ? 4'b1111 : node20749;
														assign node20749 = (inp[14]) ? 4'b1111 : 4'b1110;
											assign node20753 = (inp[7]) ? node20769 : node20754;
												assign node20754 = (inp[14]) ? node20758 : node20755;
													assign node20755 = (inp[1]) ? 4'b1110 : 4'b0110;
													assign node20758 = (inp[1]) ? node20764 : node20759;
														assign node20759 = (inp[9]) ? 4'b1011 : node20760;
															assign node20760 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node20764 = (inp[4]) ? node20766 : 4'b1111;
															assign node20766 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node20769 = (inp[14]) ? node20773 : node20770;
													assign node20770 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node20773 = (inp[2]) ? node20777 : node20774;
														assign node20774 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node20777 = (inp[9]) ? node20779 : 4'b1010;
															assign node20779 = (inp[4]) ? 4'b1010 : 4'b1110;
										assign node20782 = (inp[1]) ? node20810 : node20783;
											assign node20783 = (inp[2]) ? node20803 : node20784;
												assign node20784 = (inp[14]) ? node20796 : node20785;
													assign node20785 = (inp[8]) ? node20789 : node20786;
														assign node20786 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node20789 = (inp[4]) ? node20793 : node20790;
															assign node20790 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node20793 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node20796 = (inp[7]) ? 4'b0011 : node20797;
														assign node20797 = (inp[8]) ? 4'b0111 : node20798;
															assign node20798 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node20803 = (inp[4]) ? 4'b0111 : node20804;
													assign node20804 = (inp[14]) ? 4'b1010 : node20805;
														assign node20805 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node20810 = (inp[7]) ? node20830 : node20811;
												assign node20811 = (inp[14]) ? node20823 : node20812;
													assign node20812 = (inp[8]) ? node20818 : node20813;
														assign node20813 = (inp[4]) ? 4'b0011 : node20814;
															assign node20814 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node20818 = (inp[2]) ? 4'b0011 : node20819;
															assign node20819 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node20823 = (inp[8]) ? node20827 : node20824;
														assign node20824 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node20827 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node20830 = (inp[4]) ? node20836 : node20831;
													assign node20831 = (inp[2]) ? node20833 : 4'b0110;
														assign node20833 = (inp[14]) ? 4'b0111 : 4'b0011;
													assign node20836 = (inp[2]) ? 4'b0110 : node20837;
														assign node20837 = (inp[14]) ? 4'b0110 : 4'b0111;
								assign node20841 = (inp[6]) ? node20939 : node20842;
									assign node20842 = (inp[11]) ? node20896 : node20843;
										assign node20843 = (inp[8]) ? node20867 : node20844;
											assign node20844 = (inp[7]) ? node20850 : node20845;
												assign node20845 = (inp[1]) ? 4'b0111 : node20846;
													assign node20846 = (inp[4]) ? 4'b1011 : 4'b1010;
												assign node20850 = (inp[2]) ? node20856 : node20851;
													assign node20851 = (inp[14]) ? node20853 : 4'b1010;
														assign node20853 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node20856 = (inp[1]) ? node20862 : node20857;
														assign node20857 = (inp[14]) ? node20859 : 4'b0011;
															assign node20859 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node20862 = (inp[14]) ? node20864 : 4'b0111;
															assign node20864 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node20867 = (inp[7]) ? node20881 : node20868;
												assign node20868 = (inp[2]) ? node20874 : node20869;
													assign node20869 = (inp[14]) ? 4'b0111 : node20870;
														assign node20870 = (inp[4]) ? 4'b1010 : 4'b0010;
													assign node20874 = (inp[1]) ? 4'b0111 : node20875;
														assign node20875 = (inp[14]) ? 4'b0111 : node20876;
															assign node20876 = (inp[4]) ? 4'b0011 : 4'b0011;
												assign node20881 = (inp[14]) ? node20889 : node20882;
													assign node20882 = (inp[2]) ? 4'b0010 : node20883;
														assign node20883 = (inp[4]) ? node20885 : 4'b0011;
															assign node20885 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node20889 = (inp[1]) ? 4'b0010 : node20890;
														assign node20890 = (inp[2]) ? 4'b0110 : node20891;
															assign node20891 = (inp[4]) ? 4'b0010 : 4'b0010;
										assign node20896 = (inp[1]) ? node20924 : node20897;
											assign node20897 = (inp[14]) ? node20915 : node20898;
												assign node20898 = (inp[8]) ? node20904 : node20899;
													assign node20899 = (inp[2]) ? 4'b0110 : node20900;
														assign node20900 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node20904 = (inp[7]) ? node20910 : node20905;
														assign node20905 = (inp[2]) ? 4'b1111 : node20906;
															assign node20906 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node20910 = (inp[2]) ? node20912 : 4'b1111;
															assign node20912 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node20915 = (inp[2]) ? node20919 : node20916;
													assign node20916 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node20919 = (inp[7]) ? node20921 : 4'b1011;
														assign node20921 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node20924 = (inp[14]) ? node20932 : node20925;
												assign node20925 = (inp[9]) ? node20929 : node20926;
													assign node20926 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node20929 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node20932 = (inp[4]) ? node20934 : 4'b1011;
													assign node20934 = (inp[7]) ? 4'b1010 : node20935;
														assign node20935 = (inp[8]) ? 4'b1011 : 4'b1010;
									assign node20939 = (inp[11]) ? node20983 : node20940;
										assign node20940 = (inp[8]) ? node20964 : node20941;
											assign node20941 = (inp[7]) ? node20949 : node20942;
												assign node20942 = (inp[1]) ? node20944 : 4'b0010;
													assign node20944 = (inp[14]) ? node20946 : 4'b1010;
														assign node20946 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node20949 = (inp[14]) ? node20957 : node20950;
													assign node20950 = (inp[2]) ? node20952 : 4'b1010;
														assign node20952 = (inp[4]) ? node20954 : 4'b1111;
															assign node20954 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node20957 = (inp[1]) ? node20959 : 4'b1011;
														assign node20959 = (inp[4]) ? 4'b1011 : node20960;
															assign node20960 = (inp[9]) ? 4'b1111 : 4'b1011;
											assign node20964 = (inp[7]) ? node20976 : node20965;
												assign node20965 = (inp[14]) ? node20971 : node20966;
													assign node20966 = (inp[2]) ? node20968 : 4'b1010;
														assign node20968 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node20971 = (inp[4]) ? node20973 : 4'b1111;
														assign node20973 = (inp[1]) ? 4'b1111 : 4'b1011;
												assign node20976 = (inp[2]) ? node20978 : 4'b1111;
													assign node20978 = (inp[4]) ? 4'b1110 : node20979;
														assign node20979 = (inp[9]) ? 4'b1110 : 4'b1010;
										assign node20983 = (inp[7]) ? node21007 : node20984;
											assign node20984 = (inp[8]) ? node20998 : node20985;
												assign node20985 = (inp[1]) ? node20989 : node20986;
													assign node20986 = (inp[14]) ? 4'b1110 : 4'b1010;
													assign node20989 = (inp[2]) ? node20991 : 4'b0110;
														assign node20991 = (inp[14]) ? node20995 : node20992;
															assign node20992 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node20995 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node20998 = (inp[14]) ? node21004 : node20999;
													assign node20999 = (inp[2]) ? 4'b0011 : node21000;
														assign node21000 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node21004 = (inp[2]) ? 4'b0111 : 4'b0011;
											assign node21007 = (inp[8]) ? node21015 : node21008;
												assign node21008 = (inp[2]) ? 4'b0011 : node21009;
													assign node21009 = (inp[9]) ? node21011 : 4'b0110;
														assign node21011 = (inp[14]) ? 4'b0011 : 4'b0010;
												assign node21015 = (inp[2]) ? node21021 : node21016;
													assign node21016 = (inp[14]) ? node21018 : 4'b0011;
														assign node21018 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node21021 = (inp[1]) ? node21023 : 4'b0010;
														assign node21023 = (inp[4]) ? node21027 : node21024;
															assign node21024 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node21027 = (inp[9]) ? 4'b0010 : 4'b0110;
					assign node21030 = (inp[3]) ? node21774 : node21031;
						assign node21031 = (inp[5]) ? node21411 : node21032;
							assign node21032 = (inp[4]) ? node21208 : node21033;
								assign node21033 = (inp[9]) ? node21131 : node21034;
									assign node21034 = (inp[7]) ? node21086 : node21035;
										assign node21035 = (inp[8]) ? node21055 : node21036;
											assign node21036 = (inp[12]) ? node21050 : node21037;
												assign node21037 = (inp[6]) ? node21047 : node21038;
													assign node21038 = (inp[2]) ? node21042 : node21039;
														assign node21039 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node21042 = (inp[11]) ? node21044 : 4'b0110;
															assign node21044 = (inp[14]) ? 4'b1010 : 4'b0110;
													assign node21047 = (inp[1]) ? 4'b0010 : 4'b1010;
												assign node21050 = (inp[1]) ? node21052 : 4'b0010;
													assign node21052 = (inp[6]) ? 4'b0010 : 4'b0011;
											assign node21055 = (inp[12]) ? node21071 : node21056;
												assign node21056 = (inp[11]) ? node21064 : node21057;
													assign node21057 = (inp[2]) ? node21061 : node21058;
														assign node21058 = (inp[1]) ? 4'b1010 : 4'b0110;
														assign node21061 = (inp[6]) ? 4'b1011 : 4'b0111;
													assign node21064 = (inp[6]) ? 4'b0011 : node21065;
														assign node21065 = (inp[2]) ? 4'b1011 : node21066;
															assign node21066 = (inp[14]) ? 4'b1011 : 4'b1010;
												assign node21071 = (inp[14]) ? node21075 : node21072;
													assign node21072 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node21075 = (inp[1]) ? node21081 : node21076;
														assign node21076 = (inp[11]) ? node21078 : 4'b0011;
															assign node21078 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node21081 = (inp[11]) ? 4'b0011 : node21082;
															assign node21082 = (inp[6]) ? 4'b1011 : 4'b0011;
										assign node21086 = (inp[8]) ? node21114 : node21087;
											assign node21087 = (inp[2]) ? node21099 : node21088;
												assign node21088 = (inp[14]) ? node21096 : node21089;
													assign node21089 = (inp[11]) ? 4'b1010 : node21090;
														assign node21090 = (inp[6]) ? 4'b1010 : node21091;
															assign node21091 = (inp[1]) ? 4'b0110 : 4'b1010;
													assign node21096 = (inp[6]) ? 4'b1011 : 4'b0011;
												assign node21099 = (inp[1]) ? node21105 : node21100;
													assign node21100 = (inp[6]) ? node21102 : 4'b1011;
														assign node21102 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node21105 = (inp[14]) ? node21111 : node21106;
														assign node21106 = (inp[6]) ? node21108 : 4'b1011;
															assign node21108 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node21111 = (inp[6]) ? 4'b1011 : 4'b0011;
											assign node21114 = (inp[2]) ? node21126 : node21115;
												assign node21115 = (inp[14]) ? node21123 : node21116;
													assign node21116 = (inp[6]) ? node21120 : node21117;
														assign node21117 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node21120 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node21123 = (inp[6]) ? 4'b1010 : 4'b0110;
												assign node21126 = (inp[6]) ? node21128 : 4'b1010;
													assign node21128 = (inp[11]) ? 4'b0010 : 4'b1010;
									assign node21131 = (inp[6]) ? node21177 : node21132;
										assign node21132 = (inp[12]) ? node21146 : node21133;
											assign node21133 = (inp[11]) ? node21139 : node21134;
												assign node21134 = (inp[7]) ? node21136 : 4'b0011;
													assign node21136 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node21139 = (inp[2]) ? node21141 : 4'b0010;
													assign node21141 = (inp[7]) ? 4'b1111 : node21142;
														assign node21142 = (inp[8]) ? 4'b1111 : 4'b0010;
											assign node21146 = (inp[11]) ? node21164 : node21147;
												assign node21147 = (inp[8]) ? node21155 : node21148;
													assign node21148 = (inp[7]) ? 4'b0111 : node21149;
														assign node21149 = (inp[1]) ? 4'b0110 : node21150;
															assign node21150 = (inp[14]) ? 4'b1110 : 4'b1110;
													assign node21155 = (inp[7]) ? node21159 : node21156;
														assign node21156 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node21159 = (inp[14]) ? 4'b0110 : node21160;
															assign node21160 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node21164 = (inp[7]) ? node21172 : node21165;
													assign node21165 = (inp[1]) ? 4'b1111 : node21166;
														assign node21166 = (inp[2]) ? 4'b1111 : node21167;
															assign node21167 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node21172 = (inp[8]) ? node21174 : 4'b1111;
														assign node21174 = (inp[2]) ? 4'b1110 : 4'b1111;
										assign node21177 = (inp[11]) ? node21201 : node21178;
											assign node21178 = (inp[1]) ? node21194 : node21179;
												assign node21179 = (inp[2]) ? node21187 : node21180;
													assign node21180 = (inp[7]) ? node21182 : 4'b1111;
														assign node21182 = (inp[12]) ? node21184 : 4'b1111;
															assign node21184 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node21187 = (inp[12]) ? 4'b0110 : node21188;
														assign node21188 = (inp[8]) ? node21190 : 4'b1111;
															assign node21190 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node21194 = (inp[14]) ? 4'b1110 : node21195;
													assign node21195 = (inp[8]) ? 4'b1111 : node21196;
														assign node21196 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node21201 = (inp[8]) ? 4'b0111 : node21202;
												assign node21202 = (inp[1]) ? 4'b0111 : node21203;
													assign node21203 = (inp[2]) ? 4'b1110 : 4'b1111;
								assign node21208 = (inp[9]) ? node21312 : node21209;
									assign node21209 = (inp[12]) ? node21259 : node21210;
										assign node21210 = (inp[6]) ? node21232 : node21211;
											assign node21211 = (inp[11]) ? node21225 : node21212;
												assign node21212 = (inp[8]) ? node21220 : node21213;
													assign node21213 = (inp[7]) ? node21215 : 4'b1010;
														assign node21215 = (inp[2]) ? 4'b0011 : node21216;
															assign node21216 = (inp[14]) ? 4'b0011 : 4'b1010;
													assign node21220 = (inp[7]) ? 4'b0010 : node21221;
														assign node21221 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node21225 = (inp[2]) ? node21229 : node21226;
													assign node21226 = (inp[7]) ? 4'b1110 : 4'b0010;
													assign node21229 = (inp[7]) ? 4'b1111 : 4'b1110;
											assign node21232 = (inp[11]) ? node21246 : node21233;
												assign node21233 = (inp[7]) ? node21239 : node21234;
													assign node21234 = (inp[1]) ? node21236 : 4'b0010;
														assign node21236 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node21239 = (inp[14]) ? 4'b1110 : node21240;
														assign node21240 = (inp[2]) ? 4'b1110 : node21241;
															assign node21241 = (inp[1]) ? 4'b1110 : 4'b1111;
												assign node21246 = (inp[14]) ? node21252 : node21247;
													assign node21247 = (inp[1]) ? 4'b0110 : node21248;
														assign node21248 = (inp[7]) ? 4'b0111 : 4'b1110;
													assign node21252 = (inp[1]) ? 4'b0111 : node21253;
														assign node21253 = (inp[2]) ? node21255 : 4'b0111;
															assign node21255 = (inp[8]) ? 4'b0110 : 4'b0110;
										assign node21259 = (inp[14]) ? node21291 : node21260;
											assign node21260 = (inp[11]) ? node21274 : node21261;
												assign node21261 = (inp[8]) ? node21269 : node21262;
													assign node21262 = (inp[7]) ? 4'b0111 : node21263;
														assign node21263 = (inp[2]) ? 4'b1110 : node21264;
															assign node21264 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node21269 = (inp[2]) ? node21271 : 4'b0110;
														assign node21271 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node21274 = (inp[6]) ? node21284 : node21275;
													assign node21275 = (inp[1]) ? node21279 : node21276;
														assign node21276 = (inp[7]) ? 4'b1111 : 4'b0111;
														assign node21279 = (inp[2]) ? 4'b1110 : node21280;
															assign node21280 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node21284 = (inp[1]) ? node21288 : node21285;
														assign node21285 = (inp[8]) ? 4'b0110 : 4'b1110;
														assign node21288 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node21291 = (inp[8]) ? node21303 : node21292;
												assign node21292 = (inp[7]) ? 4'b1111 : node21293;
													assign node21293 = (inp[1]) ? 4'b1110 : node21294;
														assign node21294 = (inp[2]) ? node21298 : node21295;
															assign node21295 = (inp[6]) ? 4'b0110 : 4'b1110;
															assign node21298 = (inp[6]) ? 4'b1110 : 4'b0110;
												assign node21303 = (inp[7]) ? node21307 : node21304;
													assign node21304 = (inp[2]) ? 4'b1111 : 4'b0111;
													assign node21307 = (inp[6]) ? 4'b0110 : node21308;
														assign node21308 = (inp[11]) ? 4'b1110 : 4'b0110;
									assign node21312 = (inp[12]) ? node21372 : node21313;
										assign node21313 = (inp[6]) ? node21339 : node21314;
											assign node21314 = (inp[11]) ? node21326 : node21315;
												assign node21315 = (inp[2]) ? node21319 : node21316;
													assign node21316 = (inp[7]) ? 4'b0110 : 4'b1110;
													assign node21319 = (inp[7]) ? 4'b0111 : node21320;
														assign node21320 = (inp[1]) ? node21322 : 4'b1110;
															assign node21322 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node21326 = (inp[14]) ? node21334 : node21327;
													assign node21327 = (inp[2]) ? node21331 : node21328;
														assign node21328 = (inp[1]) ? 4'b1010 : 4'b0110;
														assign node21331 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node21334 = (inp[7]) ? node21336 : 4'b1011;
														assign node21336 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node21339 = (inp[11]) ? node21361 : node21340;
												assign node21340 = (inp[1]) ? node21348 : node21341;
													assign node21341 = (inp[8]) ? 4'b1011 : node21342;
														assign node21342 = (inp[14]) ? 4'b0110 : node21343;
															assign node21343 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node21348 = (inp[2]) ? node21354 : node21349;
														assign node21349 = (inp[8]) ? node21351 : 4'b1011;
															assign node21351 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node21354 = (inp[7]) ? node21358 : node21355;
															assign node21355 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node21358 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node21361 = (inp[14]) ? node21369 : node21362;
													assign node21362 = (inp[7]) ? node21364 : 4'b0011;
														assign node21364 = (inp[1]) ? 4'b0010 : node21365;
															assign node21365 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node21369 = (inp[8]) ? 4'b0010 : 4'b1010;
										assign node21372 = (inp[7]) ? node21394 : node21373;
											assign node21373 = (inp[8]) ? node21387 : node21374;
												assign node21374 = (inp[2]) ? node21376 : 4'b0011;
													assign node21376 = (inp[1]) ? node21382 : node21377;
														assign node21377 = (inp[6]) ? node21379 : 4'b0010;
															assign node21379 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node21382 = (inp[6]) ? node21384 : 4'b1010;
															assign node21384 = (inp[11]) ? 4'b0010 : 4'b1010;
												assign node21387 = (inp[2]) ? node21391 : node21388;
													assign node21388 = (inp[6]) ? 4'b1010 : 4'b0011;
													assign node21391 = (inp[14]) ? 4'b1011 : 4'b0011;
											assign node21394 = (inp[8]) ? node21404 : node21395;
												assign node21395 = (inp[2]) ? node21399 : node21396;
													assign node21396 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node21399 = (inp[11]) ? 4'b0011 : node21400;
														assign node21400 = (inp[6]) ? 4'b1011 : 4'b0011;
												assign node21404 = (inp[2]) ? node21406 : 4'b1011;
													assign node21406 = (inp[11]) ? node21408 : 4'b1010;
														assign node21408 = (inp[6]) ? 4'b0010 : 4'b1010;
							assign node21411 = (inp[9]) ? node21583 : node21412;
								assign node21412 = (inp[4]) ? node21500 : node21413;
									assign node21413 = (inp[6]) ? node21457 : node21414;
										assign node21414 = (inp[11]) ? node21438 : node21415;
											assign node21415 = (inp[12]) ? node21423 : node21416;
												assign node21416 = (inp[1]) ? 4'b0111 : node21417;
													assign node21417 = (inp[8]) ? 4'b0110 : node21418;
														assign node21418 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node21423 = (inp[7]) ? node21433 : node21424;
													assign node21424 = (inp[1]) ? node21430 : node21425;
														assign node21425 = (inp[14]) ? 4'b1010 : node21426;
															assign node21426 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node21430 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node21433 = (inp[1]) ? node21435 : 4'b0011;
														assign node21435 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node21438 = (inp[12]) ? node21446 : node21439;
												assign node21439 = (inp[1]) ? 4'b1010 : node21440;
													assign node21440 = (inp[2]) ? 4'b1011 : node21441;
														assign node21441 = (inp[8]) ? 4'b1011 : 4'b0110;
												assign node21446 = (inp[2]) ? 4'b1011 : node21447;
													assign node21447 = (inp[1]) ? node21453 : node21448;
														assign node21448 = (inp[7]) ? node21450 : 4'b0010;
															assign node21450 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node21453 = (inp[7]) ? 4'b1010 : 4'b1011;
										assign node21457 = (inp[11]) ? node21481 : node21458;
											assign node21458 = (inp[12]) ? node21474 : node21459;
												assign node21459 = (inp[1]) ? node21467 : node21460;
													assign node21460 = (inp[7]) ? node21462 : 4'b1011;
														assign node21462 = (inp[8]) ? node21464 : 4'b1011;
															assign node21464 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node21467 = (inp[14]) ? node21469 : 4'b1010;
														assign node21469 = (inp[8]) ? node21471 : 4'b1011;
															assign node21471 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node21474 = (inp[8]) ? node21478 : node21475;
													assign node21475 = (inp[2]) ? 4'b0010 : 4'b1010;
													assign node21478 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node21481 = (inp[1]) ? node21493 : node21482;
												assign node21482 = (inp[8]) ? node21484 : 4'b1010;
													assign node21484 = (inp[14]) ? 4'b0011 : node21485;
														assign node21485 = (inp[7]) ? node21489 : node21486;
															assign node21486 = (inp[2]) ? 4'b0011 : 4'b1010;
															assign node21489 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node21493 = (inp[14]) ? node21495 : 4'b0010;
													assign node21495 = (inp[8]) ? 4'b0010 : node21496;
														assign node21496 = (inp[7]) ? 4'b0011 : 4'b0010;
									assign node21500 = (inp[12]) ? node21548 : node21501;
										assign node21501 = (inp[11]) ? node21523 : node21502;
											assign node21502 = (inp[6]) ? node21510 : node21503;
												assign node21503 = (inp[8]) ? 4'b0011 : node21504;
													assign node21504 = (inp[2]) ? node21506 : 4'b0010;
														assign node21506 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node21510 = (inp[8]) ? node21518 : node21511;
													assign node21511 = (inp[7]) ? 4'b1101 : node21512;
														assign node21512 = (inp[2]) ? 4'b0010 : node21513;
															assign node21513 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node21518 = (inp[7]) ? node21520 : 4'b1101;
														assign node21520 = (inp[1]) ? 4'b1101 : 4'b1100;
											assign node21523 = (inp[6]) ? node21533 : node21524;
												assign node21524 = (inp[2]) ? node21526 : 4'b0011;
													assign node21526 = (inp[8]) ? node21530 : node21527;
														assign node21527 = (inp[7]) ? 4'b1101 : 4'b0010;
														assign node21530 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node21533 = (inp[1]) ? node21543 : node21534;
													assign node21534 = (inp[8]) ? node21536 : 4'b1100;
														assign node21536 = (inp[7]) ? node21540 : node21537;
															assign node21537 = (inp[14]) ? 4'b0101 : 4'b1100;
															assign node21540 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node21543 = (inp[8]) ? 4'b0100 : node21544;
														assign node21544 = (inp[14]) ? 4'b0100 : 4'b0101;
										assign node21548 = (inp[14]) ? node21566 : node21549;
											assign node21549 = (inp[11]) ? node21557 : node21550;
												assign node21550 = (inp[7]) ? node21554 : node21551;
													assign node21551 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node21554 = (inp[6]) ? 4'b1101 : 4'b0101;
												assign node21557 = (inp[6]) ? 4'b0100 : node21558;
													assign node21558 = (inp[7]) ? node21560 : 4'b1100;
														assign node21560 = (inp[1]) ? 4'b1101 : node21561;
															assign node21561 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node21566 = (inp[2]) ? node21572 : node21567;
												assign node21567 = (inp[1]) ? node21569 : 4'b0101;
													assign node21569 = (inp[8]) ? 4'b0101 : 4'b1100;
												assign node21572 = (inp[1]) ? node21576 : node21573;
													assign node21573 = (inp[7]) ? 4'b0101 : 4'b1100;
													assign node21576 = (inp[7]) ? 4'b1100 : node21577;
														assign node21577 = (inp[8]) ? 4'b0101 : node21578;
															assign node21578 = (inp[6]) ? 4'b0100 : 4'b0100;
								assign node21583 = (inp[4]) ? node21691 : node21584;
									assign node21584 = (inp[12]) ? node21634 : node21585;
										assign node21585 = (inp[6]) ? node21607 : node21586;
											assign node21586 = (inp[11]) ? node21596 : node21587;
												assign node21587 = (inp[8]) ? node21591 : node21588;
													assign node21588 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node21591 = (inp[7]) ? node21593 : 4'b0011;
														assign node21593 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node21596 = (inp[7]) ? node21602 : node21597;
													assign node21597 = (inp[2]) ? 4'b1101 : node21598;
														assign node21598 = (inp[1]) ? 4'b1100 : 4'b0010;
													assign node21602 = (inp[1]) ? 4'b1101 : node21603;
														assign node21603 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node21607 = (inp[11]) ? node21625 : node21608;
												assign node21608 = (inp[1]) ? node21612 : node21609;
													assign node21609 = (inp[7]) ? 4'b1100 : 4'b0010;
													assign node21612 = (inp[2]) ? node21618 : node21613;
														assign node21613 = (inp[8]) ? 4'b1101 : node21614;
															assign node21614 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node21618 = (inp[14]) ? node21622 : node21619;
															assign node21619 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node21622 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node21625 = (inp[7]) ? node21627 : 4'b1100;
													assign node21627 = (inp[1]) ? node21629 : 4'b0101;
														assign node21629 = (inp[14]) ? node21631 : 4'b0100;
															assign node21631 = (inp[8]) ? 4'b0100 : 4'b0101;
										assign node21634 = (inp[14]) ? node21664 : node21635;
											assign node21635 = (inp[1]) ? node21647 : node21636;
												assign node21636 = (inp[2]) ? node21644 : node21637;
													assign node21637 = (inp[11]) ? node21641 : node21638;
														assign node21638 = (inp[6]) ? 4'b0100 : 4'b1100;
														assign node21641 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node21644 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node21647 = (inp[8]) ? node21655 : node21648;
													assign node21648 = (inp[2]) ? 4'b0100 : node21649;
														assign node21649 = (inp[7]) ? node21651 : 4'b1101;
															assign node21651 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node21655 = (inp[7]) ? node21659 : node21656;
														assign node21656 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node21659 = (inp[6]) ? node21661 : 4'b1101;
															assign node21661 = (inp[11]) ? 4'b0101 : 4'b1101;
											assign node21664 = (inp[1]) ? node21676 : node21665;
												assign node21665 = (inp[11]) ? 4'b1101 : node21666;
													assign node21666 = (inp[6]) ? node21670 : node21667;
														assign node21667 = (inp[7]) ? 4'b0101 : 4'b1100;
														assign node21670 = (inp[7]) ? node21672 : 4'b1101;
															assign node21672 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node21676 = (inp[7]) ? node21684 : node21677;
													assign node21677 = (inp[8]) ? node21679 : 4'b0100;
														assign node21679 = (inp[6]) ? 4'b1101 : node21680;
															assign node21680 = (inp[2]) ? 4'b1101 : 4'b0101;
													assign node21684 = (inp[2]) ? node21686 : 4'b1101;
														assign node21686 = (inp[11]) ? node21688 : 4'b1100;
															assign node21688 = (inp[6]) ? 4'b0100 : 4'b1100;
									assign node21691 = (inp[12]) ? node21733 : node21692;
										assign node21692 = (inp[11]) ? node21712 : node21693;
											assign node21693 = (inp[6]) ? node21701 : node21694;
												assign node21694 = (inp[2]) ? node21696 : 4'b0100;
													assign node21696 = (inp[8]) ? 4'b0101 : node21697;
														assign node21697 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node21701 = (inp[14]) ? node21709 : node21702;
													assign node21702 = (inp[1]) ? 4'b1001 : node21703;
														assign node21703 = (inp[8]) ? 4'b0100 : node21704;
															assign node21704 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node21709 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node21712 = (inp[6]) ? node21722 : node21713;
												assign node21713 = (inp[7]) ? node21717 : node21714;
													assign node21714 = (inp[1]) ? 4'b1000 : 4'b0100;
													assign node21717 = (inp[14]) ? 4'b1001 : node21718;
														assign node21718 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node21722 = (inp[8]) ? node21728 : node21723;
													assign node21723 = (inp[7]) ? 4'b1000 : node21724;
														assign node21724 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node21728 = (inp[7]) ? node21730 : 4'b0001;
														assign node21730 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node21733 = (inp[6]) ? node21753 : node21734;
											assign node21734 = (inp[11]) ? node21744 : node21735;
												assign node21735 = (inp[8]) ? node21739 : node21736;
													assign node21736 = (inp[1]) ? 4'b0001 : 4'b1000;
													assign node21739 = (inp[14]) ? node21741 : 4'b0000;
														assign node21741 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node21744 = (inp[1]) ? 4'b1000 : node21745;
													assign node21745 = (inp[2]) ? node21747 : 4'b0000;
														assign node21747 = (inp[14]) ? node21749 : 4'b1001;
															assign node21749 = (inp[8]) ? 4'b1000 : 4'b0000;
											assign node21753 = (inp[11]) ? node21765 : node21754;
												assign node21754 = (inp[8]) ? node21760 : node21755;
													assign node21755 = (inp[1]) ? node21757 : 4'b0000;
														assign node21757 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node21760 = (inp[2]) ? node21762 : 4'b1001;
														assign node21762 = (inp[1]) ? 4'b1000 : 4'b1001;
												assign node21765 = (inp[7]) ? node21771 : node21766;
													assign node21766 = (inp[1]) ? 4'b0000 : node21767;
														assign node21767 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node21771 = (inp[8]) ? 4'b0000 : 4'b0001;
						assign node21774 = (inp[5]) ? node22126 : node21775;
							assign node21775 = (inp[4]) ? node21943 : node21776;
								assign node21776 = (inp[9]) ? node21858 : node21777;
									assign node21777 = (inp[12]) ? node21815 : node21778;
										assign node21778 = (inp[6]) ? node21802 : node21779;
											assign node21779 = (inp[11]) ? node21795 : node21780;
												assign node21780 = (inp[1]) ? node21786 : node21781;
													assign node21781 = (inp[2]) ? node21783 : 4'b1110;
														assign node21783 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node21786 = (inp[14]) ? node21788 : 4'b0110;
														assign node21788 = (inp[7]) ? node21792 : node21789;
															assign node21789 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node21792 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node21795 = (inp[14]) ? node21799 : node21796;
													assign node21796 = (inp[8]) ? 4'b1010 : 4'b0110;
													assign node21799 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node21802 = (inp[11]) ? node21808 : node21803;
												assign node21803 = (inp[8]) ? 4'b1010 : node21804;
													assign node21804 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node21808 = (inp[1]) ? 4'b0010 : node21809;
													assign node21809 = (inp[8]) ? node21811 : 4'b0011;
														assign node21811 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node21815 = (inp[1]) ? node21831 : node21816;
											assign node21816 = (inp[7]) ? node21826 : node21817;
												assign node21817 = (inp[14]) ? 4'b0010 : node21818;
													assign node21818 = (inp[8]) ? node21820 : 4'b1010;
														assign node21820 = (inp[2]) ? 4'b0011 : node21821;
															assign node21821 = (inp[11]) ? 4'b0010 : 4'b0010;
												assign node21826 = (inp[8]) ? node21828 : 4'b1011;
													assign node21828 = (inp[6]) ? 4'b0010 : 4'b1010;
											assign node21831 = (inp[11]) ? node21847 : node21832;
												assign node21832 = (inp[6]) ? node21838 : node21833;
													assign node21833 = (inp[14]) ? 4'b0011 : node21834;
														assign node21834 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node21838 = (inp[7]) ? 4'b1010 : node21839;
														assign node21839 = (inp[14]) ? node21843 : node21840;
															assign node21840 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node21843 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node21847 = (inp[6]) ? node21849 : 4'b1010;
													assign node21849 = (inp[8]) ? 4'b0011 : node21850;
														assign node21850 = (inp[7]) ? node21854 : node21851;
															assign node21851 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node21854 = (inp[2]) ? 4'b0011 : 4'b0010;
									assign node21858 = (inp[12]) ? node21898 : node21859;
										assign node21859 = (inp[11]) ? node21879 : node21860;
											assign node21860 = (inp[6]) ? node21872 : node21861;
												assign node21861 = (inp[8]) ? node21865 : node21862;
													assign node21862 = (inp[14]) ? 4'b0010 : 4'b1010;
													assign node21865 = (inp[1]) ? node21867 : 4'b0011;
														assign node21867 = (inp[2]) ? 4'b0010 : node21868;
															assign node21868 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node21872 = (inp[7]) ? node21876 : node21873;
													assign node21873 = (inp[8]) ? 4'b1101 : 4'b0010;
													assign node21876 = (inp[1]) ? 4'b1100 : 4'b1101;
											assign node21879 = (inp[6]) ? node21891 : node21880;
												assign node21880 = (inp[1]) ? node21884 : node21881;
													assign node21881 = (inp[7]) ? 4'b1101 : 4'b0011;
													assign node21884 = (inp[7]) ? 4'b1100 : node21885;
														assign node21885 = (inp[14]) ? node21887 : 4'b1100;
															assign node21887 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node21891 = (inp[14]) ? node21893 : 4'b0100;
													assign node21893 = (inp[2]) ? 4'b0101 : node21894;
														assign node21894 = (inp[8]) ? 4'b0100 : 4'b0101;
										assign node21898 = (inp[1]) ? node21926 : node21899;
											assign node21899 = (inp[14]) ? node21917 : node21900;
												assign node21900 = (inp[7]) ? node21908 : node21901;
													assign node21901 = (inp[8]) ? 4'b1101 : node21902;
														assign node21902 = (inp[11]) ? 4'b0100 : node21903;
															assign node21903 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node21908 = (inp[2]) ? node21912 : node21909;
														assign node21909 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node21912 = (inp[6]) ? 4'b1101 : node21913;
															assign node21913 = (inp[11]) ? 4'b1101 : 4'b0101;
												assign node21917 = (inp[11]) ? 4'b0101 : node21918;
													assign node21918 = (inp[7]) ? node21922 : node21919;
														assign node21919 = (inp[8]) ? 4'b0101 : 4'b1100;
														assign node21922 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node21926 = (inp[8]) ? node21934 : node21927;
												assign node21927 = (inp[6]) ? node21931 : node21928;
													assign node21928 = (inp[11]) ? 4'b1100 : 4'b0101;
													assign node21931 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node21934 = (inp[7]) ? node21938 : node21935;
													assign node21935 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node21938 = (inp[6]) ? node21940 : 4'b1100;
														assign node21940 = (inp[11]) ? 4'b0100 : 4'b1100;
								assign node21943 = (inp[9]) ? node22047 : node21944;
									assign node21944 = (inp[12]) ? node21986 : node21945;
										assign node21945 = (inp[6]) ? node21969 : node21946;
											assign node21946 = (inp[11]) ? node21956 : node21947;
												assign node21947 = (inp[2]) ? node21949 : 4'b0011;
													assign node21949 = (inp[14]) ? 4'b0010 : node21950;
														assign node21950 = (inp[1]) ? 4'b0011 : node21951;
															assign node21951 = (inp[7]) ? 4'b0010 : 4'b1010;
												assign node21956 = (inp[2]) ? node21964 : node21957;
													assign node21957 = (inp[8]) ? 4'b1100 : node21958;
														assign node21958 = (inp[7]) ? 4'b0010 : node21959;
															assign node21959 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node21964 = (inp[1]) ? node21966 : 4'b1100;
														assign node21966 = (inp[8]) ? 4'b1101 : 4'b1100;
											assign node21969 = (inp[11]) ? node21975 : node21970;
												assign node21970 = (inp[7]) ? 4'b1100 : node21971;
													assign node21971 = (inp[1]) ? 4'b1100 : 4'b0010;
												assign node21975 = (inp[2]) ? node21983 : node21976;
													assign node21976 = (inp[1]) ? 4'b0101 : node21977;
														assign node21977 = (inp[14]) ? 4'b0101 : node21978;
															assign node21978 = (inp[8]) ? 4'b0101 : 4'b1100;
													assign node21983 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node21986 = (inp[1]) ? node22016 : node21987;
											assign node21987 = (inp[2]) ? node22003 : node21988;
												assign node21988 = (inp[11]) ? node21996 : node21989;
													assign node21989 = (inp[8]) ? 4'b1100 : node21990;
														assign node21990 = (inp[7]) ? node21992 : 4'b1101;
															assign node21992 = (inp[6]) ? 4'b1101 : 4'b1100;
													assign node21996 = (inp[6]) ? node21998 : 4'b1101;
														assign node21998 = (inp[14]) ? 4'b0101 : node21999;
															assign node21999 = (inp[7]) ? 4'b0101 : 4'b1100;
												assign node22003 = (inp[7]) ? node22011 : node22004;
													assign node22004 = (inp[8]) ? node22006 : 4'b0100;
														assign node22006 = (inp[14]) ? node22008 : 4'b0101;
															assign node22008 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node22011 = (inp[8]) ? 4'b1100 : node22012;
														assign node22012 = (inp[14]) ? 4'b0101 : 4'b1101;
											assign node22016 = (inp[8]) ? node22038 : node22017;
												assign node22017 = (inp[7]) ? node22029 : node22018;
													assign node22018 = (inp[14]) ? node22024 : node22019;
														assign node22019 = (inp[6]) ? 4'b1101 : node22020;
															assign node22020 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node22024 = (inp[6]) ? 4'b0100 : node22025;
															assign node22025 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node22029 = (inp[14]) ? node22033 : node22030;
														assign node22030 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node22033 = (inp[2]) ? 4'b1101 : node22034;
															assign node22034 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node22038 = (inp[2]) ? node22040 : 4'b1100;
													assign node22040 = (inp[7]) ? node22042 : 4'b0101;
														assign node22042 = (inp[11]) ? 4'b0100 : node22043;
															assign node22043 = (inp[6]) ? 4'b1100 : 4'b0100;
									assign node22047 = (inp[12]) ? node22093 : node22048;
										assign node22048 = (inp[11]) ? node22068 : node22049;
											assign node22049 = (inp[6]) ? node22057 : node22050;
												assign node22050 = (inp[1]) ? 4'b0101 : node22051;
													assign node22051 = (inp[7]) ? node22053 : 4'b1100;
														assign node22053 = (inp[8]) ? 4'b0100 : 4'b1100;
												assign node22057 = (inp[7]) ? node22063 : node22058;
													assign node22058 = (inp[1]) ? node22060 : 4'b0100;
														assign node22060 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node22063 = (inp[14]) ? 4'b1000 : node22064;
														assign node22064 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node22068 = (inp[6]) ? node22084 : node22069;
												assign node22069 = (inp[14]) ? node22077 : node22070;
													assign node22070 = (inp[2]) ? node22072 : 4'b0100;
														assign node22072 = (inp[1]) ? 4'b1000 : node22073;
															assign node22073 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node22077 = (inp[2]) ? 4'b1001 : node22078;
														assign node22078 = (inp[7]) ? node22080 : 4'b1000;
															assign node22080 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node22084 = (inp[8]) ? node22086 : 4'b0001;
													assign node22086 = (inp[2]) ? node22090 : node22087;
														assign node22087 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node22090 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node22093 = (inp[11]) ? node22111 : node22094;
											assign node22094 = (inp[6]) ? node22104 : node22095;
												assign node22095 = (inp[7]) ? 4'b0001 : node22096;
													assign node22096 = (inp[8]) ? node22100 : node22097;
														assign node22097 = (inp[14]) ? 4'b1000 : 4'b0000;
														assign node22100 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node22104 = (inp[8]) ? 4'b1001 : node22105;
													assign node22105 = (inp[7]) ? node22107 : 4'b0000;
														assign node22107 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node22111 = (inp[6]) ? node22119 : node22112;
												assign node22112 = (inp[1]) ? 4'b1001 : node22113;
													assign node22113 = (inp[7]) ? node22115 : 4'b0000;
														assign node22115 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node22119 = (inp[1]) ? 4'b0000 : node22120;
													assign node22120 = (inp[7]) ? 4'b0000 : node22121;
														assign node22121 = (inp[8]) ? 4'b0001 : 4'b1001;
							assign node22126 = (inp[8]) ? node22280 : node22127;
								assign node22127 = (inp[7]) ? node22213 : node22128;
									assign node22128 = (inp[14]) ? node22168 : node22129;
										assign node22129 = (inp[2]) ? node22151 : node22130;
											assign node22130 = (inp[6]) ? node22142 : node22131;
												assign node22131 = (inp[11]) ? node22137 : node22132;
													assign node22132 = (inp[1]) ? node22134 : 4'b1101;
														assign node22134 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node22137 = (inp[1]) ? node22139 : 4'b0001;
														assign node22139 = (inp[9]) ? 4'b1101 : 4'b1001;
												assign node22142 = (inp[12]) ? 4'b1001 : node22143;
													assign node22143 = (inp[11]) ? 4'b0101 : node22144;
														assign node22144 = (inp[4]) ? node22146 : 4'b1101;
															assign node22146 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node22151 = (inp[1]) ? node22163 : node22152;
												assign node22152 = (inp[6]) ? node22156 : node22153;
													assign node22153 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node22156 = (inp[11]) ? node22158 : 4'b0100;
														assign node22158 = (inp[4]) ? 4'b1000 : node22159;
															assign node22159 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node22163 = (inp[4]) ? node22165 : 4'b1000;
													assign node22165 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node22168 = (inp[4]) ? node22186 : node22169;
											assign node22169 = (inp[9]) ? node22175 : node22170;
												assign node22170 = (inp[12]) ? 4'b1000 : node22171;
													assign node22171 = (inp[11]) ? 4'b0000 : 4'b0100;
												assign node22175 = (inp[2]) ? node22183 : node22176;
													assign node22176 = (inp[6]) ? 4'b1100 : node22177;
														assign node22177 = (inp[11]) ? node22179 : 4'b1100;
															assign node22179 = (inp[1]) ? 4'b1100 : 4'b0100;
													assign node22183 = (inp[12]) ? 4'b0100 : 4'b1100;
											assign node22186 = (inp[9]) ? node22198 : node22187;
												assign node22187 = (inp[12]) ? node22195 : node22188;
													assign node22188 = (inp[11]) ? 4'b1100 : node22189;
														assign node22189 = (inp[6]) ? 4'b1100 : node22190;
															assign node22190 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node22195 = (inp[1]) ? 4'b1100 : 4'b0100;
												assign node22198 = (inp[12]) ? node22206 : node22199;
													assign node22199 = (inp[1]) ? node22201 : 4'b0100;
														assign node22201 = (inp[11]) ? 4'b1000 : node22202;
															assign node22202 = (inp[6]) ? 4'b1000 : 4'b0100;
													assign node22206 = (inp[2]) ? node22208 : 4'b0000;
														assign node22208 = (inp[11]) ? node22210 : 4'b1000;
															assign node22210 = (inp[1]) ? 4'b0000 : 4'b1000;
									assign node22213 = (inp[2]) ? node22255 : node22214;
										assign node22214 = (inp[14]) ? node22238 : node22215;
											assign node22215 = (inp[11]) ? node22227 : node22216;
												assign node22216 = (inp[6]) ? node22224 : node22217;
													assign node22217 = (inp[1]) ? 4'b0000 : node22218;
														assign node22218 = (inp[12]) ? 4'b1000 : node22219;
															assign node22219 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node22224 = (inp[12]) ? 4'b1100 : 4'b0100;
												assign node22227 = (inp[9]) ? node22231 : node22228;
													assign node22228 = (inp[1]) ? 4'b1100 : 4'b0100;
													assign node22231 = (inp[6]) ? node22233 : 4'b0000;
														assign node22233 = (inp[1]) ? node22235 : 4'b1100;
															assign node22235 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node22238 = (inp[4]) ? node22248 : node22239;
												assign node22239 = (inp[9]) ? node22243 : node22240;
													assign node22240 = (inp[12]) ? 4'b1001 : 4'b0001;
													assign node22243 = (inp[6]) ? 4'b0101 : node22244;
														assign node22244 = (inp[11]) ? 4'b1101 : 4'b0101;
												assign node22248 = (inp[9]) ? 4'b1001 : node22249;
													assign node22249 = (inp[11]) ? node22251 : 4'b1101;
														assign node22251 = (inp[6]) ? 4'b0101 : 4'b1101;
										assign node22255 = (inp[4]) ? node22269 : node22256;
											assign node22256 = (inp[9]) ? node22264 : node22257;
												assign node22257 = (inp[11]) ? node22261 : node22258;
													assign node22258 = (inp[6]) ? 4'b1001 : 4'b0101;
													assign node22261 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node22264 = (inp[6]) ? node22266 : 4'b0001;
													assign node22266 = (inp[11]) ? 4'b0101 : 4'b1101;
											assign node22269 = (inp[9]) ? node22275 : node22270;
												assign node22270 = (inp[6]) ? 4'b1101 : node22271;
													assign node22271 = (inp[11]) ? 4'b1101 : 4'b0001;
												assign node22275 = (inp[12]) ? 4'b1001 : node22276;
													assign node22276 = (inp[6]) ? 4'b1001 : 4'b0101;
								assign node22280 = (inp[7]) ? node22364 : node22281;
									assign node22281 = (inp[14]) ? node22327 : node22282;
										assign node22282 = (inp[2]) ? node22308 : node22283;
											assign node22283 = (inp[4]) ? node22293 : node22284;
												assign node22284 = (inp[9]) ? 4'b0100 : node22285;
													assign node22285 = (inp[11]) ? node22287 : 4'b0000;
														assign node22287 = (inp[6]) ? 4'b0000 : node22288;
															assign node22288 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node22293 = (inp[9]) ? node22301 : node22294;
													assign node22294 = (inp[11]) ? 4'b1100 : node22295;
														assign node22295 = (inp[1]) ? node22297 : 4'b0100;
															assign node22297 = (inp[6]) ? 4'b1100 : 4'b0100;
													assign node22301 = (inp[12]) ? 4'b0000 : node22302;
														assign node22302 = (inp[1]) ? 4'b0100 : node22303;
															assign node22303 = (inp[11]) ? 4'b0100 : 4'b1100;
											assign node22308 = (inp[6]) ? node22314 : node22309;
												assign node22309 = (inp[4]) ? 4'b1001 : node22310;
													assign node22310 = (inp[11]) ? 4'b1101 : 4'b0101;
												assign node22314 = (inp[11]) ? node22322 : node22315;
													assign node22315 = (inp[1]) ? 4'b1101 : node22316;
														assign node22316 = (inp[9]) ? node22318 : 4'b1001;
															assign node22318 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node22322 = (inp[9]) ? 4'b0001 : node22323;
														assign node22323 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node22327 = (inp[6]) ? node22347 : node22328;
											assign node22328 = (inp[11]) ? node22340 : node22329;
												assign node22329 = (inp[1]) ? 4'b0101 : node22330;
													assign node22330 = (inp[12]) ? node22332 : 4'b0001;
														assign node22332 = (inp[9]) ? node22336 : node22333;
															assign node22333 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node22336 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node22340 = (inp[9]) ? node22344 : node22341;
													assign node22341 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node22344 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node22347 = (inp[11]) ? node22351 : node22348;
												assign node22348 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node22351 = (inp[2]) ? node22359 : node22352;
													assign node22352 = (inp[1]) ? 4'b0101 : node22353;
														assign node22353 = (inp[4]) ? node22355 : 4'b0001;
															assign node22355 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node22359 = (inp[4]) ? 4'b0001 : node22360;
														assign node22360 = (inp[9]) ? 4'b0101 : 4'b0001;
									assign node22364 = (inp[14]) ? node22412 : node22365;
										assign node22365 = (inp[2]) ? node22397 : node22366;
											assign node22366 = (inp[1]) ? node22392 : node22367;
												assign node22367 = (inp[4]) ? node22381 : node22368;
													assign node22368 = (inp[9]) ? node22376 : node22369;
														assign node22369 = (inp[11]) ? node22373 : node22370;
															assign node22370 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node22373 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node22376 = (inp[11]) ? node22378 : 4'b0001;
															assign node22378 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node22381 = (inp[9]) ? node22389 : node22382;
														assign node22382 = (inp[12]) ? node22386 : node22383;
															assign node22383 = (inp[11]) ? 4'b0101 : 4'b0001;
															assign node22386 = (inp[6]) ? 4'b1101 : 4'b0101;
														assign node22389 = (inp[11]) ? 4'b0001 : 4'b0101;
												assign node22392 = (inp[9]) ? 4'b1001 : node22393;
													assign node22393 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node22397 = (inp[6]) ? node22407 : node22398;
												assign node22398 = (inp[11]) ? node22400 : 4'b0100;
													assign node22400 = (inp[12]) ? node22402 : 4'b1100;
														assign node22402 = (inp[9]) ? 4'b1000 : node22403;
															assign node22403 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node22407 = (inp[11]) ? 4'b0000 : node22408;
													assign node22408 = (inp[12]) ? 4'b1100 : 4'b1000;
										assign node22412 = (inp[11]) ? node22432 : node22413;
											assign node22413 = (inp[6]) ? node22421 : node22414;
												assign node22414 = (inp[12]) ? 4'b0000 : node22415;
													assign node22415 = (inp[9]) ? node22417 : 4'b0000;
														assign node22417 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node22421 = (inp[12]) ? node22427 : node22422;
													assign node22422 = (inp[4]) ? node22424 : 4'b1000;
														assign node22424 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node22427 = (inp[1]) ? 4'b1100 : node22428;
														assign node22428 = (inp[2]) ? 4'b1100 : 4'b1000;
											assign node22432 = (inp[6]) ? node22438 : node22433;
												assign node22433 = (inp[1]) ? node22435 : 4'b1100;
													assign node22435 = (inp[2]) ? 4'b1000 : 4'b1100;
												assign node22438 = (inp[4]) ? node22442 : node22439;
													assign node22439 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node22442 = (inp[9]) ? 4'b0000 : 4'b0100;

endmodule