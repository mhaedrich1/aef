module dtc_split66_bm34 (
	input  wire [9-1:0] inp,
	output wire [5-1:0] outp
);

	wire [5-1:0] node1;
	wire [5-1:0] node2;
	wire [5-1:0] node3;
	wire [5-1:0] node4;
	wire [5-1:0] node5;
	wire [5-1:0] node6;
	wire [5-1:0] node9;
	wire [5-1:0] node12;
	wire [5-1:0] node13;
	wire [5-1:0] node16;
	wire [5-1:0] node19;
	wire [5-1:0] node20;
	wire [5-1:0] node21;
	wire [5-1:0] node24;
	wire [5-1:0] node27;
	wire [5-1:0] node28;
	wire [5-1:0] node31;
	wire [5-1:0] node34;
	wire [5-1:0] node35;
	wire [5-1:0] node36;
	wire [5-1:0] node37;
	wire [5-1:0] node40;
	wire [5-1:0] node43;
	wire [5-1:0] node44;
	wire [5-1:0] node47;
	wire [5-1:0] node50;
	wire [5-1:0] node51;
	wire [5-1:0] node52;
	wire [5-1:0] node55;
	wire [5-1:0] node58;
	wire [5-1:0] node59;
	wire [5-1:0] node62;
	wire [5-1:0] node65;
	wire [5-1:0] node66;
	wire [5-1:0] node67;
	wire [5-1:0] node68;
	wire [5-1:0] node69;
	wire [5-1:0] node72;
	wire [5-1:0] node76;
	wire [5-1:0] node77;
	wire [5-1:0] node78;
	wire [5-1:0] node81;
	wire [5-1:0] node84;
	wire [5-1:0] node86;
	wire [5-1:0] node89;
	wire [5-1:0] node90;
	wire [5-1:0] node91;
	wire [5-1:0] node92;
	wire [5-1:0] node95;
	wire [5-1:0] node98;
	wire [5-1:0] node99;
	wire [5-1:0] node102;
	wire [5-1:0] node105;
	wire [5-1:0] node106;
	wire [5-1:0] node107;
	wire [5-1:0] node110;
	wire [5-1:0] node113;
	wire [5-1:0] node114;
	wire [5-1:0] node117;
	wire [5-1:0] node120;
	wire [5-1:0] node121;
	wire [5-1:0] node122;
	wire [5-1:0] node123;
	wire [5-1:0] node124;
	wire [5-1:0] node125;
	wire [5-1:0] node128;
	wire [5-1:0] node131;
	wire [5-1:0] node132;
	wire [5-1:0] node135;
	wire [5-1:0] node138;
	wire [5-1:0] node139;
	wire [5-1:0] node140;
	wire [5-1:0] node143;
	wire [5-1:0] node146;
	wire [5-1:0] node147;
	wire [5-1:0] node150;
	wire [5-1:0] node153;
	wire [5-1:0] node154;
	wire [5-1:0] node156;
	wire [5-1:0] node157;
	wire [5-1:0] node160;
	wire [5-1:0] node163;
	wire [5-1:0] node164;
	wire [5-1:0] node166;
	wire [5-1:0] node169;
	wire [5-1:0] node170;
	wire [5-1:0] node173;
	wire [5-1:0] node176;
	wire [5-1:0] node177;
	wire [5-1:0] node178;
	wire [5-1:0] node179;
	wire [5-1:0] node180;
	wire [5-1:0] node183;
	wire [5-1:0] node186;
	wire [5-1:0] node187;
	wire [5-1:0] node190;
	wire [5-1:0] node193;
	wire [5-1:0] node194;
	wire [5-1:0] node195;
	wire [5-1:0] node198;
	wire [5-1:0] node201;
	wire [5-1:0] node202;
	wire [5-1:0] node205;
	wire [5-1:0] node208;
	wire [5-1:0] node209;
	wire [5-1:0] node210;
	wire [5-1:0] node211;
	wire [5-1:0] node214;
	wire [5-1:0] node217;
	wire [5-1:0] node218;
	wire [5-1:0] node221;
	wire [5-1:0] node224;
	wire [5-1:0] node225;
	wire [5-1:0] node226;
	wire [5-1:0] node229;
	wire [5-1:0] node232;
	wire [5-1:0] node233;
	wire [5-1:0] node236;

	assign outp = (inp[2]) ? node120 : node1;
		assign node1 = (inp[0]) ? node65 : node2;
			assign node2 = (inp[7]) ? node34 : node3;
				assign node3 = (inp[8]) ? node19 : node4;
					assign node4 = (inp[5]) ? node12 : node5;
						assign node5 = (inp[3]) ? node9 : node6;
							assign node6 = (inp[4]) ? 5'b01011 : 5'b00110;
							assign node9 = (inp[4]) ? 5'b00110 : 5'b10111;
						assign node12 = (inp[3]) ? node16 : node13;
							assign node13 = (inp[4]) ? 5'b00011 : 5'b11010;
							assign node16 = (inp[4]) ? 5'b11010 : 5'b01011;
					assign node19 = (inp[5]) ? node27 : node20;
						assign node20 = (inp[3]) ? node24 : node21;
							assign node21 = (inp[6]) ? 5'b11000 : 5'b01000;
							assign node24 = (inp[4]) ? 5'b10000 : 5'b10001;
						assign node27 = (inp[6]) ? node31 : node28;
							assign node28 = (inp[1]) ? 5'b11111 : 5'b00000;
							assign node31 = (inp[1]) ? 5'b01110 : 5'b11111;
				assign node34 = (inp[5]) ? node50 : node35;
					assign node35 = (inp[8]) ? node43 : node36;
						assign node36 = (inp[4]) ? node40 : node37;
							assign node37 = (inp[3]) ? 5'b01111 : 5'b01110;
							assign node40 = (inp[3]) ? 5'b10111 : 5'b00111;
						assign node43 = (inp[3]) ? node47 : node44;
							assign node44 = (inp[4]) ? 5'b01111 : 5'b00000;
							assign node47 = (inp[4]) ? 5'b01110 : 5'b01111;
					assign node50 = (inp[3]) ? node58 : node51;
						assign node51 = (inp[4]) ? node55 : node52;
							assign node52 = (inp[6]) ? 5'b00110 : 5'b11111;
							assign node55 = (inp[8]) ? 5'b10111 : 5'b11011;
						assign node58 = (inp[4]) ? node62 : node59;
							assign node59 = (inp[6]) ? 5'b00111 : 5'b10111;
							assign node62 = (inp[8]) ? 5'b10110 : 5'b00110;
			assign node65 = (inp[8]) ? node89 : node66;
				assign node66 = (inp[7]) ? node76 : node67;
					assign node67 = (inp[5]) ? 5'b00010 : node68;
						assign node68 = (inp[3]) ? node72 : node69;
							assign node69 = (inp[1]) ? 5'b00010 : 5'b00010;
							assign node72 = (inp[4]) ? 5'b00010 : 5'b10011;
					assign node76 = (inp[5]) ? node84 : node77;
						assign node77 = (inp[4]) ? node81 : node78;
							assign node78 = (inp[3]) ? 5'b11011 : 5'b01010;
							assign node81 = (inp[3]) ? 5'b01010 : 5'b00011;
						assign node84 = (inp[4]) ? node86 : 5'b00011;
							assign node86 = (inp[6]) ? 5'b00010 : 5'b00010;
				assign node89 = (inp[5]) ? node105 : node90;
					assign node90 = (inp[7]) ? node98 : node91;
						assign node91 = (inp[4]) ? node95 : node92;
							assign node92 = (inp[3]) ? 5'b00111 : 5'b01110;
							assign node95 = (inp[1]) ? 5'b10110 : 5'b00111;
						assign node98 = (inp[4]) ? node102 : node99;
							assign node99 = (inp[3]) ? 5'b11011 : 5'b00110;
							assign node102 = (inp[3]) ? 5'b01010 : 5'b11011;
					assign node105 = (inp[3]) ? node113 : node106;
						assign node106 = (inp[7]) ? node110 : node107;
							assign node107 = (inp[6]) ? 5'b00110 : 5'b00111;
							assign node110 = (inp[4]) ? 5'b00011 : 5'b11010;
						assign node113 = (inp[7]) ? node117 : node114;
							assign node114 = (inp[4]) ? 5'b01010 : 5'b11011;
							assign node117 = (inp[4]) ? 5'b00010 : 5'b00011;
		assign node120 = (inp[0]) ? node176 : node121;
			assign node121 = (inp[8]) ? node153 : node122;
				assign node122 = (inp[5]) ? node138 : node123;
					assign node123 = (inp[7]) ? node131 : node124;
						assign node124 = (inp[4]) ? node128 : node125;
							assign node125 = (inp[3]) ? 5'b00101 : 5'b00100;
							assign node128 = (inp[3]) ? 5'b00100 : 5'b11001;
						assign node131 = (inp[3]) ? node135 : node132;
							assign node132 = (inp[4]) ? 5'b00101 : 5'b01100;
							assign node135 = (inp[4]) ? 5'b01100 : 5'b01101;
					assign node138 = (inp[7]) ? node146 : node139;
						assign node139 = (inp[4]) ? node143 : node140;
							assign node140 = (inp[3]) ? 5'b01001 : 5'b01000;
							assign node143 = (inp[3]) ? 5'b10000 : 5'b00001;
						assign node146 = (inp[4]) ? node150 : node147;
							assign node147 = (inp[3]) ? 5'b00101 : 5'b00100;
							assign node150 = (inp[3]) ? 5'b10000 : 5'b01001;
				assign node153 = (inp[5]) ? node163 : node154;
					assign node154 = (inp[4]) ? node156 : 5'b11101;
						assign node156 = (inp[3]) ? node160 : node157;
							assign node157 = (inp[6]) ? 5'b11101 : 5'b11101;
							assign node160 = (inp[6]) ? 5'b01100 : 5'b01101;
					assign node163 = (inp[7]) ? node169 : node164;
						assign node164 = (inp[1]) ? node166 : 5'b11101;
							assign node166 = (inp[4]) ? 5'b11100 : 5'b11101;
						assign node169 = (inp[3]) ? node173 : node170;
							assign node170 = (inp[6]) ? 5'b10101 : 5'b01100;
							assign node173 = (inp[4]) ? 5'b00100 : 5'b00101;
			assign node176 = (inp[7]) ? node208 : node177;
				assign node177 = (inp[8]) ? node193 : node178;
					assign node178 = (inp[5]) ? node186 : node179;
						assign node179 = (inp[3]) ? node183 : node180;
							assign node180 = (inp[1]) ? 5'b11111 : 5'b00000;
							assign node183 = (inp[4]) ? 5'b00000 : 5'b00001;
						assign node186 = (inp[4]) ? node190 : node187;
							assign node187 = (inp[1]) ? 5'b01110 : 5'b01110;
							assign node190 = (inp[3]) ? 5'b00110 : 5'b00111;
					assign node193 = (inp[5]) ? node201 : node194;
						assign node194 = (inp[6]) ? node198 : node195;
							assign node195 = (inp[4]) ? 5'b00100 : 5'b01100;
							assign node198 = (inp[1]) ? 5'b00100 : 5'b10101;
						assign node201 = (inp[3]) ? node205 : node202;
							assign node202 = (inp[1]) ? 5'b01001 : 5'b00100;
							assign node205 = (inp[4]) ? 5'b01000 : 5'b11001;
				assign node208 = (inp[5]) ? node224 : node209;
					assign node209 = (inp[3]) ? node217 : node210;
						assign node210 = (inp[4]) ? node214 : node211;
							assign node211 = (inp[8]) ? 5'b00100 : 5'b01000;
							assign node214 = (inp[8]) ? 5'b11001 : 5'b10001;
						assign node217 = (inp[4]) ? node221 : node218;
							assign node218 = (inp[8]) ? 5'b11001 : 5'b01001;
							assign node221 = (inp[6]) ? 5'b01000 : 5'b01001;
					assign node224 = (inp[8]) ? node232 : node225;
						assign node225 = (inp[4]) ? node229 : node226;
							assign node226 = (inp[3]) ? 5'b10001 : 5'b00000;
							assign node229 = (inp[3]) ? 5'b00000 : 5'b11111;
						assign node232 = (inp[4]) ? node236 : node233;
							assign node233 = (inp[3]) ? 5'b00001 : 5'b11000;
							assign node236 = (inp[3]) ? 5'b00000 : 5'b00001;

endmodule