module dtc_split66_bm98 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node187;
	wire [3-1:0] node189;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node231;
	wire [3-1:0] node233;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node243;
	wire [3-1:0] node247;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node283;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node302;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node317;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node330;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node341;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node357;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node365;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node374;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node385;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node393;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node402;
	wire [3-1:0] node404;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node411;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node422;
	wire [3-1:0] node425;
	wire [3-1:0] node427;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node446;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node459;
	wire [3-1:0] node461;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node471;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node488;
	wire [3-1:0] node490;
	wire [3-1:0] node493;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node510;
	wire [3-1:0] node513;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node537;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node544;
	wire [3-1:0] node546;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node552;
	wire [3-1:0] node554;
	wire [3-1:0] node557;
	wire [3-1:0] node559;
	wire [3-1:0] node561;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node569;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node591;
	wire [3-1:0] node595;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node608;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node634;
	wire [3-1:0] node638;
	wire [3-1:0] node640;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node646;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node660;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node671;
	wire [3-1:0] node674;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node681;
	wire [3-1:0] node684;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node690;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node702;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node709;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node715;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node724;
	wire [3-1:0] node726;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node745;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node765;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node776;
	wire [3-1:0] node779;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node785;
	wire [3-1:0] node788;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node794;
	wire [3-1:0] node796;

	assign outp = (inp[0]) ? node288 : node1;
		assign node1 = (inp[6]) ? node3 : 3'b111;
			assign node3 = (inp[9]) ? node101 : node4;
				assign node4 = (inp[3]) ? node66 : node5;
					assign node5 = (inp[4]) ? node7 : 3'b100;
						assign node7 = (inp[1]) ? node41 : node8;
							assign node8 = (inp[7]) ? node10 : 3'b100;
								assign node10 = (inp[2]) ? node22 : node11;
									assign node11 = (inp[11]) ? node17 : node12;
										assign node12 = (inp[5]) ? node14 : 3'b000;
											assign node14 = (inp[10]) ? 3'b100 : 3'b000;
										assign node17 = (inp[5]) ? node19 : 3'b100;
											assign node19 = (inp[10]) ? 3'b000 : 3'b100;
									assign node22 = (inp[5]) ? node28 : node23;
										assign node23 = (inp[11]) ? node25 : 3'b100;
											assign node25 = (inp[10]) ? 3'b000 : 3'b100;
										assign node28 = (inp[8]) ? node34 : node29;
											assign node29 = (inp[11]) ? 3'b100 : node30;
												assign node30 = (inp[10]) ? 3'b000 : 3'b100;
											assign node34 = (inp[10]) ? node38 : node35;
												assign node35 = (inp[11]) ? 3'b000 : 3'b100;
												assign node38 = (inp[11]) ? 3'b100 : 3'b000;
							assign node41 = (inp[7]) ? node43 : 3'b000;
								assign node43 = (inp[2]) ? node53 : node44;
									assign node44 = (inp[10]) ? node46 : 3'b101;
										assign node46 = (inp[5]) ? node50 : node47;
											assign node47 = (inp[11]) ? 3'b100 : 3'b101;
											assign node50 = (inp[11]) ? 3'b101 : 3'b100;
									assign node53 = (inp[8]) ? node61 : node54;
										assign node54 = (inp[5]) ? node56 : 3'b100;
											assign node56 = (inp[10]) ? 3'b100 : node57;
												assign node57 = (inp[11]) ? 3'b101 : 3'b100;
										assign node61 = (inp[10]) ? 3'b101 : node62;
											assign node62 = (inp[5]) ? 3'b101 : 3'b100;
					assign node66 = (inp[1]) ? node68 : 3'b010;
						assign node68 = (inp[4]) ? node70 : 3'b010;
							assign node70 = (inp[7]) ? node72 : 3'b010;
								assign node72 = (inp[2]) ? node80 : node73;
									assign node73 = (inp[11]) ? node75 : 3'b110;
										assign node75 = (inp[5]) ? node77 : 3'b010;
											assign node77 = (inp[8]) ? 3'b110 : 3'b010;
									assign node80 = (inp[5]) ? node86 : node81;
										assign node81 = (inp[11]) ? node83 : 3'b010;
											assign node83 = (inp[10]) ? 3'b110 : 3'b010;
										assign node86 = (inp[8]) ? node94 : node87;
											assign node87 = (inp[10]) ? node91 : node88;
												assign node88 = (inp[11]) ? 3'b110 : 3'b010;
												assign node91 = (inp[11]) ? 3'b010 : 3'b110;
											assign node94 = (inp[11]) ? node98 : node95;
												assign node95 = (inp[10]) ? 3'b110 : 3'b010;
												assign node98 = (inp[10]) ? 3'b010 : 3'b110;
				assign node101 = (inp[3]) ? node247 : node102;
					assign node102 = (inp[1]) ? node172 : node103;
						assign node103 = (inp[4]) ? node125 : node104;
							assign node104 = (inp[2]) ? node114 : node105;
								assign node105 = (inp[7]) ? 3'b001 : node106;
									assign node106 = (inp[5]) ? node110 : node107;
										assign node107 = (inp[11]) ? 3'b101 : 3'b001;
										assign node110 = (inp[11]) ? 3'b001 : 3'b101;
								assign node114 = (inp[7]) ? 3'b101 : node115;
									assign node115 = (inp[10]) ? node117 : 3'b101;
										assign node117 = (inp[5]) ? node121 : node118;
											assign node118 = (inp[11]) ? 3'b101 : 3'b001;
											assign node121 = (inp[11]) ? 3'b001 : 3'b101;
							assign node125 = (inp[2]) ? node147 : node126;
								assign node126 = (inp[7]) ? node142 : node127;
									assign node127 = (inp[5]) ? node133 : node128;
										assign node128 = (inp[10]) ? node130 : 3'b101;
											assign node130 = (inp[11]) ? 3'b111 : 3'b101;
										assign node133 = (inp[8]) ? node137 : node134;
											assign node134 = (inp[11]) ? 3'b101 : 3'b111;
											assign node137 = (inp[10]) ? 3'b101 : node138;
												assign node138 = (inp[11]) ? 3'b111 : 3'b101;
									assign node142 = (inp[5]) ? node144 : 3'b111;
										assign node144 = (inp[11]) ? 3'b011 : 3'b111;
								assign node147 = (inp[7]) ? node161 : node148;
									assign node148 = (inp[5]) ? node154 : node149;
										assign node149 = (inp[11]) ? 3'b111 : node150;
											assign node150 = (inp[10]) ? 3'b011 : 3'b111;
										assign node154 = (inp[8]) ? node156 : 3'b011;
											assign node156 = (inp[10]) ? node158 : 3'b101;
												assign node158 = (inp[11]) ? 3'b011 : 3'b001;
									assign node161 = (inp[10]) ? node163 : 3'b101;
										assign node163 = (inp[8]) ? node165 : 3'b001;
											assign node165 = (inp[11]) ? node169 : node166;
												assign node166 = (inp[5]) ? 3'b001 : 3'b101;
												assign node169 = (inp[5]) ? 3'b101 : 3'b001;
						assign node172 = (inp[4]) ? node202 : node173;
							assign node173 = (inp[2]) ? node193 : node174;
								assign node174 = (inp[7]) ? 3'b001 : node175;
									assign node175 = (inp[8]) ? node181 : node176;
										assign node176 = (inp[11]) ? node178 : 3'b100;
											assign node178 = (inp[5]) ? 3'b001 : 3'b100;
										assign node181 = (inp[10]) ? node187 : node182;
											assign node182 = (inp[11]) ? 3'b100 : node183;
												assign node183 = (inp[5]) ? 3'b100 : 3'b001;
											assign node187 = (inp[11]) ? node189 : 3'b001;
												assign node189 = (inp[5]) ? 3'b001 : 3'b100;
								assign node193 = (inp[7]) ? 3'b100 : node194;
									assign node194 = (inp[5]) ? node198 : node195;
										assign node195 = (inp[11]) ? 3'b100 : 3'b001;
										assign node198 = (inp[11]) ? 3'b001 : 3'b100;
							assign node202 = (inp[2]) ? node224 : node203;
								assign node203 = (inp[7]) ? node215 : node204;
									assign node204 = (inp[5]) ? node210 : node205;
										assign node205 = (inp[8]) ? 3'b100 : node206;
											assign node206 = (inp[11]) ? 3'b100 : 3'b110;
										assign node210 = (inp[8]) ? 3'b110 : node211;
											assign node211 = (inp[11]) ? 3'b100 : 3'b110;
									assign node215 = (inp[10]) ? 3'b110 : node216;
										assign node216 = (inp[5]) ? node220 : node217;
											assign node217 = (inp[11]) ? 3'b110 : 3'b001;
											assign node220 = (inp[11]) ? 3'b001 : 3'b110;
								assign node224 = (inp[11]) ? node236 : node225;
									assign node225 = (inp[8]) ? node231 : node226;
										assign node226 = (inp[7]) ? 3'b001 : node227;
											assign node227 = (inp[10]) ? 3'b100 : 3'b001;
										assign node231 = (inp[10]) ? node233 : 3'b110;
											assign node233 = (inp[5]) ? 3'b001 : 3'b011;
									assign node236 = (inp[7]) ? 3'b110 : node237;
										assign node237 = (inp[8]) ? node239 : 3'b011;
											assign node239 = (inp[10]) ? node243 : node240;
												assign node240 = (inp[5]) ? 3'b100 : 3'b110;
												assign node243 = (inp[5]) ? 3'b011 : 3'b001;
					assign node247 = (inp[1]) ? node249 : 3'b111;
						assign node249 = (inp[7]) ? node267 : node250;
							assign node250 = (inp[4]) ? node258 : node251;
								assign node251 = (inp[5]) ? node255 : node252;
									assign node252 = (inp[11]) ? 3'b011 : 3'b111;
									assign node255 = (inp[11]) ? 3'b111 : 3'b011;
								assign node258 = (inp[2]) ? node260 : 3'b001;
									assign node260 = (inp[8]) ? node264 : node261;
										assign node261 = (inp[10]) ? 3'b001 : 3'b111;
										assign node264 = (inp[10]) ? 3'b111 : 3'b011;
							assign node267 = (inp[4]) ? node271 : node268;
								assign node268 = (inp[2]) ? 3'b001 : 3'b101;
								assign node271 = (inp[2]) ? node279 : node272;
									assign node272 = (inp[11]) ? node276 : node273;
										assign node273 = (inp[5]) ? 3'b011 : 3'b111;
										assign node276 = (inp[5]) ? 3'b111 : 3'b011;
									assign node279 = (inp[11]) ? node283 : node280;
										assign node280 = (inp[10]) ? 3'b101 : 3'b001;
										assign node283 = (inp[8]) ? node285 : 3'b011;
											assign node285 = (inp[10]) ? 3'b011 : 3'b101;
		assign node288 = (inp[3]) ? node474 : node289;
			assign node289 = (inp[6]) ? node425 : node290;
				assign node290 = (inp[9]) ? node334 : node291;
					assign node291 = (inp[4]) ? node293 : 3'b010;
						assign node293 = (inp[7]) ? node297 : node294;
							assign node294 = (inp[1]) ? 3'b000 : 3'b010;
							assign node297 = (inp[1]) ? 3'b010 : node298;
								assign node298 = (inp[2]) ? node314 : node299;
									assign node299 = (inp[11]) ? node305 : node300;
										assign node300 = (inp[5]) ? node302 : 3'b000;
											assign node302 = (inp[10]) ? 3'b010 : 3'b000;
										assign node305 = (inp[8]) ? 3'b010 : node306;
											assign node306 = (inp[10]) ? node310 : node307;
												assign node307 = (inp[5]) ? 3'b010 : 3'b000;
												assign node310 = (inp[5]) ? 3'b000 : 3'b010;
									assign node314 = (inp[5]) ? node320 : node315;
										assign node315 = (inp[11]) ? node317 : 3'b010;
											assign node317 = (inp[10]) ? 3'b000 : 3'b010;
										assign node320 = (inp[8]) ? node326 : node321;
											assign node321 = (inp[10]) ? node323 : 3'b010;
												assign node323 = (inp[11]) ? 3'b010 : 3'b000;
											assign node326 = (inp[11]) ? node330 : node327;
												assign node327 = (inp[10]) ? 3'b000 : 3'b010;
												assign node330 = (inp[10]) ? 3'b010 : 3'b000;
					assign node334 = (inp[4]) ? node378 : node335;
						assign node335 = (inp[2]) ? node345 : node336;
							assign node336 = (inp[7]) ? 3'b000 : node337;
								assign node337 = (inp[5]) ? node341 : node338;
									assign node338 = (inp[11]) ? 3'b010 : 3'b000;
									assign node341 = (inp[11]) ? 3'b000 : 3'b010;
							assign node345 = (inp[7]) ? 3'b010 : node346;
								assign node346 = (inp[1]) ? node360 : node347;
									assign node347 = (inp[10]) ? node353 : node348;
										assign node348 = (inp[5]) ? 3'b000 : node349;
											assign node349 = (inp[11]) ? 3'b010 : 3'b000;
										assign node353 = (inp[11]) ? node357 : node354;
											assign node354 = (inp[5]) ? 3'b010 : 3'b000;
											assign node357 = (inp[5]) ? 3'b000 : 3'b010;
									assign node360 = (inp[10]) ? node370 : node361;
										assign node361 = (inp[8]) ? node365 : node362;
											assign node362 = (inp[11]) ? 3'b010 : 3'b000;
											assign node365 = (inp[5]) ? node367 : 3'b010;
												assign node367 = (inp[11]) ? 3'b000 : 3'b010;
										assign node370 = (inp[11]) ? node374 : node371;
											assign node371 = (inp[5]) ? 3'b010 : 3'b000;
											assign node374 = (inp[5]) ? 3'b000 : 3'b010;
						assign node378 = (inp[2]) ? node388 : node379;
							assign node379 = (inp[7]) ? node381 : 3'b010;
								assign node381 = (inp[5]) ? node385 : node382;
									assign node382 = (inp[11]) ? 3'b010 : 3'b000;
									assign node385 = (inp[11]) ? 3'b000 : 3'b010;
							assign node388 = (inp[7]) ? node396 : node389;
								assign node389 = (inp[10]) ? node393 : node390;
									assign node390 = (inp[8]) ? 3'b010 : 3'b000;
									assign node393 = (inp[8]) ? 3'b000 : 3'b010;
								assign node396 = (inp[1]) ? node408 : node397;
									assign node397 = (inp[5]) ? 3'b010 : node398;
										assign node398 = (inp[8]) ? node402 : node399;
											assign node399 = (inp[11]) ? 3'b010 : 3'b000;
											assign node402 = (inp[10]) ? node404 : 3'b010;
												assign node404 = (inp[11]) ? 3'b000 : 3'b010;
									assign node408 = (inp[11]) ? node416 : node409;
										assign node409 = (inp[8]) ? node411 : 3'b100;
											assign node411 = (inp[5]) ? node413 : 3'b010;
												assign node413 = (inp[10]) ? 3'b100 : 3'b110;
										assign node416 = (inp[8]) ? node418 : 3'b110;
											assign node418 = (inp[5]) ? node422 : node419;
												assign node419 = (inp[10]) ? 3'b100 : 3'b110;
												assign node422 = (inp[10]) ? 3'b010 : 3'b000;
				assign node425 = (inp[4]) ? node427 : 3'b000;
					assign node427 = (inp[9]) ? node429 : 3'b000;
						assign node429 = (inp[1]) ? node471 : node430;
							assign node430 = (inp[11]) ? node454 : node431;
								assign node431 = (inp[8]) ? node437 : node432;
									assign node432 = (inp[2]) ? 3'b010 : node433;
										assign node433 = (inp[5]) ? 3'b100 : 3'b010;
									assign node437 = (inp[10]) ? node443 : node438;
										assign node438 = (inp[5]) ? 3'b110 : node439;
											assign node439 = (inp[2]) ? 3'b110 : 3'b010;
										assign node443 = (inp[7]) ? node449 : node444;
											assign node444 = (inp[2]) ? node446 : 3'b100;
												assign node446 = (inp[5]) ? 3'b010 : 3'b110;
											assign node449 = (inp[5]) ? 3'b010 : node450;
												assign node450 = (inp[2]) ? 3'b110 : 3'b010;
								assign node454 = (inp[5]) ? node464 : node455;
									assign node455 = (inp[10]) ? node459 : node456;
										assign node456 = (inp[2]) ? 3'b100 : 3'b110;
										assign node459 = (inp[2]) ? node461 : 3'b100;
											assign node461 = (inp[8]) ? 3'b000 : 3'b100;
									assign node464 = (inp[10]) ? 3'b010 : node465;
										assign node465 = (inp[8]) ? 3'b000 : node466;
											assign node466 = (inp[2]) ? 3'b100 : 3'b000;
							assign node471 = (inp[7]) ? 3'b000 : 3'b100;
			assign node474 = (inp[9]) ? node582 : node475;
				assign node475 = (inp[4]) ? node481 : node476;
					assign node476 = (inp[1]) ? 3'b000 : node477;
						assign node477 = (inp[6]) ? 3'b000 : 3'b001;
					assign node481 = (inp[1]) ? node531 : node482;
						assign node482 = (inp[7]) ? node502 : node483;
							assign node483 = (inp[6]) ? 3'b001 : node484;
								assign node484 = (inp[2]) ? node496 : node485;
									assign node485 = (inp[11]) ? node493 : node486;
										assign node486 = (inp[8]) ? node488 : 3'b111;
											assign node488 = (inp[10]) ? node490 : 3'b011;
												assign node490 = (inp[5]) ? 3'b111 : 3'b011;
										assign node493 = (inp[8]) ? 3'b111 : 3'b011;
									assign node496 = (inp[11]) ? 3'b101 : node497;
										assign node497 = (inp[8]) ? 3'b101 : 3'b011;
							assign node502 = (inp[6]) ? node506 : node503;
								assign node503 = (inp[2]) ? 3'b001 : 3'b101;
								assign node506 = (inp[11]) ? node516 : node507;
									assign node507 = (inp[2]) ? node513 : node508;
										assign node508 = (inp[5]) ? node510 : 3'b100;
											assign node510 = (inp[10]) ? 3'b010 : 3'b100;
										assign node513 = (inp[5]) ? 3'b100 : 3'b000;
									assign node516 = (inp[2]) ? node524 : node517;
										assign node517 = (inp[5]) ? node521 : node518;
											assign node518 = (inp[10]) ? 3'b010 : 3'b100;
											assign node521 = (inp[10]) ? 3'b100 : 3'b010;
										assign node524 = (inp[10]) ? node528 : node525;
											assign node525 = (inp[5]) ? 3'b110 : 3'b010;
											assign node528 = (inp[5]) ? 3'b010 : 3'b110;
						assign node531 = (inp[6]) ? node579 : node532;
							assign node532 = (inp[7]) ? node564 : node533;
								assign node533 = (inp[2]) ? node549 : node534;
									assign node534 = (inp[5]) ? node540 : node535;
										assign node535 = (inp[10]) ? node537 : 3'b001;
											assign node537 = (inp[11]) ? 3'b101 : 3'b001;
										assign node540 = (inp[11]) ? node544 : node541;
											assign node541 = (inp[8]) ? 3'b001 : 3'b101;
											assign node544 = (inp[8]) ? node546 : 3'b001;
												assign node546 = (inp[10]) ? 3'b001 : 3'b101;
									assign node549 = (inp[11]) ? node557 : node550;
										assign node550 = (inp[8]) ? node552 : 3'b001;
											assign node552 = (inp[5]) ? node554 : 3'b110;
												assign node554 = (inp[10]) ? 3'b001 : 3'b110;
										assign node557 = (inp[8]) ? node559 : 3'b110;
											assign node559 = (inp[5]) ? node561 : 3'b001;
												assign node561 = (inp[10]) ? 3'b110 : 3'b001;
								assign node564 = (inp[11]) ? node574 : node565;
									assign node565 = (inp[10]) ? 3'b010 : node566;
										assign node566 = (inp[5]) ? 3'b110 : node567;
											assign node567 = (inp[8]) ? node569 : 3'b010;
												assign node569 = (inp[2]) ? 3'b100 : 3'b010;
									assign node574 = (inp[2]) ? 3'b100 : node575;
										assign node575 = (inp[5]) ? 3'b010 : 3'b110;
							assign node579 = (inp[7]) ? 3'b000 : 3'b100;
				assign node582 = (inp[6]) ? node664 : node583;
					assign node583 = (inp[1]) ? node585 : 3'b111;
						assign node585 = (inp[4]) ? node627 : node586;
							assign node586 = (inp[11]) ? node602 : node587;
								assign node587 = (inp[8]) ? node595 : node588;
									assign node588 = (inp[2]) ? 3'b110 : node589;
										assign node589 = (inp[7]) ? node591 : 3'b010;
											assign node591 = (inp[5]) ? 3'b010 : 3'b110;
									assign node595 = (inp[10]) ? node597 : 3'b001;
										assign node597 = (inp[5]) ? 3'b010 : node598;
											assign node598 = (inp[7]) ? 3'b101 : 3'b001;
								assign node602 = (inp[8]) ? node614 : node603;
									assign node603 = (inp[5]) ? node605 : 3'b001;
										assign node605 = (inp[7]) ? node611 : node606;
											assign node606 = (inp[2]) ? node608 : 3'b001;
												assign node608 = (inp[10]) ? 3'b001 : 3'b101;
											assign node611 = (inp[2]) ? 3'b001 : 3'b101;
									assign node614 = (inp[10]) ? node618 : node615;
										assign node615 = (inp[5]) ? 3'b010 : 3'b001;
										assign node618 = (inp[5]) ? node622 : node619;
											assign node619 = (inp[2]) ? 3'b110 : 3'b010;
											assign node622 = (inp[2]) ? 3'b001 : node623;
												assign node623 = (inp[7]) ? 3'b101 : 3'b001;
							assign node627 = (inp[7]) ? node649 : node628;
								assign node628 = (inp[11]) ? node638 : node629;
									assign node629 = (inp[8]) ? node631 : 3'b011;
										assign node631 = (inp[2]) ? 3'b111 : node632;
											assign node632 = (inp[5]) ? node634 : 3'b111;
												assign node634 = (inp[10]) ? 3'b011 : 3'b111;
									assign node638 = (inp[2]) ? node640 : 3'b111;
										assign node640 = (inp[8]) ? node642 : 3'b111;
											assign node642 = (inp[10]) ? node646 : node643;
												assign node643 = (inp[5]) ? 3'b011 : 3'b111;
												assign node646 = (inp[5]) ? 3'b111 : 3'b011;
								assign node649 = (inp[2]) ? node655 : node650;
									assign node650 = (inp[8]) ? 3'b001 : node651;
										assign node651 = (inp[11]) ? 3'b001 : 3'b011;
									assign node655 = (inp[8]) ? 3'b101 : node656;
										assign node656 = (inp[11]) ? node660 : node657;
											assign node657 = (inp[5]) ? 3'b101 : 3'b011;
											assign node660 = (inp[5]) ? 3'b011 : 3'b101;
					assign node664 = (inp[1]) ? node718 : node665;
						assign node665 = (inp[7]) ? node693 : node666;
							assign node666 = (inp[4]) ? node684 : node667;
								assign node667 = (inp[8]) ? node677 : node668;
									assign node668 = (inp[10]) ? node674 : node669;
										assign node669 = (inp[2]) ? node671 : 3'b001;
											assign node671 = (inp[5]) ? 3'b101 : 3'b001;
										assign node674 = (inp[5]) ? 3'b001 : 3'b101;
									assign node677 = (inp[5]) ? node681 : node678;
										assign node678 = (inp[11]) ? 3'b001 : 3'b101;
										assign node681 = (inp[11]) ? 3'b101 : 3'b001;
								assign node684 = (inp[2]) ? node686 : 3'b010;
									assign node686 = (inp[8]) ? node690 : node687;
										assign node687 = (inp[10]) ? 3'b010 : 3'b101;
										assign node690 = (inp[10]) ? 3'b101 : 3'b001;
							assign node693 = (inp[4]) ? node697 : node694;
								assign node694 = (inp[2]) ? 3'b010 : 3'b110;
								assign node697 = (inp[2]) ? node705 : node698;
									assign node698 = (inp[5]) ? node702 : node699;
										assign node699 = (inp[11]) ? 3'b001 : 3'b101;
										assign node702 = (inp[11]) ? 3'b101 : 3'b001;
									assign node705 = (inp[11]) ? node709 : node706;
										assign node706 = (inp[8]) ? 3'b010 : 3'b110;
										assign node709 = (inp[8]) ? node711 : 3'b001;
											assign node711 = (inp[5]) ? node715 : node712;
												assign node712 = (inp[10]) ? 3'b110 : 3'b010;
												assign node715 = (inp[10]) ? 3'b001 : 3'b110;
						assign node718 = (inp[7]) ? node768 : node719;
							assign node719 = (inp[4]) ? node755 : node720;
								assign node720 = (inp[2]) ? node736 : node721;
									assign node721 = (inp[8]) ? node729 : node722;
										assign node722 = (inp[10]) ? node724 : 3'b110;
											assign node724 = (inp[5]) ? node726 : 3'b110;
												assign node726 = (inp[11]) ? 3'b110 : 3'b010;
										assign node729 = (inp[10]) ? 3'b110 : node730;
											assign node730 = (inp[5]) ? 3'b010 : node731;
												assign node731 = (inp[11]) ? 3'b010 : 3'b110;
									assign node736 = (inp[8]) ? node742 : node737;
										assign node737 = (inp[5]) ? 3'b010 : node738;
											assign node738 = (inp[11]) ? 3'b010 : 3'b110;
										assign node742 = (inp[10]) ? node748 : node743;
											assign node743 = (inp[5]) ? node745 : 3'b110;
												assign node745 = (inp[11]) ? 3'b110 : 3'b010;
											assign node748 = (inp[11]) ? node752 : node749;
												assign node749 = (inp[5]) ? 3'b010 : 3'b110;
												assign node752 = (inp[5]) ? 3'b110 : 3'b010;
								assign node755 = (inp[2]) ? node761 : node756;
									assign node756 = (inp[8]) ? 3'b000 : node757;
										assign node757 = (inp[10]) ? 3'b001 : 3'b000;
									assign node761 = (inp[10]) ? node765 : node762;
										assign node762 = (inp[8]) ? 3'b010 : 3'b110;
										assign node765 = (inp[8]) ? 3'b110 : 3'b001;
							assign node768 = (inp[4]) ? node772 : node769;
								assign node769 = (inp[2]) ? 3'b000 : 3'b100;
								assign node772 = (inp[2]) ? node788 : node773;
									assign node773 = (inp[8]) ? node779 : node774;
										assign node774 = (inp[5]) ? node776 : 3'b010;
											assign node776 = (inp[11]) ? 3'b110 : 3'b010;
										assign node779 = (inp[10]) ? node781 : 3'b110;
											assign node781 = (inp[5]) ? node785 : node782;
												assign node782 = (inp[11]) ? 3'b010 : 3'b110;
												assign node785 = (inp[11]) ? 3'b110 : 3'b010;
									assign node788 = (inp[11]) ? node794 : node789;
										assign node789 = (inp[10]) ? 3'b100 : node790;
											assign node790 = (inp[8]) ? 3'b000 : 3'b100;
										assign node794 = (inp[8]) ? node796 : 3'b010;
											assign node796 = (inp[10]) ? 3'b010 : 3'b100;

endmodule