module dtc_split875_bm62 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node15;
	wire [4-1:0] node18;
	wire [4-1:0] node20;
	wire [4-1:0] node23;
	wire [4-1:0] node24;
	wire [4-1:0] node26;
	wire [4-1:0] node29;
	wire [4-1:0] node31;
	wire [4-1:0] node34;
	wire [4-1:0] node35;
	wire [4-1:0] node36;
	wire [4-1:0] node39;
	wire [4-1:0] node42;
	wire [4-1:0] node43;
	wire [4-1:0] node44;
	wire [4-1:0] node47;
	wire [4-1:0] node50;
	wire [4-1:0] node51;
	wire [4-1:0] node54;
	wire [4-1:0] node57;
	wire [4-1:0] node58;
	wire [4-1:0] node59;
	wire [4-1:0] node61;
	wire [4-1:0] node64;
	wire [4-1:0] node66;
	wire [4-1:0] node69;
	wire [4-1:0] node70;
	wire [4-1:0] node72;
	wire [4-1:0] node75;
	wire [4-1:0] node77;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node82;
	wire [4-1:0] node83;
	wire [4-1:0] node84;
	wire [4-1:0] node86;
	wire [4-1:0] node89;
	wire [4-1:0] node91;
	wire [4-1:0] node94;
	wire [4-1:0] node95;
	wire [4-1:0] node97;
	wire [4-1:0] node101;
	wire [4-1:0] node102;
	wire [4-1:0] node103;
	wire [4-1:0] node104;
	wire [4-1:0] node107;
	wire [4-1:0] node110;
	wire [4-1:0] node111;
	wire [4-1:0] node115;
	wire [4-1:0] node116;
	wire [4-1:0] node117;
	wire [4-1:0] node120;
	wire [4-1:0] node123;
	wire [4-1:0] node124;
	wire [4-1:0] node128;
	wire [4-1:0] node129;
	wire [4-1:0] node130;
	wire [4-1:0] node131;
	wire [4-1:0] node132;
	wire [4-1:0] node135;
	wire [4-1:0] node138;
	wire [4-1:0] node139;
	wire [4-1:0] node143;
	wire [4-1:0] node144;
	wire [4-1:0] node145;
	wire [4-1:0] node148;
	wire [4-1:0] node151;
	wire [4-1:0] node152;
	wire [4-1:0] node156;
	wire [4-1:0] node157;
	wire [4-1:0] node158;
	wire [4-1:0] node159;
	wire [4-1:0] node163;
	wire [4-1:0] node164;
	wire [4-1:0] node168;
	wire [4-1:0] node169;
	wire [4-1:0] node170;
	wire [4-1:0] node174;
	wire [4-1:0] node175;
	wire [4-1:0] node179;
	wire [4-1:0] node180;
	wire [4-1:0] node181;
	wire [4-1:0] node182;
	wire [4-1:0] node183;
	wire [4-1:0] node184;
	wire [4-1:0] node186;
	wire [4-1:0] node189;
	wire [4-1:0] node191;
	wire [4-1:0] node194;
	wire [4-1:0] node195;
	wire [4-1:0] node197;
	wire [4-1:0] node200;
	wire [4-1:0] node202;
	wire [4-1:0] node205;
	wire [4-1:0] node206;
	wire [4-1:0] node207;
	wire [4-1:0] node208;
	wire [4-1:0] node211;
	wire [4-1:0] node214;
	wire [4-1:0] node215;
	wire [4-1:0] node218;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node223;
	wire [4-1:0] node226;
	wire [4-1:0] node229;
	wire [4-1:0] node230;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node236;
	wire [4-1:0] node237;
	wire [4-1:0] node238;
	wire [4-1:0] node241;
	wire [4-1:0] node244;
	wire [4-1:0] node245;
	wire [4-1:0] node248;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node253;
	wire [4-1:0] node256;
	wire [4-1:0] node259;
	wire [4-1:0] node261;
	wire [4-1:0] node264;
	wire [4-1:0] node265;
	wire [4-1:0] node266;
	wire [4-1:0] node269;
	wire [4-1:0] node272;
	wire [4-1:0] node273;
	wire [4-1:0] node274;
	wire [4-1:0] node277;
	wire [4-1:0] node280;
	wire [4-1:0] node281;
	wire [4-1:0] node284;
	wire [4-1:0] node287;
	wire [4-1:0] node288;
	wire [4-1:0] node289;
	wire [4-1:0] node290;
	wire [4-1:0] node291;
	wire [4-1:0] node292;
	wire [4-1:0] node295;
	wire [4-1:0] node298;
	wire [4-1:0] node299;
	wire [4-1:0] node302;
	wire [4-1:0] node305;
	wire [4-1:0] node306;
	wire [4-1:0] node307;
	wire [4-1:0] node310;
	wire [4-1:0] node313;
	wire [4-1:0] node314;
	wire [4-1:0] node317;
	wire [4-1:0] node320;
	wire [4-1:0] node321;
	wire [4-1:0] node322;
	wire [4-1:0] node323;
	wire [4-1:0] node326;
	wire [4-1:0] node329;
	wire [4-1:0] node330;
	wire [4-1:0] node333;
	wire [4-1:0] node336;
	wire [4-1:0] node337;
	wire [4-1:0] node340;
	wire [4-1:0] node343;
	wire [4-1:0] node344;
	wire [4-1:0] node345;
	wire [4-1:0] node346;
	wire [4-1:0] node347;
	wire [4-1:0] node350;
	wire [4-1:0] node353;
	wire [4-1:0] node354;
	wire [4-1:0] node357;
	wire [4-1:0] node360;
	wire [4-1:0] node361;
	wire [4-1:0] node362;
	wire [4-1:0] node365;
	wire [4-1:0] node368;
	wire [4-1:0] node369;
	wire [4-1:0] node372;
	wire [4-1:0] node375;
	wire [4-1:0] node376;
	wire [4-1:0] node377;
	wire [4-1:0] node378;
	wire [4-1:0] node381;
	wire [4-1:0] node384;
	wire [4-1:0] node386;
	wire [4-1:0] node389;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node394;
	wire [4-1:0] node397;
	wire [4-1:0] node398;
	wire [4-1:0] node401;
	wire [4-1:0] node404;
	wire [4-1:0] node405;
	wire [4-1:0] node406;
	wire [4-1:0] node407;
	wire [4-1:0] node408;
	wire [4-1:0] node409;
	wire [4-1:0] node410;
	wire [4-1:0] node411;
	wire [4-1:0] node414;
	wire [4-1:0] node417;
	wire [4-1:0] node418;
	wire [4-1:0] node421;
	wire [4-1:0] node424;
	wire [4-1:0] node425;
	wire [4-1:0] node426;
	wire [4-1:0] node429;
	wire [4-1:0] node432;
	wire [4-1:0] node433;
	wire [4-1:0] node436;
	wire [4-1:0] node439;
	wire [4-1:0] node440;
	wire [4-1:0] node441;
	wire [4-1:0] node442;
	wire [4-1:0] node445;
	wire [4-1:0] node448;
	wire [4-1:0] node449;
	wire [4-1:0] node453;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node459;
	wire [4-1:0] node460;
	wire [4-1:0] node463;
	wire [4-1:0] node466;
	wire [4-1:0] node467;
	wire [4-1:0] node468;
	wire [4-1:0] node469;
	wire [4-1:0] node470;
	wire [4-1:0] node473;
	wire [4-1:0] node476;
	wire [4-1:0] node477;
	wire [4-1:0] node480;
	wire [4-1:0] node483;
	wire [4-1:0] node484;
	wire [4-1:0] node485;
	wire [4-1:0] node488;
	wire [4-1:0] node491;
	wire [4-1:0] node494;
	wire [4-1:0] node495;
	wire [4-1:0] node496;
	wire [4-1:0] node497;
	wire [4-1:0] node500;
	wire [4-1:0] node503;
	wire [4-1:0] node504;
	wire [4-1:0] node507;
	wire [4-1:0] node510;
	wire [4-1:0] node511;
	wire [4-1:0] node513;
	wire [4-1:0] node516;
	wire [4-1:0] node517;
	wire [4-1:0] node520;
	wire [4-1:0] node523;
	wire [4-1:0] node524;
	wire [4-1:0] node525;
	wire [4-1:0] node526;
	wire [4-1:0] node527;
	wire [4-1:0] node528;
	wire [4-1:0] node531;
	wire [4-1:0] node534;
	wire [4-1:0] node535;
	wire [4-1:0] node538;
	wire [4-1:0] node541;
	wire [4-1:0] node542;
	wire [4-1:0] node544;
	wire [4-1:0] node547;
	wire [4-1:0] node549;
	wire [4-1:0] node552;
	wire [4-1:0] node553;
	wire [4-1:0] node554;
	wire [4-1:0] node556;
	wire [4-1:0] node559;
	wire [4-1:0] node561;
	wire [4-1:0] node564;
	wire [4-1:0] node565;
	wire [4-1:0] node566;
	wire [4-1:0] node570;
	wire [4-1:0] node571;
	wire [4-1:0] node575;
	wire [4-1:0] node576;
	wire [4-1:0] node577;
	wire [4-1:0] node578;
	wire [4-1:0] node579;
	wire [4-1:0] node582;
	wire [4-1:0] node585;
	wire [4-1:0] node586;
	wire [4-1:0] node589;
	wire [4-1:0] node592;
	wire [4-1:0] node593;
	wire [4-1:0] node594;
	wire [4-1:0] node598;
	wire [4-1:0] node599;
	wire [4-1:0] node603;
	wire [4-1:0] node604;
	wire [4-1:0] node605;
	wire [4-1:0] node606;
	wire [4-1:0] node610;
	wire [4-1:0] node611;
	wire [4-1:0] node615;
	wire [4-1:0] node616;
	wire [4-1:0] node617;
	wire [4-1:0] node622;
	wire [4-1:0] node623;
	wire [4-1:0] node624;
	wire [4-1:0] node625;
	wire [4-1:0] node626;
	wire [4-1:0] node627;
	wire [4-1:0] node628;
	wire [4-1:0] node631;
	wire [4-1:0] node634;
	wire [4-1:0] node635;
	wire [4-1:0] node638;
	wire [4-1:0] node641;
	wire [4-1:0] node642;
	wire [4-1:0] node643;
	wire [4-1:0] node646;
	wire [4-1:0] node649;
	wire [4-1:0] node650;
	wire [4-1:0] node653;
	wire [4-1:0] node656;
	wire [4-1:0] node657;
	wire [4-1:0] node658;
	wire [4-1:0] node660;
	wire [4-1:0] node663;
	wire [4-1:0] node665;
	wire [4-1:0] node668;
	wire [4-1:0] node669;
	wire [4-1:0] node671;
	wire [4-1:0] node674;
	wire [4-1:0] node676;
	wire [4-1:0] node679;
	wire [4-1:0] node680;
	wire [4-1:0] node681;
	wire [4-1:0] node682;
	wire [4-1:0] node684;
	wire [4-1:0] node687;
	wire [4-1:0] node688;
	wire [4-1:0] node691;
	wire [4-1:0] node694;
	wire [4-1:0] node695;
	wire [4-1:0] node696;
	wire [4-1:0] node700;
	wire [4-1:0] node701;
	wire [4-1:0] node705;
	wire [4-1:0] node706;
	wire [4-1:0] node707;
	wire [4-1:0] node708;
	wire [4-1:0] node711;
	wire [4-1:0] node714;
	wire [4-1:0] node716;
	wire [4-1:0] node719;
	wire [4-1:0] node720;
	wire [4-1:0] node723;
	wire [4-1:0] node726;
	wire [4-1:0] node727;
	wire [4-1:0] node728;
	wire [4-1:0] node729;
	wire [4-1:0] node730;
	wire [4-1:0] node731;
	wire [4-1:0] node734;
	wire [4-1:0] node737;
	wire [4-1:0] node738;
	wire [4-1:0] node741;
	wire [4-1:0] node744;
	wire [4-1:0] node745;
	wire [4-1:0] node746;
	wire [4-1:0] node750;
	wire [4-1:0] node751;
	wire [4-1:0] node754;
	wire [4-1:0] node757;
	wire [4-1:0] node758;
	wire [4-1:0] node759;
	wire [4-1:0] node760;
	wire [4-1:0] node765;
	wire [4-1:0] node766;
	wire [4-1:0] node769;
	wire [4-1:0] node770;
	wire [4-1:0] node774;
	wire [4-1:0] node775;
	wire [4-1:0] node776;
	wire [4-1:0] node777;
	wire [4-1:0] node778;
	wire [4-1:0] node781;
	wire [4-1:0] node784;
	wire [4-1:0] node785;
	wire [4-1:0] node789;
	wire [4-1:0] node790;
	wire [4-1:0] node792;
	wire [4-1:0] node795;
	wire [4-1:0] node796;
	wire [4-1:0] node799;
	wire [4-1:0] node802;
	wire [4-1:0] node803;
	wire [4-1:0] node804;
	wire [4-1:0] node805;
	wire [4-1:0] node808;
	wire [4-1:0] node811;
	wire [4-1:0] node812;
	wire [4-1:0] node815;
	wire [4-1:0] node818;
	wire [4-1:0] node819;
	wire [4-1:0] node820;
	wire [4-1:0] node823;
	wire [4-1:0] node826;
	wire [4-1:0] node827;
	wire [4-1:0] node830;
	wire [4-1:0] node833;
	wire [4-1:0] node834;
	wire [4-1:0] node835;
	wire [4-1:0] node836;
	wire [4-1:0] node837;
	wire [4-1:0] node838;
	wire [4-1:0] node839;
	wire [4-1:0] node840;
	wire [4-1:0] node841;
	wire [4-1:0] node844;
	wire [4-1:0] node847;
	wire [4-1:0] node848;
	wire [4-1:0] node851;
	wire [4-1:0] node854;
	wire [4-1:0] node855;
	wire [4-1:0] node856;
	wire [4-1:0] node859;
	wire [4-1:0] node862;
	wire [4-1:0] node863;
	wire [4-1:0] node866;
	wire [4-1:0] node869;
	wire [4-1:0] node870;
	wire [4-1:0] node871;
	wire [4-1:0] node872;
	wire [4-1:0] node876;
	wire [4-1:0] node877;
	wire [4-1:0] node881;
	wire [4-1:0] node882;
	wire [4-1:0] node883;
	wire [4-1:0] node887;
	wire [4-1:0] node888;
	wire [4-1:0] node892;
	wire [4-1:0] node893;
	wire [4-1:0] node894;
	wire [4-1:0] node895;
	wire [4-1:0] node896;
	wire [4-1:0] node899;
	wire [4-1:0] node902;
	wire [4-1:0] node903;
	wire [4-1:0] node906;
	wire [4-1:0] node909;
	wire [4-1:0] node910;
	wire [4-1:0] node911;
	wire [4-1:0] node914;
	wire [4-1:0] node917;
	wire [4-1:0] node919;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node924;
	wire [4-1:0] node925;
	wire [4-1:0] node928;
	wire [4-1:0] node931;
	wire [4-1:0] node932;
	wire [4-1:0] node935;
	wire [4-1:0] node938;
	wire [4-1:0] node939;
	wire [4-1:0] node942;
	wire [4-1:0] node945;
	wire [4-1:0] node946;
	wire [4-1:0] node947;
	wire [4-1:0] node948;
	wire [4-1:0] node949;
	wire [4-1:0] node950;
	wire [4-1:0] node953;
	wire [4-1:0] node956;
	wire [4-1:0] node957;
	wire [4-1:0] node960;
	wire [4-1:0] node963;
	wire [4-1:0] node964;
	wire [4-1:0] node965;
	wire [4-1:0] node968;
	wire [4-1:0] node971;
	wire [4-1:0] node972;
	wire [4-1:0] node975;
	wire [4-1:0] node978;
	wire [4-1:0] node979;
	wire [4-1:0] node980;
	wire [4-1:0] node981;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node990;
	wire [4-1:0] node991;
	wire [4-1:0] node992;
	wire [4-1:0] node996;
	wire [4-1:0] node997;
	wire [4-1:0] node1001;
	wire [4-1:0] node1002;
	wire [4-1:0] node1003;
	wire [4-1:0] node1004;
	wire [4-1:0] node1005;
	wire [4-1:0] node1009;
	wire [4-1:0] node1010;
	wire [4-1:0] node1014;
	wire [4-1:0] node1015;
	wire [4-1:0] node1016;
	wire [4-1:0] node1020;
	wire [4-1:0] node1021;
	wire [4-1:0] node1025;
	wire [4-1:0] node1026;
	wire [4-1:0] node1027;
	wire [4-1:0] node1028;
	wire [4-1:0] node1032;
	wire [4-1:0] node1033;
	wire [4-1:0] node1037;
	wire [4-1:0] node1038;
	wire [4-1:0] node1039;
	wire [4-1:0] node1043;
	wire [4-1:0] node1044;
	wire [4-1:0] node1048;
	wire [4-1:0] node1049;
	wire [4-1:0] node1050;
	wire [4-1:0] node1051;
	wire [4-1:0] node1052;
	wire [4-1:0] node1053;
	wire [4-1:0] node1054;
	wire [4-1:0] node1058;
	wire [4-1:0] node1059;
	wire [4-1:0] node1063;
	wire [4-1:0] node1064;
	wire [4-1:0] node1065;
	wire [4-1:0] node1069;
	wire [4-1:0] node1070;
	wire [4-1:0] node1074;
	wire [4-1:0] node1075;
	wire [4-1:0] node1076;
	wire [4-1:0] node1077;
	wire [4-1:0] node1081;
	wire [4-1:0] node1082;
	wire [4-1:0] node1086;
	wire [4-1:0] node1087;
	wire [4-1:0] node1088;
	wire [4-1:0] node1092;
	wire [4-1:0] node1093;
	wire [4-1:0] node1097;
	wire [4-1:0] node1098;
	wire [4-1:0] node1099;
	wire [4-1:0] node1100;
	wire [4-1:0] node1101;
	wire [4-1:0] node1105;
	wire [4-1:0] node1106;
	wire [4-1:0] node1110;
	wire [4-1:0] node1111;
	wire [4-1:0] node1112;
	wire [4-1:0] node1116;
	wire [4-1:0] node1117;
	wire [4-1:0] node1121;
	wire [4-1:0] node1122;
	wire [4-1:0] node1123;
	wire [4-1:0] node1124;
	wire [4-1:0] node1127;
	wire [4-1:0] node1130;
	wire [4-1:0] node1131;
	wire [4-1:0] node1134;
	wire [4-1:0] node1137;
	wire [4-1:0] node1138;
	wire [4-1:0] node1139;
	wire [4-1:0] node1143;
	wire [4-1:0] node1144;
	wire [4-1:0] node1147;
	wire [4-1:0] node1150;
	wire [4-1:0] node1151;
	wire [4-1:0] node1152;
	wire [4-1:0] node1153;
	wire [4-1:0] node1154;
	wire [4-1:0] node1155;
	wire [4-1:0] node1159;
	wire [4-1:0] node1160;
	wire [4-1:0] node1164;
	wire [4-1:0] node1165;
	wire [4-1:0] node1166;
	wire [4-1:0] node1170;
	wire [4-1:0] node1171;
	wire [4-1:0] node1175;
	wire [4-1:0] node1176;
	wire [4-1:0] node1177;
	wire [4-1:0] node1178;
	wire [4-1:0] node1181;
	wire [4-1:0] node1184;
	wire [4-1:0] node1185;
	wire [4-1:0] node1188;
	wire [4-1:0] node1191;
	wire [4-1:0] node1192;
	wire [4-1:0] node1193;
	wire [4-1:0] node1197;
	wire [4-1:0] node1198;
	wire [4-1:0] node1201;
	wire [4-1:0] node1204;
	wire [4-1:0] node1205;
	wire [4-1:0] node1206;
	wire [4-1:0] node1207;
	wire [4-1:0] node1208;
	wire [4-1:0] node1212;
	wire [4-1:0] node1213;
	wire [4-1:0] node1217;
	wire [4-1:0] node1218;
	wire [4-1:0] node1219;
	wire [4-1:0] node1223;
	wire [4-1:0] node1224;
	wire [4-1:0] node1228;
	wire [4-1:0] node1229;
	wire [4-1:0] node1230;
	wire [4-1:0] node1231;
	wire [4-1:0] node1234;
	wire [4-1:0] node1237;
	wire [4-1:0] node1238;
	wire [4-1:0] node1241;
	wire [4-1:0] node1244;
	wire [4-1:0] node1245;
	wire [4-1:0] node1246;
	wire [4-1:0] node1249;
	wire [4-1:0] node1252;
	wire [4-1:0] node1253;
	wire [4-1:0] node1256;
	wire [4-1:0] node1259;
	wire [4-1:0] node1260;
	wire [4-1:0] node1261;
	wire [4-1:0] node1262;
	wire [4-1:0] node1263;
	wire [4-1:0] node1264;
	wire [4-1:0] node1265;
	wire [4-1:0] node1267;
	wire [4-1:0] node1270;
	wire [4-1:0] node1271;
	wire [4-1:0] node1274;
	wire [4-1:0] node1277;
	wire [4-1:0] node1278;
	wire [4-1:0] node1279;
	wire [4-1:0] node1282;
	wire [4-1:0] node1285;
	wire [4-1:0] node1287;
	wire [4-1:0] node1290;
	wire [4-1:0] node1291;
	wire [4-1:0] node1292;
	wire [4-1:0] node1293;
	wire [4-1:0] node1296;
	wire [4-1:0] node1299;
	wire [4-1:0] node1300;
	wire [4-1:0] node1303;
	wire [4-1:0] node1306;
	wire [4-1:0] node1307;
	wire [4-1:0] node1308;
	wire [4-1:0] node1311;
	wire [4-1:0] node1314;
	wire [4-1:0] node1315;
	wire [4-1:0] node1318;
	wire [4-1:0] node1321;
	wire [4-1:0] node1322;
	wire [4-1:0] node1323;
	wire [4-1:0] node1324;
	wire [4-1:0] node1325;
	wire [4-1:0] node1329;
	wire [4-1:0] node1330;
	wire [4-1:0] node1334;
	wire [4-1:0] node1335;
	wire [4-1:0] node1336;
	wire [4-1:0] node1339;
	wire [4-1:0] node1342;
	wire [4-1:0] node1344;
	wire [4-1:0] node1347;
	wire [4-1:0] node1348;
	wire [4-1:0] node1349;
	wire [4-1:0] node1350;
	wire [4-1:0] node1353;
	wire [4-1:0] node1356;
	wire [4-1:0] node1357;
	wire [4-1:0] node1360;
	wire [4-1:0] node1363;
	wire [4-1:0] node1364;
	wire [4-1:0] node1365;
	wire [4-1:0] node1368;
	wire [4-1:0] node1371;
	wire [4-1:0] node1372;
	wire [4-1:0] node1375;
	wire [4-1:0] node1378;
	wire [4-1:0] node1379;
	wire [4-1:0] node1380;
	wire [4-1:0] node1381;
	wire [4-1:0] node1382;
	wire [4-1:0] node1383;
	wire [4-1:0] node1386;
	wire [4-1:0] node1389;
	wire [4-1:0] node1391;
	wire [4-1:0] node1394;
	wire [4-1:0] node1395;
	wire [4-1:0] node1396;
	wire [4-1:0] node1399;
	wire [4-1:0] node1402;
	wire [4-1:0] node1404;
	wire [4-1:0] node1407;
	wire [4-1:0] node1408;
	wire [4-1:0] node1409;
	wire [4-1:0] node1410;
	wire [4-1:0] node1413;
	wire [4-1:0] node1416;
	wire [4-1:0] node1417;
	wire [4-1:0] node1420;
	wire [4-1:0] node1423;
	wire [4-1:0] node1424;
	wire [4-1:0] node1425;
	wire [4-1:0] node1428;
	wire [4-1:0] node1431;
	wire [4-1:0] node1432;
	wire [4-1:0] node1435;
	wire [4-1:0] node1438;
	wire [4-1:0] node1439;
	wire [4-1:0] node1440;
	wire [4-1:0] node1441;
	wire [4-1:0] node1442;
	wire [4-1:0] node1445;
	wire [4-1:0] node1448;
	wire [4-1:0] node1449;
	wire [4-1:0] node1452;
	wire [4-1:0] node1455;
	wire [4-1:0] node1456;
	wire [4-1:0] node1457;
	wire [4-1:0] node1460;
	wire [4-1:0] node1463;
	wire [4-1:0] node1464;
	wire [4-1:0] node1467;
	wire [4-1:0] node1470;
	wire [4-1:0] node1471;
	wire [4-1:0] node1472;
	wire [4-1:0] node1474;
	wire [4-1:0] node1477;
	wire [4-1:0] node1478;
	wire [4-1:0] node1481;
	wire [4-1:0] node1484;
	wire [4-1:0] node1485;
	wire [4-1:0] node1487;
	wire [4-1:0] node1490;
	wire [4-1:0] node1491;
	wire [4-1:0] node1494;
	wire [4-1:0] node1497;
	wire [4-1:0] node1498;
	wire [4-1:0] node1499;
	wire [4-1:0] node1500;
	wire [4-1:0] node1501;
	wire [4-1:0] node1502;
	wire [4-1:0] node1503;
	wire [4-1:0] node1506;
	wire [4-1:0] node1509;
	wire [4-1:0] node1511;
	wire [4-1:0] node1514;
	wire [4-1:0] node1515;
	wire [4-1:0] node1516;
	wire [4-1:0] node1519;
	wire [4-1:0] node1522;
	wire [4-1:0] node1523;
	wire [4-1:0] node1526;
	wire [4-1:0] node1529;
	wire [4-1:0] node1530;
	wire [4-1:0] node1531;
	wire [4-1:0] node1534;
	wire [4-1:0] node1537;
	wire [4-1:0] node1538;
	wire [4-1:0] node1539;
	wire [4-1:0] node1542;
	wire [4-1:0] node1545;
	wire [4-1:0] node1546;
	wire [4-1:0] node1549;
	wire [4-1:0] node1552;
	wire [4-1:0] node1553;
	wire [4-1:0] node1554;
	wire [4-1:0] node1555;
	wire [4-1:0] node1558;
	wire [4-1:0] node1559;
	wire [4-1:0] node1562;
	wire [4-1:0] node1565;
	wire [4-1:0] node1566;
	wire [4-1:0] node1568;
	wire [4-1:0] node1571;
	wire [4-1:0] node1572;
	wire [4-1:0] node1575;
	wire [4-1:0] node1578;
	wire [4-1:0] node1579;
	wire [4-1:0] node1580;
	wire [4-1:0] node1581;
	wire [4-1:0] node1585;
	wire [4-1:0] node1586;
	wire [4-1:0] node1590;
	wire [4-1:0] node1591;
	wire [4-1:0] node1592;
	wire [4-1:0] node1596;
	wire [4-1:0] node1597;
	wire [4-1:0] node1601;
	wire [4-1:0] node1602;
	wire [4-1:0] node1603;
	wire [4-1:0] node1604;
	wire [4-1:0] node1605;
	wire [4-1:0] node1607;
	wire [4-1:0] node1610;
	wire [4-1:0] node1611;
	wire [4-1:0] node1614;
	wire [4-1:0] node1617;
	wire [4-1:0] node1618;
	wire [4-1:0] node1619;
	wire [4-1:0] node1622;
	wire [4-1:0] node1625;
	wire [4-1:0] node1626;
	wire [4-1:0] node1629;
	wire [4-1:0] node1632;
	wire [4-1:0] node1633;
	wire [4-1:0] node1634;
	wire [4-1:0] node1635;
	wire [4-1:0] node1639;
	wire [4-1:0] node1640;
	wire [4-1:0] node1644;
	wire [4-1:0] node1645;
	wire [4-1:0] node1646;
	wire [4-1:0] node1650;
	wire [4-1:0] node1651;
	wire [4-1:0] node1655;
	wire [4-1:0] node1656;
	wire [4-1:0] node1657;
	wire [4-1:0] node1658;
	wire [4-1:0] node1659;
	wire [4-1:0] node1662;
	wire [4-1:0] node1665;
	wire [4-1:0] node1666;
	wire [4-1:0] node1669;
	wire [4-1:0] node1672;
	wire [4-1:0] node1673;
	wire [4-1:0] node1674;
	wire [4-1:0] node1677;
	wire [4-1:0] node1680;
	wire [4-1:0] node1681;
	wire [4-1:0] node1684;
	wire [4-1:0] node1687;
	wire [4-1:0] node1688;
	wire [4-1:0] node1689;
	wire [4-1:0] node1690;
	wire [4-1:0] node1694;
	wire [4-1:0] node1695;
	wire [4-1:0] node1699;
	wire [4-1:0] node1700;
	wire [4-1:0] node1701;
	wire [4-1:0] node1705;
	wire [4-1:0] node1706;
	wire [4-1:0] node1710;
	wire [4-1:0] node1711;
	wire [4-1:0] node1712;
	wire [4-1:0] node1713;
	wire [4-1:0] node1714;
	wire [4-1:0] node1715;
	wire [4-1:0] node1716;
	wire [4-1:0] node1717;
	wire [4-1:0] node1718;
	wire [4-1:0] node1719;
	wire [4-1:0] node1722;
	wire [4-1:0] node1725;
	wire [4-1:0] node1726;
	wire [4-1:0] node1730;
	wire [4-1:0] node1731;
	wire [4-1:0] node1732;
	wire [4-1:0] node1735;
	wire [4-1:0] node1738;
	wire [4-1:0] node1739;
	wire [4-1:0] node1742;
	wire [4-1:0] node1745;
	wire [4-1:0] node1746;
	wire [4-1:0] node1747;
	wire [4-1:0] node1748;
	wire [4-1:0] node1751;
	wire [4-1:0] node1754;
	wire [4-1:0] node1755;
	wire [4-1:0] node1758;
	wire [4-1:0] node1761;
	wire [4-1:0] node1762;
	wire [4-1:0] node1763;
	wire [4-1:0] node1766;
	wire [4-1:0] node1769;
	wire [4-1:0] node1770;
	wire [4-1:0] node1774;
	wire [4-1:0] node1775;
	wire [4-1:0] node1776;
	wire [4-1:0] node1777;
	wire [4-1:0] node1778;
	wire [4-1:0] node1781;
	wire [4-1:0] node1784;
	wire [4-1:0] node1785;
	wire [4-1:0] node1788;
	wire [4-1:0] node1791;
	wire [4-1:0] node1792;
	wire [4-1:0] node1793;
	wire [4-1:0] node1796;
	wire [4-1:0] node1799;
	wire [4-1:0] node1800;
	wire [4-1:0] node1803;
	wire [4-1:0] node1806;
	wire [4-1:0] node1807;
	wire [4-1:0] node1808;
	wire [4-1:0] node1809;
	wire [4-1:0] node1812;
	wire [4-1:0] node1815;
	wire [4-1:0] node1816;
	wire [4-1:0] node1819;
	wire [4-1:0] node1822;
	wire [4-1:0] node1823;
	wire [4-1:0] node1824;
	wire [4-1:0] node1827;
	wire [4-1:0] node1830;
	wire [4-1:0] node1831;
	wire [4-1:0] node1834;
	wire [4-1:0] node1837;
	wire [4-1:0] node1838;
	wire [4-1:0] node1839;
	wire [4-1:0] node1840;
	wire [4-1:0] node1841;
	wire [4-1:0] node1842;
	wire [4-1:0] node1845;
	wire [4-1:0] node1848;
	wire [4-1:0] node1849;
	wire [4-1:0] node1852;
	wire [4-1:0] node1855;
	wire [4-1:0] node1856;
	wire [4-1:0] node1857;
	wire [4-1:0] node1860;
	wire [4-1:0] node1863;
	wire [4-1:0] node1865;
	wire [4-1:0] node1868;
	wire [4-1:0] node1869;
	wire [4-1:0] node1870;
	wire [4-1:0] node1871;
	wire [4-1:0] node1874;
	wire [4-1:0] node1877;
	wire [4-1:0] node1878;
	wire [4-1:0] node1881;
	wire [4-1:0] node1884;
	wire [4-1:0] node1885;
	wire [4-1:0] node1886;
	wire [4-1:0] node1889;
	wire [4-1:0] node1892;
	wire [4-1:0] node1893;
	wire [4-1:0] node1896;
	wire [4-1:0] node1899;
	wire [4-1:0] node1900;
	wire [4-1:0] node1901;
	wire [4-1:0] node1902;
	wire [4-1:0] node1903;
	wire [4-1:0] node1906;
	wire [4-1:0] node1909;
	wire [4-1:0] node1910;
	wire [4-1:0] node1913;
	wire [4-1:0] node1916;
	wire [4-1:0] node1917;
	wire [4-1:0] node1918;
	wire [4-1:0] node1921;
	wire [4-1:0] node1924;
	wire [4-1:0] node1925;
	wire [4-1:0] node1928;
	wire [4-1:0] node1931;
	wire [4-1:0] node1932;
	wire [4-1:0] node1933;
	wire [4-1:0] node1934;
	wire [4-1:0] node1937;
	wire [4-1:0] node1940;
	wire [4-1:0] node1941;
	wire [4-1:0] node1944;
	wire [4-1:0] node1947;
	wire [4-1:0] node1948;
	wire [4-1:0] node1949;
	wire [4-1:0] node1952;
	wire [4-1:0] node1955;
	wire [4-1:0] node1956;
	wire [4-1:0] node1959;
	wire [4-1:0] node1962;
	wire [4-1:0] node1963;
	wire [4-1:0] node1964;
	wire [4-1:0] node1965;
	wire [4-1:0] node1966;
	wire [4-1:0] node1967;
	wire [4-1:0] node1968;
	wire [4-1:0] node1971;
	wire [4-1:0] node1974;
	wire [4-1:0] node1975;
	wire [4-1:0] node1978;
	wire [4-1:0] node1981;
	wire [4-1:0] node1982;
	wire [4-1:0] node1983;
	wire [4-1:0] node1986;
	wire [4-1:0] node1989;
	wire [4-1:0] node1990;
	wire [4-1:0] node1993;
	wire [4-1:0] node1996;
	wire [4-1:0] node1997;
	wire [4-1:0] node1998;
	wire [4-1:0] node1999;
	wire [4-1:0] node2002;
	wire [4-1:0] node2005;
	wire [4-1:0] node2006;
	wire [4-1:0] node2009;
	wire [4-1:0] node2012;
	wire [4-1:0] node2013;
	wire [4-1:0] node2014;
	wire [4-1:0] node2017;
	wire [4-1:0] node2020;
	wire [4-1:0] node2021;
	wire [4-1:0] node2024;
	wire [4-1:0] node2027;
	wire [4-1:0] node2028;
	wire [4-1:0] node2029;
	wire [4-1:0] node2030;
	wire [4-1:0] node2031;
	wire [4-1:0] node2034;
	wire [4-1:0] node2037;
	wire [4-1:0] node2038;
	wire [4-1:0] node2041;
	wire [4-1:0] node2044;
	wire [4-1:0] node2045;
	wire [4-1:0] node2046;
	wire [4-1:0] node2049;
	wire [4-1:0] node2052;
	wire [4-1:0] node2053;
	wire [4-1:0] node2056;
	wire [4-1:0] node2059;
	wire [4-1:0] node2060;
	wire [4-1:0] node2061;
	wire [4-1:0] node2064;
	wire [4-1:0] node2067;
	wire [4-1:0] node2068;
	wire [4-1:0] node2069;
	wire [4-1:0] node2072;
	wire [4-1:0] node2075;
	wire [4-1:0] node2076;
	wire [4-1:0] node2079;
	wire [4-1:0] node2082;
	wire [4-1:0] node2083;
	wire [4-1:0] node2084;
	wire [4-1:0] node2085;
	wire [4-1:0] node2086;
	wire [4-1:0] node2087;
	wire [4-1:0] node2090;
	wire [4-1:0] node2093;
	wire [4-1:0] node2094;
	wire [4-1:0] node2097;
	wire [4-1:0] node2100;
	wire [4-1:0] node2101;
	wire [4-1:0] node2104;
	wire [4-1:0] node2107;
	wire [4-1:0] node2108;
	wire [4-1:0] node2111;
	wire [4-1:0] node2114;
	wire [4-1:0] node2115;
	wire [4-1:0] node2116;
	wire [4-1:0] node2117;
	wire [4-1:0] node2120;
	wire [4-1:0] node2123;
	wire [4-1:0] node2124;
	wire [4-1:0] node2127;
	wire [4-1:0] node2130;
	wire [4-1:0] node2131;
	wire [4-1:0] node2134;
	wire [4-1:0] node2137;
	wire [4-1:0] node2138;
	wire [4-1:0] node2139;
	wire [4-1:0] node2140;
	wire [4-1:0] node2141;
	wire [4-1:0] node2142;
	wire [4-1:0] node2143;
	wire [4-1:0] node2144;
	wire [4-1:0] node2147;
	wire [4-1:0] node2150;
	wire [4-1:0] node2151;
	wire [4-1:0] node2154;
	wire [4-1:0] node2157;
	wire [4-1:0] node2158;
	wire [4-1:0] node2159;
	wire [4-1:0] node2162;
	wire [4-1:0] node2165;
	wire [4-1:0] node2166;
	wire [4-1:0] node2169;
	wire [4-1:0] node2172;
	wire [4-1:0] node2173;
	wire [4-1:0] node2174;
	wire [4-1:0] node2175;
	wire [4-1:0] node2178;
	wire [4-1:0] node2181;
	wire [4-1:0] node2182;
	wire [4-1:0] node2185;
	wire [4-1:0] node2188;
	wire [4-1:0] node2189;
	wire [4-1:0] node2190;
	wire [4-1:0] node2193;
	wire [4-1:0] node2196;
	wire [4-1:0] node2197;
	wire [4-1:0] node2201;
	wire [4-1:0] node2202;
	wire [4-1:0] node2203;
	wire [4-1:0] node2204;
	wire [4-1:0] node2205;
	wire [4-1:0] node2208;
	wire [4-1:0] node2211;
	wire [4-1:0] node2212;
	wire [4-1:0] node2215;
	wire [4-1:0] node2218;
	wire [4-1:0] node2219;
	wire [4-1:0] node2220;
	wire [4-1:0] node2223;
	wire [4-1:0] node2226;
	wire [4-1:0] node2227;
	wire [4-1:0] node2230;
	wire [4-1:0] node2233;
	wire [4-1:0] node2234;
	wire [4-1:0] node2235;
	wire [4-1:0] node2236;
	wire [4-1:0] node2239;
	wire [4-1:0] node2242;
	wire [4-1:0] node2244;
	wire [4-1:0] node2247;
	wire [4-1:0] node2248;
	wire [4-1:0] node2249;
	wire [4-1:0] node2252;
	wire [4-1:0] node2255;
	wire [4-1:0] node2256;
	wire [4-1:0] node2260;
	wire [4-1:0] node2261;
	wire [4-1:0] node2262;
	wire [4-1:0] node2263;
	wire [4-1:0] node2264;
	wire [4-1:0] node2265;
	wire [4-1:0] node2268;
	wire [4-1:0] node2271;
	wire [4-1:0] node2272;
	wire [4-1:0] node2275;
	wire [4-1:0] node2278;
	wire [4-1:0] node2279;
	wire [4-1:0] node2280;
	wire [4-1:0] node2283;
	wire [4-1:0] node2286;
	wire [4-1:0] node2287;
	wire [4-1:0] node2291;
	wire [4-1:0] node2292;
	wire [4-1:0] node2293;
	wire [4-1:0] node2294;
	wire [4-1:0] node2297;
	wire [4-1:0] node2300;
	wire [4-1:0] node2301;
	wire [4-1:0] node2304;
	wire [4-1:0] node2307;
	wire [4-1:0] node2308;
	wire [4-1:0] node2310;
	wire [4-1:0] node2313;
	wire [4-1:0] node2314;
	wire [4-1:0] node2317;
	wire [4-1:0] node2320;
	wire [4-1:0] node2321;
	wire [4-1:0] node2322;
	wire [4-1:0] node2323;
	wire [4-1:0] node2325;
	wire [4-1:0] node2328;
	wire [4-1:0] node2330;
	wire [4-1:0] node2333;
	wire [4-1:0] node2334;
	wire [4-1:0] node2335;
	wire [4-1:0] node2338;
	wire [4-1:0] node2341;
	wire [4-1:0] node2342;
	wire [4-1:0] node2345;
	wire [4-1:0] node2348;
	wire [4-1:0] node2349;
	wire [4-1:0] node2350;
	wire [4-1:0] node2351;
	wire [4-1:0] node2354;
	wire [4-1:0] node2357;
	wire [4-1:0] node2359;
	wire [4-1:0] node2362;
	wire [4-1:0] node2363;
	wire [4-1:0] node2364;
	wire [4-1:0] node2367;
	wire [4-1:0] node2370;
	wire [4-1:0] node2372;
	wire [4-1:0] node2375;
	wire [4-1:0] node2376;
	wire [4-1:0] node2377;
	wire [4-1:0] node2378;
	wire [4-1:0] node2379;
	wire [4-1:0] node2380;
	wire [4-1:0] node2381;
	wire [4-1:0] node2385;
	wire [4-1:0] node2386;
	wire [4-1:0] node2389;
	wire [4-1:0] node2392;
	wire [4-1:0] node2393;
	wire [4-1:0] node2394;
	wire [4-1:0] node2397;
	wire [4-1:0] node2400;
	wire [4-1:0] node2401;
	wire [4-1:0] node2404;
	wire [4-1:0] node2407;
	wire [4-1:0] node2408;
	wire [4-1:0] node2409;
	wire [4-1:0] node2410;
	wire [4-1:0] node2413;
	wire [4-1:0] node2416;
	wire [4-1:0] node2417;
	wire [4-1:0] node2420;
	wire [4-1:0] node2423;
	wire [4-1:0] node2424;
	wire [4-1:0] node2425;
	wire [4-1:0] node2428;
	wire [4-1:0] node2431;
	wire [4-1:0] node2432;
	wire [4-1:0] node2435;
	wire [4-1:0] node2438;
	wire [4-1:0] node2439;
	wire [4-1:0] node2440;
	wire [4-1:0] node2441;
	wire [4-1:0] node2442;
	wire [4-1:0] node2445;
	wire [4-1:0] node2448;
	wire [4-1:0] node2449;
	wire [4-1:0] node2452;
	wire [4-1:0] node2455;
	wire [4-1:0] node2456;
	wire [4-1:0] node2457;
	wire [4-1:0] node2460;
	wire [4-1:0] node2463;
	wire [4-1:0] node2465;
	wire [4-1:0] node2468;
	wire [4-1:0] node2469;
	wire [4-1:0] node2470;
	wire [4-1:0] node2471;
	wire [4-1:0] node2474;
	wire [4-1:0] node2477;
	wire [4-1:0] node2478;
	wire [4-1:0] node2481;
	wire [4-1:0] node2484;
	wire [4-1:0] node2485;
	wire [4-1:0] node2486;
	wire [4-1:0] node2489;
	wire [4-1:0] node2492;
	wire [4-1:0] node2494;
	wire [4-1:0] node2497;
	wire [4-1:0] node2498;
	wire [4-1:0] node2499;
	wire [4-1:0] node2500;
	wire [4-1:0] node2501;
	wire [4-1:0] node2502;
	wire [4-1:0] node2505;
	wire [4-1:0] node2508;
	wire [4-1:0] node2509;
	wire [4-1:0] node2512;
	wire [4-1:0] node2515;
	wire [4-1:0] node2516;
	wire [4-1:0] node2517;
	wire [4-1:0] node2520;
	wire [4-1:0] node2523;
	wire [4-1:0] node2524;
	wire [4-1:0] node2527;
	wire [4-1:0] node2530;
	wire [4-1:0] node2531;
	wire [4-1:0] node2532;
	wire [4-1:0] node2533;
	wire [4-1:0] node2536;
	wire [4-1:0] node2539;
	wire [4-1:0] node2540;
	wire [4-1:0] node2543;
	wire [4-1:0] node2546;
	wire [4-1:0] node2547;
	wire [4-1:0] node2549;
	wire [4-1:0] node2552;
	wire [4-1:0] node2553;
	wire [4-1:0] node2556;
	wire [4-1:0] node2559;
	wire [4-1:0] node2560;
	wire [4-1:0] node2561;
	wire [4-1:0] node2562;
	wire [4-1:0] node2564;
	wire [4-1:0] node2567;
	wire [4-1:0] node2568;
	wire [4-1:0] node2571;
	wire [4-1:0] node2574;
	wire [4-1:0] node2575;
	wire [4-1:0] node2576;
	wire [4-1:0] node2579;
	wire [4-1:0] node2582;
	wire [4-1:0] node2583;
	wire [4-1:0] node2586;
	wire [4-1:0] node2589;
	wire [4-1:0] node2590;
	wire [4-1:0] node2591;
	wire [4-1:0] node2592;
	wire [4-1:0] node2595;
	wire [4-1:0] node2598;
	wire [4-1:0] node2599;
	wire [4-1:0] node2602;
	wire [4-1:0] node2605;
	wire [4-1:0] node2606;
	wire [4-1:0] node2607;
	wire [4-1:0] node2611;
	wire [4-1:0] node2612;
	wire [4-1:0] node2615;
	wire [4-1:0] node2618;
	wire [4-1:0] node2619;
	wire [4-1:0] node2620;
	wire [4-1:0] node2621;
	wire [4-1:0] node2622;
	wire [4-1:0] node2623;
	wire [4-1:0] node2624;
	wire [4-1:0] node2625;
	wire [4-1:0] node2626;
	wire [4-1:0] node2629;
	wire [4-1:0] node2632;
	wire [4-1:0] node2633;
	wire [4-1:0] node2636;
	wire [4-1:0] node2639;
	wire [4-1:0] node2640;
	wire [4-1:0] node2641;
	wire [4-1:0] node2644;
	wire [4-1:0] node2647;
	wire [4-1:0] node2648;
	wire [4-1:0] node2651;
	wire [4-1:0] node2654;
	wire [4-1:0] node2655;
	wire [4-1:0] node2656;
	wire [4-1:0] node2657;
	wire [4-1:0] node2661;
	wire [4-1:0] node2662;
	wire [4-1:0] node2666;
	wire [4-1:0] node2667;
	wire [4-1:0] node2668;
	wire [4-1:0] node2672;
	wire [4-1:0] node2673;
	wire [4-1:0] node2677;
	wire [4-1:0] node2678;
	wire [4-1:0] node2679;
	wire [4-1:0] node2680;
	wire [4-1:0] node2681;
	wire [4-1:0] node2685;
	wire [4-1:0] node2686;
	wire [4-1:0] node2690;
	wire [4-1:0] node2691;
	wire [4-1:0] node2692;
	wire [4-1:0] node2696;
	wire [4-1:0] node2697;
	wire [4-1:0] node2701;
	wire [4-1:0] node2702;
	wire [4-1:0] node2703;
	wire [4-1:0] node2704;
	wire [4-1:0] node2707;
	wire [4-1:0] node2710;
	wire [4-1:0] node2711;
	wire [4-1:0] node2714;
	wire [4-1:0] node2717;
	wire [4-1:0] node2718;
	wire [4-1:0] node2719;
	wire [4-1:0] node2722;
	wire [4-1:0] node2725;
	wire [4-1:0] node2726;
	wire [4-1:0] node2729;
	wire [4-1:0] node2732;
	wire [4-1:0] node2733;
	wire [4-1:0] node2734;
	wire [4-1:0] node2735;
	wire [4-1:0] node2736;
	wire [4-1:0] node2737;
	wire [4-1:0] node2740;
	wire [4-1:0] node2744;
	wire [4-1:0] node2745;
	wire [4-1:0] node2746;
	wire [4-1:0] node2750;
	wire [4-1:0] node2751;
	wire [4-1:0] node2755;
	wire [4-1:0] node2756;
	wire [4-1:0] node2757;
	wire [4-1:0] node2758;
	wire [4-1:0] node2762;
	wire [4-1:0] node2763;
	wire [4-1:0] node2767;
	wire [4-1:0] node2768;
	wire [4-1:0] node2769;
	wire [4-1:0] node2773;
	wire [4-1:0] node2774;
	wire [4-1:0] node2778;
	wire [4-1:0] node2779;
	wire [4-1:0] node2780;
	wire [4-1:0] node2781;
	wire [4-1:0] node2782;
	wire [4-1:0] node2786;
	wire [4-1:0] node2787;
	wire [4-1:0] node2791;
	wire [4-1:0] node2792;
	wire [4-1:0] node2793;
	wire [4-1:0] node2797;
	wire [4-1:0] node2798;
	wire [4-1:0] node2802;
	wire [4-1:0] node2803;
	wire [4-1:0] node2804;
	wire [4-1:0] node2805;
	wire [4-1:0] node2809;
	wire [4-1:0] node2810;
	wire [4-1:0] node2814;
	wire [4-1:0] node2815;
	wire [4-1:0] node2816;
	wire [4-1:0] node2820;
	wire [4-1:0] node2821;
	wire [4-1:0] node2825;
	wire [4-1:0] node2826;
	wire [4-1:0] node2827;
	wire [4-1:0] node2828;
	wire [4-1:0] node2829;
	wire [4-1:0] node2830;
	wire [4-1:0] node2831;
	wire [4-1:0] node2834;
	wire [4-1:0] node2837;
	wire [4-1:0] node2838;
	wire [4-1:0] node2841;
	wire [4-1:0] node2844;
	wire [4-1:0] node2845;
	wire [4-1:0] node2846;
	wire [4-1:0] node2849;
	wire [4-1:0] node2852;
	wire [4-1:0] node2853;
	wire [4-1:0] node2856;
	wire [4-1:0] node2859;
	wire [4-1:0] node2860;
	wire [4-1:0] node2861;
	wire [4-1:0] node2862;
	wire [4-1:0] node2866;
	wire [4-1:0] node2867;
	wire [4-1:0] node2871;
	wire [4-1:0] node2872;
	wire [4-1:0] node2873;
	wire [4-1:0] node2877;
	wire [4-1:0] node2878;
	wire [4-1:0] node2882;
	wire [4-1:0] node2883;
	wire [4-1:0] node2884;
	wire [4-1:0] node2885;
	wire [4-1:0] node2886;
	wire [4-1:0] node2890;
	wire [4-1:0] node2891;
	wire [4-1:0] node2895;
	wire [4-1:0] node2896;
	wire [4-1:0] node2897;
	wire [4-1:0] node2901;
	wire [4-1:0] node2902;
	wire [4-1:0] node2906;
	wire [4-1:0] node2907;
	wire [4-1:0] node2908;
	wire [4-1:0] node2909;
	wire [4-1:0] node2912;
	wire [4-1:0] node2915;
	wire [4-1:0] node2916;
	wire [4-1:0] node2920;
	wire [4-1:0] node2921;
	wire [4-1:0] node2922;
	wire [4-1:0] node2926;
	wire [4-1:0] node2928;
	wire [4-1:0] node2931;
	wire [4-1:0] node2932;
	wire [4-1:0] node2933;
	wire [4-1:0] node2934;
	wire [4-1:0] node2935;
	wire [4-1:0] node2936;
	wire [4-1:0] node2941;
	wire [4-1:0] node2942;
	wire [4-1:0] node2943;
	wire [4-1:0] node2947;
	wire [4-1:0] node2948;
	wire [4-1:0] node2952;
	wire [4-1:0] node2953;
	wire [4-1:0] node2954;
	wire [4-1:0] node2955;
	wire [4-1:0] node2959;
	wire [4-1:0] node2960;
	wire [4-1:0] node2964;
	wire [4-1:0] node2965;
	wire [4-1:0] node2966;
	wire [4-1:0] node2970;
	wire [4-1:0] node2971;
	wire [4-1:0] node2975;
	wire [4-1:0] node2976;
	wire [4-1:0] node2977;
	wire [4-1:0] node2978;
	wire [4-1:0] node2979;
	wire [4-1:0] node2983;
	wire [4-1:0] node2984;
	wire [4-1:0] node2988;
	wire [4-1:0] node2989;
	wire [4-1:0] node2990;
	wire [4-1:0] node2994;
	wire [4-1:0] node2995;
	wire [4-1:0] node2999;
	wire [4-1:0] node3000;
	wire [4-1:0] node3001;
	wire [4-1:0] node3002;
	wire [4-1:0] node3005;
	wire [4-1:0] node3008;
	wire [4-1:0] node3009;
	wire [4-1:0] node3012;
	wire [4-1:0] node3015;
	wire [4-1:0] node3016;
	wire [4-1:0] node3017;
	wire [4-1:0] node3020;
	wire [4-1:0] node3023;
	wire [4-1:0] node3024;
	wire [4-1:0] node3027;
	wire [4-1:0] node3030;
	wire [4-1:0] node3031;
	wire [4-1:0] node3032;
	wire [4-1:0] node3033;
	wire [4-1:0] node3034;
	wire [4-1:0] node3035;
	wire [4-1:0] node3036;
	wire [4-1:0] node3037;
	wire [4-1:0] node3040;
	wire [4-1:0] node3043;
	wire [4-1:0] node3044;
	wire [4-1:0] node3047;
	wire [4-1:0] node3050;
	wire [4-1:0] node3051;
	wire [4-1:0] node3052;
	wire [4-1:0] node3055;
	wire [4-1:0] node3058;
	wire [4-1:0] node3059;
	wire [4-1:0] node3062;
	wire [4-1:0] node3065;
	wire [4-1:0] node3066;
	wire [4-1:0] node3067;
	wire [4-1:0] node3068;
	wire [4-1:0] node3071;
	wire [4-1:0] node3074;
	wire [4-1:0] node3075;
	wire [4-1:0] node3078;
	wire [4-1:0] node3081;
	wire [4-1:0] node3082;
	wire [4-1:0] node3083;
	wire [4-1:0] node3086;
	wire [4-1:0] node3089;
	wire [4-1:0] node3090;
	wire [4-1:0] node3093;
	wire [4-1:0] node3096;
	wire [4-1:0] node3097;
	wire [4-1:0] node3098;
	wire [4-1:0] node3099;
	wire [4-1:0] node3100;
	wire [4-1:0] node3103;
	wire [4-1:0] node3106;
	wire [4-1:0] node3108;
	wire [4-1:0] node3111;
	wire [4-1:0] node3112;
	wire [4-1:0] node3113;
	wire [4-1:0] node3116;
	wire [4-1:0] node3119;
	wire [4-1:0] node3120;
	wire [4-1:0] node3123;
	wire [4-1:0] node3126;
	wire [4-1:0] node3127;
	wire [4-1:0] node3128;
	wire [4-1:0] node3129;
	wire [4-1:0] node3132;
	wire [4-1:0] node3135;
	wire [4-1:0] node3136;
	wire [4-1:0] node3139;
	wire [4-1:0] node3142;
	wire [4-1:0] node3143;
	wire [4-1:0] node3144;
	wire [4-1:0] node3147;
	wire [4-1:0] node3150;
	wire [4-1:0] node3151;
	wire [4-1:0] node3154;
	wire [4-1:0] node3157;
	wire [4-1:0] node3158;
	wire [4-1:0] node3159;
	wire [4-1:0] node3160;
	wire [4-1:0] node3161;
	wire [4-1:0] node3162;
	wire [4-1:0] node3166;
	wire [4-1:0] node3167;
	wire [4-1:0] node3171;
	wire [4-1:0] node3172;
	wire [4-1:0] node3174;
	wire [4-1:0] node3177;
	wire [4-1:0] node3178;
	wire [4-1:0] node3181;
	wire [4-1:0] node3184;
	wire [4-1:0] node3185;
	wire [4-1:0] node3186;
	wire [4-1:0] node3187;
	wire [4-1:0] node3190;
	wire [4-1:0] node3193;
	wire [4-1:0] node3195;
	wire [4-1:0] node3198;
	wire [4-1:0] node3199;
	wire [4-1:0] node3200;
	wire [4-1:0] node3203;
	wire [4-1:0] node3206;
	wire [4-1:0] node3207;
	wire [4-1:0] node3211;
	wire [4-1:0] node3212;
	wire [4-1:0] node3213;
	wire [4-1:0] node3214;
	wire [4-1:0] node3215;
	wire [4-1:0] node3218;
	wire [4-1:0] node3221;
	wire [4-1:0] node3222;
	wire [4-1:0] node3225;
	wire [4-1:0] node3228;
	wire [4-1:0] node3229;
	wire [4-1:0] node3230;
	wire [4-1:0] node3233;
	wire [4-1:0] node3236;
	wire [4-1:0] node3237;
	wire [4-1:0] node3240;
	wire [4-1:0] node3243;
	wire [4-1:0] node3244;
	wire [4-1:0] node3245;
	wire [4-1:0] node3247;
	wire [4-1:0] node3250;
	wire [4-1:0] node3251;
	wire [4-1:0] node3254;
	wire [4-1:0] node3257;
	wire [4-1:0] node3258;
	wire [4-1:0] node3259;
	wire [4-1:0] node3263;
	wire [4-1:0] node3264;
	wire [4-1:0] node3267;
	wire [4-1:0] node3270;
	wire [4-1:0] node3271;
	wire [4-1:0] node3272;
	wire [4-1:0] node3273;
	wire [4-1:0] node3274;
	wire [4-1:0] node3275;
	wire [4-1:0] node3276;
	wire [4-1:0] node3279;
	wire [4-1:0] node3282;
	wire [4-1:0] node3284;
	wire [4-1:0] node3287;
	wire [4-1:0] node3288;
	wire [4-1:0] node3289;
	wire [4-1:0] node3292;
	wire [4-1:0] node3295;
	wire [4-1:0] node3296;
	wire [4-1:0] node3299;
	wire [4-1:0] node3302;
	wire [4-1:0] node3303;
	wire [4-1:0] node3304;
	wire [4-1:0] node3305;
	wire [4-1:0] node3308;
	wire [4-1:0] node3311;
	wire [4-1:0] node3312;
	wire [4-1:0] node3315;
	wire [4-1:0] node3318;
	wire [4-1:0] node3319;
	wire [4-1:0] node3321;
	wire [4-1:0] node3324;
	wire [4-1:0] node3325;
	wire [4-1:0] node3328;
	wire [4-1:0] node3331;
	wire [4-1:0] node3332;
	wire [4-1:0] node3333;
	wire [4-1:0] node3334;
	wire [4-1:0] node3335;
	wire [4-1:0] node3338;
	wire [4-1:0] node3341;
	wire [4-1:0] node3344;
	wire [4-1:0] node3345;
	wire [4-1:0] node3346;
	wire [4-1:0] node3349;
	wire [4-1:0] node3352;
	wire [4-1:0] node3353;
	wire [4-1:0] node3357;
	wire [4-1:0] node3358;
	wire [4-1:0] node3359;
	wire [4-1:0] node3360;
	wire [4-1:0] node3363;
	wire [4-1:0] node3366;
	wire [4-1:0] node3367;
	wire [4-1:0] node3370;
	wire [4-1:0] node3373;
	wire [4-1:0] node3374;
	wire [4-1:0] node3375;
	wire [4-1:0] node3378;
	wire [4-1:0] node3381;
	wire [4-1:0] node3382;
	wire [4-1:0] node3385;
	wire [4-1:0] node3388;
	wire [4-1:0] node3389;
	wire [4-1:0] node3390;
	wire [4-1:0] node3391;
	wire [4-1:0] node3392;
	wire [4-1:0] node3393;
	wire [4-1:0] node3396;
	wire [4-1:0] node3399;
	wire [4-1:0] node3400;
	wire [4-1:0] node3403;
	wire [4-1:0] node3406;
	wire [4-1:0] node3407;
	wire [4-1:0] node3408;
	wire [4-1:0] node3411;
	wire [4-1:0] node3414;
	wire [4-1:0] node3415;
	wire [4-1:0] node3418;
	wire [4-1:0] node3421;
	wire [4-1:0] node3422;
	wire [4-1:0] node3423;
	wire [4-1:0] node3425;
	wire [4-1:0] node3428;
	wire [4-1:0] node3429;
	wire [4-1:0] node3432;
	wire [4-1:0] node3435;
	wire [4-1:0] node3436;
	wire [4-1:0] node3437;
	wire [4-1:0] node3440;
	wire [4-1:0] node3443;
	wire [4-1:0] node3444;
	wire [4-1:0] node3447;
	wire [4-1:0] node3450;
	wire [4-1:0] node3451;
	wire [4-1:0] node3452;
	wire [4-1:0] node3453;
	wire [4-1:0] node3454;
	wire [4-1:0] node3457;
	wire [4-1:0] node3460;
	wire [4-1:0] node3461;
	wire [4-1:0] node3464;
	wire [4-1:0] node3467;
	wire [4-1:0] node3468;
	wire [4-1:0] node3469;
	wire [4-1:0] node3472;
	wire [4-1:0] node3475;
	wire [4-1:0] node3476;
	wire [4-1:0] node3479;
	wire [4-1:0] node3482;
	wire [4-1:0] node3483;
	wire [4-1:0] node3484;
	wire [4-1:0] node3485;
	wire [4-1:0] node3488;
	wire [4-1:0] node3491;
	wire [4-1:0] node3492;
	wire [4-1:0] node3495;
	wire [4-1:0] node3498;
	wire [4-1:0] node3499;
	wire [4-1:0] node3500;
	wire [4-1:0] node3503;
	wire [4-1:0] node3506;
	wire [4-1:0] node3507;
	wire [4-1:0] node3511;
	wire [4-1:0] node3512;
	wire [4-1:0] node3513;
	wire [4-1:0] node3514;
	wire [4-1:0] node3515;
	wire [4-1:0] node3516;
	wire [4-1:0] node3517;
	wire [4-1:0] node3518;
	wire [4-1:0] node3519;
	wire [4-1:0] node3520;
	wire [4-1:0] node3521;
	wire [4-1:0] node3524;
	wire [4-1:0] node3527;
	wire [4-1:0] node3528;
	wire [4-1:0] node3531;
	wire [4-1:0] node3534;
	wire [4-1:0] node3535;
	wire [4-1:0] node3538;
	wire [4-1:0] node3541;
	wire [4-1:0] node3542;
	wire [4-1:0] node3543;
	wire [4-1:0] node3544;
	wire [4-1:0] node3547;
	wire [4-1:0] node3550;
	wire [4-1:0] node3551;
	wire [4-1:0] node3554;
	wire [4-1:0] node3557;
	wire [4-1:0] node3558;
	wire [4-1:0] node3559;
	wire [4-1:0] node3562;
	wire [4-1:0] node3565;
	wire [4-1:0] node3566;
	wire [4-1:0] node3569;
	wire [4-1:0] node3572;
	wire [4-1:0] node3573;
	wire [4-1:0] node3574;
	wire [4-1:0] node3575;
	wire [4-1:0] node3576;
	wire [4-1:0] node3580;
	wire [4-1:0] node3582;
	wire [4-1:0] node3585;
	wire [4-1:0] node3586;
	wire [4-1:0] node3589;
	wire [4-1:0] node3592;
	wire [4-1:0] node3593;
	wire [4-1:0] node3594;
	wire [4-1:0] node3595;
	wire [4-1:0] node3598;
	wire [4-1:0] node3601;
	wire [4-1:0] node3602;
	wire [4-1:0] node3605;
	wire [4-1:0] node3608;
	wire [4-1:0] node3609;
	wire [4-1:0] node3610;
	wire [4-1:0] node3613;
	wire [4-1:0] node3616;
	wire [4-1:0] node3617;
	wire [4-1:0] node3620;
	wire [4-1:0] node3623;
	wire [4-1:0] node3624;
	wire [4-1:0] node3625;
	wire [4-1:0] node3626;
	wire [4-1:0] node3627;
	wire [4-1:0] node3628;
	wire [4-1:0] node3631;
	wire [4-1:0] node3634;
	wire [4-1:0] node3635;
	wire [4-1:0] node3638;
	wire [4-1:0] node3641;
	wire [4-1:0] node3642;
	wire [4-1:0] node3643;
	wire [4-1:0] node3646;
	wire [4-1:0] node3649;
	wire [4-1:0] node3651;
	wire [4-1:0] node3654;
	wire [4-1:0] node3655;
	wire [4-1:0] node3656;
	wire [4-1:0] node3657;
	wire [4-1:0] node3660;
	wire [4-1:0] node3663;
	wire [4-1:0] node3664;
	wire [4-1:0] node3667;
	wire [4-1:0] node3670;
	wire [4-1:0] node3671;
	wire [4-1:0] node3672;
	wire [4-1:0] node3675;
	wire [4-1:0] node3678;
	wire [4-1:0] node3679;
	wire [4-1:0] node3682;
	wire [4-1:0] node3685;
	wire [4-1:0] node3686;
	wire [4-1:0] node3687;
	wire [4-1:0] node3688;
	wire [4-1:0] node3689;
	wire [4-1:0] node3692;
	wire [4-1:0] node3695;
	wire [4-1:0] node3696;
	wire [4-1:0] node3699;
	wire [4-1:0] node3702;
	wire [4-1:0] node3703;
	wire [4-1:0] node3704;
	wire [4-1:0] node3707;
	wire [4-1:0] node3710;
	wire [4-1:0] node3711;
	wire [4-1:0] node3714;
	wire [4-1:0] node3717;
	wire [4-1:0] node3718;
	wire [4-1:0] node3719;
	wire [4-1:0] node3721;
	wire [4-1:0] node3724;
	wire [4-1:0] node3725;
	wire [4-1:0] node3728;
	wire [4-1:0] node3731;
	wire [4-1:0] node3732;
	wire [4-1:0] node3733;
	wire [4-1:0] node3736;
	wire [4-1:0] node3739;
	wire [4-1:0] node3740;
	wire [4-1:0] node3743;
	wire [4-1:0] node3746;
	wire [4-1:0] node3747;
	wire [4-1:0] node3748;
	wire [4-1:0] node3749;
	wire [4-1:0] node3750;
	wire [4-1:0] node3751;
	wire [4-1:0] node3752;
	wire [4-1:0] node3755;
	wire [4-1:0] node3758;
	wire [4-1:0] node3759;
	wire [4-1:0] node3762;
	wire [4-1:0] node3765;
	wire [4-1:0] node3766;
	wire [4-1:0] node3768;
	wire [4-1:0] node3771;
	wire [4-1:0] node3772;
	wire [4-1:0] node3775;
	wire [4-1:0] node3778;
	wire [4-1:0] node3779;
	wire [4-1:0] node3780;
	wire [4-1:0] node3781;
	wire [4-1:0] node3784;
	wire [4-1:0] node3787;
	wire [4-1:0] node3788;
	wire [4-1:0] node3791;
	wire [4-1:0] node3794;
	wire [4-1:0] node3795;
	wire [4-1:0] node3796;
	wire [4-1:0] node3799;
	wire [4-1:0] node3802;
	wire [4-1:0] node3803;
	wire [4-1:0] node3806;
	wire [4-1:0] node3809;
	wire [4-1:0] node3810;
	wire [4-1:0] node3811;
	wire [4-1:0] node3812;
	wire [4-1:0] node3813;
	wire [4-1:0] node3816;
	wire [4-1:0] node3819;
	wire [4-1:0] node3820;
	wire [4-1:0] node3823;
	wire [4-1:0] node3826;
	wire [4-1:0] node3827;
	wire [4-1:0] node3828;
	wire [4-1:0] node3831;
	wire [4-1:0] node3834;
	wire [4-1:0] node3835;
	wire [4-1:0] node3838;
	wire [4-1:0] node3841;
	wire [4-1:0] node3842;
	wire [4-1:0] node3843;
	wire [4-1:0] node3844;
	wire [4-1:0] node3847;
	wire [4-1:0] node3850;
	wire [4-1:0] node3851;
	wire [4-1:0] node3854;
	wire [4-1:0] node3857;
	wire [4-1:0] node3858;
	wire [4-1:0] node3859;
	wire [4-1:0] node3862;
	wire [4-1:0] node3865;
	wire [4-1:0] node3866;
	wire [4-1:0] node3869;
	wire [4-1:0] node3872;
	wire [4-1:0] node3873;
	wire [4-1:0] node3874;
	wire [4-1:0] node3875;
	wire [4-1:0] node3876;
	wire [4-1:0] node3877;
	wire [4-1:0] node3880;
	wire [4-1:0] node3883;
	wire [4-1:0] node3884;
	wire [4-1:0] node3887;
	wire [4-1:0] node3890;
	wire [4-1:0] node3891;
	wire [4-1:0] node3892;
	wire [4-1:0] node3895;
	wire [4-1:0] node3898;
	wire [4-1:0] node3899;
	wire [4-1:0] node3902;
	wire [4-1:0] node3905;
	wire [4-1:0] node3906;
	wire [4-1:0] node3907;
	wire [4-1:0] node3910;
	wire [4-1:0] node3913;
	wire [4-1:0] node3914;
	wire [4-1:0] node3915;
	wire [4-1:0] node3918;
	wire [4-1:0] node3921;
	wire [4-1:0] node3922;
	wire [4-1:0] node3925;
	wire [4-1:0] node3928;
	wire [4-1:0] node3929;
	wire [4-1:0] node3930;
	wire [4-1:0] node3931;
	wire [4-1:0] node3932;
	wire [4-1:0] node3935;
	wire [4-1:0] node3938;
	wire [4-1:0] node3939;
	wire [4-1:0] node3942;
	wire [4-1:0] node3945;
	wire [4-1:0] node3946;
	wire [4-1:0] node3947;
	wire [4-1:0] node3950;
	wire [4-1:0] node3953;
	wire [4-1:0] node3954;
	wire [4-1:0] node3957;
	wire [4-1:0] node3960;
	wire [4-1:0] node3961;
	wire [4-1:0] node3962;
	wire [4-1:0] node3964;
	wire [4-1:0] node3967;
	wire [4-1:0] node3969;
	wire [4-1:0] node3972;
	wire [4-1:0] node3973;
	wire [4-1:0] node3975;
	wire [4-1:0] node3978;
	wire [4-1:0] node3981;
	wire [4-1:0] node3982;
	wire [4-1:0] node3983;
	wire [4-1:0] node3984;
	wire [4-1:0] node3985;
	wire [4-1:0] node3986;
	wire [4-1:0] node3987;
	wire [4-1:0] node3988;
	wire [4-1:0] node3991;
	wire [4-1:0] node3994;
	wire [4-1:0] node3995;
	wire [4-1:0] node3998;
	wire [4-1:0] node4001;
	wire [4-1:0] node4002;
	wire [4-1:0] node4003;
	wire [4-1:0] node4006;
	wire [4-1:0] node4009;
	wire [4-1:0] node4010;
	wire [4-1:0] node4013;
	wire [4-1:0] node4016;
	wire [4-1:0] node4017;
	wire [4-1:0] node4018;
	wire [4-1:0] node4019;
	wire [4-1:0] node4022;
	wire [4-1:0] node4025;
	wire [4-1:0] node4026;
	wire [4-1:0] node4029;
	wire [4-1:0] node4032;
	wire [4-1:0] node4033;
	wire [4-1:0] node4034;
	wire [4-1:0] node4037;
	wire [4-1:0] node4040;
	wire [4-1:0] node4041;
	wire [4-1:0] node4044;
	wire [4-1:0] node4047;
	wire [4-1:0] node4048;
	wire [4-1:0] node4049;
	wire [4-1:0] node4050;
	wire [4-1:0] node4051;
	wire [4-1:0] node4054;
	wire [4-1:0] node4057;
	wire [4-1:0] node4058;
	wire [4-1:0] node4061;
	wire [4-1:0] node4064;
	wire [4-1:0] node4065;
	wire [4-1:0] node4066;
	wire [4-1:0] node4070;
	wire [4-1:0] node4071;
	wire [4-1:0] node4074;
	wire [4-1:0] node4077;
	wire [4-1:0] node4078;
	wire [4-1:0] node4079;
	wire [4-1:0] node4082;
	wire [4-1:0] node4085;
	wire [4-1:0] node4086;
	wire [4-1:0] node4087;
	wire [4-1:0] node4090;
	wire [4-1:0] node4093;
	wire [4-1:0] node4094;
	wire [4-1:0] node4097;
	wire [4-1:0] node4100;
	wire [4-1:0] node4101;
	wire [4-1:0] node4102;
	wire [4-1:0] node4103;
	wire [4-1:0] node4104;
	wire [4-1:0] node4105;
	wire [4-1:0] node4108;
	wire [4-1:0] node4111;
	wire [4-1:0] node4112;
	wire [4-1:0] node4116;
	wire [4-1:0] node4117;
	wire [4-1:0] node4118;
	wire [4-1:0] node4121;
	wire [4-1:0] node4124;
	wire [4-1:0] node4125;
	wire [4-1:0] node4129;
	wire [4-1:0] node4130;
	wire [4-1:0] node4131;
	wire [4-1:0] node4133;
	wire [4-1:0] node4136;
	wire [4-1:0] node4138;
	wire [4-1:0] node4141;
	wire [4-1:0] node4142;
	wire [4-1:0] node4144;
	wire [4-1:0] node4147;
	wire [4-1:0] node4149;
	wire [4-1:0] node4152;
	wire [4-1:0] node4153;
	wire [4-1:0] node4154;
	wire [4-1:0] node4155;
	wire [4-1:0] node4156;
	wire [4-1:0] node4159;
	wire [4-1:0] node4162;
	wire [4-1:0] node4163;
	wire [4-1:0] node4167;
	wire [4-1:0] node4168;
	wire [4-1:0] node4169;
	wire [4-1:0] node4172;
	wire [4-1:0] node4175;
	wire [4-1:0] node4176;
	wire [4-1:0] node4179;
	wire [4-1:0] node4182;
	wire [4-1:0] node4183;
	wire [4-1:0] node4184;
	wire [4-1:0] node4185;
	wire [4-1:0] node4188;
	wire [4-1:0] node4191;
	wire [4-1:0] node4192;
	wire [4-1:0] node4195;
	wire [4-1:0] node4198;
	wire [4-1:0] node4199;
	wire [4-1:0] node4200;
	wire [4-1:0] node4203;
	wire [4-1:0] node4206;
	wire [4-1:0] node4208;
	wire [4-1:0] node4211;
	wire [4-1:0] node4212;
	wire [4-1:0] node4213;
	wire [4-1:0] node4214;
	wire [4-1:0] node4215;
	wire [4-1:0] node4216;
	wire [4-1:0] node4217;
	wire [4-1:0] node4220;
	wire [4-1:0] node4223;
	wire [4-1:0] node4224;
	wire [4-1:0] node4227;
	wire [4-1:0] node4230;
	wire [4-1:0] node4231;
	wire [4-1:0] node4232;
	wire [4-1:0] node4235;
	wire [4-1:0] node4238;
	wire [4-1:0] node4239;
	wire [4-1:0] node4242;
	wire [4-1:0] node4245;
	wire [4-1:0] node4246;
	wire [4-1:0] node4247;
	wire [4-1:0] node4248;
	wire [4-1:0] node4251;
	wire [4-1:0] node4254;
	wire [4-1:0] node4255;
	wire [4-1:0] node4258;
	wire [4-1:0] node4261;
	wire [4-1:0] node4262;
	wire [4-1:0] node4263;
	wire [4-1:0] node4266;
	wire [4-1:0] node4269;
	wire [4-1:0] node4270;
	wire [4-1:0] node4273;
	wire [4-1:0] node4276;
	wire [4-1:0] node4277;
	wire [4-1:0] node4278;
	wire [4-1:0] node4279;
	wire [4-1:0] node4280;
	wire [4-1:0] node4284;
	wire [4-1:0] node4285;
	wire [4-1:0] node4288;
	wire [4-1:0] node4291;
	wire [4-1:0] node4292;
	wire [4-1:0] node4293;
	wire [4-1:0] node4296;
	wire [4-1:0] node4299;
	wire [4-1:0] node4300;
	wire [4-1:0] node4304;
	wire [4-1:0] node4305;
	wire [4-1:0] node4306;
	wire [4-1:0] node4309;
	wire [4-1:0] node4312;
	wire [4-1:0] node4313;
	wire [4-1:0] node4316;
	wire [4-1:0] node4319;
	wire [4-1:0] node4320;
	wire [4-1:0] node4321;
	wire [4-1:0] node4322;
	wire [4-1:0] node4323;
	wire [4-1:0] node4324;
	wire [4-1:0] node4327;
	wire [4-1:0] node4330;
	wire [4-1:0] node4331;
	wire [4-1:0] node4335;
	wire [4-1:0] node4336;
	wire [4-1:0] node4337;
	wire [4-1:0] node4341;
	wire [4-1:0] node4342;
	wire [4-1:0] node4345;
	wire [4-1:0] node4348;
	wire [4-1:0] node4349;
	wire [4-1:0] node4350;
	wire [4-1:0] node4351;
	wire [4-1:0] node4355;
	wire [4-1:0] node4356;
	wire [4-1:0] node4359;
	wire [4-1:0] node4362;
	wire [4-1:0] node4363;
	wire [4-1:0] node4364;
	wire [4-1:0] node4367;
	wire [4-1:0] node4370;
	wire [4-1:0] node4371;
	wire [4-1:0] node4374;
	wire [4-1:0] node4377;
	wire [4-1:0] node4378;
	wire [4-1:0] node4379;
	wire [4-1:0] node4380;
	wire [4-1:0] node4381;
	wire [4-1:0] node4384;
	wire [4-1:0] node4387;
	wire [4-1:0] node4388;
	wire [4-1:0] node4391;
	wire [4-1:0] node4394;
	wire [4-1:0] node4395;
	wire [4-1:0] node4396;
	wire [4-1:0] node4399;
	wire [4-1:0] node4402;
	wire [4-1:0] node4403;
	wire [4-1:0] node4406;
	wire [4-1:0] node4409;
	wire [4-1:0] node4410;
	wire [4-1:0] node4411;
	wire [4-1:0] node4412;
	wire [4-1:0] node4415;
	wire [4-1:0] node4418;
	wire [4-1:0] node4419;
	wire [4-1:0] node4422;
	wire [4-1:0] node4425;
	wire [4-1:0] node4426;
	wire [4-1:0] node4427;
	wire [4-1:0] node4430;
	wire [4-1:0] node4433;
	wire [4-1:0] node4434;
	wire [4-1:0] node4437;
	wire [4-1:0] node4440;
	wire [4-1:0] node4441;
	wire [4-1:0] node4442;
	wire [4-1:0] node4443;
	wire [4-1:0] node4444;
	wire [4-1:0] node4445;
	wire [4-1:0] node4446;
	wire [4-1:0] node4447;
	wire [4-1:0] node4448;
	wire [4-1:0] node4451;
	wire [4-1:0] node4454;
	wire [4-1:0] node4455;
	wire [4-1:0] node4458;
	wire [4-1:0] node4461;
	wire [4-1:0] node4462;
	wire [4-1:0] node4463;
	wire [4-1:0] node4466;
	wire [4-1:0] node4469;
	wire [4-1:0] node4470;
	wire [4-1:0] node4473;
	wire [4-1:0] node4476;
	wire [4-1:0] node4477;
	wire [4-1:0] node4478;
	wire [4-1:0] node4480;
	wire [4-1:0] node4483;
	wire [4-1:0] node4485;
	wire [4-1:0] node4488;
	wire [4-1:0] node4489;
	wire [4-1:0] node4491;
	wire [4-1:0] node4494;
	wire [4-1:0] node4496;
	wire [4-1:0] node4499;
	wire [4-1:0] node4500;
	wire [4-1:0] node4501;
	wire [4-1:0] node4502;
	wire [4-1:0] node4503;
	wire [4-1:0] node4506;
	wire [4-1:0] node4509;
	wire [4-1:0] node4510;
	wire [4-1:0] node4513;
	wire [4-1:0] node4516;
	wire [4-1:0] node4517;
	wire [4-1:0] node4518;
	wire [4-1:0] node4521;
	wire [4-1:0] node4524;
	wire [4-1:0] node4525;
	wire [4-1:0] node4528;
	wire [4-1:0] node4531;
	wire [4-1:0] node4532;
	wire [4-1:0] node4533;
	wire [4-1:0] node4534;
	wire [4-1:0] node4537;
	wire [4-1:0] node4540;
	wire [4-1:0] node4541;
	wire [4-1:0] node4544;
	wire [4-1:0] node4547;
	wire [4-1:0] node4548;
	wire [4-1:0] node4549;
	wire [4-1:0] node4552;
	wire [4-1:0] node4555;
	wire [4-1:0] node4556;
	wire [4-1:0] node4559;
	wire [4-1:0] node4562;
	wire [4-1:0] node4563;
	wire [4-1:0] node4564;
	wire [4-1:0] node4565;
	wire [4-1:0] node4566;
	wire [4-1:0] node4567;
	wire [4-1:0] node4570;
	wire [4-1:0] node4573;
	wire [4-1:0] node4574;
	wire [4-1:0] node4577;
	wire [4-1:0] node4580;
	wire [4-1:0] node4581;
	wire [4-1:0] node4584;
	wire [4-1:0] node4585;
	wire [4-1:0] node4589;
	wire [4-1:0] node4590;
	wire [4-1:0] node4591;
	wire [4-1:0] node4594;
	wire [4-1:0] node4597;
	wire [4-1:0] node4598;
	wire [4-1:0] node4599;
	wire [4-1:0] node4602;
	wire [4-1:0] node4605;
	wire [4-1:0] node4606;
	wire [4-1:0] node4609;
	wire [4-1:0] node4612;
	wire [4-1:0] node4613;
	wire [4-1:0] node4614;
	wire [4-1:0] node4615;
	wire [4-1:0] node4616;
	wire [4-1:0] node4619;
	wire [4-1:0] node4622;
	wire [4-1:0] node4623;
	wire [4-1:0] node4626;
	wire [4-1:0] node4629;
	wire [4-1:0] node4630;
	wire [4-1:0] node4631;
	wire [4-1:0] node4634;
	wire [4-1:0] node4637;
	wire [4-1:0] node4640;
	wire [4-1:0] node4641;
	wire [4-1:0] node4642;
	wire [4-1:0] node4644;
	wire [4-1:0] node4647;
	wire [4-1:0] node4649;
	wire [4-1:0] node4652;
	wire [4-1:0] node4653;
	wire [4-1:0] node4655;
	wire [4-1:0] node4658;
	wire [4-1:0] node4660;
	wire [4-1:0] node4663;
	wire [4-1:0] node4664;
	wire [4-1:0] node4665;
	wire [4-1:0] node4666;
	wire [4-1:0] node4667;
	wire [4-1:0] node4668;
	wire [4-1:0] node4669;
	wire [4-1:0] node4672;
	wire [4-1:0] node4675;
	wire [4-1:0] node4676;
	wire [4-1:0] node4679;
	wire [4-1:0] node4682;
	wire [4-1:0] node4683;
	wire [4-1:0] node4684;
	wire [4-1:0] node4687;
	wire [4-1:0] node4690;
	wire [4-1:0] node4691;
	wire [4-1:0] node4694;
	wire [4-1:0] node4697;
	wire [4-1:0] node4698;
	wire [4-1:0] node4699;
	wire [4-1:0] node4701;
	wire [4-1:0] node4704;
	wire [4-1:0] node4706;
	wire [4-1:0] node4709;
	wire [4-1:0] node4710;
	wire [4-1:0] node4712;
	wire [4-1:0] node4715;
	wire [4-1:0] node4717;
	wire [4-1:0] node4720;
	wire [4-1:0] node4721;
	wire [4-1:0] node4722;
	wire [4-1:0] node4723;
	wire [4-1:0] node4724;
	wire [4-1:0] node4727;
	wire [4-1:0] node4730;
	wire [4-1:0] node4731;
	wire [4-1:0] node4734;
	wire [4-1:0] node4737;
	wire [4-1:0] node4738;
	wire [4-1:0] node4739;
	wire [4-1:0] node4742;
	wire [4-1:0] node4745;
	wire [4-1:0] node4746;
	wire [4-1:0] node4750;
	wire [4-1:0] node4751;
	wire [4-1:0] node4752;
	wire [4-1:0] node4754;
	wire [4-1:0] node4757;
	wire [4-1:0] node4759;
	wire [4-1:0] node4762;
	wire [4-1:0] node4763;
	wire [4-1:0] node4765;
	wire [4-1:0] node4768;
	wire [4-1:0] node4770;
	wire [4-1:0] node4773;
	wire [4-1:0] node4774;
	wire [4-1:0] node4775;
	wire [4-1:0] node4776;
	wire [4-1:0] node4777;
	wire [4-1:0] node4778;
	wire [4-1:0] node4781;
	wire [4-1:0] node4784;
	wire [4-1:0] node4785;
	wire [4-1:0] node4788;
	wire [4-1:0] node4791;
	wire [4-1:0] node4792;
	wire [4-1:0] node4793;
	wire [4-1:0] node4797;
	wire [4-1:0] node4798;
	wire [4-1:0] node4801;
	wire [4-1:0] node4804;
	wire [4-1:0] node4805;
	wire [4-1:0] node4806;
	wire [4-1:0] node4808;
	wire [4-1:0] node4811;
	wire [4-1:0] node4813;
	wire [4-1:0] node4816;
	wire [4-1:0] node4817;
	wire [4-1:0] node4819;
	wire [4-1:0] node4822;
	wire [4-1:0] node4824;
	wire [4-1:0] node4827;
	wire [4-1:0] node4828;
	wire [4-1:0] node4829;
	wire [4-1:0] node4830;
	wire [4-1:0] node4831;
	wire [4-1:0] node4834;
	wire [4-1:0] node4837;
	wire [4-1:0] node4838;
	wire [4-1:0] node4842;
	wire [4-1:0] node4843;
	wire [4-1:0] node4844;
	wire [4-1:0] node4847;
	wire [4-1:0] node4850;
	wire [4-1:0] node4851;
	wire [4-1:0] node4854;
	wire [4-1:0] node4857;
	wire [4-1:0] node4858;
	wire [4-1:0] node4859;
	wire [4-1:0] node4862;
	wire [4-1:0] node4865;
	wire [4-1:0] node4866;
	wire [4-1:0] node4867;
	wire [4-1:0] node4870;
	wire [4-1:0] node4873;
	wire [4-1:0] node4874;
	wire [4-1:0] node4877;
	wire [4-1:0] node4880;
	wire [4-1:0] node4881;
	wire [4-1:0] node4882;
	wire [4-1:0] node4883;
	wire [4-1:0] node4884;
	wire [4-1:0] node4885;
	wire [4-1:0] node4886;
	wire [4-1:0] node4887;
	wire [4-1:0] node4890;
	wire [4-1:0] node4893;
	wire [4-1:0] node4895;
	wire [4-1:0] node4898;
	wire [4-1:0] node4899;
	wire [4-1:0] node4900;
	wire [4-1:0] node4904;
	wire [4-1:0] node4905;
	wire [4-1:0] node4908;
	wire [4-1:0] node4911;
	wire [4-1:0] node4912;
	wire [4-1:0] node4913;
	wire [4-1:0] node4914;
	wire [4-1:0] node4917;
	wire [4-1:0] node4920;
	wire [4-1:0] node4921;
	wire [4-1:0] node4924;
	wire [4-1:0] node4927;
	wire [4-1:0] node4928;
	wire [4-1:0] node4929;
	wire [4-1:0] node4932;
	wire [4-1:0] node4935;
	wire [4-1:0] node4936;
	wire [4-1:0] node4939;
	wire [4-1:0] node4942;
	wire [4-1:0] node4943;
	wire [4-1:0] node4944;
	wire [4-1:0] node4945;
	wire [4-1:0] node4946;
	wire [4-1:0] node4949;
	wire [4-1:0] node4952;
	wire [4-1:0] node4953;
	wire [4-1:0] node4957;
	wire [4-1:0] node4958;
	wire [4-1:0] node4959;
	wire [4-1:0] node4962;
	wire [4-1:0] node4965;
	wire [4-1:0] node4966;
	wire [4-1:0] node4969;
	wire [4-1:0] node4972;
	wire [4-1:0] node4973;
	wire [4-1:0] node4974;
	wire [4-1:0] node4976;
	wire [4-1:0] node4979;
	wire [4-1:0] node4981;
	wire [4-1:0] node4984;
	wire [4-1:0] node4985;
	wire [4-1:0] node4987;
	wire [4-1:0] node4990;
	wire [4-1:0] node4992;
	wire [4-1:0] node4995;
	wire [4-1:0] node4996;
	wire [4-1:0] node4997;
	wire [4-1:0] node4998;
	wire [4-1:0] node4999;
	wire [4-1:0] node5000;
	wire [4-1:0] node5003;
	wire [4-1:0] node5006;
	wire [4-1:0] node5007;
	wire [4-1:0] node5010;
	wire [4-1:0] node5013;
	wire [4-1:0] node5014;
	wire [4-1:0] node5016;
	wire [4-1:0] node5019;
	wire [4-1:0] node5020;
	wire [4-1:0] node5023;
	wire [4-1:0] node5026;
	wire [4-1:0] node5027;
	wire [4-1:0] node5028;
	wire [4-1:0] node5030;
	wire [4-1:0] node5033;
	wire [4-1:0] node5035;
	wire [4-1:0] node5038;
	wire [4-1:0] node5039;
	wire [4-1:0] node5041;
	wire [4-1:0] node5044;
	wire [4-1:0] node5046;
	wire [4-1:0] node5049;
	wire [4-1:0] node5050;
	wire [4-1:0] node5051;
	wire [4-1:0] node5052;
	wire [4-1:0] node5053;
	wire [4-1:0] node5056;
	wire [4-1:0] node5059;
	wire [4-1:0] node5060;
	wire [4-1:0] node5063;
	wire [4-1:0] node5066;
	wire [4-1:0] node5067;
	wire [4-1:0] node5069;
	wire [4-1:0] node5072;
	wire [4-1:0] node5073;
	wire [4-1:0] node5076;
	wire [4-1:0] node5079;
	wire [4-1:0] node5080;
	wire [4-1:0] node5081;
	wire [4-1:0] node5084;
	wire [4-1:0] node5087;
	wire [4-1:0] node5088;
	wire [4-1:0] node5089;
	wire [4-1:0] node5093;
	wire [4-1:0] node5094;
	wire [4-1:0] node5097;
	wire [4-1:0] node5100;
	wire [4-1:0] node5101;
	wire [4-1:0] node5102;
	wire [4-1:0] node5103;
	wire [4-1:0] node5104;
	wire [4-1:0] node5105;
	wire [4-1:0] node5106;
	wire [4-1:0] node5109;
	wire [4-1:0] node5112;
	wire [4-1:0] node5113;
	wire [4-1:0] node5116;
	wire [4-1:0] node5119;
	wire [4-1:0] node5120;
	wire [4-1:0] node5121;
	wire [4-1:0] node5124;
	wire [4-1:0] node5127;
	wire [4-1:0] node5128;
	wire [4-1:0] node5132;
	wire [4-1:0] node5133;
	wire [4-1:0] node5134;
	wire [4-1:0] node5135;
	wire [4-1:0] node5138;
	wire [4-1:0] node5141;
	wire [4-1:0] node5142;
	wire [4-1:0] node5145;
	wire [4-1:0] node5148;
	wire [4-1:0] node5149;
	wire [4-1:0] node5152;
	wire [4-1:0] node5155;
	wire [4-1:0] node5156;
	wire [4-1:0] node5157;
	wire [4-1:0] node5158;
	wire [4-1:0] node5159;
	wire [4-1:0] node5162;
	wire [4-1:0] node5165;
	wire [4-1:0] node5166;
	wire [4-1:0] node5169;
	wire [4-1:0] node5172;
	wire [4-1:0] node5173;
	wire [4-1:0] node5176;
	wire [4-1:0] node5179;
	wire [4-1:0] node5180;
	wire [4-1:0] node5181;
	wire [4-1:0] node5182;
	wire [4-1:0] node5185;
	wire [4-1:0] node5188;
	wire [4-1:0] node5189;
	wire [4-1:0] node5193;
	wire [4-1:0] node5194;
	wire [4-1:0] node5195;
	wire [4-1:0] node5198;
	wire [4-1:0] node5201;
	wire [4-1:0] node5202;
	wire [4-1:0] node5205;
	wire [4-1:0] node5208;
	wire [4-1:0] node5209;
	wire [4-1:0] node5210;
	wire [4-1:0] node5211;
	wire [4-1:0] node5212;
	wire [4-1:0] node5213;
	wire [4-1:0] node5216;
	wire [4-1:0] node5219;
	wire [4-1:0] node5220;
	wire [4-1:0] node5223;
	wire [4-1:0] node5226;
	wire [4-1:0] node5227;
	wire [4-1:0] node5228;
	wire [4-1:0] node5231;
	wire [4-1:0] node5234;
	wire [4-1:0] node5235;
	wire [4-1:0] node5239;
	wire [4-1:0] node5240;
	wire [4-1:0] node5241;
	wire [4-1:0] node5243;
	wire [4-1:0] node5246;
	wire [4-1:0] node5247;
	wire [4-1:0] node5250;
	wire [4-1:0] node5253;
	wire [4-1:0] node5254;
	wire [4-1:0] node5255;
	wire [4-1:0] node5258;
	wire [4-1:0] node5261;
	wire [4-1:0] node5262;
	wire [4-1:0] node5265;
	wire [4-1:0] node5268;
	wire [4-1:0] node5269;
	wire [4-1:0] node5270;
	wire [4-1:0] node5271;
	wire [4-1:0] node5272;
	wire [4-1:0] node5275;
	wire [4-1:0] node5278;
	wire [4-1:0] node5280;
	wire [4-1:0] node5283;
	wire [4-1:0] node5284;
	wire [4-1:0] node5285;
	wire [4-1:0] node5288;
	wire [4-1:0] node5291;
	wire [4-1:0] node5293;
	wire [4-1:0] node5296;
	wire [4-1:0] node5297;
	wire [4-1:0] node5298;
	wire [4-1:0] node5299;
	wire [4-1:0] node5302;
	wire [4-1:0] node5305;
	wire [4-1:0] node5306;
	wire [4-1:0] node5309;
	wire [4-1:0] node5312;
	wire [4-1:0] node5313;
	wire [4-1:0] node5314;
	wire [4-1:0] node5317;
	wire [4-1:0] node5320;
	wire [4-1:0] node5321;
	wire [4-1:0] node5324;
	wire [4-1:0] node5327;
	wire [4-1:0] node5328;
	wire [4-1:0] node5329;
	wire [4-1:0] node5330;
	wire [4-1:0] node5331;
	wire [4-1:0] node5332;
	wire [4-1:0] node5333;
	wire [4-1:0] node5334;
	wire [4-1:0] node5336;
	wire [4-1:0] node5337;
	wire [4-1:0] node5340;
	wire [4-1:0] node5343;
	wire [4-1:0] node5344;
	wire [4-1:0] node5345;
	wire [4-1:0] node5348;
	wire [4-1:0] node5351;
	wire [4-1:0] node5352;
	wire [4-1:0] node5355;
	wire [4-1:0] node5358;
	wire [4-1:0] node5359;
	wire [4-1:0] node5360;
	wire [4-1:0] node5361;
	wire [4-1:0] node5365;
	wire [4-1:0] node5366;
	wire [4-1:0] node5369;
	wire [4-1:0] node5372;
	wire [4-1:0] node5373;
	wire [4-1:0] node5374;
	wire [4-1:0] node5377;
	wire [4-1:0] node5380;
	wire [4-1:0] node5381;
	wire [4-1:0] node5384;
	wire [4-1:0] node5387;
	wire [4-1:0] node5388;
	wire [4-1:0] node5389;
	wire [4-1:0] node5390;
	wire [4-1:0] node5391;
	wire [4-1:0] node5395;
	wire [4-1:0] node5396;
	wire [4-1:0] node5400;
	wire [4-1:0] node5401;
	wire [4-1:0] node5402;
	wire [4-1:0] node5406;
	wire [4-1:0] node5407;
	wire [4-1:0] node5411;
	wire [4-1:0] node5412;
	wire [4-1:0] node5413;
	wire [4-1:0] node5414;
	wire [4-1:0] node5417;
	wire [4-1:0] node5420;
	wire [4-1:0] node5421;
	wire [4-1:0] node5424;
	wire [4-1:0] node5427;
	wire [4-1:0] node5428;
	wire [4-1:0] node5429;
	wire [4-1:0] node5432;
	wire [4-1:0] node5435;
	wire [4-1:0] node5436;
	wire [4-1:0] node5439;
	wire [4-1:0] node5442;
	wire [4-1:0] node5443;
	wire [4-1:0] node5444;
	wire [4-1:0] node5445;
	wire [4-1:0] node5446;
	wire [4-1:0] node5447;
	wire [4-1:0] node5451;
	wire [4-1:0] node5452;
	wire [4-1:0] node5456;
	wire [4-1:0] node5457;
	wire [4-1:0] node5458;
	wire [4-1:0] node5462;
	wire [4-1:0] node5463;
	wire [4-1:0] node5467;
	wire [4-1:0] node5468;
	wire [4-1:0] node5469;
	wire [4-1:0] node5470;
	wire [4-1:0] node5473;
	wire [4-1:0] node5476;
	wire [4-1:0] node5478;
	wire [4-1:0] node5481;
	wire [4-1:0] node5482;
	wire [4-1:0] node5483;
	wire [4-1:0] node5486;
	wire [4-1:0] node5489;
	wire [4-1:0] node5490;
	wire [4-1:0] node5493;
	wire [4-1:0] node5496;
	wire [4-1:0] node5497;
	wire [4-1:0] node5498;
	wire [4-1:0] node5499;
	wire [4-1:0] node5500;
	wire [4-1:0] node5503;
	wire [4-1:0] node5506;
	wire [4-1:0] node5507;
	wire [4-1:0] node5510;
	wire [4-1:0] node5513;
	wire [4-1:0] node5514;
	wire [4-1:0] node5517;
	wire [4-1:0] node5520;
	wire [4-1:0] node5521;
	wire [4-1:0] node5522;
	wire [4-1:0] node5523;
	wire [4-1:0] node5526;
	wire [4-1:0] node5529;
	wire [4-1:0] node5530;
	wire [4-1:0] node5533;
	wire [4-1:0] node5536;
	wire [4-1:0] node5537;
	wire [4-1:0] node5538;
	wire [4-1:0] node5542;
	wire [4-1:0] node5543;
	wire [4-1:0] node5546;
	wire [4-1:0] node5549;
	wire [4-1:0] node5550;
	wire [4-1:0] node5551;
	wire [4-1:0] node5552;
	wire [4-1:0] node5553;
	wire [4-1:0] node5554;
	wire [4-1:0] node5556;
	wire [4-1:0] node5559;
	wire [4-1:0] node5561;
	wire [4-1:0] node5564;
	wire [4-1:0] node5565;
	wire [4-1:0] node5566;
	wire [4-1:0] node5569;
	wire [4-1:0] node5572;
	wire [4-1:0] node5573;
	wire [4-1:0] node5576;
	wire [4-1:0] node5579;
	wire [4-1:0] node5580;
	wire [4-1:0] node5581;
	wire [4-1:0] node5583;
	wire [4-1:0] node5586;
	wire [4-1:0] node5588;
	wire [4-1:0] node5591;
	wire [4-1:0] node5592;
	wire [4-1:0] node5594;
	wire [4-1:0] node5597;
	wire [4-1:0] node5599;
	wire [4-1:0] node5602;
	wire [4-1:0] node5603;
	wire [4-1:0] node5604;
	wire [4-1:0] node5605;
	wire [4-1:0] node5606;
	wire [4-1:0] node5609;
	wire [4-1:0] node5612;
	wire [4-1:0] node5613;
	wire [4-1:0] node5616;
	wire [4-1:0] node5619;
	wire [4-1:0] node5620;
	wire [4-1:0] node5621;
	wire [4-1:0] node5624;
	wire [4-1:0] node5627;
	wire [4-1:0] node5629;
	wire [4-1:0] node5632;
	wire [4-1:0] node5633;
	wire [4-1:0] node5634;
	wire [4-1:0] node5637;
	wire [4-1:0] node5640;
	wire [4-1:0] node5641;
	wire [4-1:0] node5642;
	wire [4-1:0] node5645;
	wire [4-1:0] node5648;
	wire [4-1:0] node5649;
	wire [4-1:0] node5652;
	wire [4-1:0] node5655;
	wire [4-1:0] node5656;
	wire [4-1:0] node5657;
	wire [4-1:0] node5658;
	wire [4-1:0] node5659;
	wire [4-1:0] node5660;
	wire [4-1:0] node5663;
	wire [4-1:0] node5666;
	wire [4-1:0] node5667;
	wire [4-1:0] node5670;
	wire [4-1:0] node5673;
	wire [4-1:0] node5674;
	wire [4-1:0] node5675;
	wire [4-1:0] node5678;
	wire [4-1:0] node5681;
	wire [4-1:0] node5683;
	wire [4-1:0] node5686;
	wire [4-1:0] node5687;
	wire [4-1:0] node5688;
	wire [4-1:0] node5690;
	wire [4-1:0] node5693;
	wire [4-1:0] node5695;
	wire [4-1:0] node5698;
	wire [4-1:0] node5699;
	wire [4-1:0] node5701;
	wire [4-1:0] node5704;
	wire [4-1:0] node5706;
	wire [4-1:0] node5709;
	wire [4-1:0] node5710;
	wire [4-1:0] node5711;
	wire [4-1:0] node5712;
	wire [4-1:0] node5714;
	wire [4-1:0] node5717;
	wire [4-1:0] node5718;
	wire [4-1:0] node5721;
	wire [4-1:0] node5724;
	wire [4-1:0] node5725;
	wire [4-1:0] node5726;
	wire [4-1:0] node5729;
	wire [4-1:0] node5732;
	wire [4-1:0] node5733;
	wire [4-1:0] node5736;
	wire [4-1:0] node5739;
	wire [4-1:0] node5740;
	wire [4-1:0] node5741;
	wire [4-1:0] node5742;
	wire [4-1:0] node5745;
	wire [4-1:0] node5748;
	wire [4-1:0] node5749;
	wire [4-1:0] node5752;
	wire [4-1:0] node5755;
	wire [4-1:0] node5756;
	wire [4-1:0] node5757;
	wire [4-1:0] node5760;
	wire [4-1:0] node5763;
	wire [4-1:0] node5764;
	wire [4-1:0] node5767;
	wire [4-1:0] node5770;
	wire [4-1:0] node5771;
	wire [4-1:0] node5772;
	wire [4-1:0] node5773;
	wire [4-1:0] node5774;
	wire [4-1:0] node5775;
	wire [4-1:0] node5776;
	wire [4-1:0] node5777;
	wire [4-1:0] node5780;
	wire [4-1:0] node5783;
	wire [4-1:0] node5784;
	wire [4-1:0] node5787;
	wire [4-1:0] node5790;
	wire [4-1:0] node5791;
	wire [4-1:0] node5792;
	wire [4-1:0] node5795;
	wire [4-1:0] node5798;
	wire [4-1:0] node5799;
	wire [4-1:0] node5802;
	wire [4-1:0] node5805;
	wire [4-1:0] node5806;
	wire [4-1:0] node5807;
	wire [4-1:0] node5809;
	wire [4-1:0] node5812;
	wire [4-1:0] node5814;
	wire [4-1:0] node5817;
	wire [4-1:0] node5818;
	wire [4-1:0] node5820;
	wire [4-1:0] node5823;
	wire [4-1:0] node5825;
	wire [4-1:0] node5828;
	wire [4-1:0] node5829;
	wire [4-1:0] node5830;
	wire [4-1:0] node5831;
	wire [4-1:0] node5832;
	wire [4-1:0] node5835;
	wire [4-1:0] node5838;
	wire [4-1:0] node5839;
	wire [4-1:0] node5842;
	wire [4-1:0] node5845;
	wire [4-1:0] node5846;
	wire [4-1:0] node5848;
	wire [4-1:0] node5851;
	wire [4-1:0] node5852;
	wire [4-1:0] node5856;
	wire [4-1:0] node5857;
	wire [4-1:0] node5858;
	wire [4-1:0] node5859;
	wire [4-1:0] node5862;
	wire [4-1:0] node5865;
	wire [4-1:0] node5866;
	wire [4-1:0] node5869;
	wire [4-1:0] node5872;
	wire [4-1:0] node5873;
	wire [4-1:0] node5874;
	wire [4-1:0] node5877;
	wire [4-1:0] node5880;
	wire [4-1:0] node5881;
	wire [4-1:0] node5884;
	wire [4-1:0] node5887;
	wire [4-1:0] node5888;
	wire [4-1:0] node5889;
	wire [4-1:0] node5890;
	wire [4-1:0] node5891;
	wire [4-1:0] node5893;
	wire [4-1:0] node5896;
	wire [4-1:0] node5897;
	wire [4-1:0] node5900;
	wire [4-1:0] node5903;
	wire [4-1:0] node5904;
	wire [4-1:0] node5905;
	wire [4-1:0] node5908;
	wire [4-1:0] node5911;
	wire [4-1:0] node5912;
	wire [4-1:0] node5915;
	wire [4-1:0] node5918;
	wire [4-1:0] node5919;
	wire [4-1:0] node5920;
	wire [4-1:0] node5921;
	wire [4-1:0] node5924;
	wire [4-1:0] node5927;
	wire [4-1:0] node5928;
	wire [4-1:0] node5931;
	wire [4-1:0] node5934;
	wire [4-1:0] node5935;
	wire [4-1:0] node5936;
	wire [4-1:0] node5939;
	wire [4-1:0] node5942;
	wire [4-1:0] node5943;
	wire [4-1:0] node5946;
	wire [4-1:0] node5949;
	wire [4-1:0] node5950;
	wire [4-1:0] node5951;
	wire [4-1:0] node5952;
	wire [4-1:0] node5953;
	wire [4-1:0] node5956;
	wire [4-1:0] node5959;
	wire [4-1:0] node5960;
	wire [4-1:0] node5963;
	wire [4-1:0] node5966;
	wire [4-1:0] node5967;
	wire [4-1:0] node5968;
	wire [4-1:0] node5971;
	wire [4-1:0] node5974;
	wire [4-1:0] node5976;
	wire [4-1:0] node5979;
	wire [4-1:0] node5980;
	wire [4-1:0] node5981;
	wire [4-1:0] node5982;
	wire [4-1:0] node5985;
	wire [4-1:0] node5988;
	wire [4-1:0] node5989;
	wire [4-1:0] node5992;
	wire [4-1:0] node5995;
	wire [4-1:0] node5996;
	wire [4-1:0] node5997;
	wire [4-1:0] node6001;
	wire [4-1:0] node6002;
	wire [4-1:0] node6005;
	wire [4-1:0] node6008;
	wire [4-1:0] node6009;
	wire [4-1:0] node6010;
	wire [4-1:0] node6011;
	wire [4-1:0] node6012;
	wire [4-1:0] node6013;
	wire [4-1:0] node6015;
	wire [4-1:0] node6018;
	wire [4-1:0] node6019;
	wire [4-1:0] node6022;
	wire [4-1:0] node6025;
	wire [4-1:0] node6026;
	wire [4-1:0] node6029;
	wire [4-1:0] node6030;
	wire [4-1:0] node6033;
	wire [4-1:0] node6036;
	wire [4-1:0] node6037;
	wire [4-1:0] node6038;
	wire [4-1:0] node6041;
	wire [4-1:0] node6043;
	wire [4-1:0] node6046;
	wire [4-1:0] node6047;
	wire [4-1:0] node6048;
	wire [4-1:0] node6051;
	wire [4-1:0] node6054;
	wire [4-1:0] node6056;
	wire [4-1:0] node6059;
	wire [4-1:0] node6060;
	wire [4-1:0] node6061;
	wire [4-1:0] node6062;
	wire [4-1:0] node6064;
	wire [4-1:0] node6067;
	wire [4-1:0] node6068;
	wire [4-1:0] node6071;
	wire [4-1:0] node6074;
	wire [4-1:0] node6075;
	wire [4-1:0] node6077;
	wire [4-1:0] node6080;
	wire [4-1:0] node6081;
	wire [4-1:0] node6084;
	wire [4-1:0] node6087;
	wire [4-1:0] node6088;
	wire [4-1:0] node6089;
	wire [4-1:0] node6090;
	wire [4-1:0] node6093;
	wire [4-1:0] node6096;
	wire [4-1:0] node6097;
	wire [4-1:0] node6100;
	wire [4-1:0] node6103;
	wire [4-1:0] node6104;
	wire [4-1:0] node6105;
	wire [4-1:0] node6108;
	wire [4-1:0] node6111;
	wire [4-1:0] node6112;
	wire [4-1:0] node6115;
	wire [4-1:0] node6118;
	wire [4-1:0] node6119;
	wire [4-1:0] node6120;
	wire [4-1:0] node6121;
	wire [4-1:0] node6122;
	wire [4-1:0] node6123;
	wire [4-1:0] node6126;
	wire [4-1:0] node6129;
	wire [4-1:0] node6130;
	wire [4-1:0] node6133;
	wire [4-1:0] node6136;
	wire [4-1:0] node6137;
	wire [4-1:0] node6138;
	wire [4-1:0] node6142;
	wire [4-1:0] node6143;
	wire [4-1:0] node6146;
	wire [4-1:0] node6149;
	wire [4-1:0] node6150;
	wire [4-1:0] node6151;
	wire [4-1:0] node6153;
	wire [4-1:0] node6156;
	wire [4-1:0] node6158;
	wire [4-1:0] node6161;
	wire [4-1:0] node6162;
	wire [4-1:0] node6164;
	wire [4-1:0] node6167;
	wire [4-1:0] node6169;
	wire [4-1:0] node6172;
	wire [4-1:0] node6173;
	wire [4-1:0] node6174;
	wire [4-1:0] node6175;
	wire [4-1:0] node6176;
	wire [4-1:0] node6179;
	wire [4-1:0] node6182;
	wire [4-1:0] node6183;
	wire [4-1:0] node6186;
	wire [4-1:0] node6189;
	wire [4-1:0] node6190;
	wire [4-1:0] node6191;
	wire [4-1:0] node6194;
	wire [4-1:0] node6197;
	wire [4-1:0] node6198;
	wire [4-1:0] node6201;
	wire [4-1:0] node6204;
	wire [4-1:0] node6205;
	wire [4-1:0] node6206;
	wire [4-1:0] node6207;
	wire [4-1:0] node6210;
	wire [4-1:0] node6213;
	wire [4-1:0] node6214;
	wire [4-1:0] node6217;
	wire [4-1:0] node6220;
	wire [4-1:0] node6221;
	wire [4-1:0] node6222;
	wire [4-1:0] node6225;
	wire [4-1:0] node6228;
	wire [4-1:0] node6229;
	wire [4-1:0] node6233;
	wire [4-1:0] node6234;
	wire [4-1:0] node6235;
	wire [4-1:0] node6236;
	wire [4-1:0] node6237;
	wire [4-1:0] node6238;
	wire [4-1:0] node6239;
	wire [4-1:0] node6240;
	wire [4-1:0] node6241;
	wire [4-1:0] node6244;
	wire [4-1:0] node6247;
	wire [4-1:0] node6248;
	wire [4-1:0] node6251;
	wire [4-1:0] node6254;
	wire [4-1:0] node6255;
	wire [4-1:0] node6256;
	wire [4-1:0] node6259;
	wire [4-1:0] node6262;
	wire [4-1:0] node6263;
	wire [4-1:0] node6266;
	wire [4-1:0] node6269;
	wire [4-1:0] node6270;
	wire [4-1:0] node6271;
	wire [4-1:0] node6272;
	wire [4-1:0] node6275;
	wire [4-1:0] node6278;
	wire [4-1:0] node6279;
	wire [4-1:0] node6282;
	wire [4-1:0] node6285;
	wire [4-1:0] node6286;
	wire [4-1:0] node6287;
	wire [4-1:0] node6290;
	wire [4-1:0] node6293;
	wire [4-1:0] node6294;
	wire [4-1:0] node6297;
	wire [4-1:0] node6300;
	wire [4-1:0] node6301;
	wire [4-1:0] node6302;
	wire [4-1:0] node6303;
	wire [4-1:0] node6306;
	wire [4-1:0] node6309;
	wire [4-1:0] node6310;
	wire [4-1:0] node6313;
	wire [4-1:0] node6316;
	wire [4-1:0] node6317;
	wire [4-1:0] node6318;
	wire [4-1:0] node6321;
	wire [4-1:0] node6324;
	wire [4-1:0] node6325;
	wire [4-1:0] node6328;
	wire [4-1:0] node6331;
	wire [4-1:0] node6332;
	wire [4-1:0] node6333;
	wire [4-1:0] node6334;
	wire [4-1:0] node6335;
	wire [4-1:0] node6336;
	wire [4-1:0] node6339;
	wire [4-1:0] node6342;
	wire [4-1:0] node6343;
	wire [4-1:0] node6346;
	wire [4-1:0] node6349;
	wire [4-1:0] node6350;
	wire [4-1:0] node6351;
	wire [4-1:0] node6354;
	wire [4-1:0] node6357;
	wire [4-1:0] node6358;
	wire [4-1:0] node6361;
	wire [4-1:0] node6364;
	wire [4-1:0] node6365;
	wire [4-1:0] node6366;
	wire [4-1:0] node6367;
	wire [4-1:0] node6370;
	wire [4-1:0] node6373;
	wire [4-1:0] node6374;
	wire [4-1:0] node6377;
	wire [4-1:0] node6380;
	wire [4-1:0] node6381;
	wire [4-1:0] node6382;
	wire [4-1:0] node6385;
	wire [4-1:0] node6388;
	wire [4-1:0] node6389;
	wire [4-1:0] node6393;
	wire [4-1:0] node6394;
	wire [4-1:0] node6395;
	wire [4-1:0] node6396;
	wire [4-1:0] node6397;
	wire [4-1:0] node6400;
	wire [4-1:0] node6403;
	wire [4-1:0] node6404;
	wire [4-1:0] node6407;
	wire [4-1:0] node6410;
	wire [4-1:0] node6411;
	wire [4-1:0] node6412;
	wire [4-1:0] node6415;
	wire [4-1:0] node6418;
	wire [4-1:0] node6419;
	wire [4-1:0] node6423;
	wire [4-1:0] node6424;
	wire [4-1:0] node6425;
	wire [4-1:0] node6426;
	wire [4-1:0] node6429;
	wire [4-1:0] node6432;
	wire [4-1:0] node6433;
	wire [4-1:0] node6436;
	wire [4-1:0] node6439;
	wire [4-1:0] node6440;
	wire [4-1:0] node6441;
	wire [4-1:0] node6444;
	wire [4-1:0] node6447;
	wire [4-1:0] node6448;
	wire [4-1:0] node6451;
	wire [4-1:0] node6454;
	wire [4-1:0] node6455;
	wire [4-1:0] node6456;
	wire [4-1:0] node6457;
	wire [4-1:0] node6458;
	wire [4-1:0] node6459;
	wire [4-1:0] node6461;
	wire [4-1:0] node6464;
	wire [4-1:0] node6465;
	wire [4-1:0] node6468;
	wire [4-1:0] node6471;
	wire [4-1:0] node6472;
	wire [4-1:0] node6473;
	wire [4-1:0] node6476;
	wire [4-1:0] node6479;
	wire [4-1:0] node6480;
	wire [4-1:0] node6483;
	wire [4-1:0] node6486;
	wire [4-1:0] node6487;
	wire [4-1:0] node6488;
	wire [4-1:0] node6489;
	wire [4-1:0] node6492;
	wire [4-1:0] node6495;
	wire [4-1:0] node6496;
	wire [4-1:0] node6500;
	wire [4-1:0] node6501;
	wire [4-1:0] node6502;
	wire [4-1:0] node6505;
	wire [4-1:0] node6508;
	wire [4-1:0] node6509;
	wire [4-1:0] node6512;
	wire [4-1:0] node6515;
	wire [4-1:0] node6516;
	wire [4-1:0] node6517;
	wire [4-1:0] node6518;
	wire [4-1:0] node6519;
	wire [4-1:0] node6522;
	wire [4-1:0] node6525;
	wire [4-1:0] node6526;
	wire [4-1:0] node6529;
	wire [4-1:0] node6532;
	wire [4-1:0] node6533;
	wire [4-1:0] node6535;
	wire [4-1:0] node6538;
	wire [4-1:0] node6540;
	wire [4-1:0] node6543;
	wire [4-1:0] node6544;
	wire [4-1:0] node6545;
	wire [4-1:0] node6546;
	wire [4-1:0] node6549;
	wire [4-1:0] node6552;
	wire [4-1:0] node6553;
	wire [4-1:0] node6557;
	wire [4-1:0] node6558;
	wire [4-1:0] node6559;
	wire [4-1:0] node6562;
	wire [4-1:0] node6565;
	wire [4-1:0] node6566;
	wire [4-1:0] node6569;
	wire [4-1:0] node6572;
	wire [4-1:0] node6573;
	wire [4-1:0] node6574;
	wire [4-1:0] node6575;
	wire [4-1:0] node6576;
	wire [4-1:0] node6577;
	wire [4-1:0] node6580;
	wire [4-1:0] node6583;
	wire [4-1:0] node6584;
	wire [4-1:0] node6587;
	wire [4-1:0] node6590;
	wire [4-1:0] node6591;
	wire [4-1:0] node6592;
	wire [4-1:0] node6595;
	wire [4-1:0] node6598;
	wire [4-1:0] node6600;
	wire [4-1:0] node6603;
	wire [4-1:0] node6604;
	wire [4-1:0] node6605;
	wire [4-1:0] node6606;
	wire [4-1:0] node6609;
	wire [4-1:0] node6612;
	wire [4-1:0] node6613;
	wire [4-1:0] node6616;
	wire [4-1:0] node6619;
	wire [4-1:0] node6620;
	wire [4-1:0] node6621;
	wire [4-1:0] node6624;
	wire [4-1:0] node6627;
	wire [4-1:0] node6628;
	wire [4-1:0] node6631;
	wire [4-1:0] node6634;
	wire [4-1:0] node6635;
	wire [4-1:0] node6636;
	wire [4-1:0] node6637;
	wire [4-1:0] node6638;
	wire [4-1:0] node6641;
	wire [4-1:0] node6644;
	wire [4-1:0] node6645;
	wire [4-1:0] node6649;
	wire [4-1:0] node6650;
	wire [4-1:0] node6651;
	wire [4-1:0] node6654;
	wire [4-1:0] node6657;
	wire [4-1:0] node6658;
	wire [4-1:0] node6661;
	wire [4-1:0] node6664;
	wire [4-1:0] node6665;
	wire [4-1:0] node6666;
	wire [4-1:0] node6667;
	wire [4-1:0] node6670;
	wire [4-1:0] node6673;
	wire [4-1:0] node6674;
	wire [4-1:0] node6677;
	wire [4-1:0] node6680;
	wire [4-1:0] node6681;
	wire [4-1:0] node6682;
	wire [4-1:0] node6685;
	wire [4-1:0] node6688;
	wire [4-1:0] node6690;
	wire [4-1:0] node6693;
	wire [4-1:0] node6694;
	wire [4-1:0] node6695;
	wire [4-1:0] node6696;
	wire [4-1:0] node6697;
	wire [4-1:0] node6698;
	wire [4-1:0] node6699;
	wire [4-1:0] node6700;
	wire [4-1:0] node6703;
	wire [4-1:0] node6706;
	wire [4-1:0] node6707;
	wire [4-1:0] node6710;
	wire [4-1:0] node6713;
	wire [4-1:0] node6714;
	wire [4-1:0] node6715;
	wire [4-1:0] node6718;
	wire [4-1:0] node6721;
	wire [4-1:0] node6722;
	wire [4-1:0] node6725;
	wire [4-1:0] node6728;
	wire [4-1:0] node6729;
	wire [4-1:0] node6730;
	wire [4-1:0] node6733;
	wire [4-1:0] node6736;
	wire [4-1:0] node6737;
	wire [4-1:0] node6739;
	wire [4-1:0] node6742;
	wire [4-1:0] node6743;
	wire [4-1:0] node6746;
	wire [4-1:0] node6749;
	wire [4-1:0] node6750;
	wire [4-1:0] node6751;
	wire [4-1:0] node6752;
	wire [4-1:0] node6753;
	wire [4-1:0] node6757;
	wire [4-1:0] node6758;
	wire [4-1:0] node6762;
	wire [4-1:0] node6763;
	wire [4-1:0] node6764;
	wire [4-1:0] node6768;
	wire [4-1:0] node6769;
	wire [4-1:0] node6772;
	wire [4-1:0] node6775;
	wire [4-1:0] node6776;
	wire [4-1:0] node6777;
	wire [4-1:0] node6778;
	wire [4-1:0] node6781;
	wire [4-1:0] node6784;
	wire [4-1:0] node6785;
	wire [4-1:0] node6788;
	wire [4-1:0] node6791;
	wire [4-1:0] node6792;
	wire [4-1:0] node6794;
	wire [4-1:0] node6797;
	wire [4-1:0] node6798;
	wire [4-1:0] node6801;
	wire [4-1:0] node6804;
	wire [4-1:0] node6805;
	wire [4-1:0] node6806;
	wire [4-1:0] node6807;
	wire [4-1:0] node6808;
	wire [4-1:0] node6809;
	wire [4-1:0] node6812;
	wire [4-1:0] node6815;
	wire [4-1:0] node6816;
	wire [4-1:0] node6819;
	wire [4-1:0] node6822;
	wire [4-1:0] node6823;
	wire [4-1:0] node6824;
	wire [4-1:0] node6827;
	wire [4-1:0] node6830;
	wire [4-1:0] node6831;
	wire [4-1:0] node6834;
	wire [4-1:0] node6837;
	wire [4-1:0] node6838;
	wire [4-1:0] node6839;
	wire [4-1:0] node6841;
	wire [4-1:0] node6844;
	wire [4-1:0] node6846;
	wire [4-1:0] node6849;
	wire [4-1:0] node6850;
	wire [4-1:0] node6852;
	wire [4-1:0] node6855;
	wire [4-1:0] node6857;
	wire [4-1:0] node6860;
	wire [4-1:0] node6861;
	wire [4-1:0] node6862;
	wire [4-1:0] node6863;
	wire [4-1:0] node6864;
	wire [4-1:0] node6867;
	wire [4-1:0] node6870;
	wire [4-1:0] node6871;
	wire [4-1:0] node6874;
	wire [4-1:0] node6877;
	wire [4-1:0] node6878;
	wire [4-1:0] node6879;
	wire [4-1:0] node6882;
	wire [4-1:0] node6885;
	wire [4-1:0] node6886;
	wire [4-1:0] node6889;
	wire [4-1:0] node6892;
	wire [4-1:0] node6893;
	wire [4-1:0] node6894;
	wire [4-1:0] node6895;
	wire [4-1:0] node6898;
	wire [4-1:0] node6901;
	wire [4-1:0] node6902;
	wire [4-1:0] node6905;
	wire [4-1:0] node6908;
	wire [4-1:0] node6909;
	wire [4-1:0] node6910;
	wire [4-1:0] node6913;
	wire [4-1:0] node6916;
	wire [4-1:0] node6917;
	wire [4-1:0] node6920;
	wire [4-1:0] node6923;
	wire [4-1:0] node6924;
	wire [4-1:0] node6925;
	wire [4-1:0] node6926;
	wire [4-1:0] node6927;
	wire [4-1:0] node6928;
	wire [4-1:0] node6929;
	wire [4-1:0] node6933;
	wire [4-1:0] node6934;
	wire [4-1:0] node6937;
	wire [4-1:0] node6940;
	wire [4-1:0] node6941;
	wire [4-1:0] node6942;
	wire [4-1:0] node6945;
	wire [4-1:0] node6948;
	wire [4-1:0] node6949;
	wire [4-1:0] node6952;
	wire [4-1:0] node6955;
	wire [4-1:0] node6956;
	wire [4-1:0] node6957;
	wire [4-1:0] node6958;
	wire [4-1:0] node6961;
	wire [4-1:0] node6964;
	wire [4-1:0] node6965;
	wire [4-1:0] node6968;
	wire [4-1:0] node6971;
	wire [4-1:0] node6972;
	wire [4-1:0] node6973;
	wire [4-1:0] node6976;
	wire [4-1:0] node6979;
	wire [4-1:0] node6980;
	wire [4-1:0] node6983;
	wire [4-1:0] node6986;
	wire [4-1:0] node6987;
	wire [4-1:0] node6988;
	wire [4-1:0] node6989;
	wire [4-1:0] node6990;
	wire [4-1:0] node6993;
	wire [4-1:0] node6996;
	wire [4-1:0] node6997;
	wire [4-1:0] node7000;
	wire [4-1:0] node7003;
	wire [4-1:0] node7004;
	wire [4-1:0] node7005;
	wire [4-1:0] node7008;
	wire [4-1:0] node7011;
	wire [4-1:0] node7013;
	wire [4-1:0] node7016;
	wire [4-1:0] node7017;
	wire [4-1:0] node7018;
	wire [4-1:0] node7019;
	wire [4-1:0] node7022;
	wire [4-1:0] node7025;
	wire [4-1:0] node7026;
	wire [4-1:0] node7029;
	wire [4-1:0] node7032;
	wire [4-1:0] node7033;
	wire [4-1:0] node7035;
	wire [4-1:0] node7038;
	wire [4-1:0] node7039;
	wire [4-1:0] node7042;
	wire [4-1:0] node7045;
	wire [4-1:0] node7046;
	wire [4-1:0] node7047;
	wire [4-1:0] node7048;
	wire [4-1:0] node7049;
	wire [4-1:0] node7050;
	wire [4-1:0] node7053;
	wire [4-1:0] node7056;
	wire [4-1:0] node7057;
	wire [4-1:0] node7060;
	wire [4-1:0] node7063;
	wire [4-1:0] node7064;
	wire [4-1:0] node7066;
	wire [4-1:0] node7069;
	wire [4-1:0] node7070;
	wire [4-1:0] node7073;
	wire [4-1:0] node7076;
	wire [4-1:0] node7077;
	wire [4-1:0] node7078;
	wire [4-1:0] node7079;
	wire [4-1:0] node7082;
	wire [4-1:0] node7085;
	wire [4-1:0] node7086;
	wire [4-1:0] node7089;
	wire [4-1:0] node7092;
	wire [4-1:0] node7093;
	wire [4-1:0] node7094;
	wire [4-1:0] node7097;
	wire [4-1:0] node7100;
	wire [4-1:0] node7101;
	wire [4-1:0] node7104;
	wire [4-1:0] node7107;
	wire [4-1:0] node7108;
	wire [4-1:0] node7109;
	wire [4-1:0] node7110;
	wire [4-1:0] node7111;
	wire [4-1:0] node7114;
	wire [4-1:0] node7117;
	wire [4-1:0] node7118;
	wire [4-1:0] node7121;
	wire [4-1:0] node7124;
	wire [4-1:0] node7125;
	wire [4-1:0] node7126;
	wire [4-1:0] node7129;
	wire [4-1:0] node7132;
	wire [4-1:0] node7133;
	wire [4-1:0] node7136;
	wire [4-1:0] node7139;
	wire [4-1:0] node7140;
	wire [4-1:0] node7141;
	wire [4-1:0] node7143;
	wire [4-1:0] node7146;
	wire [4-1:0] node7147;
	wire [4-1:0] node7150;
	wire [4-1:0] node7153;
	wire [4-1:0] node7154;
	wire [4-1:0] node7155;
	wire [4-1:0] node7158;
	wire [4-1:0] node7161;
	wire [4-1:0] node7162;
	wire [4-1:0] node7166;
	wire [4-1:0] node7167;
	wire [4-1:0] node7168;
	wire [4-1:0] node7169;
	wire [4-1:0] node7170;
	wire [4-1:0] node7171;
	wire [4-1:0] node7172;
	wire [4-1:0] node7173;
	wire [4-1:0] node7174;
	wire [4-1:0] node7175;
	wire [4-1:0] node7176;
	wire [4-1:0] node7177;
	wire [4-1:0] node7180;
	wire [4-1:0] node7183;
	wire [4-1:0] node7185;
	wire [4-1:0] node7188;
	wire [4-1:0] node7189;
	wire [4-1:0] node7190;
	wire [4-1:0] node7193;
	wire [4-1:0] node7196;
	wire [4-1:0] node7197;
	wire [4-1:0] node7200;
	wire [4-1:0] node7203;
	wire [4-1:0] node7204;
	wire [4-1:0] node7205;
	wire [4-1:0] node7206;
	wire [4-1:0] node7209;
	wire [4-1:0] node7212;
	wire [4-1:0] node7213;
	wire [4-1:0] node7216;
	wire [4-1:0] node7219;
	wire [4-1:0] node7220;
	wire [4-1:0] node7221;
	wire [4-1:0] node7224;
	wire [4-1:0] node7227;
	wire [4-1:0] node7229;
	wire [4-1:0] node7232;
	wire [4-1:0] node7233;
	wire [4-1:0] node7234;
	wire [4-1:0] node7236;
	wire [4-1:0] node7237;
	wire [4-1:0] node7240;
	wire [4-1:0] node7243;
	wire [4-1:0] node7244;
	wire [4-1:0] node7245;
	wire [4-1:0] node7248;
	wire [4-1:0] node7251;
	wire [4-1:0] node7253;
	wire [4-1:0] node7256;
	wire [4-1:0] node7257;
	wire [4-1:0] node7258;
	wire [4-1:0] node7261;
	wire [4-1:0] node7264;
	wire [4-1:0] node7265;
	wire [4-1:0] node7266;
	wire [4-1:0] node7269;
	wire [4-1:0] node7272;
	wire [4-1:0] node7274;
	wire [4-1:0] node7277;
	wire [4-1:0] node7278;
	wire [4-1:0] node7279;
	wire [4-1:0] node7280;
	wire [4-1:0] node7281;
	wire [4-1:0] node7282;
	wire [4-1:0] node7285;
	wire [4-1:0] node7288;
	wire [4-1:0] node7289;
	wire [4-1:0] node7292;
	wire [4-1:0] node7295;
	wire [4-1:0] node7296;
	wire [4-1:0] node7297;
	wire [4-1:0] node7300;
	wire [4-1:0] node7303;
	wire [4-1:0] node7304;
	wire [4-1:0] node7307;
	wire [4-1:0] node7310;
	wire [4-1:0] node7311;
	wire [4-1:0] node7312;
	wire [4-1:0] node7313;
	wire [4-1:0] node7316;
	wire [4-1:0] node7319;
	wire [4-1:0] node7321;
	wire [4-1:0] node7324;
	wire [4-1:0] node7325;
	wire [4-1:0] node7326;
	wire [4-1:0] node7329;
	wire [4-1:0] node7332;
	wire [4-1:0] node7333;
	wire [4-1:0] node7336;
	wire [4-1:0] node7339;
	wire [4-1:0] node7340;
	wire [4-1:0] node7341;
	wire [4-1:0] node7342;
	wire [4-1:0] node7343;
	wire [4-1:0] node7346;
	wire [4-1:0] node7349;
	wire [4-1:0] node7350;
	wire [4-1:0] node7353;
	wire [4-1:0] node7356;
	wire [4-1:0] node7357;
	wire [4-1:0] node7358;
	wire [4-1:0] node7361;
	wire [4-1:0] node7364;
	wire [4-1:0] node7365;
	wire [4-1:0] node7368;
	wire [4-1:0] node7371;
	wire [4-1:0] node7372;
	wire [4-1:0] node7373;
	wire [4-1:0] node7374;
	wire [4-1:0] node7378;
	wire [4-1:0] node7379;
	wire [4-1:0] node7382;
	wire [4-1:0] node7385;
	wire [4-1:0] node7386;
	wire [4-1:0] node7387;
	wire [4-1:0] node7390;
	wire [4-1:0] node7393;
	wire [4-1:0] node7394;
	wire [4-1:0] node7397;
	wire [4-1:0] node7400;
	wire [4-1:0] node7401;
	wire [4-1:0] node7402;
	wire [4-1:0] node7403;
	wire [4-1:0] node7404;
	wire [4-1:0] node7405;
	wire [4-1:0] node7406;
	wire [4-1:0] node7410;
	wire [4-1:0] node7411;
	wire [4-1:0] node7414;
	wire [4-1:0] node7417;
	wire [4-1:0] node7418;
	wire [4-1:0] node7419;
	wire [4-1:0] node7422;
	wire [4-1:0] node7425;
	wire [4-1:0] node7427;
	wire [4-1:0] node7430;
	wire [4-1:0] node7431;
	wire [4-1:0] node7432;
	wire [4-1:0] node7434;
	wire [4-1:0] node7437;
	wire [4-1:0] node7439;
	wire [4-1:0] node7442;
	wire [4-1:0] node7443;
	wire [4-1:0] node7445;
	wire [4-1:0] node7448;
	wire [4-1:0] node7450;
	wire [4-1:0] node7453;
	wire [4-1:0] node7454;
	wire [4-1:0] node7455;
	wire [4-1:0] node7456;
	wire [4-1:0] node7457;
	wire [4-1:0] node7460;
	wire [4-1:0] node7463;
	wire [4-1:0] node7464;
	wire [4-1:0] node7467;
	wire [4-1:0] node7470;
	wire [4-1:0] node7471;
	wire [4-1:0] node7472;
	wire [4-1:0] node7475;
	wire [4-1:0] node7478;
	wire [4-1:0] node7480;
	wire [4-1:0] node7483;
	wire [4-1:0] node7484;
	wire [4-1:0] node7485;
	wire [4-1:0] node7488;
	wire [4-1:0] node7491;
	wire [4-1:0] node7492;
	wire [4-1:0] node7493;
	wire [4-1:0] node7496;
	wire [4-1:0] node7499;
	wire [4-1:0] node7500;
	wire [4-1:0] node7503;
	wire [4-1:0] node7506;
	wire [4-1:0] node7507;
	wire [4-1:0] node7508;
	wire [4-1:0] node7509;
	wire [4-1:0] node7510;
	wire [4-1:0] node7511;
	wire [4-1:0] node7514;
	wire [4-1:0] node7517;
	wire [4-1:0] node7518;
	wire [4-1:0] node7521;
	wire [4-1:0] node7524;
	wire [4-1:0] node7525;
	wire [4-1:0] node7526;
	wire [4-1:0] node7530;
	wire [4-1:0] node7531;
	wire [4-1:0] node7534;
	wire [4-1:0] node7537;
	wire [4-1:0] node7538;
	wire [4-1:0] node7539;
	wire [4-1:0] node7541;
	wire [4-1:0] node7544;
	wire [4-1:0] node7546;
	wire [4-1:0] node7549;
	wire [4-1:0] node7550;
	wire [4-1:0] node7552;
	wire [4-1:0] node7555;
	wire [4-1:0] node7557;
	wire [4-1:0] node7560;
	wire [4-1:0] node7561;
	wire [4-1:0] node7562;
	wire [4-1:0] node7563;
	wire [4-1:0] node7564;
	wire [4-1:0] node7567;
	wire [4-1:0] node7570;
	wire [4-1:0] node7571;
	wire [4-1:0] node7574;
	wire [4-1:0] node7577;
	wire [4-1:0] node7578;
	wire [4-1:0] node7580;
	wire [4-1:0] node7583;
	wire [4-1:0] node7585;
	wire [4-1:0] node7588;
	wire [4-1:0] node7589;
	wire [4-1:0] node7590;
	wire [4-1:0] node7592;
	wire [4-1:0] node7595;
	wire [4-1:0] node7597;
	wire [4-1:0] node7600;
	wire [4-1:0] node7601;
	wire [4-1:0] node7603;
	wire [4-1:0] node7606;
	wire [4-1:0] node7608;
	wire [4-1:0] node7611;
	wire [4-1:0] node7612;
	wire [4-1:0] node7613;
	wire [4-1:0] node7614;
	wire [4-1:0] node7615;
	wire [4-1:0] node7616;
	wire [4-1:0] node7617;
	wire [4-1:0] node7618;
	wire [4-1:0] node7621;
	wire [4-1:0] node7624;
	wire [4-1:0] node7625;
	wire [4-1:0] node7628;
	wire [4-1:0] node7631;
	wire [4-1:0] node7632;
	wire [4-1:0] node7634;
	wire [4-1:0] node7637;
	wire [4-1:0] node7638;
	wire [4-1:0] node7641;
	wire [4-1:0] node7644;
	wire [4-1:0] node7645;
	wire [4-1:0] node7646;
	wire [4-1:0] node7647;
	wire [4-1:0] node7650;
	wire [4-1:0] node7653;
	wire [4-1:0] node7655;
	wire [4-1:0] node7658;
	wire [4-1:0] node7659;
	wire [4-1:0] node7660;
	wire [4-1:0] node7663;
	wire [4-1:0] node7666;
	wire [4-1:0] node7667;
	wire [4-1:0] node7670;
	wire [4-1:0] node7673;
	wire [4-1:0] node7674;
	wire [4-1:0] node7675;
	wire [4-1:0] node7676;
	wire [4-1:0] node7677;
	wire [4-1:0] node7680;
	wire [4-1:0] node7683;
	wire [4-1:0] node7684;
	wire [4-1:0] node7687;
	wire [4-1:0] node7690;
	wire [4-1:0] node7691;
	wire [4-1:0] node7692;
	wire [4-1:0] node7695;
	wire [4-1:0] node7698;
	wire [4-1:0] node7699;
	wire [4-1:0] node7702;
	wire [4-1:0] node7705;
	wire [4-1:0] node7706;
	wire [4-1:0] node7707;
	wire [4-1:0] node7708;
	wire [4-1:0] node7711;
	wire [4-1:0] node7714;
	wire [4-1:0] node7715;
	wire [4-1:0] node7718;
	wire [4-1:0] node7721;
	wire [4-1:0] node7722;
	wire [4-1:0] node7723;
	wire [4-1:0] node7726;
	wire [4-1:0] node7729;
	wire [4-1:0] node7730;
	wire [4-1:0] node7734;
	wire [4-1:0] node7735;
	wire [4-1:0] node7736;
	wire [4-1:0] node7737;
	wire [4-1:0] node7738;
	wire [4-1:0] node7739;
	wire [4-1:0] node7742;
	wire [4-1:0] node7745;
	wire [4-1:0] node7746;
	wire [4-1:0] node7750;
	wire [4-1:0] node7751;
	wire [4-1:0] node7753;
	wire [4-1:0] node7756;
	wire [4-1:0] node7757;
	wire [4-1:0] node7760;
	wire [4-1:0] node7763;
	wire [4-1:0] node7764;
	wire [4-1:0] node7765;
	wire [4-1:0] node7768;
	wire [4-1:0] node7771;
	wire [4-1:0] node7772;
	wire [4-1:0] node7773;
	wire [4-1:0] node7776;
	wire [4-1:0] node7779;
	wire [4-1:0] node7780;
	wire [4-1:0] node7783;
	wire [4-1:0] node7786;
	wire [4-1:0] node7787;
	wire [4-1:0] node7788;
	wire [4-1:0] node7789;
	wire [4-1:0] node7790;
	wire [4-1:0] node7793;
	wire [4-1:0] node7796;
	wire [4-1:0] node7797;
	wire [4-1:0] node7800;
	wire [4-1:0] node7803;
	wire [4-1:0] node7804;
	wire [4-1:0] node7805;
	wire [4-1:0] node7809;
	wire [4-1:0] node7810;
	wire [4-1:0] node7813;
	wire [4-1:0] node7816;
	wire [4-1:0] node7817;
	wire [4-1:0] node7818;
	wire [4-1:0] node7819;
	wire [4-1:0] node7822;
	wire [4-1:0] node7825;
	wire [4-1:0] node7826;
	wire [4-1:0] node7829;
	wire [4-1:0] node7832;
	wire [4-1:0] node7833;
	wire [4-1:0] node7834;
	wire [4-1:0] node7837;
	wire [4-1:0] node7840;
	wire [4-1:0] node7841;
	wire [4-1:0] node7844;
	wire [4-1:0] node7847;
	wire [4-1:0] node7848;
	wire [4-1:0] node7849;
	wire [4-1:0] node7850;
	wire [4-1:0] node7851;
	wire [4-1:0] node7852;
	wire [4-1:0] node7854;
	wire [4-1:0] node7857;
	wire [4-1:0] node7858;
	wire [4-1:0] node7861;
	wire [4-1:0] node7864;
	wire [4-1:0] node7865;
	wire [4-1:0] node7866;
	wire [4-1:0] node7869;
	wire [4-1:0] node7872;
	wire [4-1:0] node7873;
	wire [4-1:0] node7876;
	wire [4-1:0] node7879;
	wire [4-1:0] node7880;
	wire [4-1:0] node7881;
	wire [4-1:0] node7882;
	wire [4-1:0] node7885;
	wire [4-1:0] node7888;
	wire [4-1:0] node7889;
	wire [4-1:0] node7892;
	wire [4-1:0] node7895;
	wire [4-1:0] node7896;
	wire [4-1:0] node7897;
	wire [4-1:0] node7900;
	wire [4-1:0] node7903;
	wire [4-1:0] node7904;
	wire [4-1:0] node7907;
	wire [4-1:0] node7910;
	wire [4-1:0] node7911;
	wire [4-1:0] node7912;
	wire [4-1:0] node7913;
	wire [4-1:0] node7914;
	wire [4-1:0] node7917;
	wire [4-1:0] node7920;
	wire [4-1:0] node7921;
	wire [4-1:0] node7924;
	wire [4-1:0] node7927;
	wire [4-1:0] node7928;
	wire [4-1:0] node7931;
	wire [4-1:0] node7934;
	wire [4-1:0] node7935;
	wire [4-1:0] node7936;
	wire [4-1:0] node7937;
	wire [4-1:0] node7940;
	wire [4-1:0] node7943;
	wire [4-1:0] node7944;
	wire [4-1:0] node7947;
	wire [4-1:0] node7950;
	wire [4-1:0] node7951;
	wire [4-1:0] node7953;
	wire [4-1:0] node7956;
	wire [4-1:0] node7957;
	wire [4-1:0] node7960;
	wire [4-1:0] node7963;
	wire [4-1:0] node7964;
	wire [4-1:0] node7965;
	wire [4-1:0] node7966;
	wire [4-1:0] node7967;
	wire [4-1:0] node7968;
	wire [4-1:0] node7971;
	wire [4-1:0] node7974;
	wire [4-1:0] node7975;
	wire [4-1:0] node7978;
	wire [4-1:0] node7981;
	wire [4-1:0] node7982;
	wire [4-1:0] node7985;
	wire [4-1:0] node7988;
	wire [4-1:0] node7989;
	wire [4-1:0] node7990;
	wire [4-1:0] node7991;
	wire [4-1:0] node7994;
	wire [4-1:0] node7997;
	wire [4-1:0] node7999;
	wire [4-1:0] node8002;
	wire [4-1:0] node8003;
	wire [4-1:0] node8004;
	wire [4-1:0] node8007;
	wire [4-1:0] node8010;
	wire [4-1:0] node8011;
	wire [4-1:0] node8014;
	wire [4-1:0] node8017;
	wire [4-1:0] node8018;
	wire [4-1:0] node8019;
	wire [4-1:0] node8020;
	wire [4-1:0] node8021;
	wire [4-1:0] node8024;
	wire [4-1:0] node8027;
	wire [4-1:0] node8028;
	wire [4-1:0] node8031;
	wire [4-1:0] node8034;
	wire [4-1:0] node8035;
	wire [4-1:0] node8036;
	wire [4-1:0] node8039;
	wire [4-1:0] node8042;
	wire [4-1:0] node8043;
	wire [4-1:0] node8046;
	wire [4-1:0] node8049;
	wire [4-1:0] node8050;
	wire [4-1:0] node8051;
	wire [4-1:0] node8052;
	wire [4-1:0] node8055;
	wire [4-1:0] node8058;
	wire [4-1:0] node8059;
	wire [4-1:0] node8063;
	wire [4-1:0] node8064;
	wire [4-1:0] node8065;
	wire [4-1:0] node8069;
	wire [4-1:0] node8070;
	wire [4-1:0] node8073;
	wire [4-1:0] node8076;
	wire [4-1:0] node8077;
	wire [4-1:0] node8078;
	wire [4-1:0] node8079;
	wire [4-1:0] node8080;
	wire [4-1:0] node8081;
	wire [4-1:0] node8082;
	wire [4-1:0] node8083;
	wire [4-1:0] node8084;
	wire [4-1:0] node8087;
	wire [4-1:0] node8090;
	wire [4-1:0] node8091;
	wire [4-1:0] node8094;
	wire [4-1:0] node8097;
	wire [4-1:0] node8098;
	wire [4-1:0] node8099;
	wire [4-1:0] node8102;
	wire [4-1:0] node8105;
	wire [4-1:0] node8106;
	wire [4-1:0] node8109;
	wire [4-1:0] node8112;
	wire [4-1:0] node8113;
	wire [4-1:0] node8114;
	wire [4-1:0] node8115;
	wire [4-1:0] node8118;
	wire [4-1:0] node8121;
	wire [4-1:0] node8123;
	wire [4-1:0] node8126;
	wire [4-1:0] node8127;
	wire [4-1:0] node8128;
	wire [4-1:0] node8131;
	wire [4-1:0] node8134;
	wire [4-1:0] node8135;
	wire [4-1:0] node8138;
	wire [4-1:0] node8141;
	wire [4-1:0] node8142;
	wire [4-1:0] node8143;
	wire [4-1:0] node8144;
	wire [4-1:0] node8145;
	wire [4-1:0] node8148;
	wire [4-1:0] node8151;
	wire [4-1:0] node8152;
	wire [4-1:0] node8155;
	wire [4-1:0] node8158;
	wire [4-1:0] node8159;
	wire [4-1:0] node8162;
	wire [4-1:0] node8165;
	wire [4-1:0] node8166;
	wire [4-1:0] node8167;
	wire [4-1:0] node8169;
	wire [4-1:0] node8172;
	wire [4-1:0] node8173;
	wire [4-1:0] node8176;
	wire [4-1:0] node8179;
	wire [4-1:0] node8180;
	wire [4-1:0] node8181;
	wire [4-1:0] node8185;
	wire [4-1:0] node8186;
	wire [4-1:0] node8189;
	wire [4-1:0] node8192;
	wire [4-1:0] node8193;
	wire [4-1:0] node8194;
	wire [4-1:0] node8195;
	wire [4-1:0] node8196;
	wire [4-1:0] node8197;
	wire [4-1:0] node8201;
	wire [4-1:0] node8202;
	wire [4-1:0] node8206;
	wire [4-1:0] node8207;
	wire [4-1:0] node8208;
	wire [4-1:0] node8212;
	wire [4-1:0] node8213;
	wire [4-1:0] node8217;
	wire [4-1:0] node8218;
	wire [4-1:0] node8219;
	wire [4-1:0] node8220;
	wire [4-1:0] node8224;
	wire [4-1:0] node8225;
	wire [4-1:0] node8228;
	wire [4-1:0] node8231;
	wire [4-1:0] node8232;
	wire [4-1:0] node8233;
	wire [4-1:0] node8236;
	wire [4-1:0] node8239;
	wire [4-1:0] node8240;
	wire [4-1:0] node8243;
	wire [4-1:0] node8246;
	wire [4-1:0] node8247;
	wire [4-1:0] node8248;
	wire [4-1:0] node8249;
	wire [4-1:0] node8250;
	wire [4-1:0] node8254;
	wire [4-1:0] node8255;
	wire [4-1:0] node8259;
	wire [4-1:0] node8260;
	wire [4-1:0] node8261;
	wire [4-1:0] node8265;
	wire [4-1:0] node8266;
	wire [4-1:0] node8270;
	wire [4-1:0] node8271;
	wire [4-1:0] node8272;
	wire [4-1:0] node8273;
	wire [4-1:0] node8276;
	wire [4-1:0] node8279;
	wire [4-1:0] node8280;
	wire [4-1:0] node8284;
	wire [4-1:0] node8285;
	wire [4-1:0] node8286;
	wire [4-1:0] node8289;
	wire [4-1:0] node8292;
	wire [4-1:0] node8293;
	wire [4-1:0] node8297;
	wire [4-1:0] node8298;
	wire [4-1:0] node8299;
	wire [4-1:0] node8300;
	wire [4-1:0] node8301;
	wire [4-1:0] node8302;
	wire [4-1:0] node8303;
	wire [4-1:0] node8306;
	wire [4-1:0] node8309;
	wire [4-1:0] node8311;
	wire [4-1:0] node8314;
	wire [4-1:0] node8315;
	wire [4-1:0] node8317;
	wire [4-1:0] node8320;
	wire [4-1:0] node8321;
	wire [4-1:0] node8324;
	wire [4-1:0] node8327;
	wire [4-1:0] node8328;
	wire [4-1:0] node8329;
	wire [4-1:0] node8330;
	wire [4-1:0] node8333;
	wire [4-1:0] node8336;
	wire [4-1:0] node8337;
	wire [4-1:0] node8340;
	wire [4-1:0] node8343;
	wire [4-1:0] node8344;
	wire [4-1:0] node8345;
	wire [4-1:0] node8349;
	wire [4-1:0] node8350;
	wire [4-1:0] node8353;
	wire [4-1:0] node8356;
	wire [4-1:0] node8357;
	wire [4-1:0] node8358;
	wire [4-1:0] node8359;
	wire [4-1:0] node8360;
	wire [4-1:0] node8363;
	wire [4-1:0] node8366;
	wire [4-1:0] node8367;
	wire [4-1:0] node8370;
	wire [4-1:0] node8373;
	wire [4-1:0] node8374;
	wire [4-1:0] node8376;
	wire [4-1:0] node8379;
	wire [4-1:0] node8381;
	wire [4-1:0] node8384;
	wire [4-1:0] node8385;
	wire [4-1:0] node8386;
	wire [4-1:0] node8388;
	wire [4-1:0] node8391;
	wire [4-1:0] node8393;
	wire [4-1:0] node8396;
	wire [4-1:0] node8397;
	wire [4-1:0] node8399;
	wire [4-1:0] node8402;
	wire [4-1:0] node8404;
	wire [4-1:0] node8407;
	wire [4-1:0] node8408;
	wire [4-1:0] node8409;
	wire [4-1:0] node8410;
	wire [4-1:0] node8411;
	wire [4-1:0] node8413;
	wire [4-1:0] node8416;
	wire [4-1:0] node8417;
	wire [4-1:0] node8420;
	wire [4-1:0] node8423;
	wire [4-1:0] node8424;
	wire [4-1:0] node8426;
	wire [4-1:0] node8429;
	wire [4-1:0] node8430;
	wire [4-1:0] node8433;
	wire [4-1:0] node8436;
	wire [4-1:0] node8437;
	wire [4-1:0] node8438;
	wire [4-1:0] node8439;
	wire [4-1:0] node8442;
	wire [4-1:0] node8445;
	wire [4-1:0] node8446;
	wire [4-1:0] node8449;
	wire [4-1:0] node8452;
	wire [4-1:0] node8453;
	wire [4-1:0] node8454;
	wire [4-1:0] node8457;
	wire [4-1:0] node8460;
	wire [4-1:0] node8461;
	wire [4-1:0] node8464;
	wire [4-1:0] node8467;
	wire [4-1:0] node8468;
	wire [4-1:0] node8469;
	wire [4-1:0] node8470;
	wire [4-1:0] node8471;
	wire [4-1:0] node8474;
	wire [4-1:0] node8477;
	wire [4-1:0] node8478;
	wire [4-1:0] node8482;
	wire [4-1:0] node8483;
	wire [4-1:0] node8484;
	wire [4-1:0] node8487;
	wire [4-1:0] node8490;
	wire [4-1:0] node8491;
	wire [4-1:0] node8495;
	wire [4-1:0] node8496;
	wire [4-1:0] node8497;
	wire [4-1:0] node8499;
	wire [4-1:0] node8502;
	wire [4-1:0] node8504;
	wire [4-1:0] node8507;
	wire [4-1:0] node8508;
	wire [4-1:0] node8510;
	wire [4-1:0] node8513;
	wire [4-1:0] node8515;
	wire [4-1:0] node8518;
	wire [4-1:0] node8519;
	wire [4-1:0] node8520;
	wire [4-1:0] node8521;
	wire [4-1:0] node8522;
	wire [4-1:0] node8523;
	wire [4-1:0] node8524;
	wire [4-1:0] node8525;
	wire [4-1:0] node8528;
	wire [4-1:0] node8531;
	wire [4-1:0] node8532;
	wire [4-1:0] node8535;
	wire [4-1:0] node8538;
	wire [4-1:0] node8539;
	wire [4-1:0] node8541;
	wire [4-1:0] node8544;
	wire [4-1:0] node8545;
	wire [4-1:0] node8548;
	wire [4-1:0] node8551;
	wire [4-1:0] node8552;
	wire [4-1:0] node8553;
	wire [4-1:0] node8554;
	wire [4-1:0] node8557;
	wire [4-1:0] node8560;
	wire [4-1:0] node8561;
	wire [4-1:0] node8564;
	wire [4-1:0] node8567;
	wire [4-1:0] node8568;
	wire [4-1:0] node8569;
	wire [4-1:0] node8572;
	wire [4-1:0] node8575;
	wire [4-1:0] node8576;
	wire [4-1:0] node8580;
	wire [4-1:0] node8581;
	wire [4-1:0] node8582;
	wire [4-1:0] node8583;
	wire [4-1:0] node8584;
	wire [4-1:0] node8587;
	wire [4-1:0] node8590;
	wire [4-1:0] node8592;
	wire [4-1:0] node8595;
	wire [4-1:0] node8596;
	wire [4-1:0] node8597;
	wire [4-1:0] node8600;
	wire [4-1:0] node8603;
	wire [4-1:0] node8605;
	wire [4-1:0] node8608;
	wire [4-1:0] node8609;
	wire [4-1:0] node8610;
	wire [4-1:0] node8612;
	wire [4-1:0] node8615;
	wire [4-1:0] node8617;
	wire [4-1:0] node8620;
	wire [4-1:0] node8621;
	wire [4-1:0] node8623;
	wire [4-1:0] node8626;
	wire [4-1:0] node8628;
	wire [4-1:0] node8631;
	wire [4-1:0] node8632;
	wire [4-1:0] node8633;
	wire [4-1:0] node8634;
	wire [4-1:0] node8635;
	wire [4-1:0] node8636;
	wire [4-1:0] node8639;
	wire [4-1:0] node8642;
	wire [4-1:0] node8643;
	wire [4-1:0] node8647;
	wire [4-1:0] node8648;
	wire [4-1:0] node8649;
	wire [4-1:0] node8652;
	wire [4-1:0] node8655;
	wire [4-1:0] node8656;
	wire [4-1:0] node8659;
	wire [4-1:0] node8662;
	wire [4-1:0] node8663;
	wire [4-1:0] node8664;
	wire [4-1:0] node8666;
	wire [4-1:0] node8669;
	wire [4-1:0] node8671;
	wire [4-1:0] node8674;
	wire [4-1:0] node8675;
	wire [4-1:0] node8677;
	wire [4-1:0] node8680;
	wire [4-1:0] node8682;
	wire [4-1:0] node8685;
	wire [4-1:0] node8686;
	wire [4-1:0] node8687;
	wire [4-1:0] node8688;
	wire [4-1:0] node8689;
	wire [4-1:0] node8692;
	wire [4-1:0] node8695;
	wire [4-1:0] node8696;
	wire [4-1:0] node8699;
	wire [4-1:0] node8702;
	wire [4-1:0] node8703;
	wire [4-1:0] node8704;
	wire [4-1:0] node8707;
	wire [4-1:0] node8710;
	wire [4-1:0] node8711;
	wire [4-1:0] node8714;
	wire [4-1:0] node8717;
	wire [4-1:0] node8718;
	wire [4-1:0] node8719;
	wire [4-1:0] node8721;
	wire [4-1:0] node8724;
	wire [4-1:0] node8726;
	wire [4-1:0] node8729;
	wire [4-1:0] node8730;
	wire [4-1:0] node8732;
	wire [4-1:0] node8735;
	wire [4-1:0] node8737;
	wire [4-1:0] node8740;
	wire [4-1:0] node8741;
	wire [4-1:0] node8742;
	wire [4-1:0] node8743;
	wire [4-1:0] node8744;
	wire [4-1:0] node8745;
	wire [4-1:0] node8746;
	wire [4-1:0] node8749;
	wire [4-1:0] node8752;
	wire [4-1:0] node8754;
	wire [4-1:0] node8757;
	wire [4-1:0] node8758;
	wire [4-1:0] node8759;
	wire [4-1:0] node8762;
	wire [4-1:0] node8765;
	wire [4-1:0] node8766;
	wire [4-1:0] node8769;
	wire [4-1:0] node8772;
	wire [4-1:0] node8773;
	wire [4-1:0] node8774;
	wire [4-1:0] node8775;
	wire [4-1:0] node8778;
	wire [4-1:0] node8781;
	wire [4-1:0] node8782;
	wire [4-1:0] node8785;
	wire [4-1:0] node8788;
	wire [4-1:0] node8789;
	wire [4-1:0] node8790;
	wire [4-1:0] node8793;
	wire [4-1:0] node8796;
	wire [4-1:0] node8798;
	wire [4-1:0] node8801;
	wire [4-1:0] node8802;
	wire [4-1:0] node8803;
	wire [4-1:0] node8804;
	wire [4-1:0] node8805;
	wire [4-1:0] node8808;
	wire [4-1:0] node8811;
	wire [4-1:0] node8812;
	wire [4-1:0] node8815;
	wire [4-1:0] node8818;
	wire [4-1:0] node8819;
	wire [4-1:0] node8820;
	wire [4-1:0] node8823;
	wire [4-1:0] node8826;
	wire [4-1:0] node8827;
	wire [4-1:0] node8831;
	wire [4-1:0] node8832;
	wire [4-1:0] node8833;
	wire [4-1:0] node8834;
	wire [4-1:0] node8837;
	wire [4-1:0] node8840;
	wire [4-1:0] node8841;
	wire [4-1:0] node8844;
	wire [4-1:0] node8847;
	wire [4-1:0] node8848;
	wire [4-1:0] node8849;
	wire [4-1:0] node8852;
	wire [4-1:0] node8855;
	wire [4-1:0] node8857;
	wire [4-1:0] node8860;
	wire [4-1:0] node8861;
	wire [4-1:0] node8862;
	wire [4-1:0] node8863;
	wire [4-1:0] node8864;
	wire [4-1:0] node8865;
	wire [4-1:0] node8869;
	wire [4-1:0] node8870;
	wire [4-1:0] node8874;
	wire [4-1:0] node8875;
	wire [4-1:0] node8876;
	wire [4-1:0] node8880;
	wire [4-1:0] node8881;
	wire [4-1:0] node8884;
	wire [4-1:0] node8887;
	wire [4-1:0] node8888;
	wire [4-1:0] node8889;
	wire [4-1:0] node8892;
	wire [4-1:0] node8895;
	wire [4-1:0] node8896;
	wire [4-1:0] node8897;
	wire [4-1:0] node8900;
	wire [4-1:0] node8903;
	wire [4-1:0] node8904;
	wire [4-1:0] node8908;
	wire [4-1:0] node8909;
	wire [4-1:0] node8910;
	wire [4-1:0] node8911;
	wire [4-1:0] node8912;
	wire [4-1:0] node8915;
	wire [4-1:0] node8918;
	wire [4-1:0] node8919;
	wire [4-1:0] node8922;
	wire [4-1:0] node8925;
	wire [4-1:0] node8926;
	wire [4-1:0] node8928;
	wire [4-1:0] node8931;
	wire [4-1:0] node8932;
	wire [4-1:0] node8935;
	wire [4-1:0] node8938;
	wire [4-1:0] node8939;
	wire [4-1:0] node8940;
	wire [4-1:0] node8942;
	wire [4-1:0] node8945;
	wire [4-1:0] node8946;
	wire [4-1:0] node8949;
	wire [4-1:0] node8952;
	wire [4-1:0] node8953;
	wire [4-1:0] node8954;
	wire [4-1:0] node8957;
	wire [4-1:0] node8960;
	wire [4-1:0] node8961;
	wire [4-1:0] node8964;
	wire [4-1:0] node8967;
	wire [4-1:0] node8968;
	wire [4-1:0] node8969;
	wire [4-1:0] node8970;
	wire [4-1:0] node8971;
	wire [4-1:0] node8972;
	wire [4-1:0] node8973;
	wire [4-1:0] node8974;
	wire [4-1:0] node8975;
	wire [4-1:0] node8976;
	wire [4-1:0] node8979;
	wire [4-1:0] node8982;
	wire [4-1:0] node8983;
	wire [4-1:0] node8986;
	wire [4-1:0] node8989;
	wire [4-1:0] node8990;
	wire [4-1:0] node8991;
	wire [4-1:0] node8995;
	wire [4-1:0] node8996;
	wire [4-1:0] node8999;
	wire [4-1:0] node9002;
	wire [4-1:0] node9003;
	wire [4-1:0] node9004;
	wire [4-1:0] node9005;
	wire [4-1:0] node9008;
	wire [4-1:0] node9011;
	wire [4-1:0] node9013;
	wire [4-1:0] node9016;
	wire [4-1:0] node9017;
	wire [4-1:0] node9018;
	wire [4-1:0] node9021;
	wire [4-1:0] node9024;
	wire [4-1:0] node9025;
	wire [4-1:0] node9028;
	wire [4-1:0] node9031;
	wire [4-1:0] node9032;
	wire [4-1:0] node9033;
	wire [4-1:0] node9034;
	wire [4-1:0] node9037;
	wire [4-1:0] node9040;
	wire [4-1:0] node9041;
	wire [4-1:0] node9042;
	wire [4-1:0] node9045;
	wire [4-1:0] node9048;
	wire [4-1:0] node9049;
	wire [4-1:0] node9052;
	wire [4-1:0] node9055;
	wire [4-1:0] node9056;
	wire [4-1:0] node9057;
	wire [4-1:0] node9058;
	wire [4-1:0] node9061;
	wire [4-1:0] node9064;
	wire [4-1:0] node9065;
	wire [4-1:0] node9068;
	wire [4-1:0] node9071;
	wire [4-1:0] node9072;
	wire [4-1:0] node9075;
	wire [4-1:0] node9078;
	wire [4-1:0] node9079;
	wire [4-1:0] node9080;
	wire [4-1:0] node9081;
	wire [4-1:0] node9082;
	wire [4-1:0] node9083;
	wire [4-1:0] node9086;
	wire [4-1:0] node9089;
	wire [4-1:0] node9090;
	wire [4-1:0] node9093;
	wire [4-1:0] node9096;
	wire [4-1:0] node9097;
	wire [4-1:0] node9098;
	wire [4-1:0] node9101;
	wire [4-1:0] node9104;
	wire [4-1:0] node9105;
	wire [4-1:0] node9108;
	wire [4-1:0] node9111;
	wire [4-1:0] node9112;
	wire [4-1:0] node9113;
	wire [4-1:0] node9115;
	wire [4-1:0] node9118;
	wire [4-1:0] node9119;
	wire [4-1:0] node9122;
	wire [4-1:0] node9125;
	wire [4-1:0] node9126;
	wire [4-1:0] node9127;
	wire [4-1:0] node9130;
	wire [4-1:0] node9133;
	wire [4-1:0] node9134;
	wire [4-1:0] node9137;
	wire [4-1:0] node9140;
	wire [4-1:0] node9141;
	wire [4-1:0] node9142;
	wire [4-1:0] node9143;
	wire [4-1:0] node9144;
	wire [4-1:0] node9147;
	wire [4-1:0] node9150;
	wire [4-1:0] node9151;
	wire [4-1:0] node9154;
	wire [4-1:0] node9157;
	wire [4-1:0] node9158;
	wire [4-1:0] node9159;
	wire [4-1:0] node9162;
	wire [4-1:0] node9165;
	wire [4-1:0] node9166;
	wire [4-1:0] node9169;
	wire [4-1:0] node9172;
	wire [4-1:0] node9173;
	wire [4-1:0] node9174;
	wire [4-1:0] node9175;
	wire [4-1:0] node9178;
	wire [4-1:0] node9181;
	wire [4-1:0] node9182;
	wire [4-1:0] node9185;
	wire [4-1:0] node9188;
	wire [4-1:0] node9189;
	wire [4-1:0] node9190;
	wire [4-1:0] node9193;
	wire [4-1:0] node9196;
	wire [4-1:0] node9197;
	wire [4-1:0] node9200;
	wire [4-1:0] node9203;
	wire [4-1:0] node9204;
	wire [4-1:0] node9205;
	wire [4-1:0] node9206;
	wire [4-1:0] node9207;
	wire [4-1:0] node9208;
	wire [4-1:0] node9209;
	wire [4-1:0] node9212;
	wire [4-1:0] node9215;
	wire [4-1:0] node9216;
	wire [4-1:0] node9219;
	wire [4-1:0] node9222;
	wire [4-1:0] node9223;
	wire [4-1:0] node9224;
	wire [4-1:0] node9227;
	wire [4-1:0] node9230;
	wire [4-1:0] node9231;
	wire [4-1:0] node9234;
	wire [4-1:0] node9237;
	wire [4-1:0] node9238;
	wire [4-1:0] node9239;
	wire [4-1:0] node9240;
	wire [4-1:0] node9243;
	wire [4-1:0] node9246;
	wire [4-1:0] node9247;
	wire [4-1:0] node9250;
	wire [4-1:0] node9253;
	wire [4-1:0] node9254;
	wire [4-1:0] node9255;
	wire [4-1:0] node9258;
	wire [4-1:0] node9261;
	wire [4-1:0] node9262;
	wire [4-1:0] node9265;
	wire [4-1:0] node9268;
	wire [4-1:0] node9269;
	wire [4-1:0] node9270;
	wire [4-1:0] node9271;
	wire [4-1:0] node9273;
	wire [4-1:0] node9276;
	wire [4-1:0] node9277;
	wire [4-1:0] node9280;
	wire [4-1:0] node9283;
	wire [4-1:0] node9284;
	wire [4-1:0] node9285;
	wire [4-1:0] node9288;
	wire [4-1:0] node9291;
	wire [4-1:0] node9292;
	wire [4-1:0] node9295;
	wire [4-1:0] node9298;
	wire [4-1:0] node9299;
	wire [4-1:0] node9300;
	wire [4-1:0] node9302;
	wire [4-1:0] node9305;
	wire [4-1:0] node9307;
	wire [4-1:0] node9310;
	wire [4-1:0] node9311;
	wire [4-1:0] node9313;
	wire [4-1:0] node9316;
	wire [4-1:0] node9318;
	wire [4-1:0] node9321;
	wire [4-1:0] node9322;
	wire [4-1:0] node9323;
	wire [4-1:0] node9324;
	wire [4-1:0] node9325;
	wire [4-1:0] node9327;
	wire [4-1:0] node9330;
	wire [4-1:0] node9331;
	wire [4-1:0] node9334;
	wire [4-1:0] node9337;
	wire [4-1:0] node9338;
	wire [4-1:0] node9339;
	wire [4-1:0] node9343;
	wire [4-1:0] node9344;
	wire [4-1:0] node9347;
	wire [4-1:0] node9350;
	wire [4-1:0] node9351;
	wire [4-1:0] node9352;
	wire [4-1:0] node9353;
	wire [4-1:0] node9356;
	wire [4-1:0] node9359;
	wire [4-1:0] node9360;
	wire [4-1:0] node9363;
	wire [4-1:0] node9366;
	wire [4-1:0] node9367;
	wire [4-1:0] node9368;
	wire [4-1:0] node9371;
	wire [4-1:0] node9374;
	wire [4-1:0] node9375;
	wire [4-1:0] node9379;
	wire [4-1:0] node9380;
	wire [4-1:0] node9381;
	wire [4-1:0] node9382;
	wire [4-1:0] node9383;
	wire [4-1:0] node9386;
	wire [4-1:0] node9389;
	wire [4-1:0] node9390;
	wire [4-1:0] node9393;
	wire [4-1:0] node9396;
	wire [4-1:0] node9397;
	wire [4-1:0] node9398;
	wire [4-1:0] node9402;
	wire [4-1:0] node9403;
	wire [4-1:0] node9406;
	wire [4-1:0] node9409;
	wire [4-1:0] node9410;
	wire [4-1:0] node9411;
	wire [4-1:0] node9412;
	wire [4-1:0] node9415;
	wire [4-1:0] node9418;
	wire [4-1:0] node9419;
	wire [4-1:0] node9422;
	wire [4-1:0] node9425;
	wire [4-1:0] node9426;
	wire [4-1:0] node9427;
	wire [4-1:0] node9430;
	wire [4-1:0] node9433;
	wire [4-1:0] node9434;
	wire [4-1:0] node9437;
	wire [4-1:0] node9440;
	wire [4-1:0] node9441;
	wire [4-1:0] node9442;
	wire [4-1:0] node9443;
	wire [4-1:0] node9444;
	wire [4-1:0] node9445;
	wire [4-1:0] node9446;
	wire [4-1:0] node9448;
	wire [4-1:0] node9451;
	wire [4-1:0] node9452;
	wire [4-1:0] node9455;
	wire [4-1:0] node9458;
	wire [4-1:0] node9459;
	wire [4-1:0] node9460;
	wire [4-1:0] node9464;
	wire [4-1:0] node9465;
	wire [4-1:0] node9468;
	wire [4-1:0] node9471;
	wire [4-1:0] node9472;
	wire [4-1:0] node9473;
	wire [4-1:0] node9475;
	wire [4-1:0] node9478;
	wire [4-1:0] node9479;
	wire [4-1:0] node9482;
	wire [4-1:0] node9485;
	wire [4-1:0] node9486;
	wire [4-1:0] node9487;
	wire [4-1:0] node9491;
	wire [4-1:0] node9492;
	wire [4-1:0] node9495;
	wire [4-1:0] node9498;
	wire [4-1:0] node9499;
	wire [4-1:0] node9500;
	wire [4-1:0] node9501;
	wire [4-1:0] node9502;
	wire [4-1:0] node9505;
	wire [4-1:0] node9508;
	wire [4-1:0] node9509;
	wire [4-1:0] node9512;
	wire [4-1:0] node9515;
	wire [4-1:0] node9516;
	wire [4-1:0] node9517;
	wire [4-1:0] node9520;
	wire [4-1:0] node9523;
	wire [4-1:0] node9524;
	wire [4-1:0] node9527;
	wire [4-1:0] node9530;
	wire [4-1:0] node9531;
	wire [4-1:0] node9532;
	wire [4-1:0] node9533;
	wire [4-1:0] node9536;
	wire [4-1:0] node9539;
	wire [4-1:0] node9540;
	wire [4-1:0] node9543;
	wire [4-1:0] node9546;
	wire [4-1:0] node9547;
	wire [4-1:0] node9548;
	wire [4-1:0] node9551;
	wire [4-1:0] node9555;
	wire [4-1:0] node9556;
	wire [4-1:0] node9557;
	wire [4-1:0] node9558;
	wire [4-1:0] node9559;
	wire [4-1:0] node9560;
	wire [4-1:0] node9563;
	wire [4-1:0] node9566;
	wire [4-1:0] node9567;
	wire [4-1:0] node9571;
	wire [4-1:0] node9572;
	wire [4-1:0] node9574;
	wire [4-1:0] node9577;
	wire [4-1:0] node9579;
	wire [4-1:0] node9582;
	wire [4-1:0] node9583;
	wire [4-1:0] node9584;
	wire [4-1:0] node9585;
	wire [4-1:0] node9588;
	wire [4-1:0] node9591;
	wire [4-1:0] node9592;
	wire [4-1:0] node9595;
	wire [4-1:0] node9598;
	wire [4-1:0] node9599;
	wire [4-1:0] node9600;
	wire [4-1:0] node9603;
	wire [4-1:0] node9606;
	wire [4-1:0] node9607;
	wire [4-1:0] node9610;
	wire [4-1:0] node9613;
	wire [4-1:0] node9614;
	wire [4-1:0] node9615;
	wire [4-1:0] node9616;
	wire [4-1:0] node9617;
	wire [4-1:0] node9620;
	wire [4-1:0] node9623;
	wire [4-1:0] node9624;
	wire [4-1:0] node9627;
	wire [4-1:0] node9630;
	wire [4-1:0] node9631;
	wire [4-1:0] node9632;
	wire [4-1:0] node9635;
	wire [4-1:0] node9638;
	wire [4-1:0] node9640;
	wire [4-1:0] node9643;
	wire [4-1:0] node9644;
	wire [4-1:0] node9645;
	wire [4-1:0] node9646;
	wire [4-1:0] node9649;
	wire [4-1:0] node9652;
	wire [4-1:0] node9653;
	wire [4-1:0] node9656;
	wire [4-1:0] node9659;
	wire [4-1:0] node9660;
	wire [4-1:0] node9661;
	wire [4-1:0] node9664;
	wire [4-1:0] node9667;
	wire [4-1:0] node9668;
	wire [4-1:0] node9672;
	wire [4-1:0] node9673;
	wire [4-1:0] node9674;
	wire [4-1:0] node9675;
	wire [4-1:0] node9676;
	wire [4-1:0] node9677;
	wire [4-1:0] node9678;
	wire [4-1:0] node9682;
	wire [4-1:0] node9683;
	wire [4-1:0] node9687;
	wire [4-1:0] node9688;
	wire [4-1:0] node9689;
	wire [4-1:0] node9693;
	wire [4-1:0] node9694;
	wire [4-1:0] node9698;
	wire [4-1:0] node9699;
	wire [4-1:0] node9700;
	wire [4-1:0] node9701;
	wire [4-1:0] node9704;
	wire [4-1:0] node9707;
	wire [4-1:0] node9708;
	wire [4-1:0] node9711;
	wire [4-1:0] node9714;
	wire [4-1:0] node9715;
	wire [4-1:0] node9716;
	wire [4-1:0] node9719;
	wire [4-1:0] node9722;
	wire [4-1:0] node9724;
	wire [4-1:0] node9727;
	wire [4-1:0] node9728;
	wire [4-1:0] node9729;
	wire [4-1:0] node9730;
	wire [4-1:0] node9731;
	wire [4-1:0] node9735;
	wire [4-1:0] node9736;
	wire [4-1:0] node9740;
	wire [4-1:0] node9742;
	wire [4-1:0] node9743;
	wire [4-1:0] node9747;
	wire [4-1:0] node9748;
	wire [4-1:0] node9749;
	wire [4-1:0] node9750;
	wire [4-1:0] node9754;
	wire [4-1:0] node9755;
	wire [4-1:0] node9758;
	wire [4-1:0] node9761;
	wire [4-1:0] node9762;
	wire [4-1:0] node9763;
	wire [4-1:0] node9766;
	wire [4-1:0] node9769;
	wire [4-1:0] node9770;
	wire [4-1:0] node9773;
	wire [4-1:0] node9776;
	wire [4-1:0] node9777;
	wire [4-1:0] node9778;
	wire [4-1:0] node9779;
	wire [4-1:0] node9780;
	wire [4-1:0] node9781;
	wire [4-1:0] node9784;
	wire [4-1:0] node9787;
	wire [4-1:0] node9788;
	wire [4-1:0] node9791;
	wire [4-1:0] node9794;
	wire [4-1:0] node9795;
	wire [4-1:0] node9796;
	wire [4-1:0] node9799;
	wire [4-1:0] node9802;
	wire [4-1:0] node9803;
	wire [4-1:0] node9806;
	wire [4-1:0] node9809;
	wire [4-1:0] node9810;
	wire [4-1:0] node9811;
	wire [4-1:0] node9813;
	wire [4-1:0] node9816;
	wire [4-1:0] node9817;
	wire [4-1:0] node9820;
	wire [4-1:0] node9823;
	wire [4-1:0] node9824;
	wire [4-1:0] node9825;
	wire [4-1:0] node9828;
	wire [4-1:0] node9831;
	wire [4-1:0] node9832;
	wire [4-1:0] node9835;
	wire [4-1:0] node9838;
	wire [4-1:0] node9839;
	wire [4-1:0] node9840;
	wire [4-1:0] node9841;
	wire [4-1:0] node9842;
	wire [4-1:0] node9846;
	wire [4-1:0] node9847;
	wire [4-1:0] node9851;
	wire [4-1:0] node9852;
	wire [4-1:0] node9853;
	wire [4-1:0] node9857;
	wire [4-1:0] node9858;
	wire [4-1:0] node9862;
	wire [4-1:0] node9863;
	wire [4-1:0] node9864;
	wire [4-1:0] node9865;
	wire [4-1:0] node9868;
	wire [4-1:0] node9871;
	wire [4-1:0] node9872;
	wire [4-1:0] node9876;
	wire [4-1:0] node9877;
	wire [4-1:0] node9878;
	wire [4-1:0] node9881;
	wire [4-1:0] node9884;
	wire [4-1:0] node9885;
	wire [4-1:0] node9888;
	wire [4-1:0] node9891;
	wire [4-1:0] node9892;
	wire [4-1:0] node9893;
	wire [4-1:0] node9894;
	wire [4-1:0] node9895;
	wire [4-1:0] node9896;
	wire [4-1:0] node9897;
	wire [4-1:0] node9898;
	wire [4-1:0] node9900;
	wire [4-1:0] node9903;
	wire [4-1:0] node9904;
	wire [4-1:0] node9907;
	wire [4-1:0] node9910;
	wire [4-1:0] node9911;
	wire [4-1:0] node9912;
	wire [4-1:0] node9915;
	wire [4-1:0] node9918;
	wire [4-1:0] node9919;
	wire [4-1:0] node9922;
	wire [4-1:0] node9925;
	wire [4-1:0] node9926;
	wire [4-1:0] node9927;
	wire [4-1:0] node9929;
	wire [4-1:0] node9932;
	wire [4-1:0] node9934;
	wire [4-1:0] node9937;
	wire [4-1:0] node9938;
	wire [4-1:0] node9940;
	wire [4-1:0] node9943;
	wire [4-1:0] node9945;
	wire [4-1:0] node9948;
	wire [4-1:0] node9949;
	wire [4-1:0] node9950;
	wire [4-1:0] node9951;
	wire [4-1:0] node9952;
	wire [4-1:0] node9955;
	wire [4-1:0] node9958;
	wire [4-1:0] node9959;
	wire [4-1:0] node9962;
	wire [4-1:0] node9965;
	wire [4-1:0] node9966;
	wire [4-1:0] node9967;
	wire [4-1:0] node9970;
	wire [4-1:0] node9973;
	wire [4-1:0] node9974;
	wire [4-1:0] node9977;
	wire [4-1:0] node9980;
	wire [4-1:0] node9981;
	wire [4-1:0] node9982;
	wire [4-1:0] node9983;
	wire [4-1:0] node9986;
	wire [4-1:0] node9989;
	wire [4-1:0] node9990;
	wire [4-1:0] node9993;
	wire [4-1:0] node9996;
	wire [4-1:0] node9997;
	wire [4-1:0] node9998;
	wire [4-1:0] node10001;
	wire [4-1:0] node10004;
	wire [4-1:0] node10005;
	wire [4-1:0] node10008;
	wire [4-1:0] node10011;
	wire [4-1:0] node10012;
	wire [4-1:0] node10013;
	wire [4-1:0] node10014;
	wire [4-1:0] node10015;
	wire [4-1:0] node10016;
	wire [4-1:0] node10019;
	wire [4-1:0] node10022;
	wire [4-1:0] node10023;
	wire [4-1:0] node10026;
	wire [4-1:0] node10029;
	wire [4-1:0] node10030;
	wire [4-1:0] node10031;
	wire [4-1:0] node10034;
	wire [4-1:0] node10037;
	wire [4-1:0] node10038;
	wire [4-1:0] node10041;
	wire [4-1:0] node10044;
	wire [4-1:0] node10045;
	wire [4-1:0] node10046;
	wire [4-1:0] node10049;
	wire [4-1:0] node10052;
	wire [4-1:0] node10053;
	wire [4-1:0] node10054;
	wire [4-1:0] node10057;
	wire [4-1:0] node10060;
	wire [4-1:0] node10061;
	wire [4-1:0] node10064;
	wire [4-1:0] node10067;
	wire [4-1:0] node10068;
	wire [4-1:0] node10069;
	wire [4-1:0] node10070;
	wire [4-1:0] node10071;
	wire [4-1:0] node10074;
	wire [4-1:0] node10077;
	wire [4-1:0] node10079;
	wire [4-1:0] node10082;
	wire [4-1:0] node10083;
	wire [4-1:0] node10085;
	wire [4-1:0] node10088;
	wire [4-1:0] node10089;
	wire [4-1:0] node10092;
	wire [4-1:0] node10095;
	wire [4-1:0] node10096;
	wire [4-1:0] node10097;
	wire [4-1:0] node10098;
	wire [4-1:0] node10101;
	wire [4-1:0] node10104;
	wire [4-1:0] node10105;
	wire [4-1:0] node10108;
	wire [4-1:0] node10111;
	wire [4-1:0] node10112;
	wire [4-1:0] node10113;
	wire [4-1:0] node10116;
	wire [4-1:0] node10119;
	wire [4-1:0] node10121;
	wire [4-1:0] node10124;
	wire [4-1:0] node10125;
	wire [4-1:0] node10126;
	wire [4-1:0] node10127;
	wire [4-1:0] node10128;
	wire [4-1:0] node10129;
	wire [4-1:0] node10130;
	wire [4-1:0] node10133;
	wire [4-1:0] node10136;
	wire [4-1:0] node10137;
	wire [4-1:0] node10140;
	wire [4-1:0] node10143;
	wire [4-1:0] node10144;
	wire [4-1:0] node10146;
	wire [4-1:0] node10149;
	wire [4-1:0] node10150;
	wire [4-1:0] node10153;
	wire [4-1:0] node10156;
	wire [4-1:0] node10157;
	wire [4-1:0] node10158;
	wire [4-1:0] node10160;
	wire [4-1:0] node10163;
	wire [4-1:0] node10165;
	wire [4-1:0] node10168;
	wire [4-1:0] node10169;
	wire [4-1:0] node10171;
	wire [4-1:0] node10174;
	wire [4-1:0] node10176;
	wire [4-1:0] node10179;
	wire [4-1:0] node10180;
	wire [4-1:0] node10181;
	wire [4-1:0] node10182;
	wire [4-1:0] node10184;
	wire [4-1:0] node10187;
	wire [4-1:0] node10188;
	wire [4-1:0] node10191;
	wire [4-1:0] node10194;
	wire [4-1:0] node10195;
	wire [4-1:0] node10196;
	wire [4-1:0] node10199;
	wire [4-1:0] node10202;
	wire [4-1:0] node10203;
	wire [4-1:0] node10206;
	wire [4-1:0] node10209;
	wire [4-1:0] node10210;
	wire [4-1:0] node10211;
	wire [4-1:0] node10214;
	wire [4-1:0] node10217;
	wire [4-1:0] node10218;
	wire [4-1:0] node10219;
	wire [4-1:0] node10222;
	wire [4-1:0] node10225;
	wire [4-1:0] node10226;
	wire [4-1:0] node10230;
	wire [4-1:0] node10231;
	wire [4-1:0] node10232;
	wire [4-1:0] node10233;
	wire [4-1:0] node10234;
	wire [4-1:0] node10235;
	wire [4-1:0] node10238;
	wire [4-1:0] node10241;
	wire [4-1:0] node10243;
	wire [4-1:0] node10246;
	wire [4-1:0] node10247;
	wire [4-1:0] node10248;
	wire [4-1:0] node10252;
	wire [4-1:0] node10253;
	wire [4-1:0] node10256;
	wire [4-1:0] node10259;
	wire [4-1:0] node10260;
	wire [4-1:0] node10261;
	wire [4-1:0] node10262;
	wire [4-1:0] node10265;
	wire [4-1:0] node10268;
	wire [4-1:0] node10269;
	wire [4-1:0] node10272;
	wire [4-1:0] node10275;
	wire [4-1:0] node10276;
	wire [4-1:0] node10278;
	wire [4-1:0] node10281;
	wire [4-1:0] node10282;
	wire [4-1:0] node10285;
	wire [4-1:0] node10288;
	wire [4-1:0] node10289;
	wire [4-1:0] node10290;
	wire [4-1:0] node10291;
	wire [4-1:0] node10292;
	wire [4-1:0] node10295;
	wire [4-1:0] node10298;
	wire [4-1:0] node10299;
	wire [4-1:0] node10303;
	wire [4-1:0] node10304;
	wire [4-1:0] node10305;
	wire [4-1:0] node10309;
	wire [4-1:0] node10310;
	wire [4-1:0] node10313;
	wire [4-1:0] node10316;
	wire [4-1:0] node10317;
	wire [4-1:0] node10318;
	wire [4-1:0] node10319;
	wire [4-1:0] node10322;
	wire [4-1:0] node10325;
	wire [4-1:0] node10326;
	wire [4-1:0] node10329;
	wire [4-1:0] node10332;
	wire [4-1:0] node10333;
	wire [4-1:0] node10334;
	wire [4-1:0] node10337;
	wire [4-1:0] node10340;
	wire [4-1:0] node10341;
	wire [4-1:0] node10345;
	wire [4-1:0] node10346;
	wire [4-1:0] node10347;
	wire [4-1:0] node10348;
	wire [4-1:0] node10349;
	wire [4-1:0] node10350;
	wire [4-1:0] node10351;
	wire [4-1:0] node10352;
	wire [4-1:0] node10356;
	wire [4-1:0] node10357;
	wire [4-1:0] node10361;
	wire [4-1:0] node10362;
	wire [4-1:0] node10364;
	wire [4-1:0] node10367;
	wire [4-1:0] node10369;
	wire [4-1:0] node10372;
	wire [4-1:0] node10373;
	wire [4-1:0] node10375;
	wire [4-1:0] node10377;
	wire [4-1:0] node10380;
	wire [4-1:0] node10381;
	wire [4-1:0] node10383;
	wire [4-1:0] node10386;
	wire [4-1:0] node10388;
	wire [4-1:0] node10391;
	wire [4-1:0] node10392;
	wire [4-1:0] node10393;
	wire [4-1:0] node10394;
	wire [4-1:0] node10395;
	wire [4-1:0] node10398;
	wire [4-1:0] node10401;
	wire [4-1:0] node10402;
	wire [4-1:0] node10405;
	wire [4-1:0] node10408;
	wire [4-1:0] node10409;
	wire [4-1:0] node10410;
	wire [4-1:0] node10413;
	wire [4-1:0] node10416;
	wire [4-1:0] node10417;
	wire [4-1:0] node10420;
	wire [4-1:0] node10423;
	wire [4-1:0] node10424;
	wire [4-1:0] node10425;
	wire [4-1:0] node10426;
	wire [4-1:0] node10429;
	wire [4-1:0] node10432;
	wire [4-1:0] node10433;
	wire [4-1:0] node10436;
	wire [4-1:0] node10439;
	wire [4-1:0] node10440;
	wire [4-1:0] node10441;
	wire [4-1:0] node10444;
	wire [4-1:0] node10447;
	wire [4-1:0] node10449;
	wire [4-1:0] node10452;
	wire [4-1:0] node10453;
	wire [4-1:0] node10454;
	wire [4-1:0] node10455;
	wire [4-1:0] node10456;
	wire [4-1:0] node10457;
	wire [4-1:0] node10460;
	wire [4-1:0] node10463;
	wire [4-1:0] node10464;
	wire [4-1:0] node10467;
	wire [4-1:0] node10470;
	wire [4-1:0] node10471;
	wire [4-1:0] node10472;
	wire [4-1:0] node10476;
	wire [4-1:0] node10477;
	wire [4-1:0] node10481;
	wire [4-1:0] node10482;
	wire [4-1:0] node10483;
	wire [4-1:0] node10485;
	wire [4-1:0] node10488;
	wire [4-1:0] node10490;
	wire [4-1:0] node10493;
	wire [4-1:0] node10494;
	wire [4-1:0] node10496;
	wire [4-1:0] node10499;
	wire [4-1:0] node10501;
	wire [4-1:0] node10504;
	wire [4-1:0] node10505;
	wire [4-1:0] node10506;
	wire [4-1:0] node10507;
	wire [4-1:0] node10508;
	wire [4-1:0] node10511;
	wire [4-1:0] node10514;
	wire [4-1:0] node10515;
	wire [4-1:0] node10518;
	wire [4-1:0] node10521;
	wire [4-1:0] node10522;
	wire [4-1:0] node10523;
	wire [4-1:0] node10527;
	wire [4-1:0] node10528;
	wire [4-1:0] node10532;
	wire [4-1:0] node10533;
	wire [4-1:0] node10534;
	wire [4-1:0] node10535;
	wire [4-1:0] node10539;
	wire [4-1:0] node10540;
	wire [4-1:0] node10543;
	wire [4-1:0] node10546;
	wire [4-1:0] node10547;
	wire [4-1:0] node10548;
	wire [4-1:0] node10551;
	wire [4-1:0] node10554;
	wire [4-1:0] node10556;
	wire [4-1:0] node10559;
	wire [4-1:0] node10560;
	wire [4-1:0] node10561;
	wire [4-1:0] node10562;
	wire [4-1:0] node10563;
	wire [4-1:0] node10564;
	wire [4-1:0] node10565;
	wire [4-1:0] node10568;
	wire [4-1:0] node10571;
	wire [4-1:0] node10572;
	wire [4-1:0] node10575;
	wire [4-1:0] node10578;
	wire [4-1:0] node10579;
	wire [4-1:0] node10580;
	wire [4-1:0] node10583;
	wire [4-1:0] node10586;
	wire [4-1:0] node10587;
	wire [4-1:0] node10590;
	wire [4-1:0] node10593;
	wire [4-1:0] node10594;
	wire [4-1:0] node10595;
	wire [4-1:0] node10596;
	wire [4-1:0] node10599;
	wire [4-1:0] node10602;
	wire [4-1:0] node10603;
	wire [4-1:0] node10606;
	wire [4-1:0] node10609;
	wire [4-1:0] node10610;
	wire [4-1:0] node10611;
	wire [4-1:0] node10614;
	wire [4-1:0] node10617;
	wire [4-1:0] node10618;
	wire [4-1:0] node10621;
	wire [4-1:0] node10624;
	wire [4-1:0] node10625;
	wire [4-1:0] node10626;
	wire [4-1:0] node10627;
	wire [4-1:0] node10628;
	wire [4-1:0] node10631;
	wire [4-1:0] node10634;
	wire [4-1:0] node10635;
	wire [4-1:0] node10638;
	wire [4-1:0] node10641;
	wire [4-1:0] node10642;
	wire [4-1:0] node10643;
	wire [4-1:0] node10646;
	wire [4-1:0] node10649;
	wire [4-1:0] node10650;
	wire [4-1:0] node10653;
	wire [4-1:0] node10656;
	wire [4-1:0] node10657;
	wire [4-1:0] node10658;
	wire [4-1:0] node10659;
	wire [4-1:0] node10662;
	wire [4-1:0] node10665;
	wire [4-1:0] node10666;
	wire [4-1:0] node10669;
	wire [4-1:0] node10672;
	wire [4-1:0] node10673;
	wire [4-1:0] node10674;
	wire [4-1:0] node10677;
	wire [4-1:0] node10680;
	wire [4-1:0] node10681;
	wire [4-1:0] node10684;
	wire [4-1:0] node10687;
	wire [4-1:0] node10688;
	wire [4-1:0] node10689;
	wire [4-1:0] node10690;
	wire [4-1:0] node10691;
	wire [4-1:0] node10694;
	wire [4-1:0] node10697;
	wire [4-1:0] node10698;
	wire [4-1:0] node10700;
	wire [4-1:0] node10703;
	wire [4-1:0] node10704;
	wire [4-1:0] node10707;
	wire [4-1:0] node10710;
	wire [4-1:0] node10711;
	wire [4-1:0] node10712;
	wire [4-1:0] node10715;
	wire [4-1:0] node10718;
	wire [4-1:0] node10719;
	wire [4-1:0] node10720;
	wire [4-1:0] node10723;
	wire [4-1:0] node10726;
	wire [4-1:0] node10728;
	wire [4-1:0] node10731;
	wire [4-1:0] node10732;
	wire [4-1:0] node10733;
	wire [4-1:0] node10734;
	wire [4-1:0] node10737;
	wire [4-1:0] node10740;
	wire [4-1:0] node10741;
	wire [4-1:0] node10742;
	wire [4-1:0] node10745;
	wire [4-1:0] node10748;
	wire [4-1:0] node10749;
	wire [4-1:0] node10752;
	wire [4-1:0] node10755;
	wire [4-1:0] node10756;
	wire [4-1:0] node10757;
	wire [4-1:0] node10760;
	wire [4-1:0] node10763;
	wire [4-1:0] node10764;
	wire [4-1:0] node10765;
	wire [4-1:0] node10768;
	wire [4-1:0] node10771;
	wire [4-1:0] node10772;
	wire [4-1:0] node10775;
	wire [4-1:0] node10778;
	wire [4-1:0] node10779;
	wire [4-1:0] node10780;
	wire [4-1:0] node10781;
	wire [4-1:0] node10782;
	wire [4-1:0] node10783;
	wire [4-1:0] node10784;
	wire [4-1:0] node10785;
	wire [4-1:0] node10786;
	wire [4-1:0] node10787;
	wire [4-1:0] node10788;
	wire [4-1:0] node10791;
	wire [4-1:0] node10794;
	wire [4-1:0] node10795;
	wire [4-1:0] node10798;
	wire [4-1:0] node10801;
	wire [4-1:0] node10802;
	wire [4-1:0] node10803;
	wire [4-1:0] node10806;
	wire [4-1:0] node10809;
	wire [4-1:0] node10810;
	wire [4-1:0] node10813;
	wire [4-1:0] node10816;
	wire [4-1:0] node10817;
	wire [4-1:0] node10818;
	wire [4-1:0] node10819;
	wire [4-1:0] node10822;
	wire [4-1:0] node10825;
	wire [4-1:0] node10826;
	wire [4-1:0] node10829;
	wire [4-1:0] node10832;
	wire [4-1:0] node10833;
	wire [4-1:0] node10835;
	wire [4-1:0] node10838;
	wire [4-1:0] node10839;
	wire [4-1:0] node10842;
	wire [4-1:0] node10845;
	wire [4-1:0] node10846;
	wire [4-1:0] node10847;
	wire [4-1:0] node10848;
	wire [4-1:0] node10850;
	wire [4-1:0] node10853;
	wire [4-1:0] node10855;
	wire [4-1:0] node10858;
	wire [4-1:0] node10859;
	wire [4-1:0] node10862;
	wire [4-1:0] node10865;
	wire [4-1:0] node10866;
	wire [4-1:0] node10867;
	wire [4-1:0] node10870;
	wire [4-1:0] node10873;
	wire [4-1:0] node10874;
	wire [4-1:0] node10875;
	wire [4-1:0] node10878;
	wire [4-1:0] node10881;
	wire [4-1:0] node10882;
	wire [4-1:0] node10885;
	wire [4-1:0] node10888;
	wire [4-1:0] node10889;
	wire [4-1:0] node10890;
	wire [4-1:0] node10891;
	wire [4-1:0] node10892;
	wire [4-1:0] node10895;
	wire [4-1:0] node10898;
	wire [4-1:0] node10899;
	wire [4-1:0] node10902;
	wire [4-1:0] node10905;
	wire [4-1:0] node10906;
	wire [4-1:0] node10907;
	wire [4-1:0] node10910;
	wire [4-1:0] node10913;
	wire [4-1:0] node10914;
	wire [4-1:0] node10915;
	wire [4-1:0] node10918;
	wire [4-1:0] node10921;
	wire [4-1:0] node10923;
	wire [4-1:0] node10926;
	wire [4-1:0] node10927;
	wire [4-1:0] node10928;
	wire [4-1:0] node10929;
	wire [4-1:0] node10930;
	wire [4-1:0] node10933;
	wire [4-1:0] node10936;
	wire [4-1:0] node10938;
	wire [4-1:0] node10941;
	wire [4-1:0] node10942;
	wire [4-1:0] node10943;
	wire [4-1:0] node10946;
	wire [4-1:0] node10949;
	wire [4-1:0] node10950;
	wire [4-1:0] node10953;
	wire [4-1:0] node10956;
	wire [4-1:0] node10957;
	wire [4-1:0] node10958;
	wire [4-1:0] node10961;
	wire [4-1:0] node10964;
	wire [4-1:0] node10965;
	wire [4-1:0] node10966;
	wire [4-1:0] node10969;
	wire [4-1:0] node10972;
	wire [4-1:0] node10973;
	wire [4-1:0] node10976;
	wire [4-1:0] node10979;
	wire [4-1:0] node10980;
	wire [4-1:0] node10981;
	wire [4-1:0] node10982;
	wire [4-1:0] node10983;
	wire [4-1:0] node10984;
	wire [4-1:0] node10985;
	wire [4-1:0] node10988;
	wire [4-1:0] node10991;
	wire [4-1:0] node10992;
	wire [4-1:0] node10995;
	wire [4-1:0] node10998;
	wire [4-1:0] node10999;
	wire [4-1:0] node11000;
	wire [4-1:0] node11003;
	wire [4-1:0] node11006;
	wire [4-1:0] node11007;
	wire [4-1:0] node11010;
	wire [4-1:0] node11013;
	wire [4-1:0] node11014;
	wire [4-1:0] node11015;
	wire [4-1:0] node11016;
	wire [4-1:0] node11019;
	wire [4-1:0] node11022;
	wire [4-1:0] node11023;
	wire [4-1:0] node11026;
	wire [4-1:0] node11029;
	wire [4-1:0] node11030;
	wire [4-1:0] node11031;
	wire [4-1:0] node11034;
	wire [4-1:0] node11037;
	wire [4-1:0] node11038;
	wire [4-1:0] node11041;
	wire [4-1:0] node11044;
	wire [4-1:0] node11045;
	wire [4-1:0] node11046;
	wire [4-1:0] node11047;
	wire [4-1:0] node11048;
	wire [4-1:0] node11051;
	wire [4-1:0] node11054;
	wire [4-1:0] node11055;
	wire [4-1:0] node11059;
	wire [4-1:0] node11060;
	wire [4-1:0] node11061;
	wire [4-1:0] node11064;
	wire [4-1:0] node11067;
	wire [4-1:0] node11068;
	wire [4-1:0] node11071;
	wire [4-1:0] node11074;
	wire [4-1:0] node11075;
	wire [4-1:0] node11076;
	wire [4-1:0] node11077;
	wire [4-1:0] node11080;
	wire [4-1:0] node11083;
	wire [4-1:0] node11084;
	wire [4-1:0] node11087;
	wire [4-1:0] node11090;
	wire [4-1:0] node11091;
	wire [4-1:0] node11092;
	wire [4-1:0] node11095;
	wire [4-1:0] node11098;
	wire [4-1:0] node11100;
	wire [4-1:0] node11103;
	wire [4-1:0] node11104;
	wire [4-1:0] node11105;
	wire [4-1:0] node11106;
	wire [4-1:0] node11107;
	wire [4-1:0] node11109;
	wire [4-1:0] node11112;
	wire [4-1:0] node11113;
	wire [4-1:0] node11116;
	wire [4-1:0] node11119;
	wire [4-1:0] node11120;
	wire [4-1:0] node11121;
	wire [4-1:0] node11124;
	wire [4-1:0] node11127;
	wire [4-1:0] node11128;
	wire [4-1:0] node11132;
	wire [4-1:0] node11133;
	wire [4-1:0] node11134;
	wire [4-1:0] node11135;
	wire [4-1:0] node11138;
	wire [4-1:0] node11141;
	wire [4-1:0] node11142;
	wire [4-1:0] node11145;
	wire [4-1:0] node11148;
	wire [4-1:0] node11149;
	wire [4-1:0] node11150;
	wire [4-1:0] node11153;
	wire [4-1:0] node11156;
	wire [4-1:0] node11157;
	wire [4-1:0] node11160;
	wire [4-1:0] node11163;
	wire [4-1:0] node11164;
	wire [4-1:0] node11165;
	wire [4-1:0] node11166;
	wire [4-1:0] node11167;
	wire [4-1:0] node11170;
	wire [4-1:0] node11173;
	wire [4-1:0] node11174;
	wire [4-1:0] node11177;
	wire [4-1:0] node11180;
	wire [4-1:0] node11181;
	wire [4-1:0] node11182;
	wire [4-1:0] node11185;
	wire [4-1:0] node11188;
	wire [4-1:0] node11189;
	wire [4-1:0] node11193;
	wire [4-1:0] node11194;
	wire [4-1:0] node11195;
	wire [4-1:0] node11196;
	wire [4-1:0] node11199;
	wire [4-1:0] node11202;
	wire [4-1:0] node11203;
	wire [4-1:0] node11206;
	wire [4-1:0] node11209;
	wire [4-1:0] node11210;
	wire [4-1:0] node11212;
	wire [4-1:0] node11215;
	wire [4-1:0] node11216;
	wire [4-1:0] node11219;
	wire [4-1:0] node11222;
	wire [4-1:0] node11223;
	wire [4-1:0] node11224;
	wire [4-1:0] node11225;
	wire [4-1:0] node11226;
	wire [4-1:0] node11227;
	wire [4-1:0] node11228;
	wire [4-1:0] node11229;
	wire [4-1:0] node11232;
	wire [4-1:0] node11235;
	wire [4-1:0] node11236;
	wire [4-1:0] node11239;
	wire [4-1:0] node11242;
	wire [4-1:0] node11243;
	wire [4-1:0] node11244;
	wire [4-1:0] node11247;
	wire [4-1:0] node11250;
	wire [4-1:0] node11251;
	wire [4-1:0] node11254;
	wire [4-1:0] node11257;
	wire [4-1:0] node11258;
	wire [4-1:0] node11259;
	wire [4-1:0] node11260;
	wire [4-1:0] node11263;
	wire [4-1:0] node11266;
	wire [4-1:0] node11267;
	wire [4-1:0] node11270;
	wire [4-1:0] node11273;
	wire [4-1:0] node11274;
	wire [4-1:0] node11275;
	wire [4-1:0] node11278;
	wire [4-1:0] node11281;
	wire [4-1:0] node11282;
	wire [4-1:0] node11285;
	wire [4-1:0] node11288;
	wire [4-1:0] node11289;
	wire [4-1:0] node11290;
	wire [4-1:0] node11291;
	wire [4-1:0] node11292;
	wire [4-1:0] node11295;
	wire [4-1:0] node11298;
	wire [4-1:0] node11299;
	wire [4-1:0] node11302;
	wire [4-1:0] node11305;
	wire [4-1:0] node11306;
	wire [4-1:0] node11307;
	wire [4-1:0] node11310;
	wire [4-1:0] node11313;
	wire [4-1:0] node11314;
	wire [4-1:0] node11317;
	wire [4-1:0] node11320;
	wire [4-1:0] node11321;
	wire [4-1:0] node11322;
	wire [4-1:0] node11323;
	wire [4-1:0] node11326;
	wire [4-1:0] node11329;
	wire [4-1:0] node11330;
	wire [4-1:0] node11333;
	wire [4-1:0] node11336;
	wire [4-1:0] node11337;
	wire [4-1:0] node11338;
	wire [4-1:0] node11341;
	wire [4-1:0] node11344;
	wire [4-1:0] node11345;
	wire [4-1:0] node11348;
	wire [4-1:0] node11351;
	wire [4-1:0] node11352;
	wire [4-1:0] node11353;
	wire [4-1:0] node11354;
	wire [4-1:0] node11355;
	wire [4-1:0] node11356;
	wire [4-1:0] node11359;
	wire [4-1:0] node11363;
	wire [4-1:0] node11364;
	wire [4-1:0] node11365;
	wire [4-1:0] node11368;
	wire [4-1:0] node11371;
	wire [4-1:0] node11372;
	wire [4-1:0] node11375;
	wire [4-1:0] node11378;
	wire [4-1:0] node11379;
	wire [4-1:0] node11380;
	wire [4-1:0] node11381;
	wire [4-1:0] node11384;
	wire [4-1:0] node11387;
	wire [4-1:0] node11388;
	wire [4-1:0] node11391;
	wire [4-1:0] node11394;
	wire [4-1:0] node11395;
	wire [4-1:0] node11396;
	wire [4-1:0] node11399;
	wire [4-1:0] node11402;
	wire [4-1:0] node11403;
	wire [4-1:0] node11406;
	wire [4-1:0] node11409;
	wire [4-1:0] node11410;
	wire [4-1:0] node11411;
	wire [4-1:0] node11412;
	wire [4-1:0] node11413;
	wire [4-1:0] node11416;
	wire [4-1:0] node11419;
	wire [4-1:0] node11420;
	wire [4-1:0] node11423;
	wire [4-1:0] node11426;
	wire [4-1:0] node11427;
	wire [4-1:0] node11428;
	wire [4-1:0] node11431;
	wire [4-1:0] node11434;
	wire [4-1:0] node11435;
	wire [4-1:0] node11438;
	wire [4-1:0] node11441;
	wire [4-1:0] node11442;
	wire [4-1:0] node11443;
	wire [4-1:0] node11444;
	wire [4-1:0] node11447;
	wire [4-1:0] node11450;
	wire [4-1:0] node11451;
	wire [4-1:0] node11454;
	wire [4-1:0] node11457;
	wire [4-1:0] node11458;
	wire [4-1:0] node11459;
	wire [4-1:0] node11462;
	wire [4-1:0] node11465;
	wire [4-1:0] node11466;
	wire [4-1:0] node11469;
	wire [4-1:0] node11472;
	wire [4-1:0] node11473;
	wire [4-1:0] node11474;
	wire [4-1:0] node11475;
	wire [4-1:0] node11476;
	wire [4-1:0] node11477;
	wire [4-1:0] node11478;
	wire [4-1:0] node11481;
	wire [4-1:0] node11484;
	wire [4-1:0] node11486;
	wire [4-1:0] node11489;
	wire [4-1:0] node11490;
	wire [4-1:0] node11491;
	wire [4-1:0] node11494;
	wire [4-1:0] node11497;
	wire [4-1:0] node11498;
	wire [4-1:0] node11501;
	wire [4-1:0] node11504;
	wire [4-1:0] node11505;
	wire [4-1:0] node11506;
	wire [4-1:0] node11507;
	wire [4-1:0] node11510;
	wire [4-1:0] node11513;
	wire [4-1:0] node11514;
	wire [4-1:0] node11517;
	wire [4-1:0] node11520;
	wire [4-1:0] node11521;
	wire [4-1:0] node11522;
	wire [4-1:0] node11526;
	wire [4-1:0] node11527;
	wire [4-1:0] node11530;
	wire [4-1:0] node11533;
	wire [4-1:0] node11534;
	wire [4-1:0] node11535;
	wire [4-1:0] node11536;
	wire [4-1:0] node11537;
	wire [4-1:0] node11540;
	wire [4-1:0] node11543;
	wire [4-1:0] node11544;
	wire [4-1:0] node11547;
	wire [4-1:0] node11550;
	wire [4-1:0] node11551;
	wire [4-1:0] node11552;
	wire [4-1:0] node11555;
	wire [4-1:0] node11558;
	wire [4-1:0] node11559;
	wire [4-1:0] node11562;
	wire [4-1:0] node11565;
	wire [4-1:0] node11566;
	wire [4-1:0] node11567;
	wire [4-1:0] node11568;
	wire [4-1:0] node11571;
	wire [4-1:0] node11574;
	wire [4-1:0] node11575;
	wire [4-1:0] node11578;
	wire [4-1:0] node11581;
	wire [4-1:0] node11582;
	wire [4-1:0] node11583;
	wire [4-1:0] node11586;
	wire [4-1:0] node11589;
	wire [4-1:0] node11590;
	wire [4-1:0] node11593;
	wire [4-1:0] node11596;
	wire [4-1:0] node11597;
	wire [4-1:0] node11598;
	wire [4-1:0] node11599;
	wire [4-1:0] node11600;
	wire [4-1:0] node11601;
	wire [4-1:0] node11604;
	wire [4-1:0] node11607;
	wire [4-1:0] node11608;
	wire [4-1:0] node11612;
	wire [4-1:0] node11613;
	wire [4-1:0] node11614;
	wire [4-1:0] node11617;
	wire [4-1:0] node11620;
	wire [4-1:0] node11622;
	wire [4-1:0] node11625;
	wire [4-1:0] node11626;
	wire [4-1:0] node11627;
	wire [4-1:0] node11628;
	wire [4-1:0] node11631;
	wire [4-1:0] node11634;
	wire [4-1:0] node11635;
	wire [4-1:0] node11638;
	wire [4-1:0] node11641;
	wire [4-1:0] node11642;
	wire [4-1:0] node11643;
	wire [4-1:0] node11646;
	wire [4-1:0] node11649;
	wire [4-1:0] node11650;
	wire [4-1:0] node11653;
	wire [4-1:0] node11656;
	wire [4-1:0] node11657;
	wire [4-1:0] node11658;
	wire [4-1:0] node11659;
	wire [4-1:0] node11660;
	wire [4-1:0] node11663;
	wire [4-1:0] node11666;
	wire [4-1:0] node11667;
	wire [4-1:0] node11670;
	wire [4-1:0] node11673;
	wire [4-1:0] node11674;
	wire [4-1:0] node11675;
	wire [4-1:0] node11678;
	wire [4-1:0] node11681;
	wire [4-1:0] node11682;
	wire [4-1:0] node11685;
	wire [4-1:0] node11688;
	wire [4-1:0] node11689;
	wire [4-1:0] node11690;
	wire [4-1:0] node11691;
	wire [4-1:0] node11694;
	wire [4-1:0] node11697;
	wire [4-1:0] node11699;
	wire [4-1:0] node11702;
	wire [4-1:0] node11703;
	wire [4-1:0] node11704;
	wire [4-1:0] node11707;
	wire [4-1:0] node11710;
	wire [4-1:0] node11711;
	wire [4-1:0] node11714;
	wire [4-1:0] node11717;
	wire [4-1:0] node11718;
	wire [4-1:0] node11719;
	wire [4-1:0] node11720;
	wire [4-1:0] node11721;
	wire [4-1:0] node11722;
	wire [4-1:0] node11723;
	wire [4-1:0] node11726;
	wire [4-1:0] node11729;
	wire [4-1:0] node11730;
	wire [4-1:0] node11731;
	wire [4-1:0] node11732;
	wire [4-1:0] node11735;
	wire [4-1:0] node11738;
	wire [4-1:0] node11739;
	wire [4-1:0] node11742;
	wire [4-1:0] node11745;
	wire [4-1:0] node11746;
	wire [4-1:0] node11747;
	wire [4-1:0] node11750;
	wire [4-1:0] node11753;
	wire [4-1:0] node11754;
	wire [4-1:0] node11757;
	wire [4-1:0] node11760;
	wire [4-1:0] node11761;
	wire [4-1:0] node11762;
	wire [4-1:0] node11763;
	wire [4-1:0] node11766;
	wire [4-1:0] node11769;
	wire [4-1:0] node11770;
	wire [4-1:0] node11773;
	wire [4-1:0] node11776;
	wire [4-1:0] node11777;
	wire [4-1:0] node11778;
	wire [4-1:0] node11781;
	wire [4-1:0] node11784;
	wire [4-1:0] node11785;
	wire [4-1:0] node11786;
	wire [4-1:0] node11789;
	wire [4-1:0] node11792;
	wire [4-1:0] node11793;
	wire [4-1:0] node11796;
	wire [4-1:0] node11799;
	wire [4-1:0] node11800;
	wire [4-1:0] node11801;
	wire [4-1:0] node11802;
	wire [4-1:0] node11803;
	wire [4-1:0] node11804;
	wire [4-1:0] node11808;
	wire [4-1:0] node11809;
	wire [4-1:0] node11813;
	wire [4-1:0] node11814;
	wire [4-1:0] node11815;
	wire [4-1:0] node11819;
	wire [4-1:0] node11820;
	wire [4-1:0] node11824;
	wire [4-1:0] node11825;
	wire [4-1:0] node11826;
	wire [4-1:0] node11827;
	wire [4-1:0] node11831;
	wire [4-1:0] node11832;
	wire [4-1:0] node11836;
	wire [4-1:0] node11837;
	wire [4-1:0] node11838;
	wire [4-1:0] node11842;
	wire [4-1:0] node11843;
	wire [4-1:0] node11847;
	wire [4-1:0] node11848;
	wire [4-1:0] node11849;
	wire [4-1:0] node11850;
	wire [4-1:0] node11854;
	wire [4-1:0] node11855;
	wire [4-1:0] node11859;
	wire [4-1:0] node11860;
	wire [4-1:0] node11861;
	wire [4-1:0] node11865;
	wire [4-1:0] node11866;
	wire [4-1:0] node11870;
	wire [4-1:0] node11871;
	wire [4-1:0] node11872;
	wire [4-1:0] node11873;
	wire [4-1:0] node11874;
	wire [4-1:0] node11875;
	wire [4-1:0] node11876;
	wire [4-1:0] node11879;
	wire [4-1:0] node11882;
	wire [4-1:0] node11883;
	wire [4-1:0] node11886;
	wire [4-1:0] node11889;
	wire [4-1:0] node11890;
	wire [4-1:0] node11891;
	wire [4-1:0] node11894;
	wire [4-1:0] node11897;
	wire [4-1:0] node11898;
	wire [4-1:0] node11901;
	wire [4-1:0] node11904;
	wire [4-1:0] node11905;
	wire [4-1:0] node11906;
	wire [4-1:0] node11907;
	wire [4-1:0] node11910;
	wire [4-1:0] node11913;
	wire [4-1:0] node11914;
	wire [4-1:0] node11917;
	wire [4-1:0] node11920;
	wire [4-1:0] node11921;
	wire [4-1:0] node11923;
	wire [4-1:0] node11926;
	wire [4-1:0] node11928;
	wire [4-1:0] node11931;
	wire [4-1:0] node11932;
	wire [4-1:0] node11933;
	wire [4-1:0] node11934;
	wire [4-1:0] node11935;
	wire [4-1:0] node11938;
	wire [4-1:0] node11941;
	wire [4-1:0] node11942;
	wire [4-1:0] node11945;
	wire [4-1:0] node11948;
	wire [4-1:0] node11949;
	wire [4-1:0] node11950;
	wire [4-1:0] node11953;
	wire [4-1:0] node11956;
	wire [4-1:0] node11957;
	wire [4-1:0] node11960;
	wire [4-1:0] node11963;
	wire [4-1:0] node11964;
	wire [4-1:0] node11965;
	wire [4-1:0] node11966;
	wire [4-1:0] node11969;
	wire [4-1:0] node11972;
	wire [4-1:0] node11973;
	wire [4-1:0] node11976;
	wire [4-1:0] node11979;
	wire [4-1:0] node11980;
	wire [4-1:0] node11981;
	wire [4-1:0] node11984;
	wire [4-1:0] node11987;
	wire [4-1:0] node11988;
	wire [4-1:0] node11991;
	wire [4-1:0] node11994;
	wire [4-1:0] node11995;
	wire [4-1:0] node11996;
	wire [4-1:0] node11997;
	wire [4-1:0] node11998;
	wire [4-1:0] node11999;
	wire [4-1:0] node12002;
	wire [4-1:0] node12005;
	wire [4-1:0] node12006;
	wire [4-1:0] node12009;
	wire [4-1:0] node12012;
	wire [4-1:0] node12013;
	wire [4-1:0] node12014;
	wire [4-1:0] node12018;
	wire [4-1:0] node12021;
	wire [4-1:0] node12022;
	wire [4-1:0] node12023;
	wire [4-1:0] node12024;
	wire [4-1:0] node12027;
	wire [4-1:0] node12030;
	wire [4-1:0] node12031;
	wire [4-1:0] node12034;
	wire [4-1:0] node12037;
	wire [4-1:0] node12038;
	wire [4-1:0] node12039;
	wire [4-1:0] node12043;
	wire [4-1:0] node12046;
	wire [4-1:0] node12047;
	wire [4-1:0] node12048;
	wire [4-1:0] node12049;
	wire [4-1:0] node12050;
	wire [4-1:0] node12053;
	wire [4-1:0] node12056;
	wire [4-1:0] node12057;
	wire [4-1:0] node12060;
	wire [4-1:0] node12063;
	wire [4-1:0] node12064;
	wire [4-1:0] node12065;
	wire [4-1:0] node12069;
	wire [4-1:0] node12072;
	wire [4-1:0] node12073;
	wire [4-1:0] node12074;
	wire [4-1:0] node12075;
	wire [4-1:0] node12078;
	wire [4-1:0] node12081;
	wire [4-1:0] node12082;
	wire [4-1:0] node12085;
	wire [4-1:0] node12088;
	wire [4-1:0] node12089;
	wire [4-1:0] node12090;
	wire [4-1:0] node12094;
	wire [4-1:0] node12097;
	wire [4-1:0] node12098;
	wire [4-1:0] node12099;
	wire [4-1:0] node12100;
	wire [4-1:0] node12101;
	wire [4-1:0] node12102;
	wire [4-1:0] node12103;
	wire [4-1:0] node12106;
	wire [4-1:0] node12109;
	wire [4-1:0] node12110;
	wire [4-1:0] node12113;
	wire [4-1:0] node12116;
	wire [4-1:0] node12117;
	wire [4-1:0] node12118;
	wire [4-1:0] node12119;
	wire [4-1:0] node12123;
	wire [4-1:0] node12124;
	wire [4-1:0] node12127;
	wire [4-1:0] node12130;
	wire [4-1:0] node12131;
	wire [4-1:0] node12134;
	wire [4-1:0] node12137;
	wire [4-1:0] node12138;
	wire [4-1:0] node12139;
	wire [4-1:0] node12140;
	wire [4-1:0] node12143;
	wire [4-1:0] node12146;
	wire [4-1:0] node12147;
	wire [4-1:0] node12150;
	wire [4-1:0] node12153;
	wire [4-1:0] node12154;
	wire [4-1:0] node12155;
	wire [4-1:0] node12158;
	wire [4-1:0] node12161;
	wire [4-1:0] node12162;
	wire [4-1:0] node12165;
	wire [4-1:0] node12168;
	wire [4-1:0] node12169;
	wire [4-1:0] node12170;
	wire [4-1:0] node12171;
	wire [4-1:0] node12172;
	wire [4-1:0] node12176;
	wire [4-1:0] node12179;
	wire [4-1:0] node12180;
	wire [4-1:0] node12181;
	wire [4-1:0] node12184;
	wire [4-1:0] node12187;
	wire [4-1:0] node12188;
	wire [4-1:0] node12189;
	wire [4-1:0] node12193;
	wire [4-1:0] node12194;
	wire [4-1:0] node12197;
	wire [4-1:0] node12200;
	wire [4-1:0] node12201;
	wire [4-1:0] node12202;
	wire [4-1:0] node12203;
	wire [4-1:0] node12207;
	wire [4-1:0] node12210;
	wire [4-1:0] node12211;
	wire [4-1:0] node12212;
	wire [4-1:0] node12216;
	wire [4-1:0] node12219;
	wire [4-1:0] node12220;
	wire [4-1:0] node12221;
	wire [4-1:0] node12222;
	wire [4-1:0] node12223;
	wire [4-1:0] node12224;
	wire [4-1:0] node12225;
	wire [4-1:0] node12228;
	wire [4-1:0] node12231;
	wire [4-1:0] node12232;
	wire [4-1:0] node12235;
	wire [4-1:0] node12238;
	wire [4-1:0] node12239;
	wire [4-1:0] node12242;
	wire [4-1:0] node12245;
	wire [4-1:0] node12246;
	wire [4-1:0] node12247;
	wire [4-1:0] node12251;
	wire [4-1:0] node12254;
	wire [4-1:0] node12255;
	wire [4-1:0] node12256;
	wire [4-1:0] node12257;
	wire [4-1:0] node12260;
	wire [4-1:0] node12263;
	wire [4-1:0] node12264;
	wire [4-1:0] node12267;
	wire [4-1:0] node12270;
	wire [4-1:0] node12271;
	wire [4-1:0] node12272;
	wire [4-1:0] node12276;
	wire [4-1:0] node12279;
	wire [4-1:0] node12280;
	wire [4-1:0] node12281;
	wire [4-1:0] node12282;
	wire [4-1:0] node12283;
	wire [4-1:0] node12284;
	wire [4-1:0] node12287;
	wire [4-1:0] node12290;
	wire [4-1:0] node12291;
	wire [4-1:0] node12294;
	wire [4-1:0] node12297;
	wire [4-1:0] node12298;
	wire [4-1:0] node12301;
	wire [4-1:0] node12304;
	wire [4-1:0] node12305;
	wire [4-1:0] node12306;
	wire [4-1:0] node12310;
	wire [4-1:0] node12313;
	wire [4-1:0] node12314;
	wire [4-1:0] node12315;
	wire [4-1:0] node12316;
	wire [4-1:0] node12319;
	wire [4-1:0] node12322;
	wire [4-1:0] node12323;
	wire [4-1:0] node12326;
	wire [4-1:0] node12329;
	wire [4-1:0] node12330;
	wire [4-1:0] node12331;
	wire [4-1:0] node12335;
	wire [4-1:0] node12338;
	wire [4-1:0] node12339;
	wire [4-1:0] node12340;
	wire [4-1:0] node12341;
	wire [4-1:0] node12342;
	wire [4-1:0] node12343;
	wire [4-1:0] node12344;
	wire [4-1:0] node12345;
	wire [4-1:0] node12346;
	wire [4-1:0] node12347;
	wire [4-1:0] node12350;
	wire [4-1:0] node12353;
	wire [4-1:0] node12354;
	wire [4-1:0] node12358;
	wire [4-1:0] node12359;
	wire [4-1:0] node12360;
	wire [4-1:0] node12363;
	wire [4-1:0] node12366;
	wire [4-1:0] node12367;
	wire [4-1:0] node12370;
	wire [4-1:0] node12373;
	wire [4-1:0] node12374;
	wire [4-1:0] node12375;
	wire [4-1:0] node12376;
	wire [4-1:0] node12379;
	wire [4-1:0] node12382;
	wire [4-1:0] node12383;
	wire [4-1:0] node12386;
	wire [4-1:0] node12389;
	wire [4-1:0] node12390;
	wire [4-1:0] node12391;
	wire [4-1:0] node12394;
	wire [4-1:0] node12397;
	wire [4-1:0] node12398;
	wire [4-1:0] node12401;
	wire [4-1:0] node12404;
	wire [4-1:0] node12405;
	wire [4-1:0] node12406;
	wire [4-1:0] node12407;
	wire [4-1:0] node12408;
	wire [4-1:0] node12411;
	wire [4-1:0] node12414;
	wire [4-1:0] node12415;
	wire [4-1:0] node12418;
	wire [4-1:0] node12421;
	wire [4-1:0] node12422;
	wire [4-1:0] node12423;
	wire [4-1:0] node12426;
	wire [4-1:0] node12429;
	wire [4-1:0] node12430;
	wire [4-1:0] node12433;
	wire [4-1:0] node12436;
	wire [4-1:0] node12437;
	wire [4-1:0] node12438;
	wire [4-1:0] node12439;
	wire [4-1:0] node12442;
	wire [4-1:0] node12445;
	wire [4-1:0] node12446;
	wire [4-1:0] node12449;
	wire [4-1:0] node12452;
	wire [4-1:0] node12453;
	wire [4-1:0] node12454;
	wire [4-1:0] node12457;
	wire [4-1:0] node12460;
	wire [4-1:0] node12461;
	wire [4-1:0] node12464;
	wire [4-1:0] node12467;
	wire [4-1:0] node12468;
	wire [4-1:0] node12469;
	wire [4-1:0] node12470;
	wire [4-1:0] node12471;
	wire [4-1:0] node12472;
	wire [4-1:0] node12475;
	wire [4-1:0] node12478;
	wire [4-1:0] node12479;
	wire [4-1:0] node12482;
	wire [4-1:0] node12485;
	wire [4-1:0] node12486;
	wire [4-1:0] node12487;
	wire [4-1:0] node12490;
	wire [4-1:0] node12493;
	wire [4-1:0] node12494;
	wire [4-1:0] node12498;
	wire [4-1:0] node12499;
	wire [4-1:0] node12500;
	wire [4-1:0] node12501;
	wire [4-1:0] node12504;
	wire [4-1:0] node12507;
	wire [4-1:0] node12508;
	wire [4-1:0] node12511;
	wire [4-1:0] node12514;
	wire [4-1:0] node12515;
	wire [4-1:0] node12516;
	wire [4-1:0] node12519;
	wire [4-1:0] node12522;
	wire [4-1:0] node12523;
	wire [4-1:0] node12526;
	wire [4-1:0] node12529;
	wire [4-1:0] node12530;
	wire [4-1:0] node12531;
	wire [4-1:0] node12532;
	wire [4-1:0] node12533;
	wire [4-1:0] node12536;
	wire [4-1:0] node12539;
	wire [4-1:0] node12540;
	wire [4-1:0] node12543;
	wire [4-1:0] node12546;
	wire [4-1:0] node12547;
	wire [4-1:0] node12549;
	wire [4-1:0] node12552;
	wire [4-1:0] node12554;
	wire [4-1:0] node12557;
	wire [4-1:0] node12558;
	wire [4-1:0] node12559;
	wire [4-1:0] node12560;
	wire [4-1:0] node12564;
	wire [4-1:0] node12565;
	wire [4-1:0] node12568;
	wire [4-1:0] node12571;
	wire [4-1:0] node12572;
	wire [4-1:0] node12573;
	wire [4-1:0] node12576;
	wire [4-1:0] node12579;
	wire [4-1:0] node12580;
	wire [4-1:0] node12583;
	wire [4-1:0] node12586;
	wire [4-1:0] node12587;
	wire [4-1:0] node12588;
	wire [4-1:0] node12589;
	wire [4-1:0] node12590;
	wire [4-1:0] node12591;
	wire [4-1:0] node12594;
	wire [4-1:0] node12597;
	wire [4-1:0] node12598;
	wire [4-1:0] node12599;
	wire [4-1:0] node12602;
	wire [4-1:0] node12605;
	wire [4-1:0] node12606;
	wire [4-1:0] node12609;
	wire [4-1:0] node12612;
	wire [4-1:0] node12613;
	wire [4-1:0] node12614;
	wire [4-1:0] node12615;
	wire [4-1:0] node12618;
	wire [4-1:0] node12621;
	wire [4-1:0] node12622;
	wire [4-1:0] node12625;
	wire [4-1:0] node12628;
	wire [4-1:0] node12629;
	wire [4-1:0] node12630;
	wire [4-1:0] node12633;
	wire [4-1:0] node12636;
	wire [4-1:0] node12637;
	wire [4-1:0] node12640;
	wire [4-1:0] node12643;
	wire [4-1:0] node12644;
	wire [4-1:0] node12645;
	wire [4-1:0] node12646;
	wire [4-1:0] node12647;
	wire [4-1:0] node12650;
	wire [4-1:0] node12653;
	wire [4-1:0] node12654;
	wire [4-1:0] node12658;
	wire [4-1:0] node12659;
	wire [4-1:0] node12660;
	wire [4-1:0] node12663;
	wire [4-1:0] node12666;
	wire [4-1:0] node12667;
	wire [4-1:0] node12671;
	wire [4-1:0] node12672;
	wire [4-1:0] node12673;
	wire [4-1:0] node12674;
	wire [4-1:0] node12677;
	wire [4-1:0] node12680;
	wire [4-1:0] node12681;
	wire [4-1:0] node12684;
	wire [4-1:0] node12687;
	wire [4-1:0] node12688;
	wire [4-1:0] node12689;
	wire [4-1:0] node12692;
	wire [4-1:0] node12695;
	wire [4-1:0] node12696;
	wire [4-1:0] node12699;
	wire [4-1:0] node12702;
	wire [4-1:0] node12703;
	wire [4-1:0] node12704;
	wire [4-1:0] node12705;
	wire [4-1:0] node12706;
	wire [4-1:0] node12707;
	wire [4-1:0] node12710;
	wire [4-1:0] node12713;
	wire [4-1:0] node12714;
	wire [4-1:0] node12717;
	wire [4-1:0] node12720;
	wire [4-1:0] node12721;
	wire [4-1:0] node12722;
	wire [4-1:0] node12726;
	wire [4-1:0] node12727;
	wire [4-1:0] node12730;
	wire [4-1:0] node12733;
	wire [4-1:0] node12734;
	wire [4-1:0] node12735;
	wire [4-1:0] node12736;
	wire [4-1:0] node12739;
	wire [4-1:0] node12742;
	wire [4-1:0] node12744;
	wire [4-1:0] node12747;
	wire [4-1:0] node12748;
	wire [4-1:0] node12749;
	wire [4-1:0] node12752;
	wire [4-1:0] node12755;
	wire [4-1:0] node12757;
	wire [4-1:0] node12760;
	wire [4-1:0] node12761;
	wire [4-1:0] node12762;
	wire [4-1:0] node12763;
	wire [4-1:0] node12764;
	wire [4-1:0] node12767;
	wire [4-1:0] node12770;
	wire [4-1:0] node12771;
	wire [4-1:0] node12774;
	wire [4-1:0] node12777;
	wire [4-1:0] node12778;
	wire [4-1:0] node12779;
	wire [4-1:0] node12782;
	wire [4-1:0] node12785;
	wire [4-1:0] node12786;
	wire [4-1:0] node12789;
	wire [4-1:0] node12792;
	wire [4-1:0] node12793;
	wire [4-1:0] node12794;
	wire [4-1:0] node12795;
	wire [4-1:0] node12798;
	wire [4-1:0] node12801;
	wire [4-1:0] node12802;
	wire [4-1:0] node12805;
	wire [4-1:0] node12808;
	wire [4-1:0] node12809;
	wire [4-1:0] node12810;
	wire [4-1:0] node12814;
	wire [4-1:0] node12816;
	wire [4-1:0] node12819;
	wire [4-1:0] node12820;
	wire [4-1:0] node12821;
	wire [4-1:0] node12822;
	wire [4-1:0] node12823;
	wire [4-1:0] node12824;
	wire [4-1:0] node12825;
	wire [4-1:0] node12826;
	wire [4-1:0] node12829;
	wire [4-1:0] node12832;
	wire [4-1:0] node12833;
	wire [4-1:0] node12836;
	wire [4-1:0] node12839;
	wire [4-1:0] node12840;
	wire [4-1:0] node12841;
	wire [4-1:0] node12844;
	wire [4-1:0] node12847;
	wire [4-1:0] node12848;
	wire [4-1:0] node12851;
	wire [4-1:0] node12854;
	wire [4-1:0] node12855;
	wire [4-1:0] node12856;
	wire [4-1:0] node12857;
	wire [4-1:0] node12860;
	wire [4-1:0] node12863;
	wire [4-1:0] node12864;
	wire [4-1:0] node12867;
	wire [4-1:0] node12870;
	wire [4-1:0] node12871;
	wire [4-1:0] node12872;
	wire [4-1:0] node12875;
	wire [4-1:0] node12878;
	wire [4-1:0] node12879;
	wire [4-1:0] node12882;
	wire [4-1:0] node12885;
	wire [4-1:0] node12886;
	wire [4-1:0] node12887;
	wire [4-1:0] node12888;
	wire [4-1:0] node12889;
	wire [4-1:0] node12892;
	wire [4-1:0] node12895;
	wire [4-1:0] node12897;
	wire [4-1:0] node12900;
	wire [4-1:0] node12901;
	wire [4-1:0] node12903;
	wire [4-1:0] node12906;
	wire [4-1:0] node12907;
	wire [4-1:0] node12910;
	wire [4-1:0] node12913;
	wire [4-1:0] node12914;
	wire [4-1:0] node12915;
	wire [4-1:0] node12916;
	wire [4-1:0] node12920;
	wire [4-1:0] node12921;
	wire [4-1:0] node12924;
	wire [4-1:0] node12927;
	wire [4-1:0] node12928;
	wire [4-1:0] node12929;
	wire [4-1:0] node12932;
	wire [4-1:0] node12935;
	wire [4-1:0] node12936;
	wire [4-1:0] node12939;
	wire [4-1:0] node12942;
	wire [4-1:0] node12943;
	wire [4-1:0] node12944;
	wire [4-1:0] node12945;
	wire [4-1:0] node12946;
	wire [4-1:0] node12947;
	wire [4-1:0] node12950;
	wire [4-1:0] node12953;
	wire [4-1:0] node12954;
	wire [4-1:0] node12957;
	wire [4-1:0] node12960;
	wire [4-1:0] node12961;
	wire [4-1:0] node12962;
	wire [4-1:0] node12965;
	wire [4-1:0] node12968;
	wire [4-1:0] node12969;
	wire [4-1:0] node12972;
	wire [4-1:0] node12975;
	wire [4-1:0] node12976;
	wire [4-1:0] node12977;
	wire [4-1:0] node12978;
	wire [4-1:0] node12981;
	wire [4-1:0] node12984;
	wire [4-1:0] node12985;
	wire [4-1:0] node12988;
	wire [4-1:0] node12991;
	wire [4-1:0] node12992;
	wire [4-1:0] node12993;
	wire [4-1:0] node12996;
	wire [4-1:0] node12999;
	wire [4-1:0] node13000;
	wire [4-1:0] node13003;
	wire [4-1:0] node13006;
	wire [4-1:0] node13007;
	wire [4-1:0] node13008;
	wire [4-1:0] node13009;
	wire [4-1:0] node13011;
	wire [4-1:0] node13014;
	wire [4-1:0] node13015;
	wire [4-1:0] node13018;
	wire [4-1:0] node13021;
	wire [4-1:0] node13022;
	wire [4-1:0] node13023;
	wire [4-1:0] node13026;
	wire [4-1:0] node13029;
	wire [4-1:0] node13030;
	wire [4-1:0] node13033;
	wire [4-1:0] node13036;
	wire [4-1:0] node13037;
	wire [4-1:0] node13038;
	wire [4-1:0] node13040;
	wire [4-1:0] node13043;
	wire [4-1:0] node13044;
	wire [4-1:0] node13047;
	wire [4-1:0] node13050;
	wire [4-1:0] node13051;
	wire [4-1:0] node13052;
	wire [4-1:0] node13055;
	wire [4-1:0] node13058;
	wire [4-1:0] node13059;
	wire [4-1:0] node13062;
	wire [4-1:0] node13065;
	wire [4-1:0] node13066;
	wire [4-1:0] node13067;
	wire [4-1:0] node13068;
	wire [4-1:0] node13069;
	wire [4-1:0] node13070;
	wire [4-1:0] node13072;
	wire [4-1:0] node13075;
	wire [4-1:0] node13076;
	wire [4-1:0] node13079;
	wire [4-1:0] node13082;
	wire [4-1:0] node13083;
	wire [4-1:0] node13084;
	wire [4-1:0] node13087;
	wire [4-1:0] node13090;
	wire [4-1:0] node13091;
	wire [4-1:0] node13094;
	wire [4-1:0] node13097;
	wire [4-1:0] node13098;
	wire [4-1:0] node13099;
	wire [4-1:0] node13100;
	wire [4-1:0] node13104;
	wire [4-1:0] node13105;
	wire [4-1:0] node13108;
	wire [4-1:0] node13111;
	wire [4-1:0] node13112;
	wire [4-1:0] node13113;
	wire [4-1:0] node13116;
	wire [4-1:0] node13119;
	wire [4-1:0] node13120;
	wire [4-1:0] node13123;
	wire [4-1:0] node13126;
	wire [4-1:0] node13127;
	wire [4-1:0] node13128;
	wire [4-1:0] node13129;
	wire [4-1:0] node13130;
	wire [4-1:0] node13133;
	wire [4-1:0] node13136;
	wire [4-1:0] node13137;
	wire [4-1:0] node13140;
	wire [4-1:0] node13143;
	wire [4-1:0] node13144;
	wire [4-1:0] node13145;
	wire [4-1:0] node13148;
	wire [4-1:0] node13151;
	wire [4-1:0] node13152;
	wire [4-1:0] node13155;
	wire [4-1:0] node13158;
	wire [4-1:0] node13159;
	wire [4-1:0] node13160;
	wire [4-1:0] node13161;
	wire [4-1:0] node13164;
	wire [4-1:0] node13167;
	wire [4-1:0] node13168;
	wire [4-1:0] node13171;
	wire [4-1:0] node13174;
	wire [4-1:0] node13175;
	wire [4-1:0] node13177;
	wire [4-1:0] node13180;
	wire [4-1:0] node13181;
	wire [4-1:0] node13185;
	wire [4-1:0] node13186;
	wire [4-1:0] node13187;
	wire [4-1:0] node13188;
	wire [4-1:0] node13189;
	wire [4-1:0] node13191;
	wire [4-1:0] node13194;
	wire [4-1:0] node13195;
	wire [4-1:0] node13198;
	wire [4-1:0] node13201;
	wire [4-1:0] node13202;
	wire [4-1:0] node13204;
	wire [4-1:0] node13207;
	wire [4-1:0] node13208;
	wire [4-1:0] node13211;
	wire [4-1:0] node13214;
	wire [4-1:0] node13215;
	wire [4-1:0] node13216;
	wire [4-1:0] node13217;
	wire [4-1:0] node13221;
	wire [4-1:0] node13222;
	wire [4-1:0] node13225;
	wire [4-1:0] node13228;
	wire [4-1:0] node13229;
	wire [4-1:0] node13230;
	wire [4-1:0] node13233;
	wire [4-1:0] node13236;
	wire [4-1:0] node13237;
	wire [4-1:0] node13240;
	wire [4-1:0] node13243;
	wire [4-1:0] node13244;
	wire [4-1:0] node13245;
	wire [4-1:0] node13246;
	wire [4-1:0] node13247;
	wire [4-1:0] node13250;
	wire [4-1:0] node13253;
	wire [4-1:0] node13254;
	wire [4-1:0] node13257;
	wire [4-1:0] node13260;
	wire [4-1:0] node13261;
	wire [4-1:0] node13262;
	wire [4-1:0] node13265;
	wire [4-1:0] node13268;
	wire [4-1:0] node13269;
	wire [4-1:0] node13272;
	wire [4-1:0] node13275;
	wire [4-1:0] node13276;
	wire [4-1:0] node13277;
	wire [4-1:0] node13278;
	wire [4-1:0] node13281;
	wire [4-1:0] node13284;
	wire [4-1:0] node13286;
	wire [4-1:0] node13289;
	wire [4-1:0] node13290;
	wire [4-1:0] node13291;
	wire [4-1:0] node13294;
	wire [4-1:0] node13297;
	wire [4-1:0] node13300;
	wire [4-1:0] node13301;
	wire [4-1:0] node13302;
	wire [4-1:0] node13303;
	wire [4-1:0] node13304;
	wire [4-1:0] node13305;
	wire [4-1:0] node13306;
	wire [4-1:0] node13307;
	wire [4-1:0] node13308;
	wire [4-1:0] node13311;
	wire [4-1:0] node13314;
	wire [4-1:0] node13315;
	wire [4-1:0] node13318;
	wire [4-1:0] node13321;
	wire [4-1:0] node13322;
	wire [4-1:0] node13323;
	wire [4-1:0] node13326;
	wire [4-1:0] node13329;
	wire [4-1:0] node13330;
	wire [4-1:0] node13333;
	wire [4-1:0] node13336;
	wire [4-1:0] node13337;
	wire [4-1:0] node13338;
	wire [4-1:0] node13339;
	wire [4-1:0] node13342;
	wire [4-1:0] node13345;
	wire [4-1:0] node13346;
	wire [4-1:0] node13349;
	wire [4-1:0] node13352;
	wire [4-1:0] node13353;
	wire [4-1:0] node13354;
	wire [4-1:0] node13357;
	wire [4-1:0] node13360;
	wire [4-1:0] node13362;
	wire [4-1:0] node13365;
	wire [4-1:0] node13366;
	wire [4-1:0] node13367;
	wire [4-1:0] node13368;
	wire [4-1:0] node13369;
	wire [4-1:0] node13372;
	wire [4-1:0] node13375;
	wire [4-1:0] node13376;
	wire [4-1:0] node13379;
	wire [4-1:0] node13382;
	wire [4-1:0] node13383;
	wire [4-1:0] node13384;
	wire [4-1:0] node13387;
	wire [4-1:0] node13390;
	wire [4-1:0] node13391;
	wire [4-1:0] node13394;
	wire [4-1:0] node13397;
	wire [4-1:0] node13398;
	wire [4-1:0] node13399;
	wire [4-1:0] node13400;
	wire [4-1:0] node13403;
	wire [4-1:0] node13406;
	wire [4-1:0] node13407;
	wire [4-1:0] node13410;
	wire [4-1:0] node13413;
	wire [4-1:0] node13414;
	wire [4-1:0] node13415;
	wire [4-1:0] node13418;
	wire [4-1:0] node13421;
	wire [4-1:0] node13422;
	wire [4-1:0] node13425;
	wire [4-1:0] node13428;
	wire [4-1:0] node13429;
	wire [4-1:0] node13430;
	wire [4-1:0] node13431;
	wire [4-1:0] node13432;
	wire [4-1:0] node13434;
	wire [4-1:0] node13437;
	wire [4-1:0] node13438;
	wire [4-1:0] node13441;
	wire [4-1:0] node13444;
	wire [4-1:0] node13445;
	wire [4-1:0] node13446;
	wire [4-1:0] node13449;
	wire [4-1:0] node13452;
	wire [4-1:0] node13453;
	wire [4-1:0] node13456;
	wire [4-1:0] node13459;
	wire [4-1:0] node13460;
	wire [4-1:0] node13461;
	wire [4-1:0] node13462;
	wire [4-1:0] node13465;
	wire [4-1:0] node13468;
	wire [4-1:0] node13469;
	wire [4-1:0] node13472;
	wire [4-1:0] node13475;
	wire [4-1:0] node13476;
	wire [4-1:0] node13477;
	wire [4-1:0] node13480;
	wire [4-1:0] node13483;
	wire [4-1:0] node13485;
	wire [4-1:0] node13488;
	wire [4-1:0] node13489;
	wire [4-1:0] node13490;
	wire [4-1:0] node13491;
	wire [4-1:0] node13492;
	wire [4-1:0] node13495;
	wire [4-1:0] node13498;
	wire [4-1:0] node13499;
	wire [4-1:0] node13502;
	wire [4-1:0] node13505;
	wire [4-1:0] node13506;
	wire [4-1:0] node13507;
	wire [4-1:0] node13510;
	wire [4-1:0] node13513;
	wire [4-1:0] node13514;
	wire [4-1:0] node13517;
	wire [4-1:0] node13520;
	wire [4-1:0] node13521;
	wire [4-1:0] node13522;
	wire [4-1:0] node13523;
	wire [4-1:0] node13526;
	wire [4-1:0] node13529;
	wire [4-1:0] node13530;
	wire [4-1:0] node13533;
	wire [4-1:0] node13536;
	wire [4-1:0] node13537;
	wire [4-1:0] node13539;
	wire [4-1:0] node13542;
	wire [4-1:0] node13543;
	wire [4-1:0] node13546;
	wire [4-1:0] node13549;
	wire [4-1:0] node13550;
	wire [4-1:0] node13551;
	wire [4-1:0] node13552;
	wire [4-1:0] node13553;
	wire [4-1:0] node13554;
	wire [4-1:0] node13555;
	wire [4-1:0] node13559;
	wire [4-1:0] node13560;
	wire [4-1:0] node13564;
	wire [4-1:0] node13565;
	wire [4-1:0] node13566;
	wire [4-1:0] node13569;
	wire [4-1:0] node13572;
	wire [4-1:0] node13573;
	wire [4-1:0] node13576;
	wire [4-1:0] node13579;
	wire [4-1:0] node13580;
	wire [4-1:0] node13581;
	wire [4-1:0] node13582;
	wire [4-1:0] node13585;
	wire [4-1:0] node13588;
	wire [4-1:0] node13589;
	wire [4-1:0] node13592;
	wire [4-1:0] node13595;
	wire [4-1:0] node13596;
	wire [4-1:0] node13597;
	wire [4-1:0] node13600;
	wire [4-1:0] node13603;
	wire [4-1:0] node13604;
	wire [4-1:0] node13607;
	wire [4-1:0] node13610;
	wire [4-1:0] node13611;
	wire [4-1:0] node13612;
	wire [4-1:0] node13613;
	wire [4-1:0] node13614;
	wire [4-1:0] node13617;
	wire [4-1:0] node13620;
	wire [4-1:0] node13621;
	wire [4-1:0] node13624;
	wire [4-1:0] node13627;
	wire [4-1:0] node13628;
	wire [4-1:0] node13629;
	wire [4-1:0] node13632;
	wire [4-1:0] node13635;
	wire [4-1:0] node13636;
	wire [4-1:0] node13639;
	wire [4-1:0] node13642;
	wire [4-1:0] node13643;
	wire [4-1:0] node13644;
	wire [4-1:0] node13645;
	wire [4-1:0] node13648;
	wire [4-1:0] node13651;
	wire [4-1:0] node13652;
	wire [4-1:0] node13655;
	wire [4-1:0] node13658;
	wire [4-1:0] node13659;
	wire [4-1:0] node13660;
	wire [4-1:0] node13663;
	wire [4-1:0] node13666;
	wire [4-1:0] node13667;
	wire [4-1:0] node13670;
	wire [4-1:0] node13673;
	wire [4-1:0] node13674;
	wire [4-1:0] node13675;
	wire [4-1:0] node13676;
	wire [4-1:0] node13677;
	wire [4-1:0] node13678;
	wire [4-1:0] node13681;
	wire [4-1:0] node13684;
	wire [4-1:0] node13685;
	wire [4-1:0] node13688;
	wire [4-1:0] node13691;
	wire [4-1:0] node13692;
	wire [4-1:0] node13693;
	wire [4-1:0] node13696;
	wire [4-1:0] node13699;
	wire [4-1:0] node13700;
	wire [4-1:0] node13703;
	wire [4-1:0] node13706;
	wire [4-1:0] node13707;
	wire [4-1:0] node13708;
	wire [4-1:0] node13709;
	wire [4-1:0] node13712;
	wire [4-1:0] node13715;
	wire [4-1:0] node13716;
	wire [4-1:0] node13719;
	wire [4-1:0] node13722;
	wire [4-1:0] node13723;
	wire [4-1:0] node13726;
	wire [4-1:0] node13729;
	wire [4-1:0] node13730;
	wire [4-1:0] node13731;
	wire [4-1:0] node13732;
	wire [4-1:0] node13733;
	wire [4-1:0] node13736;
	wire [4-1:0] node13739;
	wire [4-1:0] node13740;
	wire [4-1:0] node13743;
	wire [4-1:0] node13746;
	wire [4-1:0] node13747;
	wire [4-1:0] node13750;
	wire [4-1:0] node13753;
	wire [4-1:0] node13754;
	wire [4-1:0] node13755;
	wire [4-1:0] node13756;
	wire [4-1:0] node13759;
	wire [4-1:0] node13762;
	wire [4-1:0] node13763;
	wire [4-1:0] node13766;
	wire [4-1:0] node13769;
	wire [4-1:0] node13770;
	wire [4-1:0] node13771;
	wire [4-1:0] node13774;
	wire [4-1:0] node13777;
	wire [4-1:0] node13778;
	wire [4-1:0] node13781;
	wire [4-1:0] node13784;
	wire [4-1:0] node13785;
	wire [4-1:0] node13786;
	wire [4-1:0] node13787;
	wire [4-1:0] node13788;
	wire [4-1:0] node13789;
	wire [4-1:0] node13790;
	wire [4-1:0] node13791;
	wire [4-1:0] node13794;
	wire [4-1:0] node13797;
	wire [4-1:0] node13798;
	wire [4-1:0] node13801;
	wire [4-1:0] node13804;
	wire [4-1:0] node13805;
	wire [4-1:0] node13807;
	wire [4-1:0] node13810;
	wire [4-1:0] node13811;
	wire [4-1:0] node13815;
	wire [4-1:0] node13816;
	wire [4-1:0] node13817;
	wire [4-1:0] node13818;
	wire [4-1:0] node13821;
	wire [4-1:0] node13824;
	wire [4-1:0] node13825;
	wire [4-1:0] node13828;
	wire [4-1:0] node13831;
	wire [4-1:0] node13832;
	wire [4-1:0] node13833;
	wire [4-1:0] node13836;
	wire [4-1:0] node13839;
	wire [4-1:0] node13840;
	wire [4-1:0] node13844;
	wire [4-1:0] node13845;
	wire [4-1:0] node13846;
	wire [4-1:0] node13847;
	wire [4-1:0] node13848;
	wire [4-1:0] node13851;
	wire [4-1:0] node13854;
	wire [4-1:0] node13855;
	wire [4-1:0] node13858;
	wire [4-1:0] node13861;
	wire [4-1:0] node13862;
	wire [4-1:0] node13864;
	wire [4-1:0] node13867;
	wire [4-1:0] node13868;
	wire [4-1:0] node13871;
	wire [4-1:0] node13874;
	wire [4-1:0] node13875;
	wire [4-1:0] node13876;
	wire [4-1:0] node13877;
	wire [4-1:0] node13880;
	wire [4-1:0] node13883;
	wire [4-1:0] node13884;
	wire [4-1:0] node13887;
	wire [4-1:0] node13890;
	wire [4-1:0] node13891;
	wire [4-1:0] node13893;
	wire [4-1:0] node13896;
	wire [4-1:0] node13897;
	wire [4-1:0] node13901;
	wire [4-1:0] node13902;
	wire [4-1:0] node13903;
	wire [4-1:0] node13904;
	wire [4-1:0] node13905;
	wire [4-1:0] node13906;
	wire [4-1:0] node13909;
	wire [4-1:0] node13912;
	wire [4-1:0] node13914;
	wire [4-1:0] node13917;
	wire [4-1:0] node13918;
	wire [4-1:0] node13919;
	wire [4-1:0] node13923;
	wire [4-1:0] node13924;
	wire [4-1:0] node13927;
	wire [4-1:0] node13930;
	wire [4-1:0] node13931;
	wire [4-1:0] node13932;
	wire [4-1:0] node13933;
	wire [4-1:0] node13936;
	wire [4-1:0] node13939;
	wire [4-1:0] node13941;
	wire [4-1:0] node13944;
	wire [4-1:0] node13945;
	wire [4-1:0] node13946;
	wire [4-1:0] node13949;
	wire [4-1:0] node13952;
	wire [4-1:0] node13953;
	wire [4-1:0] node13956;
	wire [4-1:0] node13959;
	wire [4-1:0] node13960;
	wire [4-1:0] node13961;
	wire [4-1:0] node13962;
	wire [4-1:0] node13963;
	wire [4-1:0] node13966;
	wire [4-1:0] node13969;
	wire [4-1:0] node13970;
	wire [4-1:0] node13973;
	wire [4-1:0] node13976;
	wire [4-1:0] node13977;
	wire [4-1:0] node13978;
	wire [4-1:0] node13981;
	wire [4-1:0] node13984;
	wire [4-1:0] node13985;
	wire [4-1:0] node13988;
	wire [4-1:0] node13991;
	wire [4-1:0] node13992;
	wire [4-1:0] node13993;
	wire [4-1:0] node13994;
	wire [4-1:0] node13997;
	wire [4-1:0] node14000;
	wire [4-1:0] node14001;
	wire [4-1:0] node14004;
	wire [4-1:0] node14007;
	wire [4-1:0] node14008;
	wire [4-1:0] node14009;
	wire [4-1:0] node14012;
	wire [4-1:0] node14015;
	wire [4-1:0] node14016;
	wire [4-1:0] node14019;
	wire [4-1:0] node14022;
	wire [4-1:0] node14023;
	wire [4-1:0] node14024;
	wire [4-1:0] node14025;
	wire [4-1:0] node14026;
	wire [4-1:0] node14027;
	wire [4-1:0] node14029;
	wire [4-1:0] node14032;
	wire [4-1:0] node14033;
	wire [4-1:0] node14036;
	wire [4-1:0] node14039;
	wire [4-1:0] node14040;
	wire [4-1:0] node14041;
	wire [4-1:0] node14044;
	wire [4-1:0] node14047;
	wire [4-1:0] node14048;
	wire [4-1:0] node14052;
	wire [4-1:0] node14053;
	wire [4-1:0] node14054;
	wire [4-1:0] node14055;
	wire [4-1:0] node14058;
	wire [4-1:0] node14061;
	wire [4-1:0] node14062;
	wire [4-1:0] node14065;
	wire [4-1:0] node14068;
	wire [4-1:0] node14069;
	wire [4-1:0] node14070;
	wire [4-1:0] node14073;
	wire [4-1:0] node14076;
	wire [4-1:0] node14077;
	wire [4-1:0] node14080;
	wire [4-1:0] node14083;
	wire [4-1:0] node14084;
	wire [4-1:0] node14085;
	wire [4-1:0] node14086;
	wire [4-1:0] node14087;
	wire [4-1:0] node14090;
	wire [4-1:0] node14093;
	wire [4-1:0] node14094;
	wire [4-1:0] node14097;
	wire [4-1:0] node14100;
	wire [4-1:0] node14101;
	wire [4-1:0] node14103;
	wire [4-1:0] node14106;
	wire [4-1:0] node14107;
	wire [4-1:0] node14111;
	wire [4-1:0] node14112;
	wire [4-1:0] node14113;
	wire [4-1:0] node14114;
	wire [4-1:0] node14117;
	wire [4-1:0] node14120;
	wire [4-1:0] node14121;
	wire [4-1:0] node14124;
	wire [4-1:0] node14127;
	wire [4-1:0] node14128;
	wire [4-1:0] node14129;
	wire [4-1:0] node14132;
	wire [4-1:0] node14135;
	wire [4-1:0] node14136;
	wire [4-1:0] node14139;
	wire [4-1:0] node14142;
	wire [4-1:0] node14143;
	wire [4-1:0] node14144;
	wire [4-1:0] node14145;
	wire [4-1:0] node14146;
	wire [4-1:0] node14147;
	wire [4-1:0] node14150;
	wire [4-1:0] node14153;
	wire [4-1:0] node14154;
	wire [4-1:0] node14158;
	wire [4-1:0] node14159;
	wire [4-1:0] node14160;
	wire [4-1:0] node14163;
	wire [4-1:0] node14166;
	wire [4-1:0] node14167;
	wire [4-1:0] node14170;
	wire [4-1:0] node14173;
	wire [4-1:0] node14174;
	wire [4-1:0] node14175;
	wire [4-1:0] node14176;
	wire [4-1:0] node14179;
	wire [4-1:0] node14182;
	wire [4-1:0] node14183;
	wire [4-1:0] node14186;
	wire [4-1:0] node14189;
	wire [4-1:0] node14190;
	wire [4-1:0] node14191;
	wire [4-1:0] node14194;
	wire [4-1:0] node14197;
	wire [4-1:0] node14198;
	wire [4-1:0] node14201;
	wire [4-1:0] node14204;
	wire [4-1:0] node14205;
	wire [4-1:0] node14206;
	wire [4-1:0] node14207;
	wire [4-1:0] node14208;
	wire [4-1:0] node14211;
	wire [4-1:0] node14214;
	wire [4-1:0] node14215;
	wire [4-1:0] node14218;
	wire [4-1:0] node14221;
	wire [4-1:0] node14222;
	wire [4-1:0] node14223;
	wire [4-1:0] node14226;
	wire [4-1:0] node14229;
	wire [4-1:0] node14230;
	wire [4-1:0] node14233;
	wire [4-1:0] node14236;
	wire [4-1:0] node14237;
	wire [4-1:0] node14238;
	wire [4-1:0] node14241;
	wire [4-1:0] node14244;
	wire [4-1:0] node14245;
	wire [4-1:0] node14246;
	wire [4-1:0] node14249;
	wire [4-1:0] node14252;
	wire [4-1:0] node14253;
	wire [4-1:0] node14256;
	wire [4-1:0] node14259;
	wire [4-1:0] node14260;
	wire [4-1:0] node14261;
	wire [4-1:0] node14262;
	wire [4-1:0] node14263;
	wire [4-1:0] node14264;
	wire [4-1:0] node14265;
	wire [4-1:0] node14266;
	wire [4-1:0] node14267;
	wire [4-1:0] node14268;
	wire [4-1:0] node14269;
	wire [4-1:0] node14270;
	wire [4-1:0] node14271;
	wire [4-1:0] node14274;
	wire [4-1:0] node14277;
	wire [4-1:0] node14278;
	wire [4-1:0] node14281;
	wire [4-1:0] node14284;
	wire [4-1:0] node14285;
	wire [4-1:0] node14286;
	wire [4-1:0] node14289;
	wire [4-1:0] node14292;
	wire [4-1:0] node14293;
	wire [4-1:0] node14296;
	wire [4-1:0] node14299;
	wire [4-1:0] node14300;
	wire [4-1:0] node14301;
	wire [4-1:0] node14302;
	wire [4-1:0] node14305;
	wire [4-1:0] node14308;
	wire [4-1:0] node14309;
	wire [4-1:0] node14312;
	wire [4-1:0] node14315;
	wire [4-1:0] node14316;
	wire [4-1:0] node14317;
	wire [4-1:0] node14320;
	wire [4-1:0] node14323;
	wire [4-1:0] node14324;
	wire [4-1:0] node14327;
	wire [4-1:0] node14330;
	wire [4-1:0] node14331;
	wire [4-1:0] node14332;
	wire [4-1:0] node14333;
	wire [4-1:0] node14334;
	wire [4-1:0] node14337;
	wire [4-1:0] node14340;
	wire [4-1:0] node14341;
	wire [4-1:0] node14344;
	wire [4-1:0] node14347;
	wire [4-1:0] node14348;
	wire [4-1:0] node14349;
	wire [4-1:0] node14352;
	wire [4-1:0] node14355;
	wire [4-1:0] node14356;
	wire [4-1:0] node14359;
	wire [4-1:0] node14362;
	wire [4-1:0] node14363;
	wire [4-1:0] node14364;
	wire [4-1:0] node14365;
	wire [4-1:0] node14368;
	wire [4-1:0] node14371;
	wire [4-1:0] node14372;
	wire [4-1:0] node14375;
	wire [4-1:0] node14378;
	wire [4-1:0] node14379;
	wire [4-1:0] node14380;
	wire [4-1:0] node14383;
	wire [4-1:0] node14386;
	wire [4-1:0] node14387;
	wire [4-1:0] node14390;
	wire [4-1:0] node14393;
	wire [4-1:0] node14394;
	wire [4-1:0] node14395;
	wire [4-1:0] node14396;
	wire [4-1:0] node14397;
	wire [4-1:0] node14398;
	wire [4-1:0] node14401;
	wire [4-1:0] node14404;
	wire [4-1:0] node14405;
	wire [4-1:0] node14408;
	wire [4-1:0] node14411;
	wire [4-1:0] node14412;
	wire [4-1:0] node14413;
	wire [4-1:0] node14416;
	wire [4-1:0] node14419;
	wire [4-1:0] node14420;
	wire [4-1:0] node14423;
	wire [4-1:0] node14426;
	wire [4-1:0] node14427;
	wire [4-1:0] node14428;
	wire [4-1:0] node14429;
	wire [4-1:0] node14433;
	wire [4-1:0] node14434;
	wire [4-1:0] node14437;
	wire [4-1:0] node14440;
	wire [4-1:0] node14441;
	wire [4-1:0] node14442;
	wire [4-1:0] node14445;
	wire [4-1:0] node14448;
	wire [4-1:0] node14450;
	wire [4-1:0] node14453;
	wire [4-1:0] node14454;
	wire [4-1:0] node14455;
	wire [4-1:0] node14456;
	wire [4-1:0] node14457;
	wire [4-1:0] node14460;
	wire [4-1:0] node14463;
	wire [4-1:0] node14464;
	wire [4-1:0] node14467;
	wire [4-1:0] node14470;
	wire [4-1:0] node14471;
	wire [4-1:0] node14472;
	wire [4-1:0] node14475;
	wire [4-1:0] node14478;
	wire [4-1:0] node14479;
	wire [4-1:0] node14482;
	wire [4-1:0] node14485;
	wire [4-1:0] node14486;
	wire [4-1:0] node14487;
	wire [4-1:0] node14488;
	wire [4-1:0] node14491;
	wire [4-1:0] node14494;
	wire [4-1:0] node14495;
	wire [4-1:0] node14498;
	wire [4-1:0] node14501;
	wire [4-1:0] node14502;
	wire [4-1:0] node14503;
	wire [4-1:0] node14507;
	wire [4-1:0] node14508;
	wire [4-1:0] node14511;
	wire [4-1:0] node14514;
	wire [4-1:0] node14515;
	wire [4-1:0] node14516;
	wire [4-1:0] node14517;
	wire [4-1:0] node14518;
	wire [4-1:0] node14519;
	wire [4-1:0] node14520;
	wire [4-1:0] node14523;
	wire [4-1:0] node14526;
	wire [4-1:0] node14527;
	wire [4-1:0] node14530;
	wire [4-1:0] node14533;
	wire [4-1:0] node14534;
	wire [4-1:0] node14535;
	wire [4-1:0] node14539;
	wire [4-1:0] node14540;
	wire [4-1:0] node14543;
	wire [4-1:0] node14546;
	wire [4-1:0] node14547;
	wire [4-1:0] node14548;
	wire [4-1:0] node14550;
	wire [4-1:0] node14553;
	wire [4-1:0] node14555;
	wire [4-1:0] node14558;
	wire [4-1:0] node14559;
	wire [4-1:0] node14561;
	wire [4-1:0] node14564;
	wire [4-1:0] node14566;
	wire [4-1:0] node14569;
	wire [4-1:0] node14570;
	wire [4-1:0] node14571;
	wire [4-1:0] node14572;
	wire [4-1:0] node14574;
	wire [4-1:0] node14577;
	wire [4-1:0] node14578;
	wire [4-1:0] node14581;
	wire [4-1:0] node14584;
	wire [4-1:0] node14585;
	wire [4-1:0] node14586;
	wire [4-1:0] node14589;
	wire [4-1:0] node14592;
	wire [4-1:0] node14593;
	wire [4-1:0] node14597;
	wire [4-1:0] node14598;
	wire [4-1:0] node14599;
	wire [4-1:0] node14601;
	wire [4-1:0] node14604;
	wire [4-1:0] node14606;
	wire [4-1:0] node14609;
	wire [4-1:0] node14610;
	wire [4-1:0] node14612;
	wire [4-1:0] node14615;
	wire [4-1:0] node14617;
	wire [4-1:0] node14620;
	wire [4-1:0] node14621;
	wire [4-1:0] node14622;
	wire [4-1:0] node14623;
	wire [4-1:0] node14624;
	wire [4-1:0] node14625;
	wire [4-1:0] node14628;
	wire [4-1:0] node14631;
	wire [4-1:0] node14632;
	wire [4-1:0] node14635;
	wire [4-1:0] node14638;
	wire [4-1:0] node14639;
	wire [4-1:0] node14640;
	wire [4-1:0] node14643;
	wire [4-1:0] node14646;
	wire [4-1:0] node14647;
	wire [4-1:0] node14650;
	wire [4-1:0] node14653;
	wire [4-1:0] node14654;
	wire [4-1:0] node14655;
	wire [4-1:0] node14658;
	wire [4-1:0] node14661;
	wire [4-1:0] node14662;
	wire [4-1:0] node14663;
	wire [4-1:0] node14666;
	wire [4-1:0] node14669;
	wire [4-1:0] node14670;
	wire [4-1:0] node14673;
	wire [4-1:0] node14676;
	wire [4-1:0] node14677;
	wire [4-1:0] node14678;
	wire [4-1:0] node14679;
	wire [4-1:0] node14680;
	wire [4-1:0] node14683;
	wire [4-1:0] node14686;
	wire [4-1:0] node14687;
	wire [4-1:0] node14690;
	wire [4-1:0] node14693;
	wire [4-1:0] node14694;
	wire [4-1:0] node14695;
	wire [4-1:0] node14698;
	wire [4-1:0] node14701;
	wire [4-1:0] node14703;
	wire [4-1:0] node14706;
	wire [4-1:0] node14707;
	wire [4-1:0] node14708;
	wire [4-1:0] node14710;
	wire [4-1:0] node14713;
	wire [4-1:0] node14715;
	wire [4-1:0] node14718;
	wire [4-1:0] node14719;
	wire [4-1:0] node14721;
	wire [4-1:0] node14724;
	wire [4-1:0] node14726;
	wire [4-1:0] node14729;
	wire [4-1:0] node14730;
	wire [4-1:0] node14731;
	wire [4-1:0] node14732;
	wire [4-1:0] node14733;
	wire [4-1:0] node14734;
	wire [4-1:0] node14735;
	wire [4-1:0] node14737;
	wire [4-1:0] node14740;
	wire [4-1:0] node14741;
	wire [4-1:0] node14744;
	wire [4-1:0] node14747;
	wire [4-1:0] node14748;
	wire [4-1:0] node14749;
	wire [4-1:0] node14753;
	wire [4-1:0] node14754;
	wire [4-1:0] node14757;
	wire [4-1:0] node14760;
	wire [4-1:0] node14761;
	wire [4-1:0] node14762;
	wire [4-1:0] node14763;
	wire [4-1:0] node14766;
	wire [4-1:0] node14769;
	wire [4-1:0] node14770;
	wire [4-1:0] node14773;
	wire [4-1:0] node14776;
	wire [4-1:0] node14777;
	wire [4-1:0] node14778;
	wire [4-1:0] node14781;
	wire [4-1:0] node14784;
	wire [4-1:0] node14785;
	wire [4-1:0] node14788;
	wire [4-1:0] node14791;
	wire [4-1:0] node14792;
	wire [4-1:0] node14793;
	wire [4-1:0] node14794;
	wire [4-1:0] node14796;
	wire [4-1:0] node14799;
	wire [4-1:0] node14800;
	wire [4-1:0] node14803;
	wire [4-1:0] node14806;
	wire [4-1:0] node14807;
	wire [4-1:0] node14808;
	wire [4-1:0] node14811;
	wire [4-1:0] node14814;
	wire [4-1:0] node14816;
	wire [4-1:0] node14819;
	wire [4-1:0] node14820;
	wire [4-1:0] node14821;
	wire [4-1:0] node14822;
	wire [4-1:0] node14826;
	wire [4-1:0] node14827;
	wire [4-1:0] node14831;
	wire [4-1:0] node14832;
	wire [4-1:0] node14833;
	wire [4-1:0] node14836;
	wire [4-1:0] node14839;
	wire [4-1:0] node14841;
	wire [4-1:0] node14844;
	wire [4-1:0] node14845;
	wire [4-1:0] node14846;
	wire [4-1:0] node14847;
	wire [4-1:0] node14848;
	wire [4-1:0] node14850;
	wire [4-1:0] node14853;
	wire [4-1:0] node14854;
	wire [4-1:0] node14857;
	wire [4-1:0] node14860;
	wire [4-1:0] node14861;
	wire [4-1:0] node14862;
	wire [4-1:0] node14865;
	wire [4-1:0] node14868;
	wire [4-1:0] node14870;
	wire [4-1:0] node14873;
	wire [4-1:0] node14874;
	wire [4-1:0] node14875;
	wire [4-1:0] node14877;
	wire [4-1:0] node14880;
	wire [4-1:0] node14882;
	wire [4-1:0] node14885;
	wire [4-1:0] node14886;
	wire [4-1:0] node14888;
	wire [4-1:0] node14891;
	wire [4-1:0] node14893;
	wire [4-1:0] node14896;
	wire [4-1:0] node14897;
	wire [4-1:0] node14898;
	wire [4-1:0] node14899;
	wire [4-1:0] node14900;
	wire [4-1:0] node14903;
	wire [4-1:0] node14906;
	wire [4-1:0] node14907;
	wire [4-1:0] node14910;
	wire [4-1:0] node14913;
	wire [4-1:0] node14914;
	wire [4-1:0] node14915;
	wire [4-1:0] node14918;
	wire [4-1:0] node14921;
	wire [4-1:0] node14922;
	wire [4-1:0] node14925;
	wire [4-1:0] node14928;
	wire [4-1:0] node14929;
	wire [4-1:0] node14930;
	wire [4-1:0] node14932;
	wire [4-1:0] node14935;
	wire [4-1:0] node14937;
	wire [4-1:0] node14940;
	wire [4-1:0] node14941;
	wire [4-1:0] node14943;
	wire [4-1:0] node14946;
	wire [4-1:0] node14948;
	wire [4-1:0] node14951;
	wire [4-1:0] node14952;
	wire [4-1:0] node14953;
	wire [4-1:0] node14954;
	wire [4-1:0] node14955;
	wire [4-1:0] node14956;
	wire [4-1:0] node14957;
	wire [4-1:0] node14960;
	wire [4-1:0] node14963;
	wire [4-1:0] node14964;
	wire [4-1:0] node14967;
	wire [4-1:0] node14970;
	wire [4-1:0] node14971;
	wire [4-1:0] node14972;
	wire [4-1:0] node14975;
	wire [4-1:0] node14978;
	wire [4-1:0] node14979;
	wire [4-1:0] node14982;
	wire [4-1:0] node14985;
	wire [4-1:0] node14986;
	wire [4-1:0] node14987;
	wire [4-1:0] node14988;
	wire [4-1:0] node14991;
	wire [4-1:0] node14994;
	wire [4-1:0] node14995;
	wire [4-1:0] node14998;
	wire [4-1:0] node15001;
	wire [4-1:0] node15002;
	wire [4-1:0] node15003;
	wire [4-1:0] node15006;
	wire [4-1:0] node15009;
	wire [4-1:0] node15010;
	wire [4-1:0] node15013;
	wire [4-1:0] node15016;
	wire [4-1:0] node15017;
	wire [4-1:0] node15018;
	wire [4-1:0] node15019;
	wire [4-1:0] node15020;
	wire [4-1:0] node15024;
	wire [4-1:0] node15025;
	wire [4-1:0] node15029;
	wire [4-1:0] node15030;
	wire [4-1:0] node15031;
	wire [4-1:0] node15035;
	wire [4-1:0] node15036;
	wire [4-1:0] node15040;
	wire [4-1:0] node15041;
	wire [4-1:0] node15042;
	wire [4-1:0] node15043;
	wire [4-1:0] node15046;
	wire [4-1:0] node15049;
	wire [4-1:0] node15050;
	wire [4-1:0] node15053;
	wire [4-1:0] node15056;
	wire [4-1:0] node15057;
	wire [4-1:0] node15058;
	wire [4-1:0] node15061;
	wire [4-1:0] node15064;
	wire [4-1:0] node15066;
	wire [4-1:0] node15069;
	wire [4-1:0] node15070;
	wire [4-1:0] node15071;
	wire [4-1:0] node15072;
	wire [4-1:0] node15073;
	wire [4-1:0] node15074;
	wire [4-1:0] node15078;
	wire [4-1:0] node15079;
	wire [4-1:0] node15082;
	wire [4-1:0] node15085;
	wire [4-1:0] node15086;
	wire [4-1:0] node15087;
	wire [4-1:0] node15090;
	wire [4-1:0] node15093;
	wire [4-1:0] node15094;
	wire [4-1:0] node15097;
	wire [4-1:0] node15100;
	wire [4-1:0] node15101;
	wire [4-1:0] node15102;
	wire [4-1:0] node15103;
	wire [4-1:0] node15106;
	wire [4-1:0] node15109;
	wire [4-1:0] node15110;
	wire [4-1:0] node15113;
	wire [4-1:0] node15116;
	wire [4-1:0] node15117;
	wire [4-1:0] node15119;
	wire [4-1:0] node15122;
	wire [4-1:0] node15123;
	wire [4-1:0] node15126;
	wire [4-1:0] node15129;
	wire [4-1:0] node15130;
	wire [4-1:0] node15131;
	wire [4-1:0] node15132;
	wire [4-1:0] node15133;
	wire [4-1:0] node15137;
	wire [4-1:0] node15138;
	wire [4-1:0] node15142;
	wire [4-1:0] node15143;
	wire [4-1:0] node15144;
	wire [4-1:0] node15148;
	wire [4-1:0] node15149;
	wire [4-1:0] node15153;
	wire [4-1:0] node15154;
	wire [4-1:0] node15155;
	wire [4-1:0] node15156;
	wire [4-1:0] node15159;
	wire [4-1:0] node15162;
	wire [4-1:0] node15163;
	wire [4-1:0] node15166;
	wire [4-1:0] node15169;
	wire [4-1:0] node15170;
	wire [4-1:0] node15171;
	wire [4-1:0] node15174;
	wire [4-1:0] node15177;
	wire [4-1:0] node15179;
	wire [4-1:0] node15182;
	wire [4-1:0] node15183;
	wire [4-1:0] node15184;
	wire [4-1:0] node15185;
	wire [4-1:0] node15186;
	wire [4-1:0] node15187;
	wire [4-1:0] node15188;
	wire [4-1:0] node15189;
	wire [4-1:0] node15190;
	wire [4-1:0] node15193;
	wire [4-1:0] node15196;
	wire [4-1:0] node15198;
	wire [4-1:0] node15201;
	wire [4-1:0] node15202;
	wire [4-1:0] node15203;
	wire [4-1:0] node15206;
	wire [4-1:0] node15209;
	wire [4-1:0] node15210;
	wire [4-1:0] node15214;
	wire [4-1:0] node15215;
	wire [4-1:0] node15216;
	wire [4-1:0] node15217;
	wire [4-1:0] node15221;
	wire [4-1:0] node15222;
	wire [4-1:0] node15225;
	wire [4-1:0] node15228;
	wire [4-1:0] node15229;
	wire [4-1:0] node15230;
	wire [4-1:0] node15233;
	wire [4-1:0] node15236;
	wire [4-1:0] node15237;
	wire [4-1:0] node15240;
	wire [4-1:0] node15243;
	wire [4-1:0] node15244;
	wire [4-1:0] node15245;
	wire [4-1:0] node15246;
	wire [4-1:0] node15247;
	wire [4-1:0] node15250;
	wire [4-1:0] node15253;
	wire [4-1:0] node15254;
	wire [4-1:0] node15257;
	wire [4-1:0] node15260;
	wire [4-1:0] node15261;
	wire [4-1:0] node15263;
	wire [4-1:0] node15266;
	wire [4-1:0] node15267;
	wire [4-1:0] node15270;
	wire [4-1:0] node15273;
	wire [4-1:0] node15274;
	wire [4-1:0] node15275;
	wire [4-1:0] node15276;
	wire [4-1:0] node15280;
	wire [4-1:0] node15281;
	wire [4-1:0] node15284;
	wire [4-1:0] node15287;
	wire [4-1:0] node15288;
	wire [4-1:0] node15289;
	wire [4-1:0] node15292;
	wire [4-1:0] node15295;
	wire [4-1:0] node15296;
	wire [4-1:0] node15299;
	wire [4-1:0] node15302;
	wire [4-1:0] node15303;
	wire [4-1:0] node15304;
	wire [4-1:0] node15305;
	wire [4-1:0] node15306;
	wire [4-1:0] node15307;
	wire [4-1:0] node15310;
	wire [4-1:0] node15313;
	wire [4-1:0] node15314;
	wire [4-1:0] node15317;
	wire [4-1:0] node15320;
	wire [4-1:0] node15321;
	wire [4-1:0] node15322;
	wire [4-1:0] node15325;
	wire [4-1:0] node15328;
	wire [4-1:0] node15329;
	wire [4-1:0] node15332;
	wire [4-1:0] node15335;
	wire [4-1:0] node15336;
	wire [4-1:0] node15337;
	wire [4-1:0] node15339;
	wire [4-1:0] node15342;
	wire [4-1:0] node15344;
	wire [4-1:0] node15347;
	wire [4-1:0] node15348;
	wire [4-1:0] node15350;
	wire [4-1:0] node15353;
	wire [4-1:0] node15355;
	wire [4-1:0] node15358;
	wire [4-1:0] node15359;
	wire [4-1:0] node15360;
	wire [4-1:0] node15361;
	wire [4-1:0] node15362;
	wire [4-1:0] node15365;
	wire [4-1:0] node15368;
	wire [4-1:0] node15369;
	wire [4-1:0] node15372;
	wire [4-1:0] node15375;
	wire [4-1:0] node15376;
	wire [4-1:0] node15378;
	wire [4-1:0] node15381;
	wire [4-1:0] node15382;
	wire [4-1:0] node15385;
	wire [4-1:0] node15388;
	wire [4-1:0] node15389;
	wire [4-1:0] node15390;
	wire [4-1:0] node15393;
	wire [4-1:0] node15395;
	wire [4-1:0] node15398;
	wire [4-1:0] node15399;
	wire [4-1:0] node15401;
	wire [4-1:0] node15404;
	wire [4-1:0] node15406;
	wire [4-1:0] node15409;
	wire [4-1:0] node15410;
	wire [4-1:0] node15411;
	wire [4-1:0] node15412;
	wire [4-1:0] node15413;
	wire [4-1:0] node15414;
	wire [4-1:0] node15415;
	wire [4-1:0] node15418;
	wire [4-1:0] node15421;
	wire [4-1:0] node15422;
	wire [4-1:0] node15425;
	wire [4-1:0] node15428;
	wire [4-1:0] node15429;
	wire [4-1:0] node15430;
	wire [4-1:0] node15434;
	wire [4-1:0] node15435;
	wire [4-1:0] node15438;
	wire [4-1:0] node15441;
	wire [4-1:0] node15442;
	wire [4-1:0] node15443;
	wire [4-1:0] node15446;
	wire [4-1:0] node15449;
	wire [4-1:0] node15450;
	wire [4-1:0] node15452;
	wire [4-1:0] node15455;
	wire [4-1:0] node15456;
	wire [4-1:0] node15459;
	wire [4-1:0] node15462;
	wire [4-1:0] node15463;
	wire [4-1:0] node15464;
	wire [4-1:0] node15465;
	wire [4-1:0] node15466;
	wire [4-1:0] node15469;
	wire [4-1:0] node15472;
	wire [4-1:0] node15473;
	wire [4-1:0] node15476;
	wire [4-1:0] node15479;
	wire [4-1:0] node15480;
	wire [4-1:0] node15481;
	wire [4-1:0] node15485;
	wire [4-1:0] node15486;
	wire [4-1:0] node15489;
	wire [4-1:0] node15492;
	wire [4-1:0] node15493;
	wire [4-1:0] node15494;
	wire [4-1:0] node15497;
	wire [4-1:0] node15500;
	wire [4-1:0] node15501;
	wire [4-1:0] node15502;
	wire [4-1:0] node15505;
	wire [4-1:0] node15508;
	wire [4-1:0] node15509;
	wire [4-1:0] node15512;
	wire [4-1:0] node15515;
	wire [4-1:0] node15516;
	wire [4-1:0] node15517;
	wire [4-1:0] node15518;
	wire [4-1:0] node15519;
	wire [4-1:0] node15520;
	wire [4-1:0] node15523;
	wire [4-1:0] node15526;
	wire [4-1:0] node15527;
	wire [4-1:0] node15530;
	wire [4-1:0] node15533;
	wire [4-1:0] node15534;
	wire [4-1:0] node15535;
	wire [4-1:0] node15539;
	wire [4-1:0] node15540;
	wire [4-1:0] node15543;
	wire [4-1:0] node15546;
	wire [4-1:0] node15547;
	wire [4-1:0] node15548;
	wire [4-1:0] node15549;
	wire [4-1:0] node15552;
	wire [4-1:0] node15555;
	wire [4-1:0] node15556;
	wire [4-1:0] node15559;
	wire [4-1:0] node15562;
	wire [4-1:0] node15563;
	wire [4-1:0] node15564;
	wire [4-1:0] node15567;
	wire [4-1:0] node15570;
	wire [4-1:0] node15571;
	wire [4-1:0] node15574;
	wire [4-1:0] node15577;
	wire [4-1:0] node15578;
	wire [4-1:0] node15579;
	wire [4-1:0] node15580;
	wire [4-1:0] node15581;
	wire [4-1:0] node15584;
	wire [4-1:0] node15587;
	wire [4-1:0] node15588;
	wire [4-1:0] node15591;
	wire [4-1:0] node15594;
	wire [4-1:0] node15595;
	wire [4-1:0] node15596;
	wire [4-1:0] node15599;
	wire [4-1:0] node15602;
	wire [4-1:0] node15603;
	wire [4-1:0] node15607;
	wire [4-1:0] node15608;
	wire [4-1:0] node15609;
	wire [4-1:0] node15611;
	wire [4-1:0] node15614;
	wire [4-1:0] node15616;
	wire [4-1:0] node15619;
	wire [4-1:0] node15620;
	wire [4-1:0] node15622;
	wire [4-1:0] node15625;
	wire [4-1:0] node15627;
	wire [4-1:0] node15630;
	wire [4-1:0] node15631;
	wire [4-1:0] node15632;
	wire [4-1:0] node15633;
	wire [4-1:0] node15634;
	wire [4-1:0] node15635;
	wire [4-1:0] node15636;
	wire [4-1:0] node15638;
	wire [4-1:0] node15641;
	wire [4-1:0] node15642;
	wire [4-1:0] node15645;
	wire [4-1:0] node15648;
	wire [4-1:0] node15649;
	wire [4-1:0] node15650;
	wire [4-1:0] node15654;
	wire [4-1:0] node15655;
	wire [4-1:0] node15659;
	wire [4-1:0] node15660;
	wire [4-1:0] node15661;
	wire [4-1:0] node15663;
	wire [4-1:0] node15666;
	wire [4-1:0] node15668;
	wire [4-1:0] node15671;
	wire [4-1:0] node15672;
	wire [4-1:0] node15674;
	wire [4-1:0] node15677;
	wire [4-1:0] node15679;
	wire [4-1:0] node15682;
	wire [4-1:0] node15683;
	wire [4-1:0] node15684;
	wire [4-1:0] node15685;
	wire [4-1:0] node15686;
	wire [4-1:0] node15689;
	wire [4-1:0] node15692;
	wire [4-1:0] node15693;
	wire [4-1:0] node15697;
	wire [4-1:0] node15698;
	wire [4-1:0] node15699;
	wire [4-1:0] node15703;
	wire [4-1:0] node15704;
	wire [4-1:0] node15707;
	wire [4-1:0] node15710;
	wire [4-1:0] node15711;
	wire [4-1:0] node15712;
	wire [4-1:0] node15714;
	wire [4-1:0] node15717;
	wire [4-1:0] node15719;
	wire [4-1:0] node15722;
	wire [4-1:0] node15723;
	wire [4-1:0] node15725;
	wire [4-1:0] node15728;
	wire [4-1:0] node15730;
	wire [4-1:0] node15733;
	wire [4-1:0] node15734;
	wire [4-1:0] node15735;
	wire [4-1:0] node15736;
	wire [4-1:0] node15737;
	wire [4-1:0] node15738;
	wire [4-1:0] node15741;
	wire [4-1:0] node15744;
	wire [4-1:0] node15745;
	wire [4-1:0] node15748;
	wire [4-1:0] node15751;
	wire [4-1:0] node15752;
	wire [4-1:0] node15754;
	wire [4-1:0] node15757;
	wire [4-1:0] node15758;
	wire [4-1:0] node15761;
	wire [4-1:0] node15764;
	wire [4-1:0] node15765;
	wire [4-1:0] node15766;
	wire [4-1:0] node15767;
	wire [4-1:0] node15770;
	wire [4-1:0] node15773;
	wire [4-1:0] node15774;
	wire [4-1:0] node15777;
	wire [4-1:0] node15780;
	wire [4-1:0] node15781;
	wire [4-1:0] node15782;
	wire [4-1:0] node15785;
	wire [4-1:0] node15788;
	wire [4-1:0] node15789;
	wire [4-1:0] node15792;
	wire [4-1:0] node15795;
	wire [4-1:0] node15796;
	wire [4-1:0] node15797;
	wire [4-1:0] node15798;
	wire [4-1:0] node15799;
	wire [4-1:0] node15802;
	wire [4-1:0] node15805;
	wire [4-1:0] node15806;
	wire [4-1:0] node15809;
	wire [4-1:0] node15812;
	wire [4-1:0] node15813;
	wire [4-1:0] node15814;
	wire [4-1:0] node15817;
	wire [4-1:0] node15820;
	wire [4-1:0] node15821;
	wire [4-1:0] node15824;
	wire [4-1:0] node15827;
	wire [4-1:0] node15828;
	wire [4-1:0] node15829;
	wire [4-1:0] node15830;
	wire [4-1:0] node15833;
	wire [4-1:0] node15836;
	wire [4-1:0] node15837;
	wire [4-1:0] node15841;
	wire [4-1:0] node15842;
	wire [4-1:0] node15843;
	wire [4-1:0] node15846;
	wire [4-1:0] node15849;
	wire [4-1:0] node15850;
	wire [4-1:0] node15854;
	wire [4-1:0] node15855;
	wire [4-1:0] node15856;
	wire [4-1:0] node15857;
	wire [4-1:0] node15858;
	wire [4-1:0] node15859;
	wire [4-1:0] node15860;
	wire [4-1:0] node15864;
	wire [4-1:0] node15865;
	wire [4-1:0] node15869;
	wire [4-1:0] node15870;
	wire [4-1:0] node15871;
	wire [4-1:0] node15875;
	wire [4-1:0] node15876;
	wire [4-1:0] node15880;
	wire [4-1:0] node15881;
	wire [4-1:0] node15882;
	wire [4-1:0] node15883;
	wire [4-1:0] node15887;
	wire [4-1:0] node15888;
	wire [4-1:0] node15892;
	wire [4-1:0] node15893;
	wire [4-1:0] node15894;
	wire [4-1:0] node15898;
	wire [4-1:0] node15899;
	wire [4-1:0] node15903;
	wire [4-1:0] node15904;
	wire [4-1:0] node15905;
	wire [4-1:0] node15906;
	wire [4-1:0] node15907;
	wire [4-1:0] node15911;
	wire [4-1:0] node15912;
	wire [4-1:0] node15916;
	wire [4-1:0] node15917;
	wire [4-1:0] node15918;
	wire [4-1:0] node15922;
	wire [4-1:0] node15923;
	wire [4-1:0] node15927;
	wire [4-1:0] node15928;
	wire [4-1:0] node15929;
	wire [4-1:0] node15930;
	wire [4-1:0] node15934;
	wire [4-1:0] node15935;
	wire [4-1:0] node15939;
	wire [4-1:0] node15940;
	wire [4-1:0] node15941;
	wire [4-1:0] node15945;
	wire [4-1:0] node15946;
	wire [4-1:0] node15950;
	wire [4-1:0] node15951;
	wire [4-1:0] node15952;
	wire [4-1:0] node15953;
	wire [4-1:0] node15954;
	wire [4-1:0] node15955;
	wire [4-1:0] node15958;
	wire [4-1:0] node15961;
	wire [4-1:0] node15963;
	wire [4-1:0] node15966;
	wire [4-1:0] node15967;
	wire [4-1:0] node15969;
	wire [4-1:0] node15972;
	wire [4-1:0] node15973;
	wire [4-1:0] node15976;
	wire [4-1:0] node15979;
	wire [4-1:0] node15980;
	wire [4-1:0] node15981;
	wire [4-1:0] node15982;
	wire [4-1:0] node15986;
	wire [4-1:0] node15987;
	wire [4-1:0] node15991;
	wire [4-1:0] node15992;
	wire [4-1:0] node15993;
	wire [4-1:0] node15996;
	wire [4-1:0] node15999;
	wire [4-1:0] node16000;
	wire [4-1:0] node16003;
	wire [4-1:0] node16006;
	wire [4-1:0] node16007;
	wire [4-1:0] node16008;
	wire [4-1:0] node16009;
	wire [4-1:0] node16010;
	wire [4-1:0] node16013;
	wire [4-1:0] node16016;
	wire [4-1:0] node16017;
	wire [4-1:0] node16020;
	wire [4-1:0] node16023;
	wire [4-1:0] node16024;
	wire [4-1:0] node16025;
	wire [4-1:0] node16028;
	wire [4-1:0] node16031;
	wire [4-1:0] node16032;
	wire [4-1:0] node16035;
	wire [4-1:0] node16038;
	wire [4-1:0] node16039;
	wire [4-1:0] node16040;
	wire [4-1:0] node16041;
	wire [4-1:0] node16044;
	wire [4-1:0] node16047;
	wire [4-1:0] node16049;
	wire [4-1:0] node16052;
	wire [4-1:0] node16053;
	wire [4-1:0] node16054;
	wire [4-1:0] node16057;
	wire [4-1:0] node16060;
	wire [4-1:0] node16061;
	wire [4-1:0] node16064;
	wire [4-1:0] node16067;
	wire [4-1:0] node16068;
	wire [4-1:0] node16069;
	wire [4-1:0] node16070;
	wire [4-1:0] node16071;
	wire [4-1:0] node16072;
	wire [4-1:0] node16073;
	wire [4-1:0] node16074;
	wire [4-1:0] node16075;
	wire [4-1:0] node16076;
	wire [4-1:0] node16079;
	wire [4-1:0] node16082;
	wire [4-1:0] node16084;
	wire [4-1:0] node16087;
	wire [4-1:0] node16088;
	wire [4-1:0] node16089;
	wire [4-1:0] node16092;
	wire [4-1:0] node16095;
	wire [4-1:0] node16096;
	wire [4-1:0] node16099;
	wire [4-1:0] node16102;
	wire [4-1:0] node16103;
	wire [4-1:0] node16104;
	wire [4-1:0] node16105;
	wire [4-1:0] node16108;
	wire [4-1:0] node16111;
	wire [4-1:0] node16112;
	wire [4-1:0] node16115;
	wire [4-1:0] node16118;
	wire [4-1:0] node16119;
	wire [4-1:0] node16120;
	wire [4-1:0] node16123;
	wire [4-1:0] node16126;
	wire [4-1:0] node16127;
	wire [4-1:0] node16130;
	wire [4-1:0] node16133;
	wire [4-1:0] node16134;
	wire [4-1:0] node16135;
	wire [4-1:0] node16136;
	wire [4-1:0] node16139;
	wire [4-1:0] node16142;
	wire [4-1:0] node16143;
	wire [4-1:0] node16146;
	wire [4-1:0] node16149;
	wire [4-1:0] node16150;
	wire [4-1:0] node16151;
	wire [4-1:0] node16154;
	wire [4-1:0] node16157;
	wire [4-1:0] node16158;
	wire [4-1:0] node16159;
	wire [4-1:0] node16162;
	wire [4-1:0] node16165;
	wire [4-1:0] node16166;
	wire [4-1:0] node16169;
	wire [4-1:0] node16172;
	wire [4-1:0] node16173;
	wire [4-1:0] node16174;
	wire [4-1:0] node16175;
	wire [4-1:0] node16176;
	wire [4-1:0] node16177;
	wire [4-1:0] node16180;
	wire [4-1:0] node16183;
	wire [4-1:0] node16185;
	wire [4-1:0] node16188;
	wire [4-1:0] node16189;
	wire [4-1:0] node16190;
	wire [4-1:0] node16193;
	wire [4-1:0] node16196;
	wire [4-1:0] node16197;
	wire [4-1:0] node16200;
	wire [4-1:0] node16203;
	wire [4-1:0] node16204;
	wire [4-1:0] node16205;
	wire [4-1:0] node16206;
	wire [4-1:0] node16209;
	wire [4-1:0] node16212;
	wire [4-1:0] node16213;
	wire [4-1:0] node16216;
	wire [4-1:0] node16219;
	wire [4-1:0] node16220;
	wire [4-1:0] node16221;
	wire [4-1:0] node16224;
	wire [4-1:0] node16227;
	wire [4-1:0] node16228;
	wire [4-1:0] node16231;
	wire [4-1:0] node16234;
	wire [4-1:0] node16235;
	wire [4-1:0] node16236;
	wire [4-1:0] node16237;
	wire [4-1:0] node16238;
	wire [4-1:0] node16242;
	wire [4-1:0] node16243;
	wire [4-1:0] node16246;
	wire [4-1:0] node16249;
	wire [4-1:0] node16250;
	wire [4-1:0] node16251;
	wire [4-1:0] node16254;
	wire [4-1:0] node16257;
	wire [4-1:0] node16258;
	wire [4-1:0] node16261;
	wire [4-1:0] node16264;
	wire [4-1:0] node16265;
	wire [4-1:0] node16266;
	wire [4-1:0] node16267;
	wire [4-1:0] node16270;
	wire [4-1:0] node16273;
	wire [4-1:0] node16275;
	wire [4-1:0] node16278;
	wire [4-1:0] node16279;
	wire [4-1:0] node16280;
	wire [4-1:0] node16283;
	wire [4-1:0] node16286;
	wire [4-1:0] node16287;
	wire [4-1:0] node16290;
	wire [4-1:0] node16293;
	wire [4-1:0] node16294;
	wire [4-1:0] node16295;
	wire [4-1:0] node16296;
	wire [4-1:0] node16297;
	wire [4-1:0] node16298;
	wire [4-1:0] node16299;
	wire [4-1:0] node16302;
	wire [4-1:0] node16305;
	wire [4-1:0] node16306;
	wire [4-1:0] node16310;
	wire [4-1:0] node16311;
	wire [4-1:0] node16312;
	wire [4-1:0] node16315;
	wire [4-1:0] node16318;
	wire [4-1:0] node16319;
	wire [4-1:0] node16322;
	wire [4-1:0] node16325;
	wire [4-1:0] node16326;
	wire [4-1:0] node16327;
	wire [4-1:0] node16328;
	wire [4-1:0] node16331;
	wire [4-1:0] node16334;
	wire [4-1:0] node16335;
	wire [4-1:0] node16338;
	wire [4-1:0] node16341;
	wire [4-1:0] node16342;
	wire [4-1:0] node16343;
	wire [4-1:0] node16346;
	wire [4-1:0] node16349;
	wire [4-1:0] node16350;
	wire [4-1:0] node16353;
	wire [4-1:0] node16356;
	wire [4-1:0] node16357;
	wire [4-1:0] node16358;
	wire [4-1:0] node16359;
	wire [4-1:0] node16360;
	wire [4-1:0] node16363;
	wire [4-1:0] node16366;
	wire [4-1:0] node16367;
	wire [4-1:0] node16370;
	wire [4-1:0] node16373;
	wire [4-1:0] node16374;
	wire [4-1:0] node16375;
	wire [4-1:0] node16379;
	wire [4-1:0] node16380;
	wire [4-1:0] node16384;
	wire [4-1:0] node16385;
	wire [4-1:0] node16386;
	wire [4-1:0] node16389;
	wire [4-1:0] node16392;
	wire [4-1:0] node16393;
	wire [4-1:0] node16394;
	wire [4-1:0] node16397;
	wire [4-1:0] node16400;
	wire [4-1:0] node16401;
	wire [4-1:0] node16404;
	wire [4-1:0] node16407;
	wire [4-1:0] node16408;
	wire [4-1:0] node16409;
	wire [4-1:0] node16410;
	wire [4-1:0] node16411;
	wire [4-1:0] node16412;
	wire [4-1:0] node16415;
	wire [4-1:0] node16418;
	wire [4-1:0] node16419;
	wire [4-1:0] node16422;
	wire [4-1:0] node16425;
	wire [4-1:0] node16426;
	wire [4-1:0] node16427;
	wire [4-1:0] node16430;
	wire [4-1:0] node16434;
	wire [4-1:0] node16435;
	wire [4-1:0] node16436;
	wire [4-1:0] node16438;
	wire [4-1:0] node16441;
	wire [4-1:0] node16443;
	wire [4-1:0] node16446;
	wire [4-1:0] node16447;
	wire [4-1:0] node16449;
	wire [4-1:0] node16452;
	wire [4-1:0] node16454;
	wire [4-1:0] node16457;
	wire [4-1:0] node16458;
	wire [4-1:0] node16459;
	wire [4-1:0] node16460;
	wire [4-1:0] node16461;
	wire [4-1:0] node16464;
	wire [4-1:0] node16467;
	wire [4-1:0] node16469;
	wire [4-1:0] node16472;
	wire [4-1:0] node16473;
	wire [4-1:0] node16474;
	wire [4-1:0] node16477;
	wire [4-1:0] node16480;
	wire [4-1:0] node16481;
	wire [4-1:0] node16484;
	wire [4-1:0] node16487;
	wire [4-1:0] node16488;
	wire [4-1:0] node16489;
	wire [4-1:0] node16490;
	wire [4-1:0] node16493;
	wire [4-1:0] node16496;
	wire [4-1:0] node16497;
	wire [4-1:0] node16500;
	wire [4-1:0] node16503;
	wire [4-1:0] node16504;
	wire [4-1:0] node16505;
	wire [4-1:0] node16508;
	wire [4-1:0] node16511;
	wire [4-1:0] node16512;
	wire [4-1:0] node16515;
	wire [4-1:0] node16518;
	wire [4-1:0] node16519;
	wire [4-1:0] node16520;
	wire [4-1:0] node16521;
	wire [4-1:0] node16522;
	wire [4-1:0] node16523;
	wire [4-1:0] node16524;
	wire [4-1:0] node16525;
	wire [4-1:0] node16529;
	wire [4-1:0] node16530;
	wire [4-1:0] node16533;
	wire [4-1:0] node16536;
	wire [4-1:0] node16537;
	wire [4-1:0] node16538;
	wire [4-1:0] node16541;
	wire [4-1:0] node16544;
	wire [4-1:0] node16545;
	wire [4-1:0] node16549;
	wire [4-1:0] node16550;
	wire [4-1:0] node16551;
	wire [4-1:0] node16552;
	wire [4-1:0] node16555;
	wire [4-1:0] node16558;
	wire [4-1:0] node16559;
	wire [4-1:0] node16562;
	wire [4-1:0] node16565;
	wire [4-1:0] node16566;
	wire [4-1:0] node16567;
	wire [4-1:0] node16570;
	wire [4-1:0] node16573;
	wire [4-1:0] node16575;
	wire [4-1:0] node16578;
	wire [4-1:0] node16579;
	wire [4-1:0] node16580;
	wire [4-1:0] node16581;
	wire [4-1:0] node16582;
	wire [4-1:0] node16585;
	wire [4-1:0] node16588;
	wire [4-1:0] node16589;
	wire [4-1:0] node16592;
	wire [4-1:0] node16595;
	wire [4-1:0] node16596;
	wire [4-1:0] node16597;
	wire [4-1:0] node16601;
	wire [4-1:0] node16602;
	wire [4-1:0] node16605;
	wire [4-1:0] node16608;
	wire [4-1:0] node16609;
	wire [4-1:0] node16610;
	wire [4-1:0] node16611;
	wire [4-1:0] node16614;
	wire [4-1:0] node16617;
	wire [4-1:0] node16619;
	wire [4-1:0] node16622;
	wire [4-1:0] node16623;
	wire [4-1:0] node16624;
	wire [4-1:0] node16627;
	wire [4-1:0] node16630;
	wire [4-1:0] node16631;
	wire [4-1:0] node16634;
	wire [4-1:0] node16637;
	wire [4-1:0] node16638;
	wire [4-1:0] node16639;
	wire [4-1:0] node16640;
	wire [4-1:0] node16641;
	wire [4-1:0] node16643;
	wire [4-1:0] node16646;
	wire [4-1:0] node16647;
	wire [4-1:0] node16650;
	wire [4-1:0] node16653;
	wire [4-1:0] node16654;
	wire [4-1:0] node16655;
	wire [4-1:0] node16658;
	wire [4-1:0] node16661;
	wire [4-1:0] node16662;
	wire [4-1:0] node16665;
	wire [4-1:0] node16668;
	wire [4-1:0] node16669;
	wire [4-1:0] node16670;
	wire [4-1:0] node16672;
	wire [4-1:0] node16675;
	wire [4-1:0] node16677;
	wire [4-1:0] node16680;
	wire [4-1:0] node16681;
	wire [4-1:0] node16683;
	wire [4-1:0] node16686;
	wire [4-1:0] node16688;
	wire [4-1:0] node16691;
	wire [4-1:0] node16692;
	wire [4-1:0] node16693;
	wire [4-1:0] node16694;
	wire [4-1:0] node16695;
	wire [4-1:0] node16698;
	wire [4-1:0] node16701;
	wire [4-1:0] node16702;
	wire [4-1:0] node16705;
	wire [4-1:0] node16708;
	wire [4-1:0] node16709;
	wire [4-1:0] node16710;
	wire [4-1:0] node16713;
	wire [4-1:0] node16716;
	wire [4-1:0] node16718;
	wire [4-1:0] node16721;
	wire [4-1:0] node16722;
	wire [4-1:0] node16723;
	wire [4-1:0] node16725;
	wire [4-1:0] node16728;
	wire [4-1:0] node16730;
	wire [4-1:0] node16733;
	wire [4-1:0] node16734;
	wire [4-1:0] node16736;
	wire [4-1:0] node16739;
	wire [4-1:0] node16741;
	wire [4-1:0] node16744;
	wire [4-1:0] node16745;
	wire [4-1:0] node16746;
	wire [4-1:0] node16747;
	wire [4-1:0] node16748;
	wire [4-1:0] node16749;
	wire [4-1:0] node16750;
	wire [4-1:0] node16753;
	wire [4-1:0] node16756;
	wire [4-1:0] node16757;
	wire [4-1:0] node16760;
	wire [4-1:0] node16763;
	wire [4-1:0] node16764;
	wire [4-1:0] node16765;
	wire [4-1:0] node16768;
	wire [4-1:0] node16771;
	wire [4-1:0] node16772;
	wire [4-1:0] node16775;
	wire [4-1:0] node16778;
	wire [4-1:0] node16779;
	wire [4-1:0] node16780;
	wire [4-1:0] node16781;
	wire [4-1:0] node16784;
	wire [4-1:0] node16787;
	wire [4-1:0] node16788;
	wire [4-1:0] node16792;
	wire [4-1:0] node16793;
	wire [4-1:0] node16794;
	wire [4-1:0] node16797;
	wire [4-1:0] node16800;
	wire [4-1:0] node16801;
	wire [4-1:0] node16805;
	wire [4-1:0] node16806;
	wire [4-1:0] node16807;
	wire [4-1:0] node16808;
	wire [4-1:0] node16809;
	wire [4-1:0] node16812;
	wire [4-1:0] node16815;
	wire [4-1:0] node16817;
	wire [4-1:0] node16820;
	wire [4-1:0] node16821;
	wire [4-1:0] node16822;
	wire [4-1:0] node16825;
	wire [4-1:0] node16828;
	wire [4-1:0] node16829;
	wire [4-1:0] node16832;
	wire [4-1:0] node16835;
	wire [4-1:0] node16836;
	wire [4-1:0] node16837;
	wire [4-1:0] node16838;
	wire [4-1:0] node16842;
	wire [4-1:0] node16843;
	wire [4-1:0] node16846;
	wire [4-1:0] node16849;
	wire [4-1:0] node16850;
	wire [4-1:0] node16852;
	wire [4-1:0] node16855;
	wire [4-1:0] node16856;
	wire [4-1:0] node16859;
	wire [4-1:0] node16862;
	wire [4-1:0] node16863;
	wire [4-1:0] node16864;
	wire [4-1:0] node16865;
	wire [4-1:0] node16866;
	wire [4-1:0] node16867;
	wire [4-1:0] node16871;
	wire [4-1:0] node16872;
	wire [4-1:0] node16876;
	wire [4-1:0] node16877;
	wire [4-1:0] node16878;
	wire [4-1:0] node16882;
	wire [4-1:0] node16883;
	wire [4-1:0] node16887;
	wire [4-1:0] node16888;
	wire [4-1:0] node16889;
	wire [4-1:0] node16890;
	wire [4-1:0] node16893;
	wire [4-1:0] node16896;
	wire [4-1:0] node16897;
	wire [4-1:0] node16900;
	wire [4-1:0] node16903;
	wire [4-1:0] node16904;
	wire [4-1:0] node16905;
	wire [4-1:0] node16909;
	wire [4-1:0] node16910;
	wire [4-1:0] node16913;
	wire [4-1:0] node16916;
	wire [4-1:0] node16917;
	wire [4-1:0] node16918;
	wire [4-1:0] node16919;
	wire [4-1:0] node16920;
	wire [4-1:0] node16923;
	wire [4-1:0] node16926;
	wire [4-1:0] node16928;
	wire [4-1:0] node16931;
	wire [4-1:0] node16932;
	wire [4-1:0] node16933;
	wire [4-1:0] node16937;
	wire [4-1:0] node16938;
	wire [4-1:0] node16941;
	wire [4-1:0] node16944;
	wire [4-1:0] node16945;
	wire [4-1:0] node16946;
	wire [4-1:0] node16947;
	wire [4-1:0] node16951;
	wire [4-1:0] node16952;
	wire [4-1:0] node16955;
	wire [4-1:0] node16958;
	wire [4-1:0] node16959;
	wire [4-1:0] node16960;
	wire [4-1:0] node16963;
	wire [4-1:0] node16966;
	wire [4-1:0] node16967;
	wire [4-1:0] node16971;
	wire [4-1:0] node16972;
	wire [4-1:0] node16973;
	wire [4-1:0] node16974;
	wire [4-1:0] node16975;
	wire [4-1:0] node16976;
	wire [4-1:0] node16977;
	wire [4-1:0] node16978;
	wire [4-1:0] node16979;
	wire [4-1:0] node16982;
	wire [4-1:0] node16985;
	wire [4-1:0] node16986;
	wire [4-1:0] node16989;
	wire [4-1:0] node16992;
	wire [4-1:0] node16993;
	wire [4-1:0] node16995;
	wire [4-1:0] node16998;
	wire [4-1:0] node16999;
	wire [4-1:0] node17002;
	wire [4-1:0] node17005;
	wire [4-1:0] node17006;
	wire [4-1:0] node17007;
	wire [4-1:0] node17008;
	wire [4-1:0] node17011;
	wire [4-1:0] node17014;
	wire [4-1:0] node17015;
	wire [4-1:0] node17018;
	wire [4-1:0] node17021;
	wire [4-1:0] node17022;
	wire [4-1:0] node17023;
	wire [4-1:0] node17026;
	wire [4-1:0] node17029;
	wire [4-1:0] node17030;
	wire [4-1:0] node17033;
	wire [4-1:0] node17036;
	wire [4-1:0] node17037;
	wire [4-1:0] node17038;
	wire [4-1:0] node17039;
	wire [4-1:0] node17042;
	wire [4-1:0] node17045;
	wire [4-1:0] node17046;
	wire [4-1:0] node17049;
	wire [4-1:0] node17052;
	wire [4-1:0] node17053;
	wire [4-1:0] node17054;
	wire [4-1:0] node17056;
	wire [4-1:0] node17059;
	wire [4-1:0] node17060;
	wire [4-1:0] node17063;
	wire [4-1:0] node17066;
	wire [4-1:0] node17067;
	wire [4-1:0] node17068;
	wire [4-1:0] node17071;
	wire [4-1:0] node17074;
	wire [4-1:0] node17075;
	wire [4-1:0] node17078;
	wire [4-1:0] node17081;
	wire [4-1:0] node17082;
	wire [4-1:0] node17083;
	wire [4-1:0] node17084;
	wire [4-1:0] node17085;
	wire [4-1:0] node17086;
	wire [4-1:0] node17089;
	wire [4-1:0] node17092;
	wire [4-1:0] node17093;
	wire [4-1:0] node17096;
	wire [4-1:0] node17099;
	wire [4-1:0] node17100;
	wire [4-1:0] node17101;
	wire [4-1:0] node17104;
	wire [4-1:0] node17107;
	wire [4-1:0] node17108;
	wire [4-1:0] node17111;
	wire [4-1:0] node17114;
	wire [4-1:0] node17115;
	wire [4-1:0] node17116;
	wire [4-1:0] node17117;
	wire [4-1:0] node17121;
	wire [4-1:0] node17122;
	wire [4-1:0] node17125;
	wire [4-1:0] node17128;
	wire [4-1:0] node17129;
	wire [4-1:0] node17130;
	wire [4-1:0] node17133;
	wire [4-1:0] node17136;
	wire [4-1:0] node17137;
	wire [4-1:0] node17140;
	wire [4-1:0] node17143;
	wire [4-1:0] node17144;
	wire [4-1:0] node17145;
	wire [4-1:0] node17146;
	wire [4-1:0] node17147;
	wire [4-1:0] node17150;
	wire [4-1:0] node17153;
	wire [4-1:0] node17154;
	wire [4-1:0] node17157;
	wire [4-1:0] node17160;
	wire [4-1:0] node17161;
	wire [4-1:0] node17162;
	wire [4-1:0] node17165;
	wire [4-1:0] node17168;
	wire [4-1:0] node17170;
	wire [4-1:0] node17173;
	wire [4-1:0] node17174;
	wire [4-1:0] node17175;
	wire [4-1:0] node17177;
	wire [4-1:0] node17180;
	wire [4-1:0] node17181;
	wire [4-1:0] node17184;
	wire [4-1:0] node17187;
	wire [4-1:0] node17188;
	wire [4-1:0] node17189;
	wire [4-1:0] node17193;
	wire [4-1:0] node17194;
	wire [4-1:0] node17197;
	wire [4-1:0] node17200;
	wire [4-1:0] node17201;
	wire [4-1:0] node17202;
	wire [4-1:0] node17203;
	wire [4-1:0] node17204;
	wire [4-1:0] node17205;
	wire [4-1:0] node17206;
	wire [4-1:0] node17209;
	wire [4-1:0] node17212;
	wire [4-1:0] node17213;
	wire [4-1:0] node17216;
	wire [4-1:0] node17219;
	wire [4-1:0] node17220;
	wire [4-1:0] node17221;
	wire [4-1:0] node17224;
	wire [4-1:0] node17227;
	wire [4-1:0] node17228;
	wire [4-1:0] node17231;
	wire [4-1:0] node17234;
	wire [4-1:0] node17235;
	wire [4-1:0] node17236;
	wire [4-1:0] node17239;
	wire [4-1:0] node17242;
	wire [4-1:0] node17243;
	wire [4-1:0] node17244;
	wire [4-1:0] node17247;
	wire [4-1:0] node17250;
	wire [4-1:0] node17251;
	wire [4-1:0] node17254;
	wire [4-1:0] node17257;
	wire [4-1:0] node17258;
	wire [4-1:0] node17259;
	wire [4-1:0] node17260;
	wire [4-1:0] node17261;
	wire [4-1:0] node17264;
	wire [4-1:0] node17267;
	wire [4-1:0] node17268;
	wire [4-1:0] node17271;
	wire [4-1:0] node17274;
	wire [4-1:0] node17275;
	wire [4-1:0] node17277;
	wire [4-1:0] node17280;
	wire [4-1:0] node17281;
	wire [4-1:0] node17284;
	wire [4-1:0] node17287;
	wire [4-1:0] node17288;
	wire [4-1:0] node17289;
	wire [4-1:0] node17291;
	wire [4-1:0] node17294;
	wire [4-1:0] node17296;
	wire [4-1:0] node17299;
	wire [4-1:0] node17300;
	wire [4-1:0] node17302;
	wire [4-1:0] node17305;
	wire [4-1:0] node17307;
	wire [4-1:0] node17310;
	wire [4-1:0] node17311;
	wire [4-1:0] node17312;
	wire [4-1:0] node17313;
	wire [4-1:0] node17314;
	wire [4-1:0] node17315;
	wire [4-1:0] node17318;
	wire [4-1:0] node17321;
	wire [4-1:0] node17322;
	wire [4-1:0] node17325;
	wire [4-1:0] node17328;
	wire [4-1:0] node17329;
	wire [4-1:0] node17330;
	wire [4-1:0] node17333;
	wire [4-1:0] node17336;
	wire [4-1:0] node17337;
	wire [4-1:0] node17340;
	wire [4-1:0] node17343;
	wire [4-1:0] node17344;
	wire [4-1:0] node17345;
	wire [4-1:0] node17347;
	wire [4-1:0] node17350;
	wire [4-1:0] node17352;
	wire [4-1:0] node17355;
	wire [4-1:0] node17356;
	wire [4-1:0] node17358;
	wire [4-1:0] node17361;
	wire [4-1:0] node17363;
	wire [4-1:0] node17366;
	wire [4-1:0] node17367;
	wire [4-1:0] node17368;
	wire [4-1:0] node17369;
	wire [4-1:0] node17370;
	wire [4-1:0] node17373;
	wire [4-1:0] node17376;
	wire [4-1:0] node17377;
	wire [4-1:0] node17380;
	wire [4-1:0] node17383;
	wire [4-1:0] node17384;
	wire [4-1:0] node17385;
	wire [4-1:0] node17388;
	wire [4-1:0] node17391;
	wire [4-1:0] node17392;
	wire [4-1:0] node17395;
	wire [4-1:0] node17398;
	wire [4-1:0] node17399;
	wire [4-1:0] node17400;
	wire [4-1:0] node17401;
	wire [4-1:0] node17404;
	wire [4-1:0] node17407;
	wire [4-1:0] node17408;
	wire [4-1:0] node17411;
	wire [4-1:0] node17414;
	wire [4-1:0] node17415;
	wire [4-1:0] node17416;
	wire [4-1:0] node17420;
	wire [4-1:0] node17421;
	wire [4-1:0] node17424;
	wire [4-1:0] node17427;
	wire [4-1:0] node17428;
	wire [4-1:0] node17429;
	wire [4-1:0] node17430;
	wire [4-1:0] node17431;
	wire [4-1:0] node17432;
	wire [4-1:0] node17433;
	wire [4-1:0] node17434;
	wire [4-1:0] node17437;
	wire [4-1:0] node17440;
	wire [4-1:0] node17441;
	wire [4-1:0] node17444;
	wire [4-1:0] node17447;
	wire [4-1:0] node17448;
	wire [4-1:0] node17449;
	wire [4-1:0] node17453;
	wire [4-1:0] node17454;
	wire [4-1:0] node17457;
	wire [4-1:0] node17460;
	wire [4-1:0] node17461;
	wire [4-1:0] node17462;
	wire [4-1:0] node17463;
	wire [4-1:0] node17466;
	wire [4-1:0] node17469;
	wire [4-1:0] node17470;
	wire [4-1:0] node17473;
	wire [4-1:0] node17476;
	wire [4-1:0] node17477;
	wire [4-1:0] node17478;
	wire [4-1:0] node17481;
	wire [4-1:0] node17484;
	wire [4-1:0] node17485;
	wire [4-1:0] node17488;
	wire [4-1:0] node17491;
	wire [4-1:0] node17492;
	wire [4-1:0] node17493;
	wire [4-1:0] node17494;
	wire [4-1:0] node17495;
	wire [4-1:0] node17498;
	wire [4-1:0] node17501;
	wire [4-1:0] node17502;
	wire [4-1:0] node17506;
	wire [4-1:0] node17507;
	wire [4-1:0] node17508;
	wire [4-1:0] node17511;
	wire [4-1:0] node17514;
	wire [4-1:0] node17515;
	wire [4-1:0] node17518;
	wire [4-1:0] node17521;
	wire [4-1:0] node17522;
	wire [4-1:0] node17523;
	wire [4-1:0] node17524;
	wire [4-1:0] node17527;
	wire [4-1:0] node17530;
	wire [4-1:0] node17531;
	wire [4-1:0] node17535;
	wire [4-1:0] node17536;
	wire [4-1:0] node17537;
	wire [4-1:0] node17540;
	wire [4-1:0] node17543;
	wire [4-1:0] node17544;
	wire [4-1:0] node17547;
	wire [4-1:0] node17550;
	wire [4-1:0] node17551;
	wire [4-1:0] node17552;
	wire [4-1:0] node17553;
	wire [4-1:0] node17554;
	wire [4-1:0] node17555;
	wire [4-1:0] node17558;
	wire [4-1:0] node17561;
	wire [4-1:0] node17562;
	wire [4-1:0] node17565;
	wire [4-1:0] node17568;
	wire [4-1:0] node17569;
	wire [4-1:0] node17570;
	wire [4-1:0] node17574;
	wire [4-1:0] node17575;
	wire [4-1:0] node17578;
	wire [4-1:0] node17581;
	wire [4-1:0] node17582;
	wire [4-1:0] node17583;
	wire [4-1:0] node17585;
	wire [4-1:0] node17588;
	wire [4-1:0] node17590;
	wire [4-1:0] node17593;
	wire [4-1:0] node17594;
	wire [4-1:0] node17596;
	wire [4-1:0] node17599;
	wire [4-1:0] node17601;
	wire [4-1:0] node17604;
	wire [4-1:0] node17605;
	wire [4-1:0] node17606;
	wire [4-1:0] node17607;
	wire [4-1:0] node17608;
	wire [4-1:0] node17611;
	wire [4-1:0] node17614;
	wire [4-1:0] node17615;
	wire [4-1:0] node17618;
	wire [4-1:0] node17621;
	wire [4-1:0] node17622;
	wire [4-1:0] node17624;
	wire [4-1:0] node17627;
	wire [4-1:0] node17628;
	wire [4-1:0] node17631;
	wire [4-1:0] node17634;
	wire [4-1:0] node17635;
	wire [4-1:0] node17636;
	wire [4-1:0] node17638;
	wire [4-1:0] node17641;
	wire [4-1:0] node17643;
	wire [4-1:0] node17646;
	wire [4-1:0] node17647;
	wire [4-1:0] node17649;
	wire [4-1:0] node17652;
	wire [4-1:0] node17654;
	wire [4-1:0] node17657;
	wire [4-1:0] node17658;
	wire [4-1:0] node17659;
	wire [4-1:0] node17660;
	wire [4-1:0] node17661;
	wire [4-1:0] node17662;
	wire [4-1:0] node17663;
	wire [4-1:0] node17666;
	wire [4-1:0] node17669;
	wire [4-1:0] node17670;
	wire [4-1:0] node17673;
	wire [4-1:0] node17676;
	wire [4-1:0] node17677;
	wire [4-1:0] node17678;
	wire [4-1:0] node17681;
	wire [4-1:0] node17684;
	wire [4-1:0] node17685;
	wire [4-1:0] node17688;
	wire [4-1:0] node17691;
	wire [4-1:0] node17692;
	wire [4-1:0] node17693;
	wire [4-1:0] node17694;
	wire [4-1:0] node17698;
	wire [4-1:0] node17699;
	wire [4-1:0] node17702;
	wire [4-1:0] node17705;
	wire [4-1:0] node17706;
	wire [4-1:0] node17707;
	wire [4-1:0] node17710;
	wire [4-1:0] node17713;
	wire [4-1:0] node17715;
	wire [4-1:0] node17718;
	wire [4-1:0] node17719;
	wire [4-1:0] node17720;
	wire [4-1:0] node17721;
	wire [4-1:0] node17722;
	wire [4-1:0] node17725;
	wire [4-1:0] node17728;
	wire [4-1:0] node17729;
	wire [4-1:0] node17732;
	wire [4-1:0] node17735;
	wire [4-1:0] node17736;
	wire [4-1:0] node17737;
	wire [4-1:0] node17740;
	wire [4-1:0] node17743;
	wire [4-1:0] node17744;
	wire [4-1:0] node17747;
	wire [4-1:0] node17750;
	wire [4-1:0] node17751;
	wire [4-1:0] node17752;
	wire [4-1:0] node17753;
	wire [4-1:0] node17757;
	wire [4-1:0] node17758;
	wire [4-1:0] node17761;
	wire [4-1:0] node17764;
	wire [4-1:0] node17765;
	wire [4-1:0] node17766;
	wire [4-1:0] node17770;
	wire [4-1:0] node17772;
	wire [4-1:0] node17775;
	wire [4-1:0] node17776;
	wire [4-1:0] node17777;
	wire [4-1:0] node17778;
	wire [4-1:0] node17779;
	wire [4-1:0] node17782;
	wire [4-1:0] node17785;
	wire [4-1:0] node17786;
	wire [4-1:0] node17788;
	wire [4-1:0] node17791;
	wire [4-1:0] node17792;
	wire [4-1:0] node17795;
	wire [4-1:0] node17798;
	wire [4-1:0] node17799;
	wire [4-1:0] node17800;
	wire [4-1:0] node17803;
	wire [4-1:0] node17806;
	wire [4-1:0] node17807;
	wire [4-1:0] node17808;
	wire [4-1:0] node17811;
	wire [4-1:0] node17814;
	wire [4-1:0] node17815;
	wire [4-1:0] node17818;
	wire [4-1:0] node17821;
	wire [4-1:0] node17822;
	wire [4-1:0] node17823;
	wire [4-1:0] node17824;
	wire [4-1:0] node17825;
	wire [4-1:0] node17828;
	wire [4-1:0] node17831;
	wire [4-1:0] node17832;
	wire [4-1:0] node17835;
	wire [4-1:0] node17838;
	wire [4-1:0] node17839;
	wire [4-1:0] node17840;
	wire [4-1:0] node17844;
	wire [4-1:0] node17845;
	wire [4-1:0] node17848;
	wire [4-1:0] node17851;
	wire [4-1:0] node17852;
	wire [4-1:0] node17853;
	wire [4-1:0] node17854;
	wire [4-1:0] node17857;
	wire [4-1:0] node17860;
	wire [4-1:0] node17861;
	wire [4-1:0] node17864;
	wire [4-1:0] node17867;
	wire [4-1:0] node17868;
	wire [4-1:0] node17869;
	wire [4-1:0] node17872;
	wire [4-1:0] node17875;
	wire [4-1:0] node17876;
	wire [4-1:0] node17879;
	wire [4-1:0] node17882;
	wire [4-1:0] node17883;
	wire [4-1:0] node17884;
	wire [4-1:0] node17885;
	wire [4-1:0] node17886;
	wire [4-1:0] node17887;
	wire [4-1:0] node17888;
	wire [4-1:0] node17889;
	wire [4-1:0] node17890;
	wire [4-1:0] node17891;
	wire [4-1:0] node17892;
	wire [4-1:0] node17895;
	wire [4-1:0] node17898;
	wire [4-1:0] node17899;
	wire [4-1:0] node17902;
	wire [4-1:0] node17905;
	wire [4-1:0] node17906;
	wire [4-1:0] node17909;
	wire [4-1:0] node17912;
	wire [4-1:0] node17913;
	wire [4-1:0] node17914;
	wire [4-1:0] node17915;
	wire [4-1:0] node17919;
	wire [4-1:0] node17920;
	wire [4-1:0] node17923;
	wire [4-1:0] node17926;
	wire [4-1:0] node17927;
	wire [4-1:0] node17929;
	wire [4-1:0] node17932;
	wire [4-1:0] node17933;
	wire [4-1:0] node17937;
	wire [4-1:0] node17938;
	wire [4-1:0] node17939;
	wire [4-1:0] node17940;
	wire [4-1:0] node17941;
	wire [4-1:0] node17944;
	wire [4-1:0] node17947;
	wire [4-1:0] node17948;
	wire [4-1:0] node17951;
	wire [4-1:0] node17954;
	wire [4-1:0] node17955;
	wire [4-1:0] node17958;
	wire [4-1:0] node17961;
	wire [4-1:0] node17962;
	wire [4-1:0] node17963;
	wire [4-1:0] node17964;
	wire [4-1:0] node17967;
	wire [4-1:0] node17970;
	wire [4-1:0] node17972;
	wire [4-1:0] node17975;
	wire [4-1:0] node17976;
	wire [4-1:0] node17977;
	wire [4-1:0] node17980;
	wire [4-1:0] node17983;
	wire [4-1:0] node17984;
	wire [4-1:0] node17987;
	wire [4-1:0] node17990;
	wire [4-1:0] node17991;
	wire [4-1:0] node17992;
	wire [4-1:0] node17993;
	wire [4-1:0] node17994;
	wire [4-1:0] node17995;
	wire [4-1:0] node17998;
	wire [4-1:0] node18001;
	wire [4-1:0] node18002;
	wire [4-1:0] node18005;
	wire [4-1:0] node18008;
	wire [4-1:0] node18009;
	wire [4-1:0] node18012;
	wire [4-1:0] node18015;
	wire [4-1:0] node18016;
	wire [4-1:0] node18017;
	wire [4-1:0] node18018;
	wire [4-1:0] node18021;
	wire [4-1:0] node18024;
	wire [4-1:0] node18025;
	wire [4-1:0] node18028;
	wire [4-1:0] node18031;
	wire [4-1:0] node18032;
	wire [4-1:0] node18033;
	wire [4-1:0] node18036;
	wire [4-1:0] node18039;
	wire [4-1:0] node18040;
	wire [4-1:0] node18043;
	wire [4-1:0] node18046;
	wire [4-1:0] node18047;
	wire [4-1:0] node18048;
	wire [4-1:0] node18049;
	wire [4-1:0] node18050;
	wire [4-1:0] node18053;
	wire [4-1:0] node18056;
	wire [4-1:0] node18057;
	wire [4-1:0] node18060;
	wire [4-1:0] node18063;
	wire [4-1:0] node18064;
	wire [4-1:0] node18065;
	wire [4-1:0] node18068;
	wire [4-1:0] node18071;
	wire [4-1:0] node18072;
	wire [4-1:0] node18075;
	wire [4-1:0] node18078;
	wire [4-1:0] node18079;
	wire [4-1:0] node18080;
	wire [4-1:0] node18082;
	wire [4-1:0] node18085;
	wire [4-1:0] node18086;
	wire [4-1:0] node18089;
	wire [4-1:0] node18092;
	wire [4-1:0] node18093;
	wire [4-1:0] node18094;
	wire [4-1:0] node18097;
	wire [4-1:0] node18100;
	wire [4-1:0] node18101;
	wire [4-1:0] node18104;
	wire [4-1:0] node18107;
	wire [4-1:0] node18108;
	wire [4-1:0] node18109;
	wire [4-1:0] node18110;
	wire [4-1:0] node18111;
	wire [4-1:0] node18112;
	wire [4-1:0] node18113;
	wire [4-1:0] node18116;
	wire [4-1:0] node18119;
	wire [4-1:0] node18120;
	wire [4-1:0] node18123;
	wire [4-1:0] node18126;
	wire [4-1:0] node18127;
	wire [4-1:0] node18128;
	wire [4-1:0] node18131;
	wire [4-1:0] node18134;
	wire [4-1:0] node18135;
	wire [4-1:0] node18138;
	wire [4-1:0] node18141;
	wire [4-1:0] node18142;
	wire [4-1:0] node18143;
	wire [4-1:0] node18144;
	wire [4-1:0] node18147;
	wire [4-1:0] node18150;
	wire [4-1:0] node18151;
	wire [4-1:0] node18154;
	wire [4-1:0] node18157;
	wire [4-1:0] node18158;
	wire [4-1:0] node18159;
	wire [4-1:0] node18162;
	wire [4-1:0] node18165;
	wire [4-1:0] node18166;
	wire [4-1:0] node18169;
	wire [4-1:0] node18172;
	wire [4-1:0] node18173;
	wire [4-1:0] node18174;
	wire [4-1:0] node18175;
	wire [4-1:0] node18176;
	wire [4-1:0] node18179;
	wire [4-1:0] node18182;
	wire [4-1:0] node18183;
	wire [4-1:0] node18186;
	wire [4-1:0] node18189;
	wire [4-1:0] node18190;
	wire [4-1:0] node18191;
	wire [4-1:0] node18194;
	wire [4-1:0] node18197;
	wire [4-1:0] node18198;
	wire [4-1:0] node18201;
	wire [4-1:0] node18204;
	wire [4-1:0] node18205;
	wire [4-1:0] node18206;
	wire [4-1:0] node18208;
	wire [4-1:0] node18211;
	wire [4-1:0] node18213;
	wire [4-1:0] node18216;
	wire [4-1:0] node18217;
	wire [4-1:0] node18219;
	wire [4-1:0] node18222;
	wire [4-1:0] node18224;
	wire [4-1:0] node18227;
	wire [4-1:0] node18228;
	wire [4-1:0] node18229;
	wire [4-1:0] node18230;
	wire [4-1:0] node18231;
	wire [4-1:0] node18232;
	wire [4-1:0] node18235;
	wire [4-1:0] node18238;
	wire [4-1:0] node18240;
	wire [4-1:0] node18243;
	wire [4-1:0] node18244;
	wire [4-1:0] node18247;
	wire [4-1:0] node18248;
	wire [4-1:0] node18251;
	wire [4-1:0] node18254;
	wire [4-1:0] node18255;
	wire [4-1:0] node18256;
	wire [4-1:0] node18259;
	wire [4-1:0] node18262;
	wire [4-1:0] node18263;
	wire [4-1:0] node18264;
	wire [4-1:0] node18267;
	wire [4-1:0] node18270;
	wire [4-1:0] node18271;
	wire [4-1:0] node18274;
	wire [4-1:0] node18277;
	wire [4-1:0] node18278;
	wire [4-1:0] node18279;
	wire [4-1:0] node18280;
	wire [4-1:0] node18281;
	wire [4-1:0] node18284;
	wire [4-1:0] node18287;
	wire [4-1:0] node18289;
	wire [4-1:0] node18292;
	wire [4-1:0] node18293;
	wire [4-1:0] node18294;
	wire [4-1:0] node18298;
	wire [4-1:0] node18300;
	wire [4-1:0] node18303;
	wire [4-1:0] node18304;
	wire [4-1:0] node18305;
	wire [4-1:0] node18307;
	wire [4-1:0] node18310;
	wire [4-1:0] node18312;
	wire [4-1:0] node18315;
	wire [4-1:0] node18316;
	wire [4-1:0] node18318;
	wire [4-1:0] node18321;
	wire [4-1:0] node18323;
	wire [4-1:0] node18326;
	wire [4-1:0] node18327;
	wire [4-1:0] node18328;
	wire [4-1:0] node18329;
	wire [4-1:0] node18330;
	wire [4-1:0] node18331;
	wire [4-1:0] node18332;
	wire [4-1:0] node18333;
	wire [4-1:0] node18336;
	wire [4-1:0] node18339;
	wire [4-1:0] node18340;
	wire [4-1:0] node18343;
	wire [4-1:0] node18346;
	wire [4-1:0] node18347;
	wire [4-1:0] node18348;
	wire [4-1:0] node18351;
	wire [4-1:0] node18354;
	wire [4-1:0] node18356;
	wire [4-1:0] node18359;
	wire [4-1:0] node18360;
	wire [4-1:0] node18361;
	wire [4-1:0] node18362;
	wire [4-1:0] node18365;
	wire [4-1:0] node18368;
	wire [4-1:0] node18369;
	wire [4-1:0] node18372;
	wire [4-1:0] node18375;
	wire [4-1:0] node18376;
	wire [4-1:0] node18378;
	wire [4-1:0] node18381;
	wire [4-1:0] node18382;
	wire [4-1:0] node18386;
	wire [4-1:0] node18387;
	wire [4-1:0] node18388;
	wire [4-1:0] node18389;
	wire [4-1:0] node18390;
	wire [4-1:0] node18393;
	wire [4-1:0] node18396;
	wire [4-1:0] node18397;
	wire [4-1:0] node18400;
	wire [4-1:0] node18403;
	wire [4-1:0] node18404;
	wire [4-1:0] node18406;
	wire [4-1:0] node18409;
	wire [4-1:0] node18410;
	wire [4-1:0] node18413;
	wire [4-1:0] node18416;
	wire [4-1:0] node18417;
	wire [4-1:0] node18418;
	wire [4-1:0] node18420;
	wire [4-1:0] node18423;
	wire [4-1:0] node18425;
	wire [4-1:0] node18428;
	wire [4-1:0] node18429;
	wire [4-1:0] node18431;
	wire [4-1:0] node18434;
	wire [4-1:0] node18436;
	wire [4-1:0] node18439;
	wire [4-1:0] node18440;
	wire [4-1:0] node18441;
	wire [4-1:0] node18442;
	wire [4-1:0] node18443;
	wire [4-1:0] node18444;
	wire [4-1:0] node18447;
	wire [4-1:0] node18450;
	wire [4-1:0] node18451;
	wire [4-1:0] node18454;
	wire [4-1:0] node18457;
	wire [4-1:0] node18458;
	wire [4-1:0] node18460;
	wire [4-1:0] node18463;
	wire [4-1:0] node18464;
	wire [4-1:0] node18468;
	wire [4-1:0] node18469;
	wire [4-1:0] node18470;
	wire [4-1:0] node18473;
	wire [4-1:0] node18476;
	wire [4-1:0] node18477;
	wire [4-1:0] node18478;
	wire [4-1:0] node18481;
	wire [4-1:0] node18484;
	wire [4-1:0] node18485;
	wire [4-1:0] node18488;
	wire [4-1:0] node18491;
	wire [4-1:0] node18492;
	wire [4-1:0] node18493;
	wire [4-1:0] node18494;
	wire [4-1:0] node18495;
	wire [4-1:0] node18498;
	wire [4-1:0] node18501;
	wire [4-1:0] node18503;
	wire [4-1:0] node18506;
	wire [4-1:0] node18507;
	wire [4-1:0] node18508;
	wire [4-1:0] node18511;
	wire [4-1:0] node18514;
	wire [4-1:0] node18515;
	wire [4-1:0] node18519;
	wire [4-1:0] node18520;
	wire [4-1:0] node18521;
	wire [4-1:0] node18523;
	wire [4-1:0] node18526;
	wire [4-1:0] node18528;
	wire [4-1:0] node18531;
	wire [4-1:0] node18532;
	wire [4-1:0] node18534;
	wire [4-1:0] node18538;
	wire [4-1:0] node18539;
	wire [4-1:0] node18540;
	wire [4-1:0] node18541;
	wire [4-1:0] node18542;
	wire [4-1:0] node18543;
	wire [4-1:0] node18544;
	wire [4-1:0] node18547;
	wire [4-1:0] node18550;
	wire [4-1:0] node18551;
	wire [4-1:0] node18554;
	wire [4-1:0] node18557;
	wire [4-1:0] node18558;
	wire [4-1:0] node18559;
	wire [4-1:0] node18562;
	wire [4-1:0] node18565;
	wire [4-1:0] node18567;
	wire [4-1:0] node18570;
	wire [4-1:0] node18571;
	wire [4-1:0] node18572;
	wire [4-1:0] node18574;
	wire [4-1:0] node18577;
	wire [4-1:0] node18579;
	wire [4-1:0] node18582;
	wire [4-1:0] node18583;
	wire [4-1:0] node18584;
	wire [4-1:0] node18588;
	wire [4-1:0] node18590;
	wire [4-1:0] node18593;
	wire [4-1:0] node18594;
	wire [4-1:0] node18595;
	wire [4-1:0] node18596;
	wire [4-1:0] node18597;
	wire [4-1:0] node18600;
	wire [4-1:0] node18603;
	wire [4-1:0] node18604;
	wire [4-1:0] node18607;
	wire [4-1:0] node18610;
	wire [4-1:0] node18611;
	wire [4-1:0] node18612;
	wire [4-1:0] node18615;
	wire [4-1:0] node18618;
	wire [4-1:0] node18619;
	wire [4-1:0] node18622;
	wire [4-1:0] node18625;
	wire [4-1:0] node18626;
	wire [4-1:0] node18627;
	wire [4-1:0] node18630;
	wire [4-1:0] node18633;
	wire [4-1:0] node18634;
	wire [4-1:0] node18635;
	wire [4-1:0] node18638;
	wire [4-1:0] node18641;
	wire [4-1:0] node18643;
	wire [4-1:0] node18646;
	wire [4-1:0] node18647;
	wire [4-1:0] node18648;
	wire [4-1:0] node18649;
	wire [4-1:0] node18650;
	wire [4-1:0] node18651;
	wire [4-1:0] node18654;
	wire [4-1:0] node18657;
	wire [4-1:0] node18659;
	wire [4-1:0] node18662;
	wire [4-1:0] node18663;
	wire [4-1:0] node18665;
	wire [4-1:0] node18668;
	wire [4-1:0] node18669;
	wire [4-1:0] node18672;
	wire [4-1:0] node18675;
	wire [4-1:0] node18676;
	wire [4-1:0] node18677;
	wire [4-1:0] node18679;
	wire [4-1:0] node18682;
	wire [4-1:0] node18684;
	wire [4-1:0] node18687;
	wire [4-1:0] node18688;
	wire [4-1:0] node18690;
	wire [4-1:0] node18693;
	wire [4-1:0] node18695;
	wire [4-1:0] node18698;
	wire [4-1:0] node18699;
	wire [4-1:0] node18700;
	wire [4-1:0] node18701;
	wire [4-1:0] node18702;
	wire [4-1:0] node18705;
	wire [4-1:0] node18708;
	wire [4-1:0] node18709;
	wire [4-1:0] node18712;
	wire [4-1:0] node18715;
	wire [4-1:0] node18716;
	wire [4-1:0] node18718;
	wire [4-1:0] node18721;
	wire [4-1:0] node18722;
	wire [4-1:0] node18725;
	wire [4-1:0] node18728;
	wire [4-1:0] node18729;
	wire [4-1:0] node18730;
	wire [4-1:0] node18731;
	wire [4-1:0] node18734;
	wire [4-1:0] node18737;
	wire [4-1:0] node18738;
	wire [4-1:0] node18741;
	wire [4-1:0] node18744;
	wire [4-1:0] node18745;
	wire [4-1:0] node18746;
	wire [4-1:0] node18749;
	wire [4-1:0] node18752;
	wire [4-1:0] node18753;
	wire [4-1:0] node18756;
	wire [4-1:0] node18759;
	wire [4-1:0] node18760;
	wire [4-1:0] node18761;
	wire [4-1:0] node18762;
	wire [4-1:0] node18763;
	wire [4-1:0] node18764;
	wire [4-1:0] node18765;
	wire [4-1:0] node18766;
	wire [4-1:0] node18767;
	wire [4-1:0] node18771;
	wire [4-1:0] node18772;
	wire [4-1:0] node18776;
	wire [4-1:0] node18777;
	wire [4-1:0] node18778;
	wire [4-1:0] node18782;
	wire [4-1:0] node18783;
	wire [4-1:0] node18787;
	wire [4-1:0] node18788;
	wire [4-1:0] node18789;
	wire [4-1:0] node18790;
	wire [4-1:0] node18793;
	wire [4-1:0] node18796;
	wire [4-1:0] node18797;
	wire [4-1:0] node18800;
	wire [4-1:0] node18803;
	wire [4-1:0] node18804;
	wire [4-1:0] node18807;
	wire [4-1:0] node18808;
	wire [4-1:0] node18811;
	wire [4-1:0] node18814;
	wire [4-1:0] node18815;
	wire [4-1:0] node18816;
	wire [4-1:0] node18817;
	wire [4-1:0] node18818;
	wire [4-1:0] node18821;
	wire [4-1:0] node18824;
	wire [4-1:0] node18825;
	wire [4-1:0] node18828;
	wire [4-1:0] node18831;
	wire [4-1:0] node18832;
	wire [4-1:0] node18835;
	wire [4-1:0] node18838;
	wire [4-1:0] node18839;
	wire [4-1:0] node18840;
	wire [4-1:0] node18841;
	wire [4-1:0] node18844;
	wire [4-1:0] node18847;
	wire [4-1:0] node18848;
	wire [4-1:0] node18851;
	wire [4-1:0] node18854;
	wire [4-1:0] node18855;
	wire [4-1:0] node18856;
	wire [4-1:0] node18859;
	wire [4-1:0] node18862;
	wire [4-1:0] node18863;
	wire [4-1:0] node18866;
	wire [4-1:0] node18869;
	wire [4-1:0] node18870;
	wire [4-1:0] node18871;
	wire [4-1:0] node18872;
	wire [4-1:0] node18873;
	wire [4-1:0] node18874;
	wire [4-1:0] node18878;
	wire [4-1:0] node18879;
	wire [4-1:0] node18883;
	wire [4-1:0] node18884;
	wire [4-1:0] node18885;
	wire [4-1:0] node18889;
	wire [4-1:0] node18890;
	wire [4-1:0] node18894;
	wire [4-1:0] node18895;
	wire [4-1:0] node18896;
	wire [4-1:0] node18897;
	wire [4-1:0] node18900;
	wire [4-1:0] node18903;
	wire [4-1:0] node18904;
	wire [4-1:0] node18907;
	wire [4-1:0] node18910;
	wire [4-1:0] node18911;
	wire [4-1:0] node18912;
	wire [4-1:0] node18915;
	wire [4-1:0] node18918;
	wire [4-1:0] node18919;
	wire [4-1:0] node18922;
	wire [4-1:0] node18925;
	wire [4-1:0] node18926;
	wire [4-1:0] node18927;
	wire [4-1:0] node18928;
	wire [4-1:0] node18929;
	wire [4-1:0] node18932;
	wire [4-1:0] node18935;
	wire [4-1:0] node18936;
	wire [4-1:0] node18939;
	wire [4-1:0] node18942;
	wire [4-1:0] node18943;
	wire [4-1:0] node18945;
	wire [4-1:0] node18948;
	wire [4-1:0] node18949;
	wire [4-1:0] node18952;
	wire [4-1:0] node18955;
	wire [4-1:0] node18956;
	wire [4-1:0] node18957;
	wire [4-1:0] node18959;
	wire [4-1:0] node18962;
	wire [4-1:0] node18963;
	wire [4-1:0] node18967;
	wire [4-1:0] node18968;
	wire [4-1:0] node18969;
	wire [4-1:0] node18972;
	wire [4-1:0] node18975;
	wire [4-1:0] node18976;
	wire [4-1:0] node18979;
	wire [4-1:0] node18982;
	wire [4-1:0] node18983;
	wire [4-1:0] node18984;
	wire [4-1:0] node18985;
	wire [4-1:0] node18986;
	wire [4-1:0] node18987;
	wire [4-1:0] node18989;
	wire [4-1:0] node18992;
	wire [4-1:0] node18993;
	wire [4-1:0] node18996;
	wire [4-1:0] node18999;
	wire [4-1:0] node19000;
	wire [4-1:0] node19001;
	wire [4-1:0] node19004;
	wire [4-1:0] node19007;
	wire [4-1:0] node19008;
	wire [4-1:0] node19012;
	wire [4-1:0] node19013;
	wire [4-1:0] node19014;
	wire [4-1:0] node19017;
	wire [4-1:0] node19020;
	wire [4-1:0] node19021;
	wire [4-1:0] node19022;
	wire [4-1:0] node19025;
	wire [4-1:0] node19028;
	wire [4-1:0] node19029;
	wire [4-1:0] node19032;
	wire [4-1:0] node19035;
	wire [4-1:0] node19036;
	wire [4-1:0] node19037;
	wire [4-1:0] node19038;
	wire [4-1:0] node19039;
	wire [4-1:0] node19042;
	wire [4-1:0] node19045;
	wire [4-1:0] node19046;
	wire [4-1:0] node19049;
	wire [4-1:0] node19052;
	wire [4-1:0] node19053;
	wire [4-1:0] node19054;
	wire [4-1:0] node19057;
	wire [4-1:0] node19060;
	wire [4-1:0] node19061;
	wire [4-1:0] node19065;
	wire [4-1:0] node19066;
	wire [4-1:0] node19067;
	wire [4-1:0] node19068;
	wire [4-1:0] node19072;
	wire [4-1:0] node19073;
	wire [4-1:0] node19077;
	wire [4-1:0] node19078;
	wire [4-1:0] node19079;
	wire [4-1:0] node19083;
	wire [4-1:0] node19084;
	wire [4-1:0] node19088;
	wire [4-1:0] node19089;
	wire [4-1:0] node19090;
	wire [4-1:0] node19091;
	wire [4-1:0] node19092;
	wire [4-1:0] node19093;
	wire [4-1:0] node19096;
	wire [4-1:0] node19099;
	wire [4-1:0] node19100;
	wire [4-1:0] node19103;
	wire [4-1:0] node19106;
	wire [4-1:0] node19107;
	wire [4-1:0] node19108;
	wire [4-1:0] node19111;
	wire [4-1:0] node19114;
	wire [4-1:0] node19115;
	wire [4-1:0] node19118;
	wire [4-1:0] node19121;
	wire [4-1:0] node19122;
	wire [4-1:0] node19123;
	wire [4-1:0] node19124;
	wire [4-1:0] node19127;
	wire [4-1:0] node19130;
	wire [4-1:0] node19131;
	wire [4-1:0] node19134;
	wire [4-1:0] node19137;
	wire [4-1:0] node19138;
	wire [4-1:0] node19141;
	wire [4-1:0] node19144;
	wire [4-1:0] node19145;
	wire [4-1:0] node19146;
	wire [4-1:0] node19147;
	wire [4-1:0] node19148;
	wire [4-1:0] node19151;
	wire [4-1:0] node19154;
	wire [4-1:0] node19155;
	wire [4-1:0] node19158;
	wire [4-1:0] node19161;
	wire [4-1:0] node19162;
	wire [4-1:0] node19164;
	wire [4-1:0] node19167;
	wire [4-1:0] node19168;
	wire [4-1:0] node19171;
	wire [4-1:0] node19174;
	wire [4-1:0] node19175;
	wire [4-1:0] node19176;
	wire [4-1:0] node19177;
	wire [4-1:0] node19180;
	wire [4-1:0] node19183;
	wire [4-1:0] node19184;
	wire [4-1:0] node19187;
	wire [4-1:0] node19190;
	wire [4-1:0] node19191;
	wire [4-1:0] node19193;
	wire [4-1:0] node19196;
	wire [4-1:0] node19197;
	wire [4-1:0] node19200;
	wire [4-1:0] node19203;
	wire [4-1:0] node19204;
	wire [4-1:0] node19205;
	wire [4-1:0] node19206;
	wire [4-1:0] node19207;
	wire [4-1:0] node19208;
	wire [4-1:0] node19209;
	wire [4-1:0] node19210;
	wire [4-1:0] node19213;
	wire [4-1:0] node19216;
	wire [4-1:0] node19217;
	wire [4-1:0] node19220;
	wire [4-1:0] node19223;
	wire [4-1:0] node19225;
	wire [4-1:0] node19226;
	wire [4-1:0] node19229;
	wire [4-1:0] node19232;
	wire [4-1:0] node19233;
	wire [4-1:0] node19234;
	wire [4-1:0] node19235;
	wire [4-1:0] node19238;
	wire [4-1:0] node19241;
	wire [4-1:0] node19242;
	wire [4-1:0] node19245;
	wire [4-1:0] node19248;
	wire [4-1:0] node19249;
	wire [4-1:0] node19250;
	wire [4-1:0] node19253;
	wire [4-1:0] node19256;
	wire [4-1:0] node19257;
	wire [4-1:0] node19260;
	wire [4-1:0] node19263;
	wire [4-1:0] node19264;
	wire [4-1:0] node19265;
	wire [4-1:0] node19266;
	wire [4-1:0] node19267;
	wire [4-1:0] node19270;
	wire [4-1:0] node19273;
	wire [4-1:0] node19274;
	wire [4-1:0] node19277;
	wire [4-1:0] node19280;
	wire [4-1:0] node19281;
	wire [4-1:0] node19283;
	wire [4-1:0] node19286;
	wire [4-1:0] node19287;
	wire [4-1:0] node19290;
	wire [4-1:0] node19293;
	wire [4-1:0] node19294;
	wire [4-1:0] node19295;
	wire [4-1:0] node19296;
	wire [4-1:0] node19299;
	wire [4-1:0] node19302;
	wire [4-1:0] node19303;
	wire [4-1:0] node19306;
	wire [4-1:0] node19309;
	wire [4-1:0] node19310;
	wire [4-1:0] node19311;
	wire [4-1:0] node19315;
	wire [4-1:0] node19316;
	wire [4-1:0] node19319;
	wire [4-1:0] node19322;
	wire [4-1:0] node19323;
	wire [4-1:0] node19324;
	wire [4-1:0] node19325;
	wire [4-1:0] node19326;
	wire [4-1:0] node19327;
	wire [4-1:0] node19330;
	wire [4-1:0] node19333;
	wire [4-1:0] node19334;
	wire [4-1:0] node19337;
	wire [4-1:0] node19340;
	wire [4-1:0] node19341;
	wire [4-1:0] node19343;
	wire [4-1:0] node19346;
	wire [4-1:0] node19347;
	wire [4-1:0] node19350;
	wire [4-1:0] node19353;
	wire [4-1:0] node19354;
	wire [4-1:0] node19355;
	wire [4-1:0] node19356;
	wire [4-1:0] node19359;
	wire [4-1:0] node19362;
	wire [4-1:0] node19363;
	wire [4-1:0] node19366;
	wire [4-1:0] node19369;
	wire [4-1:0] node19370;
	wire [4-1:0] node19371;
	wire [4-1:0] node19374;
	wire [4-1:0] node19377;
	wire [4-1:0] node19378;
	wire [4-1:0] node19381;
	wire [4-1:0] node19384;
	wire [4-1:0] node19385;
	wire [4-1:0] node19386;
	wire [4-1:0] node19387;
	wire [4-1:0] node19388;
	wire [4-1:0] node19391;
	wire [4-1:0] node19394;
	wire [4-1:0] node19395;
	wire [4-1:0] node19398;
	wire [4-1:0] node19401;
	wire [4-1:0] node19402;
	wire [4-1:0] node19403;
	wire [4-1:0] node19406;
	wire [4-1:0] node19409;
	wire [4-1:0] node19410;
	wire [4-1:0] node19413;
	wire [4-1:0] node19416;
	wire [4-1:0] node19417;
	wire [4-1:0] node19418;
	wire [4-1:0] node19419;
	wire [4-1:0] node19422;
	wire [4-1:0] node19425;
	wire [4-1:0] node19426;
	wire [4-1:0] node19429;
	wire [4-1:0] node19432;
	wire [4-1:0] node19433;
	wire [4-1:0] node19434;
	wire [4-1:0] node19438;
	wire [4-1:0] node19441;
	wire [4-1:0] node19442;
	wire [4-1:0] node19443;
	wire [4-1:0] node19444;
	wire [4-1:0] node19445;
	wire [4-1:0] node19446;
	wire [4-1:0] node19447;
	wire [4-1:0] node19451;
	wire [4-1:0] node19452;
	wire [4-1:0] node19455;
	wire [4-1:0] node19458;
	wire [4-1:0] node19459;
	wire [4-1:0] node19460;
	wire [4-1:0] node19463;
	wire [4-1:0] node19466;
	wire [4-1:0] node19467;
	wire [4-1:0] node19470;
	wire [4-1:0] node19473;
	wire [4-1:0] node19474;
	wire [4-1:0] node19475;
	wire [4-1:0] node19476;
	wire [4-1:0] node19479;
	wire [4-1:0] node19482;
	wire [4-1:0] node19483;
	wire [4-1:0] node19486;
	wire [4-1:0] node19489;
	wire [4-1:0] node19490;
	wire [4-1:0] node19493;
	wire [4-1:0] node19496;
	wire [4-1:0] node19497;
	wire [4-1:0] node19498;
	wire [4-1:0] node19499;
	wire [4-1:0] node19500;
	wire [4-1:0] node19503;
	wire [4-1:0] node19506;
	wire [4-1:0] node19507;
	wire [4-1:0] node19510;
	wire [4-1:0] node19513;
	wire [4-1:0] node19514;
	wire [4-1:0] node19515;
	wire [4-1:0] node19518;
	wire [4-1:0] node19521;
	wire [4-1:0] node19522;
	wire [4-1:0] node19526;
	wire [4-1:0] node19527;
	wire [4-1:0] node19528;
	wire [4-1:0] node19529;
	wire [4-1:0] node19532;
	wire [4-1:0] node19535;
	wire [4-1:0] node19536;
	wire [4-1:0] node19539;
	wire [4-1:0] node19542;
	wire [4-1:0] node19543;
	wire [4-1:0] node19544;
	wire [4-1:0] node19547;
	wire [4-1:0] node19550;
	wire [4-1:0] node19551;
	wire [4-1:0] node19554;
	wire [4-1:0] node19557;
	wire [4-1:0] node19558;
	wire [4-1:0] node19559;
	wire [4-1:0] node19560;
	wire [4-1:0] node19561;
	wire [4-1:0] node19563;
	wire [4-1:0] node19566;
	wire [4-1:0] node19567;
	wire [4-1:0] node19570;
	wire [4-1:0] node19573;
	wire [4-1:0] node19574;
	wire [4-1:0] node19575;
	wire [4-1:0] node19579;
	wire [4-1:0] node19580;
	wire [4-1:0] node19583;
	wire [4-1:0] node19586;
	wire [4-1:0] node19587;
	wire [4-1:0] node19588;
	wire [4-1:0] node19589;
	wire [4-1:0] node19592;
	wire [4-1:0] node19595;
	wire [4-1:0] node19596;
	wire [4-1:0] node19599;
	wire [4-1:0] node19602;
	wire [4-1:0] node19603;
	wire [4-1:0] node19604;
	wire [4-1:0] node19607;
	wire [4-1:0] node19610;
	wire [4-1:0] node19611;
	wire [4-1:0] node19614;
	wire [4-1:0] node19617;
	wire [4-1:0] node19618;
	wire [4-1:0] node19619;
	wire [4-1:0] node19620;
	wire [4-1:0] node19621;
	wire [4-1:0] node19624;
	wire [4-1:0] node19627;
	wire [4-1:0] node19628;
	wire [4-1:0] node19631;
	wire [4-1:0] node19634;
	wire [4-1:0] node19635;
	wire [4-1:0] node19638;
	wire [4-1:0] node19639;
	wire [4-1:0] node19642;
	wire [4-1:0] node19645;
	wire [4-1:0] node19646;
	wire [4-1:0] node19647;
	wire [4-1:0] node19648;
	wire [4-1:0] node19651;
	wire [4-1:0] node19654;
	wire [4-1:0] node19655;
	wire [4-1:0] node19658;
	wire [4-1:0] node19661;
	wire [4-1:0] node19662;
	wire [4-1:0] node19663;
	wire [4-1:0] node19666;
	wire [4-1:0] node19669;
	wire [4-1:0] node19670;
	wire [4-1:0] node19673;
	wire [4-1:0] node19676;
	wire [4-1:0] node19677;
	wire [4-1:0] node19678;
	wire [4-1:0] node19679;
	wire [4-1:0] node19680;
	wire [4-1:0] node19681;
	wire [4-1:0] node19682;
	wire [4-1:0] node19683;
	wire [4-1:0] node19684;
	wire [4-1:0] node19685;
	wire [4-1:0] node19688;
	wire [4-1:0] node19691;
	wire [4-1:0] node19693;
	wire [4-1:0] node19696;
	wire [4-1:0] node19697;
	wire [4-1:0] node19698;
	wire [4-1:0] node19701;
	wire [4-1:0] node19704;
	wire [4-1:0] node19705;
	wire [4-1:0] node19708;
	wire [4-1:0] node19711;
	wire [4-1:0] node19712;
	wire [4-1:0] node19713;
	wire [4-1:0] node19714;
	wire [4-1:0] node19717;
	wire [4-1:0] node19720;
	wire [4-1:0] node19721;
	wire [4-1:0] node19724;
	wire [4-1:0] node19727;
	wire [4-1:0] node19728;
	wire [4-1:0] node19729;
	wire [4-1:0] node19732;
	wire [4-1:0] node19735;
	wire [4-1:0] node19736;
	wire [4-1:0] node19739;
	wire [4-1:0] node19742;
	wire [4-1:0] node19743;
	wire [4-1:0] node19744;
	wire [4-1:0] node19745;
	wire [4-1:0] node19746;
	wire [4-1:0] node19749;
	wire [4-1:0] node19752;
	wire [4-1:0] node19753;
	wire [4-1:0] node19756;
	wire [4-1:0] node19759;
	wire [4-1:0] node19760;
	wire [4-1:0] node19761;
	wire [4-1:0] node19764;
	wire [4-1:0] node19767;
	wire [4-1:0] node19768;
	wire [4-1:0] node19771;
	wire [4-1:0] node19774;
	wire [4-1:0] node19775;
	wire [4-1:0] node19776;
	wire [4-1:0] node19777;
	wire [4-1:0] node19780;
	wire [4-1:0] node19783;
	wire [4-1:0] node19784;
	wire [4-1:0] node19788;
	wire [4-1:0] node19789;
	wire [4-1:0] node19790;
	wire [4-1:0] node19793;
	wire [4-1:0] node19796;
	wire [4-1:0] node19797;
	wire [4-1:0] node19800;
	wire [4-1:0] node19803;
	wire [4-1:0] node19804;
	wire [4-1:0] node19805;
	wire [4-1:0] node19806;
	wire [4-1:0] node19807;
	wire [4-1:0] node19808;
	wire [4-1:0] node19812;
	wire [4-1:0] node19813;
	wire [4-1:0] node19816;
	wire [4-1:0] node19819;
	wire [4-1:0] node19820;
	wire [4-1:0] node19821;
	wire [4-1:0] node19824;
	wire [4-1:0] node19827;
	wire [4-1:0] node19829;
	wire [4-1:0] node19832;
	wire [4-1:0] node19833;
	wire [4-1:0] node19834;
	wire [4-1:0] node19835;
	wire [4-1:0] node19838;
	wire [4-1:0] node19841;
	wire [4-1:0] node19842;
	wire [4-1:0] node19845;
	wire [4-1:0] node19848;
	wire [4-1:0] node19849;
	wire [4-1:0] node19850;
	wire [4-1:0] node19853;
	wire [4-1:0] node19856;
	wire [4-1:0] node19857;
	wire [4-1:0] node19860;
	wire [4-1:0] node19863;
	wire [4-1:0] node19864;
	wire [4-1:0] node19865;
	wire [4-1:0] node19866;
	wire [4-1:0] node19867;
	wire [4-1:0] node19870;
	wire [4-1:0] node19873;
	wire [4-1:0] node19874;
	wire [4-1:0] node19877;
	wire [4-1:0] node19880;
	wire [4-1:0] node19881;
	wire [4-1:0] node19882;
	wire [4-1:0] node19885;
	wire [4-1:0] node19888;
	wire [4-1:0] node19889;
	wire [4-1:0] node19892;
	wire [4-1:0] node19895;
	wire [4-1:0] node19896;
	wire [4-1:0] node19897;
	wire [4-1:0] node19898;
	wire [4-1:0] node19901;
	wire [4-1:0] node19904;
	wire [4-1:0] node19905;
	wire [4-1:0] node19909;
	wire [4-1:0] node19910;
	wire [4-1:0] node19911;
	wire [4-1:0] node19914;
	wire [4-1:0] node19917;
	wire [4-1:0] node19918;
	wire [4-1:0] node19921;
	wire [4-1:0] node19924;
	wire [4-1:0] node19925;
	wire [4-1:0] node19926;
	wire [4-1:0] node19927;
	wire [4-1:0] node19928;
	wire [4-1:0] node19929;
	wire [4-1:0] node19930;
	wire [4-1:0] node19933;
	wire [4-1:0] node19936;
	wire [4-1:0] node19937;
	wire [4-1:0] node19940;
	wire [4-1:0] node19943;
	wire [4-1:0] node19944;
	wire [4-1:0] node19945;
	wire [4-1:0] node19948;
	wire [4-1:0] node19951;
	wire [4-1:0] node19953;
	wire [4-1:0] node19956;
	wire [4-1:0] node19957;
	wire [4-1:0] node19958;
	wire [4-1:0] node19960;
	wire [4-1:0] node19963;
	wire [4-1:0] node19965;
	wire [4-1:0] node19968;
	wire [4-1:0] node19969;
	wire [4-1:0] node19971;
	wire [4-1:0] node19974;
	wire [4-1:0] node19977;
	wire [4-1:0] node19978;
	wire [4-1:0] node19979;
	wire [4-1:0] node19980;
	wire [4-1:0] node19982;
	wire [4-1:0] node19985;
	wire [4-1:0] node19986;
	wire [4-1:0] node19989;
	wire [4-1:0] node19992;
	wire [4-1:0] node19993;
	wire [4-1:0] node19995;
	wire [4-1:0] node19998;
	wire [4-1:0] node19999;
	wire [4-1:0] node20002;
	wire [4-1:0] node20005;
	wire [4-1:0] node20006;
	wire [4-1:0] node20007;
	wire [4-1:0] node20008;
	wire [4-1:0] node20011;
	wire [4-1:0] node20014;
	wire [4-1:0] node20015;
	wire [4-1:0] node20018;
	wire [4-1:0] node20021;
	wire [4-1:0] node20022;
	wire [4-1:0] node20024;
	wire [4-1:0] node20027;
	wire [4-1:0] node20028;
	wire [4-1:0] node20031;
	wire [4-1:0] node20034;
	wire [4-1:0] node20035;
	wire [4-1:0] node20036;
	wire [4-1:0] node20037;
	wire [4-1:0] node20038;
	wire [4-1:0] node20039;
	wire [4-1:0] node20043;
	wire [4-1:0] node20044;
	wire [4-1:0] node20048;
	wire [4-1:0] node20049;
	wire [4-1:0] node20050;
	wire [4-1:0] node20053;
	wire [4-1:0] node20056;
	wire [4-1:0] node20057;
	wire [4-1:0] node20061;
	wire [4-1:0] node20062;
	wire [4-1:0] node20063;
	wire [4-1:0] node20064;
	wire [4-1:0] node20067;
	wire [4-1:0] node20070;
	wire [4-1:0] node20071;
	wire [4-1:0] node20075;
	wire [4-1:0] node20076;
	wire [4-1:0] node20077;
	wire [4-1:0] node20080;
	wire [4-1:0] node20083;
	wire [4-1:0] node20084;
	wire [4-1:0] node20087;
	wire [4-1:0] node20090;
	wire [4-1:0] node20091;
	wire [4-1:0] node20092;
	wire [4-1:0] node20093;
	wire [4-1:0] node20095;
	wire [4-1:0] node20098;
	wire [4-1:0] node20099;
	wire [4-1:0] node20102;
	wire [4-1:0] node20105;
	wire [4-1:0] node20106;
	wire [4-1:0] node20107;
	wire [4-1:0] node20110;
	wire [4-1:0] node20113;
	wire [4-1:0] node20114;
	wire [4-1:0] node20118;
	wire [4-1:0] node20119;
	wire [4-1:0] node20120;
	wire [4-1:0] node20121;
	wire [4-1:0] node20125;
	wire [4-1:0] node20126;
	wire [4-1:0] node20130;
	wire [4-1:0] node20131;
	wire [4-1:0] node20132;
	wire [4-1:0] node20136;
	wire [4-1:0] node20137;
	wire [4-1:0] node20141;
	wire [4-1:0] node20142;
	wire [4-1:0] node20143;
	wire [4-1:0] node20144;
	wire [4-1:0] node20145;
	wire [4-1:0] node20146;
	wire [4-1:0] node20147;
	wire [4-1:0] node20148;
	wire [4-1:0] node20151;
	wire [4-1:0] node20154;
	wire [4-1:0] node20155;
	wire [4-1:0] node20158;
	wire [4-1:0] node20161;
	wire [4-1:0] node20162;
	wire [4-1:0] node20163;
	wire [4-1:0] node20166;
	wire [4-1:0] node20169;
	wire [4-1:0] node20171;
	wire [4-1:0] node20174;
	wire [4-1:0] node20175;
	wire [4-1:0] node20176;
	wire [4-1:0] node20178;
	wire [4-1:0] node20181;
	wire [4-1:0] node20183;
	wire [4-1:0] node20186;
	wire [4-1:0] node20187;
	wire [4-1:0] node20189;
	wire [4-1:0] node20192;
	wire [4-1:0] node20194;
	wire [4-1:0] node20197;
	wire [4-1:0] node20198;
	wire [4-1:0] node20199;
	wire [4-1:0] node20200;
	wire [4-1:0] node20201;
	wire [4-1:0] node20204;
	wire [4-1:0] node20207;
	wire [4-1:0] node20208;
	wire [4-1:0] node20211;
	wire [4-1:0] node20214;
	wire [4-1:0] node20215;
	wire [4-1:0] node20218;
	wire [4-1:0] node20220;
	wire [4-1:0] node20223;
	wire [4-1:0] node20224;
	wire [4-1:0] node20225;
	wire [4-1:0] node20226;
	wire [4-1:0] node20229;
	wire [4-1:0] node20232;
	wire [4-1:0] node20233;
	wire [4-1:0] node20236;
	wire [4-1:0] node20239;
	wire [4-1:0] node20240;
	wire [4-1:0] node20241;
	wire [4-1:0] node20244;
	wire [4-1:0] node20247;
	wire [4-1:0] node20248;
	wire [4-1:0] node20251;
	wire [4-1:0] node20254;
	wire [4-1:0] node20255;
	wire [4-1:0] node20256;
	wire [4-1:0] node20257;
	wire [4-1:0] node20258;
	wire [4-1:0] node20259;
	wire [4-1:0] node20262;
	wire [4-1:0] node20265;
	wire [4-1:0] node20266;
	wire [4-1:0] node20269;
	wire [4-1:0] node20272;
	wire [4-1:0] node20273;
	wire [4-1:0] node20274;
	wire [4-1:0] node20277;
	wire [4-1:0] node20280;
	wire [4-1:0] node20281;
	wire [4-1:0] node20285;
	wire [4-1:0] node20286;
	wire [4-1:0] node20287;
	wire [4-1:0] node20288;
	wire [4-1:0] node20292;
	wire [4-1:0] node20293;
	wire [4-1:0] node20297;
	wire [4-1:0] node20298;
	wire [4-1:0] node20299;
	wire [4-1:0] node20303;
	wire [4-1:0] node20304;
	wire [4-1:0] node20308;
	wire [4-1:0] node20309;
	wire [4-1:0] node20310;
	wire [4-1:0] node20311;
	wire [4-1:0] node20312;
	wire [4-1:0] node20316;
	wire [4-1:0] node20317;
	wire [4-1:0] node20320;
	wire [4-1:0] node20323;
	wire [4-1:0] node20324;
	wire [4-1:0] node20325;
	wire [4-1:0] node20328;
	wire [4-1:0] node20331;
	wire [4-1:0] node20332;
	wire [4-1:0] node20335;
	wire [4-1:0] node20338;
	wire [4-1:0] node20339;
	wire [4-1:0] node20340;
	wire [4-1:0] node20341;
	wire [4-1:0] node20345;
	wire [4-1:0] node20346;
	wire [4-1:0] node20350;
	wire [4-1:0] node20351;
	wire [4-1:0] node20352;
	wire [4-1:0] node20356;
	wire [4-1:0] node20357;
	wire [4-1:0] node20361;
	wire [4-1:0] node20362;
	wire [4-1:0] node20363;
	wire [4-1:0] node20364;
	wire [4-1:0] node20365;
	wire [4-1:0] node20366;
	wire [4-1:0] node20367;
	wire [4-1:0] node20370;
	wire [4-1:0] node20373;
	wire [4-1:0] node20374;
	wire [4-1:0] node20378;
	wire [4-1:0] node20379;
	wire [4-1:0] node20380;
	wire [4-1:0] node20383;
	wire [4-1:0] node20386;
	wire [4-1:0] node20387;
	wire [4-1:0] node20391;
	wire [4-1:0] node20392;
	wire [4-1:0] node20393;
	wire [4-1:0] node20394;
	wire [4-1:0] node20398;
	wire [4-1:0] node20399;
	wire [4-1:0] node20403;
	wire [4-1:0] node20404;
	wire [4-1:0] node20405;
	wire [4-1:0] node20409;
	wire [4-1:0] node20410;
	wire [4-1:0] node20414;
	wire [4-1:0] node20415;
	wire [4-1:0] node20416;
	wire [4-1:0] node20417;
	wire [4-1:0] node20418;
	wire [4-1:0] node20422;
	wire [4-1:0] node20423;
	wire [4-1:0] node20426;
	wire [4-1:0] node20429;
	wire [4-1:0] node20430;
	wire [4-1:0] node20431;
	wire [4-1:0] node20435;
	wire [4-1:0] node20437;
	wire [4-1:0] node20440;
	wire [4-1:0] node20441;
	wire [4-1:0] node20442;
	wire [4-1:0] node20443;
	wire [4-1:0] node20447;
	wire [4-1:0] node20448;
	wire [4-1:0] node20452;
	wire [4-1:0] node20453;
	wire [4-1:0] node20454;
	wire [4-1:0] node20458;
	wire [4-1:0] node20459;
	wire [4-1:0] node20463;
	wire [4-1:0] node20464;
	wire [4-1:0] node20465;
	wire [4-1:0] node20466;
	wire [4-1:0] node20467;
	wire [4-1:0] node20468;
	wire [4-1:0] node20472;
	wire [4-1:0] node20473;
	wire [4-1:0] node20476;
	wire [4-1:0] node20479;
	wire [4-1:0] node20480;
	wire [4-1:0] node20481;
	wire [4-1:0] node20484;
	wire [4-1:0] node20487;
	wire [4-1:0] node20488;
	wire [4-1:0] node20491;
	wire [4-1:0] node20494;
	wire [4-1:0] node20495;
	wire [4-1:0] node20496;
	wire [4-1:0] node20497;
	wire [4-1:0] node20500;
	wire [4-1:0] node20503;
	wire [4-1:0] node20504;
	wire [4-1:0] node20507;
	wire [4-1:0] node20510;
	wire [4-1:0] node20511;
	wire [4-1:0] node20512;
	wire [4-1:0] node20515;
	wire [4-1:0] node20518;
	wire [4-1:0] node20519;
	wire [4-1:0] node20522;
	wire [4-1:0] node20525;
	wire [4-1:0] node20526;
	wire [4-1:0] node20527;
	wire [4-1:0] node20528;
	wire [4-1:0] node20529;
	wire [4-1:0] node20532;
	wire [4-1:0] node20535;
	wire [4-1:0] node20536;
	wire [4-1:0] node20539;
	wire [4-1:0] node20542;
	wire [4-1:0] node20543;
	wire [4-1:0] node20544;
	wire [4-1:0] node20547;
	wire [4-1:0] node20550;
	wire [4-1:0] node20551;
	wire [4-1:0] node20555;
	wire [4-1:0] node20556;
	wire [4-1:0] node20557;
	wire [4-1:0] node20558;
	wire [4-1:0] node20561;
	wire [4-1:0] node20564;
	wire [4-1:0] node20565;
	wire [4-1:0] node20568;
	wire [4-1:0] node20571;
	wire [4-1:0] node20572;
	wire [4-1:0] node20573;
	wire [4-1:0] node20576;
	wire [4-1:0] node20579;
	wire [4-1:0] node20580;
	wire [4-1:0] node20584;
	wire [4-1:0] node20585;
	wire [4-1:0] node20586;
	wire [4-1:0] node20587;
	wire [4-1:0] node20588;
	wire [4-1:0] node20589;
	wire [4-1:0] node20590;
	wire [4-1:0] node20591;
	wire [4-1:0] node20592;
	wire [4-1:0] node20595;
	wire [4-1:0] node20598;
	wire [4-1:0] node20599;
	wire [4-1:0] node20602;
	wire [4-1:0] node20605;
	wire [4-1:0] node20606;
	wire [4-1:0] node20607;
	wire [4-1:0] node20610;
	wire [4-1:0] node20613;
	wire [4-1:0] node20614;
	wire [4-1:0] node20617;
	wire [4-1:0] node20620;
	wire [4-1:0] node20621;
	wire [4-1:0] node20622;
	wire [4-1:0] node20623;
	wire [4-1:0] node20626;
	wire [4-1:0] node20629;
	wire [4-1:0] node20630;
	wire [4-1:0] node20633;
	wire [4-1:0] node20636;
	wire [4-1:0] node20637;
	wire [4-1:0] node20638;
	wire [4-1:0] node20641;
	wire [4-1:0] node20644;
	wire [4-1:0] node20645;
	wire [4-1:0] node20648;
	wire [4-1:0] node20651;
	wire [4-1:0] node20652;
	wire [4-1:0] node20653;
	wire [4-1:0] node20654;
	wire [4-1:0] node20655;
	wire [4-1:0] node20658;
	wire [4-1:0] node20661;
	wire [4-1:0] node20662;
	wire [4-1:0] node20665;
	wire [4-1:0] node20668;
	wire [4-1:0] node20669;
	wire [4-1:0] node20670;
	wire [4-1:0] node20673;
	wire [4-1:0] node20676;
	wire [4-1:0] node20677;
	wire [4-1:0] node20680;
	wire [4-1:0] node20683;
	wire [4-1:0] node20684;
	wire [4-1:0] node20685;
	wire [4-1:0] node20686;
	wire [4-1:0] node20689;
	wire [4-1:0] node20692;
	wire [4-1:0] node20693;
	wire [4-1:0] node20696;
	wire [4-1:0] node20699;
	wire [4-1:0] node20700;
	wire [4-1:0] node20702;
	wire [4-1:0] node20705;
	wire [4-1:0] node20706;
	wire [4-1:0] node20709;
	wire [4-1:0] node20712;
	wire [4-1:0] node20713;
	wire [4-1:0] node20714;
	wire [4-1:0] node20715;
	wire [4-1:0] node20716;
	wire [4-1:0] node20717;
	wire [4-1:0] node20720;
	wire [4-1:0] node20723;
	wire [4-1:0] node20724;
	wire [4-1:0] node20728;
	wire [4-1:0] node20729;
	wire [4-1:0] node20732;
	wire [4-1:0] node20735;
	wire [4-1:0] node20736;
	wire [4-1:0] node20737;
	wire [4-1:0] node20738;
	wire [4-1:0] node20741;
	wire [4-1:0] node20744;
	wire [4-1:0] node20745;
	wire [4-1:0] node20748;
	wire [4-1:0] node20751;
	wire [4-1:0] node20752;
	wire [4-1:0] node20753;
	wire [4-1:0] node20756;
	wire [4-1:0] node20759;
	wire [4-1:0] node20760;
	wire [4-1:0] node20763;
	wire [4-1:0] node20766;
	wire [4-1:0] node20767;
	wire [4-1:0] node20768;
	wire [4-1:0] node20769;
	wire [4-1:0] node20770;
	wire [4-1:0] node20774;
	wire [4-1:0] node20775;
	wire [4-1:0] node20779;
	wire [4-1:0] node20780;
	wire [4-1:0] node20781;
	wire [4-1:0] node20785;
	wire [4-1:0] node20786;
	wire [4-1:0] node20790;
	wire [4-1:0] node20791;
	wire [4-1:0] node20792;
	wire [4-1:0] node20793;
	wire [4-1:0] node20796;
	wire [4-1:0] node20799;
	wire [4-1:0] node20800;
	wire [4-1:0] node20803;
	wire [4-1:0] node20806;
	wire [4-1:0] node20807;
	wire [4-1:0] node20808;
	wire [4-1:0] node20811;
	wire [4-1:0] node20814;
	wire [4-1:0] node20815;
	wire [4-1:0] node20818;
	wire [4-1:0] node20821;
	wire [4-1:0] node20822;
	wire [4-1:0] node20823;
	wire [4-1:0] node20824;
	wire [4-1:0] node20825;
	wire [4-1:0] node20826;
	wire [4-1:0] node20827;
	wire [4-1:0] node20830;
	wire [4-1:0] node20833;
	wire [4-1:0] node20835;
	wire [4-1:0] node20838;
	wire [4-1:0] node20839;
	wire [4-1:0] node20840;
	wire [4-1:0] node20844;
	wire [4-1:0] node20845;
	wire [4-1:0] node20848;
	wire [4-1:0] node20851;
	wire [4-1:0] node20852;
	wire [4-1:0] node20853;
	wire [4-1:0] node20854;
	wire [4-1:0] node20857;
	wire [4-1:0] node20860;
	wire [4-1:0] node20862;
	wire [4-1:0] node20865;
	wire [4-1:0] node20866;
	wire [4-1:0] node20867;
	wire [4-1:0] node20870;
	wire [4-1:0] node20873;
	wire [4-1:0] node20874;
	wire [4-1:0] node20877;
	wire [4-1:0] node20880;
	wire [4-1:0] node20881;
	wire [4-1:0] node20882;
	wire [4-1:0] node20883;
	wire [4-1:0] node20884;
	wire [4-1:0] node20887;
	wire [4-1:0] node20890;
	wire [4-1:0] node20891;
	wire [4-1:0] node20894;
	wire [4-1:0] node20897;
	wire [4-1:0] node20898;
	wire [4-1:0] node20899;
	wire [4-1:0] node20902;
	wire [4-1:0] node20905;
	wire [4-1:0] node20906;
	wire [4-1:0] node20910;
	wire [4-1:0] node20911;
	wire [4-1:0] node20912;
	wire [4-1:0] node20913;
	wire [4-1:0] node20916;
	wire [4-1:0] node20919;
	wire [4-1:0] node20920;
	wire [4-1:0] node20924;
	wire [4-1:0] node20925;
	wire [4-1:0] node20926;
	wire [4-1:0] node20929;
	wire [4-1:0] node20932;
	wire [4-1:0] node20933;
	wire [4-1:0] node20936;
	wire [4-1:0] node20939;
	wire [4-1:0] node20940;
	wire [4-1:0] node20941;
	wire [4-1:0] node20942;
	wire [4-1:0] node20943;
	wire [4-1:0] node20944;
	wire [4-1:0] node20947;
	wire [4-1:0] node20950;
	wire [4-1:0] node20951;
	wire [4-1:0] node20954;
	wire [4-1:0] node20957;
	wire [4-1:0] node20958;
	wire [4-1:0] node20959;
	wire [4-1:0] node20963;
	wire [4-1:0] node20964;
	wire [4-1:0] node20967;
	wire [4-1:0] node20970;
	wire [4-1:0] node20971;
	wire [4-1:0] node20972;
	wire [4-1:0] node20973;
	wire [4-1:0] node20976;
	wire [4-1:0] node20979;
	wire [4-1:0] node20980;
	wire [4-1:0] node20984;
	wire [4-1:0] node20985;
	wire [4-1:0] node20988;
	wire [4-1:0] node20991;
	wire [4-1:0] node20992;
	wire [4-1:0] node20993;
	wire [4-1:0] node20994;
	wire [4-1:0] node20995;
	wire [4-1:0] node20998;
	wire [4-1:0] node21001;
	wire [4-1:0] node21003;
	wire [4-1:0] node21006;
	wire [4-1:0] node21007;
	wire [4-1:0] node21009;
	wire [4-1:0] node21012;
	wire [4-1:0] node21013;
	wire [4-1:0] node21016;
	wire [4-1:0] node21019;
	wire [4-1:0] node21020;
	wire [4-1:0] node21021;
	wire [4-1:0] node21022;
	wire [4-1:0] node21025;
	wire [4-1:0] node21028;
	wire [4-1:0] node21030;
	wire [4-1:0] node21033;
	wire [4-1:0] node21034;
	wire [4-1:0] node21037;
	wire [4-1:0] node21040;
	wire [4-1:0] node21041;
	wire [4-1:0] node21042;
	wire [4-1:0] node21043;
	wire [4-1:0] node21044;
	wire [4-1:0] node21045;
	wire [4-1:0] node21046;
	wire [4-1:0] node21047;
	wire [4-1:0] node21050;
	wire [4-1:0] node21053;
	wire [4-1:0] node21054;
	wire [4-1:0] node21058;
	wire [4-1:0] node21059;
	wire [4-1:0] node21060;
	wire [4-1:0] node21064;
	wire [4-1:0] node21065;
	wire [4-1:0] node21069;
	wire [4-1:0] node21070;
	wire [4-1:0] node21071;
	wire [4-1:0] node21072;
	wire [4-1:0] node21075;
	wire [4-1:0] node21078;
	wire [4-1:0] node21079;
	wire [4-1:0] node21082;
	wire [4-1:0] node21085;
	wire [4-1:0] node21086;
	wire [4-1:0] node21087;
	wire [4-1:0] node21090;
	wire [4-1:0] node21093;
	wire [4-1:0] node21094;
	wire [4-1:0] node21097;
	wire [4-1:0] node21100;
	wire [4-1:0] node21101;
	wire [4-1:0] node21102;
	wire [4-1:0] node21103;
	wire [4-1:0] node21104;
	wire [4-1:0] node21107;
	wire [4-1:0] node21110;
	wire [4-1:0] node21111;
	wire [4-1:0] node21114;
	wire [4-1:0] node21117;
	wire [4-1:0] node21118;
	wire [4-1:0] node21120;
	wire [4-1:0] node21123;
	wire [4-1:0] node21124;
	wire [4-1:0] node21127;
	wire [4-1:0] node21130;
	wire [4-1:0] node21131;
	wire [4-1:0] node21132;
	wire [4-1:0] node21133;
	wire [4-1:0] node21137;
	wire [4-1:0] node21138;
	wire [4-1:0] node21142;
	wire [4-1:0] node21143;
	wire [4-1:0] node21144;
	wire [4-1:0] node21148;
	wire [4-1:0] node21149;
	wire [4-1:0] node21153;
	wire [4-1:0] node21154;
	wire [4-1:0] node21155;
	wire [4-1:0] node21156;
	wire [4-1:0] node21157;
	wire [4-1:0] node21158;
	wire [4-1:0] node21161;
	wire [4-1:0] node21164;
	wire [4-1:0] node21166;
	wire [4-1:0] node21169;
	wire [4-1:0] node21170;
	wire [4-1:0] node21171;
	wire [4-1:0] node21175;
	wire [4-1:0] node21176;
	wire [4-1:0] node21179;
	wire [4-1:0] node21182;
	wire [4-1:0] node21183;
	wire [4-1:0] node21184;
	wire [4-1:0] node21185;
	wire [4-1:0] node21188;
	wire [4-1:0] node21191;
	wire [4-1:0] node21192;
	wire [4-1:0] node21195;
	wire [4-1:0] node21198;
	wire [4-1:0] node21199;
	wire [4-1:0] node21202;
	wire [4-1:0] node21205;
	wire [4-1:0] node21206;
	wire [4-1:0] node21207;
	wire [4-1:0] node21208;
	wire [4-1:0] node21209;
	wire [4-1:0] node21213;
	wire [4-1:0] node21214;
	wire [4-1:0] node21217;
	wire [4-1:0] node21220;
	wire [4-1:0] node21221;
	wire [4-1:0] node21222;
	wire [4-1:0] node21225;
	wire [4-1:0] node21228;
	wire [4-1:0] node21230;
	wire [4-1:0] node21233;
	wire [4-1:0] node21234;
	wire [4-1:0] node21235;
	wire [4-1:0] node21236;
	wire [4-1:0] node21239;
	wire [4-1:0] node21242;
	wire [4-1:0] node21243;
	wire [4-1:0] node21246;
	wire [4-1:0] node21249;
	wire [4-1:0] node21250;
	wire [4-1:0] node21251;
	wire [4-1:0] node21254;
	wire [4-1:0] node21257;
	wire [4-1:0] node21258;
	wire [4-1:0] node21261;
	wire [4-1:0] node21264;
	wire [4-1:0] node21265;
	wire [4-1:0] node21266;
	wire [4-1:0] node21267;
	wire [4-1:0] node21268;
	wire [4-1:0] node21269;
	wire [4-1:0] node21270;
	wire [4-1:0] node21273;
	wire [4-1:0] node21276;
	wire [4-1:0] node21277;
	wire [4-1:0] node21280;
	wire [4-1:0] node21283;
	wire [4-1:0] node21284;
	wire [4-1:0] node21285;
	wire [4-1:0] node21288;
	wire [4-1:0] node21291;
	wire [4-1:0] node21292;
	wire [4-1:0] node21295;
	wire [4-1:0] node21298;
	wire [4-1:0] node21299;
	wire [4-1:0] node21300;
	wire [4-1:0] node21301;
	wire [4-1:0] node21305;
	wire [4-1:0] node21306;
	wire [4-1:0] node21310;
	wire [4-1:0] node21311;
	wire [4-1:0] node21312;
	wire [4-1:0] node21316;
	wire [4-1:0] node21317;
	wire [4-1:0] node21321;
	wire [4-1:0] node21322;
	wire [4-1:0] node21323;
	wire [4-1:0] node21324;
	wire [4-1:0] node21325;
	wire [4-1:0] node21328;
	wire [4-1:0] node21331;
	wire [4-1:0] node21332;
	wire [4-1:0] node21335;
	wire [4-1:0] node21338;
	wire [4-1:0] node21339;
	wire [4-1:0] node21340;
	wire [4-1:0] node21344;
	wire [4-1:0] node21345;
	wire [4-1:0] node21348;
	wire [4-1:0] node21351;
	wire [4-1:0] node21352;
	wire [4-1:0] node21353;
	wire [4-1:0] node21354;
	wire [4-1:0] node21358;
	wire [4-1:0] node21359;
	wire [4-1:0] node21363;
	wire [4-1:0] node21364;
	wire [4-1:0] node21365;
	wire [4-1:0] node21369;
	wire [4-1:0] node21370;
	wire [4-1:0] node21374;
	wire [4-1:0] node21375;
	wire [4-1:0] node21376;
	wire [4-1:0] node21377;
	wire [4-1:0] node21378;
	wire [4-1:0] node21379;
	wire [4-1:0] node21382;
	wire [4-1:0] node21385;
	wire [4-1:0] node21386;
	wire [4-1:0] node21390;
	wire [4-1:0] node21391;
	wire [4-1:0] node21392;
	wire [4-1:0] node21395;
	wire [4-1:0] node21398;
	wire [4-1:0] node21399;
	wire [4-1:0] node21402;
	wire [4-1:0] node21405;
	wire [4-1:0] node21406;
	wire [4-1:0] node21407;
	wire [4-1:0] node21408;
	wire [4-1:0] node21411;
	wire [4-1:0] node21414;
	wire [4-1:0] node21415;
	wire [4-1:0] node21418;
	wire [4-1:0] node21421;
	wire [4-1:0] node21422;
	wire [4-1:0] node21423;
	wire [4-1:0] node21426;
	wire [4-1:0] node21429;
	wire [4-1:0] node21430;
	wire [4-1:0] node21433;
	wire [4-1:0] node21436;
	wire [4-1:0] node21437;
	wire [4-1:0] node21438;
	wire [4-1:0] node21439;
	wire [4-1:0] node21440;
	wire [4-1:0] node21443;
	wire [4-1:0] node21446;
	wire [4-1:0] node21447;
	wire [4-1:0] node21450;
	wire [4-1:0] node21453;
	wire [4-1:0] node21454;
	wire [4-1:0] node21455;
	wire [4-1:0] node21458;
	wire [4-1:0] node21461;
	wire [4-1:0] node21462;
	wire [4-1:0] node21465;
	wire [4-1:0] node21468;
	wire [4-1:0] node21469;
	wire [4-1:0] node21470;
	wire [4-1:0] node21471;
	wire [4-1:0] node21475;
	wire [4-1:0] node21476;
	wire [4-1:0] node21480;
	wire [4-1:0] node21482;
	wire [4-1:0] node21483;
	wire [4-1:0] node21487;
	wire [4-1:0] node21488;
	wire [4-1:0] node21489;
	wire [4-1:0] node21490;
	wire [4-1:0] node21491;
	wire [4-1:0] node21492;
	wire [4-1:0] node21493;
	wire [4-1:0] node21494;
	wire [4-1:0] node21495;
	wire [4-1:0] node21496;
	wire [4-1:0] node21497;
	wire [4-1:0] node21498;
	wire [4-1:0] node21502;
	wire [4-1:0] node21503;
	wire [4-1:0] node21507;
	wire [4-1:0] node21508;
	wire [4-1:0] node21509;
	wire [4-1:0] node21513;
	wire [4-1:0] node21514;
	wire [4-1:0] node21518;
	wire [4-1:0] node21519;
	wire [4-1:0] node21520;
	wire [4-1:0] node21522;
	wire [4-1:0] node21525;
	wire [4-1:0] node21526;
	wire [4-1:0] node21529;
	wire [4-1:0] node21532;
	wire [4-1:0] node21533;
	wire [4-1:0] node21534;
	wire [4-1:0] node21537;
	wire [4-1:0] node21540;
	wire [4-1:0] node21541;
	wire [4-1:0] node21544;
	wire [4-1:0] node21547;
	wire [4-1:0] node21548;
	wire [4-1:0] node21549;
	wire [4-1:0] node21550;
	wire [4-1:0] node21552;
	wire [4-1:0] node21555;
	wire [4-1:0] node21556;
	wire [4-1:0] node21559;
	wire [4-1:0] node21562;
	wire [4-1:0] node21563;
	wire [4-1:0] node21566;
	wire [4-1:0] node21569;
	wire [4-1:0] node21570;
	wire [4-1:0] node21571;
	wire [4-1:0] node21573;
	wire [4-1:0] node21576;
	wire [4-1:0] node21577;
	wire [4-1:0] node21580;
	wire [4-1:0] node21583;
	wire [4-1:0] node21584;
	wire [4-1:0] node21586;
	wire [4-1:0] node21589;
	wire [4-1:0] node21590;
	wire [4-1:0] node21593;
	wire [4-1:0] node21596;
	wire [4-1:0] node21597;
	wire [4-1:0] node21598;
	wire [4-1:0] node21599;
	wire [4-1:0] node21600;
	wire [4-1:0] node21601;
	wire [4-1:0] node21605;
	wire [4-1:0] node21606;
	wire [4-1:0] node21610;
	wire [4-1:0] node21611;
	wire [4-1:0] node21612;
	wire [4-1:0] node21616;
	wire [4-1:0] node21617;
	wire [4-1:0] node21621;
	wire [4-1:0] node21622;
	wire [4-1:0] node21623;
	wire [4-1:0] node21624;
	wire [4-1:0] node21628;
	wire [4-1:0] node21629;
	wire [4-1:0] node21632;
	wire [4-1:0] node21635;
	wire [4-1:0] node21636;
	wire [4-1:0] node21637;
	wire [4-1:0] node21641;
	wire [4-1:0] node21642;
	wire [4-1:0] node21646;
	wire [4-1:0] node21647;
	wire [4-1:0] node21648;
	wire [4-1:0] node21649;
	wire [4-1:0] node21650;
	wire [4-1:0] node21654;
	wire [4-1:0] node21655;
	wire [4-1:0] node21659;
	wire [4-1:0] node21660;
	wire [4-1:0] node21661;
	wire [4-1:0] node21665;
	wire [4-1:0] node21666;
	wire [4-1:0] node21670;
	wire [4-1:0] node21671;
	wire [4-1:0] node21672;
	wire [4-1:0] node21673;
	wire [4-1:0] node21676;
	wire [4-1:0] node21679;
	wire [4-1:0] node21680;
	wire [4-1:0] node21683;
	wire [4-1:0] node21686;
	wire [4-1:0] node21687;
	wire [4-1:0] node21689;
	wire [4-1:0] node21692;
	wire [4-1:0] node21693;
	wire [4-1:0] node21696;
	wire [4-1:0] node21699;
	wire [4-1:0] node21700;
	wire [4-1:0] node21701;
	wire [4-1:0] node21702;
	wire [4-1:0] node21703;
	wire [4-1:0] node21704;
	wire [4-1:0] node21705;
	wire [4-1:0] node21708;
	wire [4-1:0] node21711;
	wire [4-1:0] node21712;
	wire [4-1:0] node21715;
	wire [4-1:0] node21718;
	wire [4-1:0] node21719;
	wire [4-1:0] node21721;
	wire [4-1:0] node21724;
	wire [4-1:0] node21726;
	wire [4-1:0] node21729;
	wire [4-1:0] node21730;
	wire [4-1:0] node21731;
	wire [4-1:0] node21732;
	wire [4-1:0] node21735;
	wire [4-1:0] node21738;
	wire [4-1:0] node21739;
	wire [4-1:0] node21743;
	wire [4-1:0] node21744;
	wire [4-1:0] node21745;
	wire [4-1:0] node21748;
	wire [4-1:0] node21751;
	wire [4-1:0] node21752;
	wire [4-1:0] node21755;
	wire [4-1:0] node21758;
	wire [4-1:0] node21759;
	wire [4-1:0] node21760;
	wire [4-1:0] node21761;
	wire [4-1:0] node21762;
	wire [4-1:0] node21765;
	wire [4-1:0] node21768;
	wire [4-1:0] node21769;
	wire [4-1:0] node21772;
	wire [4-1:0] node21775;
	wire [4-1:0] node21776;
	wire [4-1:0] node21777;
	wire [4-1:0] node21780;
	wire [4-1:0] node21783;
	wire [4-1:0] node21784;
	wire [4-1:0] node21787;
	wire [4-1:0] node21790;
	wire [4-1:0] node21791;
	wire [4-1:0] node21792;
	wire [4-1:0] node21794;
	wire [4-1:0] node21797;
	wire [4-1:0] node21799;
	wire [4-1:0] node21802;
	wire [4-1:0] node21803;
	wire [4-1:0] node21805;
	wire [4-1:0] node21808;
	wire [4-1:0] node21810;
	wire [4-1:0] node21813;
	wire [4-1:0] node21814;
	wire [4-1:0] node21815;
	wire [4-1:0] node21816;
	wire [4-1:0] node21817;
	wire [4-1:0] node21818;
	wire [4-1:0] node21821;
	wire [4-1:0] node21824;
	wire [4-1:0] node21825;
	wire [4-1:0] node21828;
	wire [4-1:0] node21831;
	wire [4-1:0] node21832;
	wire [4-1:0] node21833;
	wire [4-1:0] node21836;
	wire [4-1:0] node21839;
	wire [4-1:0] node21841;
	wire [4-1:0] node21844;
	wire [4-1:0] node21845;
	wire [4-1:0] node21846;
	wire [4-1:0] node21847;
	wire [4-1:0] node21850;
	wire [4-1:0] node21853;
	wire [4-1:0] node21854;
	wire [4-1:0] node21857;
	wire [4-1:0] node21860;
	wire [4-1:0] node21861;
	wire [4-1:0] node21862;
	wire [4-1:0] node21865;
	wire [4-1:0] node21868;
	wire [4-1:0] node21869;
	wire [4-1:0] node21872;
	wire [4-1:0] node21875;
	wire [4-1:0] node21876;
	wire [4-1:0] node21877;
	wire [4-1:0] node21878;
	wire [4-1:0] node21879;
	wire [4-1:0] node21882;
	wire [4-1:0] node21885;
	wire [4-1:0] node21886;
	wire [4-1:0] node21889;
	wire [4-1:0] node21892;
	wire [4-1:0] node21893;
	wire [4-1:0] node21894;
	wire [4-1:0] node21897;
	wire [4-1:0] node21900;
	wire [4-1:0] node21901;
	wire [4-1:0] node21905;
	wire [4-1:0] node21906;
	wire [4-1:0] node21907;
	wire [4-1:0] node21909;
	wire [4-1:0] node21912;
	wire [4-1:0] node21914;
	wire [4-1:0] node21917;
	wire [4-1:0] node21918;
	wire [4-1:0] node21920;
	wire [4-1:0] node21923;
	wire [4-1:0] node21925;
	wire [4-1:0] node21928;
	wire [4-1:0] node21929;
	wire [4-1:0] node21930;
	wire [4-1:0] node21931;
	wire [4-1:0] node21932;
	wire [4-1:0] node21933;
	wire [4-1:0] node21934;
	wire [4-1:0] node21935;
	wire [4-1:0] node21938;
	wire [4-1:0] node21941;
	wire [4-1:0] node21942;
	wire [4-1:0] node21945;
	wire [4-1:0] node21948;
	wire [4-1:0] node21949;
	wire [4-1:0] node21950;
	wire [4-1:0] node21953;
	wire [4-1:0] node21956;
	wire [4-1:0] node21958;
	wire [4-1:0] node21961;
	wire [4-1:0] node21962;
	wire [4-1:0] node21963;
	wire [4-1:0] node21965;
	wire [4-1:0] node21968;
	wire [4-1:0] node21970;
	wire [4-1:0] node21973;
	wire [4-1:0] node21974;
	wire [4-1:0] node21976;
	wire [4-1:0] node21979;
	wire [4-1:0] node21981;
	wire [4-1:0] node21984;
	wire [4-1:0] node21985;
	wire [4-1:0] node21986;
	wire [4-1:0] node21987;
	wire [4-1:0] node21988;
	wire [4-1:0] node21992;
	wire [4-1:0] node21993;
	wire [4-1:0] node21996;
	wire [4-1:0] node21999;
	wire [4-1:0] node22000;
	wire [4-1:0] node22001;
	wire [4-1:0] node22004;
	wire [4-1:0] node22007;
	wire [4-1:0] node22008;
	wire [4-1:0] node22011;
	wire [4-1:0] node22014;
	wire [4-1:0] node22015;
	wire [4-1:0] node22016;
	wire [4-1:0] node22018;
	wire [4-1:0] node22021;
	wire [4-1:0] node22023;
	wire [4-1:0] node22026;
	wire [4-1:0] node22027;
	wire [4-1:0] node22029;
	wire [4-1:0] node22032;
	wire [4-1:0] node22035;
	wire [4-1:0] node22036;
	wire [4-1:0] node22037;
	wire [4-1:0] node22038;
	wire [4-1:0] node22039;
	wire [4-1:0] node22040;
	wire [4-1:0] node22043;
	wire [4-1:0] node22046;
	wire [4-1:0] node22047;
	wire [4-1:0] node22050;
	wire [4-1:0] node22053;
	wire [4-1:0] node22054;
	wire [4-1:0] node22055;
	wire [4-1:0] node22059;
	wire [4-1:0] node22061;
	wire [4-1:0] node22064;
	wire [4-1:0] node22065;
	wire [4-1:0] node22066;
	wire [4-1:0] node22067;
	wire [4-1:0] node22070;
	wire [4-1:0] node22073;
	wire [4-1:0] node22075;
	wire [4-1:0] node22078;
	wire [4-1:0] node22079;
	wire [4-1:0] node22080;
	wire [4-1:0] node22083;
	wire [4-1:0] node22086;
	wire [4-1:0] node22087;
	wire [4-1:0] node22090;
	wire [4-1:0] node22093;
	wire [4-1:0] node22094;
	wire [4-1:0] node22095;
	wire [4-1:0] node22096;
	wire [4-1:0] node22097;
	wire [4-1:0] node22100;
	wire [4-1:0] node22103;
	wire [4-1:0] node22104;
	wire [4-1:0] node22107;
	wire [4-1:0] node22110;
	wire [4-1:0] node22111;
	wire [4-1:0] node22112;
	wire [4-1:0] node22115;
	wire [4-1:0] node22118;
	wire [4-1:0] node22119;
	wire [4-1:0] node22122;
	wire [4-1:0] node22125;
	wire [4-1:0] node22126;
	wire [4-1:0] node22127;
	wire [4-1:0] node22129;
	wire [4-1:0] node22132;
	wire [4-1:0] node22134;
	wire [4-1:0] node22137;
	wire [4-1:0] node22138;
	wire [4-1:0] node22140;
	wire [4-1:0] node22143;
	wire [4-1:0] node22145;
	wire [4-1:0] node22148;
	wire [4-1:0] node22149;
	wire [4-1:0] node22150;
	wire [4-1:0] node22151;
	wire [4-1:0] node22152;
	wire [4-1:0] node22153;
	wire [4-1:0] node22154;
	wire [4-1:0] node22157;
	wire [4-1:0] node22160;
	wire [4-1:0] node22161;
	wire [4-1:0] node22164;
	wire [4-1:0] node22167;
	wire [4-1:0] node22168;
	wire [4-1:0] node22170;
	wire [4-1:0] node22173;
	wire [4-1:0] node22174;
	wire [4-1:0] node22177;
	wire [4-1:0] node22180;
	wire [4-1:0] node22181;
	wire [4-1:0] node22182;
	wire [4-1:0] node22184;
	wire [4-1:0] node22187;
	wire [4-1:0] node22189;
	wire [4-1:0] node22192;
	wire [4-1:0] node22193;
	wire [4-1:0] node22195;
	wire [4-1:0] node22198;
	wire [4-1:0] node22200;
	wire [4-1:0] node22203;
	wire [4-1:0] node22204;
	wire [4-1:0] node22205;
	wire [4-1:0] node22206;
	wire [4-1:0] node22208;
	wire [4-1:0] node22211;
	wire [4-1:0] node22212;
	wire [4-1:0] node22215;
	wire [4-1:0] node22218;
	wire [4-1:0] node22219;
	wire [4-1:0] node22221;
	wire [4-1:0] node22224;
	wire [4-1:0] node22225;
	wire [4-1:0] node22228;
	wire [4-1:0] node22231;
	wire [4-1:0] node22232;
	wire [4-1:0] node22233;
	wire [4-1:0] node22235;
	wire [4-1:0] node22238;
	wire [4-1:0] node22240;
	wire [4-1:0] node22243;
	wire [4-1:0] node22244;
	wire [4-1:0] node22246;
	wire [4-1:0] node22249;
	wire [4-1:0] node22251;
	wire [4-1:0] node22254;
	wire [4-1:0] node22255;
	wire [4-1:0] node22256;
	wire [4-1:0] node22257;
	wire [4-1:0] node22258;
	wire [4-1:0] node22259;
	wire [4-1:0] node22262;
	wire [4-1:0] node22265;
	wire [4-1:0] node22267;
	wire [4-1:0] node22270;
	wire [4-1:0] node22271;
	wire [4-1:0] node22272;
	wire [4-1:0] node22276;
	wire [4-1:0] node22277;
	wire [4-1:0] node22281;
	wire [4-1:0] node22282;
	wire [4-1:0] node22283;
	wire [4-1:0] node22285;
	wire [4-1:0] node22288;
	wire [4-1:0] node22290;
	wire [4-1:0] node22293;
	wire [4-1:0] node22294;
	wire [4-1:0] node22296;
	wire [4-1:0] node22299;
	wire [4-1:0] node22301;
	wire [4-1:0] node22304;
	wire [4-1:0] node22305;
	wire [4-1:0] node22306;
	wire [4-1:0] node22307;
	wire [4-1:0] node22308;
	wire [4-1:0] node22312;
	wire [4-1:0] node22313;
	wire [4-1:0] node22316;
	wire [4-1:0] node22319;
	wire [4-1:0] node22320;
	wire [4-1:0] node22321;
	wire [4-1:0] node22325;
	wire [4-1:0] node22326;
	wire [4-1:0] node22329;
	wire [4-1:0] node22332;
	wire [4-1:0] node22333;
	wire [4-1:0] node22334;
	wire [4-1:0] node22337;
	wire [4-1:0] node22340;
	wire [4-1:0] node22341;
	wire [4-1:0] node22342;
	wire [4-1:0] node22345;
	wire [4-1:0] node22348;
	wire [4-1:0] node22349;
	wire [4-1:0] node22352;
	wire [4-1:0] node22355;
	wire [4-1:0] node22356;
	wire [4-1:0] node22357;
	wire [4-1:0] node22358;
	wire [4-1:0] node22359;
	wire [4-1:0] node22360;
	wire [4-1:0] node22361;
	wire [4-1:0] node22362;
	wire [4-1:0] node22363;
	wire [4-1:0] node22366;
	wire [4-1:0] node22369;
	wire [4-1:0] node22370;
	wire [4-1:0] node22373;
	wire [4-1:0] node22376;
	wire [4-1:0] node22377;
	wire [4-1:0] node22378;
	wire [4-1:0] node22381;
	wire [4-1:0] node22384;
	wire [4-1:0] node22385;
	wire [4-1:0] node22388;
	wire [4-1:0] node22391;
	wire [4-1:0] node22392;
	wire [4-1:0] node22393;
	wire [4-1:0] node22394;
	wire [4-1:0] node22397;
	wire [4-1:0] node22400;
	wire [4-1:0] node22401;
	wire [4-1:0] node22404;
	wire [4-1:0] node22407;
	wire [4-1:0] node22408;
	wire [4-1:0] node22409;
	wire [4-1:0] node22412;
	wire [4-1:0] node22415;
	wire [4-1:0] node22417;
	wire [4-1:0] node22420;
	wire [4-1:0] node22421;
	wire [4-1:0] node22422;
	wire [4-1:0] node22423;
	wire [4-1:0] node22424;
	wire [4-1:0] node22427;
	wire [4-1:0] node22430;
	wire [4-1:0] node22431;
	wire [4-1:0] node22434;
	wire [4-1:0] node22437;
	wire [4-1:0] node22438;
	wire [4-1:0] node22439;
	wire [4-1:0] node22442;
	wire [4-1:0] node22445;
	wire [4-1:0] node22446;
	wire [4-1:0] node22449;
	wire [4-1:0] node22452;
	wire [4-1:0] node22453;
	wire [4-1:0] node22454;
	wire [4-1:0] node22455;
	wire [4-1:0] node22459;
	wire [4-1:0] node22460;
	wire [4-1:0] node22463;
	wire [4-1:0] node22466;
	wire [4-1:0] node22467;
	wire [4-1:0] node22468;
	wire [4-1:0] node22471;
	wire [4-1:0] node22474;
	wire [4-1:0] node22475;
	wire [4-1:0] node22478;
	wire [4-1:0] node22481;
	wire [4-1:0] node22482;
	wire [4-1:0] node22483;
	wire [4-1:0] node22484;
	wire [4-1:0] node22485;
	wire [4-1:0] node22486;
	wire [4-1:0] node22489;
	wire [4-1:0] node22492;
	wire [4-1:0] node22493;
	wire [4-1:0] node22496;
	wire [4-1:0] node22499;
	wire [4-1:0] node22500;
	wire [4-1:0] node22501;
	wire [4-1:0] node22504;
	wire [4-1:0] node22507;
	wire [4-1:0] node22508;
	wire [4-1:0] node22511;
	wire [4-1:0] node22514;
	wire [4-1:0] node22515;
	wire [4-1:0] node22516;
	wire [4-1:0] node22517;
	wire [4-1:0] node22520;
	wire [4-1:0] node22523;
	wire [4-1:0] node22524;
	wire [4-1:0] node22527;
	wire [4-1:0] node22530;
	wire [4-1:0] node22531;
	wire [4-1:0] node22532;
	wire [4-1:0] node22535;
	wire [4-1:0] node22538;
	wire [4-1:0] node22539;
	wire [4-1:0] node22543;
	wire [4-1:0] node22544;
	wire [4-1:0] node22545;
	wire [4-1:0] node22546;
	wire [4-1:0] node22547;
	wire [4-1:0] node22550;
	wire [4-1:0] node22553;
	wire [4-1:0] node22554;
	wire [4-1:0] node22557;
	wire [4-1:0] node22560;
	wire [4-1:0] node22561;
	wire [4-1:0] node22562;
	wire [4-1:0] node22565;
	wire [4-1:0] node22568;
	wire [4-1:0] node22569;
	wire [4-1:0] node22572;
	wire [4-1:0] node22575;
	wire [4-1:0] node22576;
	wire [4-1:0] node22577;
	wire [4-1:0] node22578;
	wire [4-1:0] node22581;
	wire [4-1:0] node22584;
	wire [4-1:0] node22585;
	wire [4-1:0] node22588;
	wire [4-1:0] node22591;
	wire [4-1:0] node22592;
	wire [4-1:0] node22593;
	wire [4-1:0] node22596;
	wire [4-1:0] node22599;
	wire [4-1:0] node22600;
	wire [4-1:0] node22603;
	wire [4-1:0] node22606;
	wire [4-1:0] node22607;
	wire [4-1:0] node22608;
	wire [4-1:0] node22609;
	wire [4-1:0] node22610;
	wire [4-1:0] node22611;
	wire [4-1:0] node22612;
	wire [4-1:0] node22615;
	wire [4-1:0] node22618;
	wire [4-1:0] node22619;
	wire [4-1:0] node22623;
	wire [4-1:0] node22624;
	wire [4-1:0] node22625;
	wire [4-1:0] node22628;
	wire [4-1:0] node22631;
	wire [4-1:0] node22632;
	wire [4-1:0] node22635;
	wire [4-1:0] node22638;
	wire [4-1:0] node22639;
	wire [4-1:0] node22640;
	wire [4-1:0] node22642;
	wire [4-1:0] node22645;
	wire [4-1:0] node22647;
	wire [4-1:0] node22650;
	wire [4-1:0] node22651;
	wire [4-1:0] node22653;
	wire [4-1:0] node22656;
	wire [4-1:0] node22658;
	wire [4-1:0] node22661;
	wire [4-1:0] node22662;
	wire [4-1:0] node22663;
	wire [4-1:0] node22664;
	wire [4-1:0] node22665;
	wire [4-1:0] node22668;
	wire [4-1:0] node22671;
	wire [4-1:0] node22672;
	wire [4-1:0] node22675;
	wire [4-1:0] node22678;
	wire [4-1:0] node22679;
	wire [4-1:0] node22680;
	wire [4-1:0] node22684;
	wire [4-1:0] node22686;
	wire [4-1:0] node22689;
	wire [4-1:0] node22690;
	wire [4-1:0] node22691;
	wire [4-1:0] node22692;
	wire [4-1:0] node22695;
	wire [4-1:0] node22698;
	wire [4-1:0] node22699;
	wire [4-1:0] node22703;
	wire [4-1:0] node22704;
	wire [4-1:0] node22705;
	wire [4-1:0] node22708;
	wire [4-1:0] node22711;
	wire [4-1:0] node22712;
	wire [4-1:0] node22715;
	wire [4-1:0] node22718;
	wire [4-1:0] node22719;
	wire [4-1:0] node22720;
	wire [4-1:0] node22721;
	wire [4-1:0] node22722;
	wire [4-1:0] node22723;
	wire [4-1:0] node22726;
	wire [4-1:0] node22729;
	wire [4-1:0] node22730;
	wire [4-1:0] node22733;
	wire [4-1:0] node22736;
	wire [4-1:0] node22737;
	wire [4-1:0] node22738;
	wire [4-1:0] node22741;
	wire [4-1:0] node22744;
	wire [4-1:0] node22746;
	wire [4-1:0] node22749;
	wire [4-1:0] node22750;
	wire [4-1:0] node22751;
	wire [4-1:0] node22752;
	wire [4-1:0] node22755;
	wire [4-1:0] node22758;
	wire [4-1:0] node22759;
	wire [4-1:0] node22762;
	wire [4-1:0] node22765;
	wire [4-1:0] node22766;
	wire [4-1:0] node22769;
	wire [4-1:0] node22772;
	wire [4-1:0] node22773;
	wire [4-1:0] node22774;
	wire [4-1:0] node22775;
	wire [4-1:0] node22776;
	wire [4-1:0] node22779;
	wire [4-1:0] node22782;
	wire [4-1:0] node22783;
	wire [4-1:0] node22786;
	wire [4-1:0] node22789;
	wire [4-1:0] node22790;
	wire [4-1:0] node22791;
	wire [4-1:0] node22795;
	wire [4-1:0] node22797;
	wire [4-1:0] node22800;
	wire [4-1:0] node22801;
	wire [4-1:0] node22802;
	wire [4-1:0] node22803;
	wire [4-1:0] node22806;
	wire [4-1:0] node22809;
	wire [4-1:0] node22810;
	wire [4-1:0] node22813;
	wire [4-1:0] node22816;
	wire [4-1:0] node22817;
	wire [4-1:0] node22820;
	wire [4-1:0] node22823;
	wire [4-1:0] node22824;
	wire [4-1:0] node22825;
	wire [4-1:0] node22826;
	wire [4-1:0] node22827;
	wire [4-1:0] node22828;
	wire [4-1:0] node22829;
	wire [4-1:0] node22830;
	wire [4-1:0] node22833;
	wire [4-1:0] node22836;
	wire [4-1:0] node22837;
	wire [4-1:0] node22840;
	wire [4-1:0] node22843;
	wire [4-1:0] node22844;
	wire [4-1:0] node22845;
	wire [4-1:0] node22848;
	wire [4-1:0] node22851;
	wire [4-1:0] node22852;
	wire [4-1:0] node22855;
	wire [4-1:0] node22858;
	wire [4-1:0] node22859;
	wire [4-1:0] node22860;
	wire [4-1:0] node22862;
	wire [4-1:0] node22865;
	wire [4-1:0] node22868;
	wire [4-1:0] node22869;
	wire [4-1:0] node22871;
	wire [4-1:0] node22874;
	wire [4-1:0] node22876;
	wire [4-1:0] node22879;
	wire [4-1:0] node22880;
	wire [4-1:0] node22881;
	wire [4-1:0] node22882;
	wire [4-1:0] node22883;
	wire [4-1:0] node22886;
	wire [4-1:0] node22889;
	wire [4-1:0] node22890;
	wire [4-1:0] node22893;
	wire [4-1:0] node22896;
	wire [4-1:0] node22897;
	wire [4-1:0] node22898;
	wire [4-1:0] node22902;
	wire [4-1:0] node22903;
	wire [4-1:0] node22906;
	wire [4-1:0] node22909;
	wire [4-1:0] node22910;
	wire [4-1:0] node22911;
	wire [4-1:0] node22912;
	wire [4-1:0] node22916;
	wire [4-1:0] node22919;
	wire [4-1:0] node22920;
	wire [4-1:0] node22921;
	wire [4-1:0] node22925;
	wire [4-1:0] node22926;
	wire [4-1:0] node22930;
	wire [4-1:0] node22931;
	wire [4-1:0] node22932;
	wire [4-1:0] node22933;
	wire [4-1:0] node22934;
	wire [4-1:0] node22935;
	wire [4-1:0] node22938;
	wire [4-1:0] node22941;
	wire [4-1:0] node22942;
	wire [4-1:0] node22945;
	wire [4-1:0] node22948;
	wire [4-1:0] node22949;
	wire [4-1:0] node22950;
	wire [4-1:0] node22954;
	wire [4-1:0] node22955;
	wire [4-1:0] node22958;
	wire [4-1:0] node22961;
	wire [4-1:0] node22962;
	wire [4-1:0] node22963;
	wire [4-1:0] node22964;
	wire [4-1:0] node22967;
	wire [4-1:0] node22970;
	wire [4-1:0] node22971;
	wire [4-1:0] node22974;
	wire [4-1:0] node22977;
	wire [4-1:0] node22978;
	wire [4-1:0] node22980;
	wire [4-1:0] node22983;
	wire [4-1:0] node22984;
	wire [4-1:0] node22987;
	wire [4-1:0] node22990;
	wire [4-1:0] node22991;
	wire [4-1:0] node22992;
	wire [4-1:0] node22993;
	wire [4-1:0] node22994;
	wire [4-1:0] node22997;
	wire [4-1:0] node23000;
	wire [4-1:0] node23001;
	wire [4-1:0] node23005;
	wire [4-1:0] node23006;
	wire [4-1:0] node23007;
	wire [4-1:0] node23010;
	wire [4-1:0] node23014;
	wire [4-1:0] node23015;
	wire [4-1:0] node23016;
	wire [4-1:0] node23017;
	wire [4-1:0] node23021;
	wire [4-1:0] node23022;
	wire [4-1:0] node23026;
	wire [4-1:0] node23027;
	wire [4-1:0] node23028;
	wire [4-1:0] node23032;
	wire [4-1:0] node23033;
	wire [4-1:0] node23037;
	wire [4-1:0] node23038;
	wire [4-1:0] node23039;
	wire [4-1:0] node23040;
	wire [4-1:0] node23041;
	wire [4-1:0] node23042;
	wire [4-1:0] node23043;
	wire [4-1:0] node23046;
	wire [4-1:0] node23049;
	wire [4-1:0] node23050;
	wire [4-1:0] node23053;
	wire [4-1:0] node23056;
	wire [4-1:0] node23057;
	wire [4-1:0] node23058;
	wire [4-1:0] node23061;
	wire [4-1:0] node23064;
	wire [4-1:0] node23065;
	wire [4-1:0] node23068;
	wire [4-1:0] node23071;
	wire [4-1:0] node23072;
	wire [4-1:0] node23073;
	wire [4-1:0] node23074;
	wire [4-1:0] node23077;
	wire [4-1:0] node23080;
	wire [4-1:0] node23081;
	wire [4-1:0] node23084;
	wire [4-1:0] node23087;
	wire [4-1:0] node23088;
	wire [4-1:0] node23089;
	wire [4-1:0] node23092;
	wire [4-1:0] node23095;
	wire [4-1:0] node23096;
	wire [4-1:0] node23099;
	wire [4-1:0] node23102;
	wire [4-1:0] node23103;
	wire [4-1:0] node23104;
	wire [4-1:0] node23105;
	wire [4-1:0] node23106;
	wire [4-1:0] node23110;
	wire [4-1:0] node23111;
	wire [4-1:0] node23114;
	wire [4-1:0] node23117;
	wire [4-1:0] node23118;
	wire [4-1:0] node23119;
	wire [4-1:0] node23122;
	wire [4-1:0] node23125;
	wire [4-1:0] node23126;
	wire [4-1:0] node23129;
	wire [4-1:0] node23132;
	wire [4-1:0] node23133;
	wire [4-1:0] node23134;
	wire [4-1:0] node23135;
	wire [4-1:0] node23138;
	wire [4-1:0] node23141;
	wire [4-1:0] node23142;
	wire [4-1:0] node23145;
	wire [4-1:0] node23148;
	wire [4-1:0] node23149;
	wire [4-1:0] node23150;
	wire [4-1:0] node23153;
	wire [4-1:0] node23156;
	wire [4-1:0] node23157;
	wire [4-1:0] node23160;
	wire [4-1:0] node23163;
	wire [4-1:0] node23164;
	wire [4-1:0] node23165;
	wire [4-1:0] node23166;
	wire [4-1:0] node23167;
	wire [4-1:0] node23168;
	wire [4-1:0] node23171;
	wire [4-1:0] node23174;
	wire [4-1:0] node23175;
	wire [4-1:0] node23179;
	wire [4-1:0] node23180;
	wire [4-1:0] node23181;
	wire [4-1:0] node23184;
	wire [4-1:0] node23187;
	wire [4-1:0] node23188;
	wire [4-1:0] node23191;
	wire [4-1:0] node23194;
	wire [4-1:0] node23195;
	wire [4-1:0] node23196;
	wire [4-1:0] node23197;
	wire [4-1:0] node23200;
	wire [4-1:0] node23203;
	wire [4-1:0] node23206;
	wire [4-1:0] node23207;
	wire [4-1:0] node23208;
	wire [4-1:0] node23211;
	wire [4-1:0] node23214;
	wire [4-1:0] node23215;
	wire [4-1:0] node23218;
	wire [4-1:0] node23221;
	wire [4-1:0] node23222;
	wire [4-1:0] node23223;
	wire [4-1:0] node23224;
	wire [4-1:0] node23225;
	wire [4-1:0] node23228;
	wire [4-1:0] node23231;
	wire [4-1:0] node23232;
	wire [4-1:0] node23235;
	wire [4-1:0] node23238;
	wire [4-1:0] node23239;
	wire [4-1:0] node23241;
	wire [4-1:0] node23244;
	wire [4-1:0] node23245;
	wire [4-1:0] node23248;
	wire [4-1:0] node23251;
	wire [4-1:0] node23252;
	wire [4-1:0] node23253;
	wire [4-1:0] node23254;
	wire [4-1:0] node23257;
	wire [4-1:0] node23260;
	wire [4-1:0] node23261;
	wire [4-1:0] node23264;
	wire [4-1:0] node23267;
	wire [4-1:0] node23268;
	wire [4-1:0] node23269;
	wire [4-1:0] node23273;
	wire [4-1:0] node23275;
	wire [4-1:0] node23278;
	wire [4-1:0] node23279;
	wire [4-1:0] node23280;
	wire [4-1:0] node23281;
	wire [4-1:0] node23282;
	wire [4-1:0] node23283;
	wire [4-1:0] node23284;
	wire [4-1:0] node23285;
	wire [4-1:0] node23286;
	wire [4-1:0] node23287;
	wire [4-1:0] node23291;
	wire [4-1:0] node23292;
	wire [4-1:0] node23296;
	wire [4-1:0] node23297;
	wire [4-1:0] node23298;
	wire [4-1:0] node23302;
	wire [4-1:0] node23303;
	wire [4-1:0] node23307;
	wire [4-1:0] node23308;
	wire [4-1:0] node23309;
	wire [4-1:0] node23311;
	wire [4-1:0] node23314;
	wire [4-1:0] node23315;
	wire [4-1:0] node23318;
	wire [4-1:0] node23321;
	wire [4-1:0] node23322;
	wire [4-1:0] node23323;
	wire [4-1:0] node23326;
	wire [4-1:0] node23329;
	wire [4-1:0] node23330;
	wire [4-1:0] node23333;
	wire [4-1:0] node23336;
	wire [4-1:0] node23337;
	wire [4-1:0] node23338;
	wire [4-1:0] node23339;
	wire [4-1:0] node23340;
	wire [4-1:0] node23343;
	wire [4-1:0] node23346;
	wire [4-1:0] node23347;
	wire [4-1:0] node23350;
	wire [4-1:0] node23353;
	wire [4-1:0] node23354;
	wire [4-1:0] node23357;
	wire [4-1:0] node23360;
	wire [4-1:0] node23361;
	wire [4-1:0] node23362;
	wire [4-1:0] node23363;
	wire [4-1:0] node23366;
	wire [4-1:0] node23369;
	wire [4-1:0] node23370;
	wire [4-1:0] node23374;
	wire [4-1:0] node23375;
	wire [4-1:0] node23376;
	wire [4-1:0] node23379;
	wire [4-1:0] node23382;
	wire [4-1:0] node23383;
	wire [4-1:0] node23386;
	wire [4-1:0] node23389;
	wire [4-1:0] node23390;
	wire [4-1:0] node23391;
	wire [4-1:0] node23392;
	wire [4-1:0] node23393;
	wire [4-1:0] node23394;
	wire [4-1:0] node23397;
	wire [4-1:0] node23400;
	wire [4-1:0] node23401;
	wire [4-1:0] node23404;
	wire [4-1:0] node23407;
	wire [4-1:0] node23408;
	wire [4-1:0] node23409;
	wire [4-1:0] node23412;
	wire [4-1:0] node23415;
	wire [4-1:0] node23416;
	wire [4-1:0] node23419;
	wire [4-1:0] node23422;
	wire [4-1:0] node23423;
	wire [4-1:0] node23424;
	wire [4-1:0] node23426;
	wire [4-1:0] node23429;
	wire [4-1:0] node23430;
	wire [4-1:0] node23433;
	wire [4-1:0] node23436;
	wire [4-1:0] node23437;
	wire [4-1:0] node23438;
	wire [4-1:0] node23441;
	wire [4-1:0] node23444;
	wire [4-1:0] node23446;
	wire [4-1:0] node23449;
	wire [4-1:0] node23450;
	wire [4-1:0] node23451;
	wire [4-1:0] node23452;
	wire [4-1:0] node23453;
	wire [4-1:0] node23457;
	wire [4-1:0] node23458;
	wire [4-1:0] node23462;
	wire [4-1:0] node23463;
	wire [4-1:0] node23466;
	wire [4-1:0] node23467;
	wire [4-1:0] node23471;
	wire [4-1:0] node23472;
	wire [4-1:0] node23473;
	wire [4-1:0] node23475;
	wire [4-1:0] node23478;
	wire [4-1:0] node23479;
	wire [4-1:0] node23482;
	wire [4-1:0] node23485;
	wire [4-1:0] node23486;
	wire [4-1:0] node23487;
	wire [4-1:0] node23490;
	wire [4-1:0] node23493;
	wire [4-1:0] node23495;
	wire [4-1:0] node23498;
	wire [4-1:0] node23499;
	wire [4-1:0] node23500;
	wire [4-1:0] node23501;
	wire [4-1:0] node23502;
	wire [4-1:0] node23503;
	wire [4-1:0] node23504;
	wire [4-1:0] node23507;
	wire [4-1:0] node23510;
	wire [4-1:0] node23512;
	wire [4-1:0] node23515;
	wire [4-1:0] node23516;
	wire [4-1:0] node23517;
	wire [4-1:0] node23520;
	wire [4-1:0] node23523;
	wire [4-1:0] node23524;
	wire [4-1:0] node23527;
	wire [4-1:0] node23530;
	wire [4-1:0] node23531;
	wire [4-1:0] node23532;
	wire [4-1:0] node23535;
	wire [4-1:0] node23538;
	wire [4-1:0] node23539;
	wire [4-1:0] node23540;
	wire [4-1:0] node23543;
	wire [4-1:0] node23546;
	wire [4-1:0] node23547;
	wire [4-1:0] node23550;
	wire [4-1:0] node23553;
	wire [4-1:0] node23554;
	wire [4-1:0] node23555;
	wire [4-1:0] node23556;
	wire [4-1:0] node23557;
	wire [4-1:0] node23560;
	wire [4-1:0] node23563;
	wire [4-1:0] node23564;
	wire [4-1:0] node23567;
	wire [4-1:0] node23570;
	wire [4-1:0] node23571;
	wire [4-1:0] node23572;
	wire [4-1:0] node23575;
	wire [4-1:0] node23578;
	wire [4-1:0] node23579;
	wire [4-1:0] node23583;
	wire [4-1:0] node23584;
	wire [4-1:0] node23585;
	wire [4-1:0] node23586;
	wire [4-1:0] node23589;
	wire [4-1:0] node23592;
	wire [4-1:0] node23593;
	wire [4-1:0] node23596;
	wire [4-1:0] node23599;
	wire [4-1:0] node23600;
	wire [4-1:0] node23601;
	wire [4-1:0] node23604;
	wire [4-1:0] node23607;
	wire [4-1:0] node23608;
	wire [4-1:0] node23611;
	wire [4-1:0] node23614;
	wire [4-1:0] node23615;
	wire [4-1:0] node23616;
	wire [4-1:0] node23617;
	wire [4-1:0] node23618;
	wire [4-1:0] node23619;
	wire [4-1:0] node23622;
	wire [4-1:0] node23625;
	wire [4-1:0] node23627;
	wire [4-1:0] node23630;
	wire [4-1:0] node23631;
	wire [4-1:0] node23632;
	wire [4-1:0] node23635;
	wire [4-1:0] node23638;
	wire [4-1:0] node23639;
	wire [4-1:0] node23642;
	wire [4-1:0] node23645;
	wire [4-1:0] node23646;
	wire [4-1:0] node23647;
	wire [4-1:0] node23648;
	wire [4-1:0] node23651;
	wire [4-1:0] node23654;
	wire [4-1:0] node23655;
	wire [4-1:0] node23658;
	wire [4-1:0] node23661;
	wire [4-1:0] node23662;
	wire [4-1:0] node23665;
	wire [4-1:0] node23668;
	wire [4-1:0] node23669;
	wire [4-1:0] node23670;
	wire [4-1:0] node23671;
	wire [4-1:0] node23673;
	wire [4-1:0] node23676;
	wire [4-1:0] node23677;
	wire [4-1:0] node23680;
	wire [4-1:0] node23683;
	wire [4-1:0] node23684;
	wire [4-1:0] node23685;
	wire [4-1:0] node23688;
	wire [4-1:0] node23691;
	wire [4-1:0] node23694;
	wire [4-1:0] node23695;
	wire [4-1:0] node23696;
	wire [4-1:0] node23697;
	wire [4-1:0] node23701;
	wire [4-1:0] node23702;
	wire [4-1:0] node23706;
	wire [4-1:0] node23707;
	wire [4-1:0] node23708;
	wire [4-1:0] node23712;
	wire [4-1:0] node23713;
	wire [4-1:0] node23717;
	wire [4-1:0] node23718;
	wire [4-1:0] node23719;
	wire [4-1:0] node23720;
	wire [4-1:0] node23721;
	wire [4-1:0] node23722;
	wire [4-1:0] node23723;
	wire [4-1:0] node23724;
	wire [4-1:0] node23728;
	wire [4-1:0] node23730;
	wire [4-1:0] node23733;
	wire [4-1:0] node23734;
	wire [4-1:0] node23735;
	wire [4-1:0] node23738;
	wire [4-1:0] node23741;
	wire [4-1:0] node23742;
	wire [4-1:0] node23746;
	wire [4-1:0] node23747;
	wire [4-1:0] node23748;
	wire [4-1:0] node23749;
	wire [4-1:0] node23752;
	wire [4-1:0] node23755;
	wire [4-1:0] node23757;
	wire [4-1:0] node23760;
	wire [4-1:0] node23761;
	wire [4-1:0] node23762;
	wire [4-1:0] node23765;
	wire [4-1:0] node23768;
	wire [4-1:0] node23769;
	wire [4-1:0] node23772;
	wire [4-1:0] node23775;
	wire [4-1:0] node23776;
	wire [4-1:0] node23777;
	wire [4-1:0] node23778;
	wire [4-1:0] node23779;
	wire [4-1:0] node23782;
	wire [4-1:0] node23785;
	wire [4-1:0] node23786;
	wire [4-1:0] node23789;
	wire [4-1:0] node23792;
	wire [4-1:0] node23793;
	wire [4-1:0] node23794;
	wire [4-1:0] node23798;
	wire [4-1:0] node23799;
	wire [4-1:0] node23802;
	wire [4-1:0] node23805;
	wire [4-1:0] node23806;
	wire [4-1:0] node23807;
	wire [4-1:0] node23808;
	wire [4-1:0] node23812;
	wire [4-1:0] node23813;
	wire [4-1:0] node23816;
	wire [4-1:0] node23819;
	wire [4-1:0] node23820;
	wire [4-1:0] node23821;
	wire [4-1:0] node23824;
	wire [4-1:0] node23827;
	wire [4-1:0] node23828;
	wire [4-1:0] node23831;
	wire [4-1:0] node23834;
	wire [4-1:0] node23835;
	wire [4-1:0] node23836;
	wire [4-1:0] node23837;
	wire [4-1:0] node23838;
	wire [4-1:0] node23839;
	wire [4-1:0] node23842;
	wire [4-1:0] node23845;
	wire [4-1:0] node23846;
	wire [4-1:0] node23850;
	wire [4-1:0] node23851;
	wire [4-1:0] node23852;
	wire [4-1:0] node23855;
	wire [4-1:0] node23858;
	wire [4-1:0] node23859;
	wire [4-1:0] node23863;
	wire [4-1:0] node23864;
	wire [4-1:0] node23865;
	wire [4-1:0] node23866;
	wire [4-1:0] node23869;
	wire [4-1:0] node23872;
	wire [4-1:0] node23873;
	wire [4-1:0] node23876;
	wire [4-1:0] node23879;
	wire [4-1:0] node23880;
	wire [4-1:0] node23882;
	wire [4-1:0] node23885;
	wire [4-1:0] node23886;
	wire [4-1:0] node23889;
	wire [4-1:0] node23892;
	wire [4-1:0] node23893;
	wire [4-1:0] node23894;
	wire [4-1:0] node23895;
	wire [4-1:0] node23896;
	wire [4-1:0] node23899;
	wire [4-1:0] node23902;
	wire [4-1:0] node23903;
	wire [4-1:0] node23906;
	wire [4-1:0] node23909;
	wire [4-1:0] node23910;
	wire [4-1:0] node23911;
	wire [4-1:0] node23915;
	wire [4-1:0] node23916;
	wire [4-1:0] node23919;
	wire [4-1:0] node23922;
	wire [4-1:0] node23923;
	wire [4-1:0] node23924;
	wire [4-1:0] node23925;
	wire [4-1:0] node23928;
	wire [4-1:0] node23931;
	wire [4-1:0] node23932;
	wire [4-1:0] node23935;
	wire [4-1:0] node23938;
	wire [4-1:0] node23939;
	wire [4-1:0] node23940;
	wire [4-1:0] node23943;
	wire [4-1:0] node23946;
	wire [4-1:0] node23947;
	wire [4-1:0] node23950;
	wire [4-1:0] node23953;
	wire [4-1:0] node23954;
	wire [4-1:0] node23955;
	wire [4-1:0] node23956;
	wire [4-1:0] node23957;
	wire [4-1:0] node23958;
	wire [4-1:0] node23959;
	wire [4-1:0] node23962;
	wire [4-1:0] node23965;
	wire [4-1:0] node23966;
	wire [4-1:0] node23969;
	wire [4-1:0] node23972;
	wire [4-1:0] node23973;
	wire [4-1:0] node23974;
	wire [4-1:0] node23977;
	wire [4-1:0] node23980;
	wire [4-1:0] node23981;
	wire [4-1:0] node23984;
	wire [4-1:0] node23987;
	wire [4-1:0] node23988;
	wire [4-1:0] node23989;
	wire [4-1:0] node23990;
	wire [4-1:0] node23993;
	wire [4-1:0] node23996;
	wire [4-1:0] node23997;
	wire [4-1:0] node24000;
	wire [4-1:0] node24003;
	wire [4-1:0] node24004;
	wire [4-1:0] node24005;
	wire [4-1:0] node24008;
	wire [4-1:0] node24011;
	wire [4-1:0] node24012;
	wire [4-1:0] node24016;
	wire [4-1:0] node24017;
	wire [4-1:0] node24018;
	wire [4-1:0] node24019;
	wire [4-1:0] node24020;
	wire [4-1:0] node24023;
	wire [4-1:0] node24026;
	wire [4-1:0] node24027;
	wire [4-1:0] node24031;
	wire [4-1:0] node24032;
	wire [4-1:0] node24033;
	wire [4-1:0] node24036;
	wire [4-1:0] node24039;
	wire [4-1:0] node24040;
	wire [4-1:0] node24043;
	wire [4-1:0] node24046;
	wire [4-1:0] node24047;
	wire [4-1:0] node24048;
	wire [4-1:0] node24049;
	wire [4-1:0] node24052;
	wire [4-1:0] node24055;
	wire [4-1:0] node24056;
	wire [4-1:0] node24059;
	wire [4-1:0] node24062;
	wire [4-1:0] node24063;
	wire [4-1:0] node24064;
	wire [4-1:0] node24067;
	wire [4-1:0] node24070;
	wire [4-1:0] node24071;
	wire [4-1:0] node24074;
	wire [4-1:0] node24077;
	wire [4-1:0] node24078;
	wire [4-1:0] node24079;
	wire [4-1:0] node24080;
	wire [4-1:0] node24081;
	wire [4-1:0] node24082;
	wire [4-1:0] node24085;
	wire [4-1:0] node24088;
	wire [4-1:0] node24089;
	wire [4-1:0] node24093;
	wire [4-1:0] node24094;
	wire [4-1:0] node24097;
	wire [4-1:0] node24100;
	wire [4-1:0] node24101;
	wire [4-1:0] node24102;
	wire [4-1:0] node24103;
	wire [4-1:0] node24107;
	wire [4-1:0] node24108;
	wire [4-1:0] node24111;
	wire [4-1:0] node24114;
	wire [4-1:0] node24115;
	wire [4-1:0] node24116;
	wire [4-1:0] node24119;
	wire [4-1:0] node24122;
	wire [4-1:0] node24123;
	wire [4-1:0] node24126;
	wire [4-1:0] node24129;
	wire [4-1:0] node24130;
	wire [4-1:0] node24131;
	wire [4-1:0] node24132;
	wire [4-1:0] node24133;
	wire [4-1:0] node24136;
	wire [4-1:0] node24139;
	wire [4-1:0] node24140;
	wire [4-1:0] node24143;
	wire [4-1:0] node24146;
	wire [4-1:0] node24147;
	wire [4-1:0] node24148;
	wire [4-1:0] node24151;
	wire [4-1:0] node24154;
	wire [4-1:0] node24155;
	wire [4-1:0] node24158;
	wire [4-1:0] node24161;
	wire [4-1:0] node24162;
	wire [4-1:0] node24163;
	wire [4-1:0] node24164;
	wire [4-1:0] node24167;
	wire [4-1:0] node24170;
	wire [4-1:0] node24171;
	wire [4-1:0] node24174;
	wire [4-1:0] node24177;
	wire [4-1:0] node24178;
	wire [4-1:0] node24179;
	wire [4-1:0] node24182;
	wire [4-1:0] node24185;
	wire [4-1:0] node24186;
	wire [4-1:0] node24189;
	wire [4-1:0] node24192;
	wire [4-1:0] node24193;
	wire [4-1:0] node24194;
	wire [4-1:0] node24195;
	wire [4-1:0] node24196;
	wire [4-1:0] node24197;
	wire [4-1:0] node24198;
	wire [4-1:0] node24199;
	wire [4-1:0] node24200;
	wire [4-1:0] node24203;
	wire [4-1:0] node24206;
	wire [4-1:0] node24207;
	wire [4-1:0] node24210;
	wire [4-1:0] node24213;
	wire [4-1:0] node24214;
	wire [4-1:0] node24215;
	wire [4-1:0] node24218;
	wire [4-1:0] node24221;
	wire [4-1:0] node24222;
	wire [4-1:0] node24225;
	wire [4-1:0] node24228;
	wire [4-1:0] node24229;
	wire [4-1:0] node24230;
	wire [4-1:0] node24231;
	wire [4-1:0] node24234;
	wire [4-1:0] node24237;
	wire [4-1:0] node24238;
	wire [4-1:0] node24241;
	wire [4-1:0] node24244;
	wire [4-1:0] node24245;
	wire [4-1:0] node24248;
	wire [4-1:0] node24251;
	wire [4-1:0] node24252;
	wire [4-1:0] node24253;
	wire [4-1:0] node24254;
	wire [4-1:0] node24255;
	wire [4-1:0] node24258;
	wire [4-1:0] node24261;
	wire [4-1:0] node24263;
	wire [4-1:0] node24266;
	wire [4-1:0] node24267;
	wire [4-1:0] node24268;
	wire [4-1:0] node24271;
	wire [4-1:0] node24274;
	wire [4-1:0] node24275;
	wire [4-1:0] node24279;
	wire [4-1:0] node24280;
	wire [4-1:0] node24281;
	wire [4-1:0] node24282;
	wire [4-1:0] node24286;
	wire [4-1:0] node24287;
	wire [4-1:0] node24291;
	wire [4-1:0] node24292;
	wire [4-1:0] node24293;
	wire [4-1:0] node24297;
	wire [4-1:0] node24298;
	wire [4-1:0] node24302;
	wire [4-1:0] node24303;
	wire [4-1:0] node24304;
	wire [4-1:0] node24305;
	wire [4-1:0] node24306;
	wire [4-1:0] node24307;
	wire [4-1:0] node24310;
	wire [4-1:0] node24313;
	wire [4-1:0] node24314;
	wire [4-1:0] node24317;
	wire [4-1:0] node24320;
	wire [4-1:0] node24321;
	wire [4-1:0] node24322;
	wire [4-1:0] node24325;
	wire [4-1:0] node24328;
	wire [4-1:0] node24329;
	wire [4-1:0] node24332;
	wire [4-1:0] node24335;
	wire [4-1:0] node24336;
	wire [4-1:0] node24337;
	wire [4-1:0] node24338;
	wire [4-1:0] node24341;
	wire [4-1:0] node24344;
	wire [4-1:0] node24345;
	wire [4-1:0] node24348;
	wire [4-1:0] node24351;
	wire [4-1:0] node24352;
	wire [4-1:0] node24353;
	wire [4-1:0] node24356;
	wire [4-1:0] node24359;
	wire [4-1:0] node24360;
	wire [4-1:0] node24363;
	wire [4-1:0] node24366;
	wire [4-1:0] node24367;
	wire [4-1:0] node24368;
	wire [4-1:0] node24369;
	wire [4-1:0] node24370;
	wire [4-1:0] node24373;
	wire [4-1:0] node24376;
	wire [4-1:0] node24377;
	wire [4-1:0] node24380;
	wire [4-1:0] node24383;
	wire [4-1:0] node24384;
	wire [4-1:0] node24385;
	wire [4-1:0] node24388;
	wire [4-1:0] node24391;
	wire [4-1:0] node24392;
	wire [4-1:0] node24395;
	wire [4-1:0] node24398;
	wire [4-1:0] node24399;
	wire [4-1:0] node24400;
	wire [4-1:0] node24401;
	wire [4-1:0] node24405;
	wire [4-1:0] node24406;
	wire [4-1:0] node24409;
	wire [4-1:0] node24412;
	wire [4-1:0] node24413;
	wire [4-1:0] node24414;
	wire [4-1:0] node24417;
	wire [4-1:0] node24420;
	wire [4-1:0] node24421;
	wire [4-1:0] node24424;
	wire [4-1:0] node24427;
	wire [4-1:0] node24428;
	wire [4-1:0] node24429;
	wire [4-1:0] node24430;
	wire [4-1:0] node24431;
	wire [4-1:0] node24432;
	wire [4-1:0] node24434;
	wire [4-1:0] node24437;
	wire [4-1:0] node24438;
	wire [4-1:0] node24441;
	wire [4-1:0] node24444;
	wire [4-1:0] node24445;
	wire [4-1:0] node24446;
	wire [4-1:0] node24449;
	wire [4-1:0] node24452;
	wire [4-1:0] node24453;
	wire [4-1:0] node24457;
	wire [4-1:0] node24458;
	wire [4-1:0] node24459;
	wire [4-1:0] node24460;
	wire [4-1:0] node24464;
	wire [4-1:0] node24465;
	wire [4-1:0] node24469;
	wire [4-1:0] node24470;
	wire [4-1:0] node24471;
	wire [4-1:0] node24475;
	wire [4-1:0] node24477;
	wire [4-1:0] node24480;
	wire [4-1:0] node24481;
	wire [4-1:0] node24482;
	wire [4-1:0] node24483;
	wire [4-1:0] node24484;
	wire [4-1:0] node24487;
	wire [4-1:0] node24490;
	wire [4-1:0] node24491;
	wire [4-1:0] node24494;
	wire [4-1:0] node24497;
	wire [4-1:0] node24498;
	wire [4-1:0] node24500;
	wire [4-1:0] node24503;
	wire [4-1:0] node24504;
	wire [4-1:0] node24507;
	wire [4-1:0] node24510;
	wire [4-1:0] node24511;
	wire [4-1:0] node24512;
	wire [4-1:0] node24513;
	wire [4-1:0] node24517;
	wire [4-1:0] node24518;
	wire [4-1:0] node24522;
	wire [4-1:0] node24523;
	wire [4-1:0] node24524;
	wire [4-1:0] node24528;
	wire [4-1:0] node24529;
	wire [4-1:0] node24533;
	wire [4-1:0] node24534;
	wire [4-1:0] node24535;
	wire [4-1:0] node24536;
	wire [4-1:0] node24537;
	wire [4-1:0] node24539;
	wire [4-1:0] node24542;
	wire [4-1:0] node24543;
	wire [4-1:0] node24546;
	wire [4-1:0] node24549;
	wire [4-1:0] node24550;
	wire [4-1:0] node24551;
	wire [4-1:0] node24554;
	wire [4-1:0] node24557;
	wire [4-1:0] node24558;
	wire [4-1:0] node24561;
	wire [4-1:0] node24564;
	wire [4-1:0] node24565;
	wire [4-1:0] node24566;
	wire [4-1:0] node24567;
	wire [4-1:0] node24570;
	wire [4-1:0] node24573;
	wire [4-1:0] node24574;
	wire [4-1:0] node24577;
	wire [4-1:0] node24580;
	wire [4-1:0] node24581;
	wire [4-1:0] node24582;
	wire [4-1:0] node24585;
	wire [4-1:0] node24588;
	wire [4-1:0] node24589;
	wire [4-1:0] node24592;
	wire [4-1:0] node24595;
	wire [4-1:0] node24596;
	wire [4-1:0] node24597;
	wire [4-1:0] node24598;
	wire [4-1:0] node24599;
	wire [4-1:0] node24602;
	wire [4-1:0] node24605;
	wire [4-1:0] node24607;
	wire [4-1:0] node24610;
	wire [4-1:0] node24611;
	wire [4-1:0] node24613;
	wire [4-1:0] node24616;
	wire [4-1:0] node24617;
	wire [4-1:0] node24620;
	wire [4-1:0] node24623;
	wire [4-1:0] node24624;
	wire [4-1:0] node24625;
	wire [4-1:0] node24627;
	wire [4-1:0] node24630;
	wire [4-1:0] node24631;
	wire [4-1:0] node24634;
	wire [4-1:0] node24637;
	wire [4-1:0] node24638;
	wire [4-1:0] node24641;
	wire [4-1:0] node24644;
	wire [4-1:0] node24645;
	wire [4-1:0] node24646;
	wire [4-1:0] node24647;
	wire [4-1:0] node24648;
	wire [4-1:0] node24649;
	wire [4-1:0] node24650;
	wire [4-1:0] node24651;
	wire [4-1:0] node24655;
	wire [4-1:0] node24656;
	wire [4-1:0] node24659;
	wire [4-1:0] node24662;
	wire [4-1:0] node24663;
	wire [4-1:0] node24664;
	wire [4-1:0] node24667;
	wire [4-1:0] node24670;
	wire [4-1:0] node24671;
	wire [4-1:0] node24674;
	wire [4-1:0] node24677;
	wire [4-1:0] node24678;
	wire [4-1:0] node24679;
	wire [4-1:0] node24682;
	wire [4-1:0] node24683;
	wire [4-1:0] node24687;
	wire [4-1:0] node24688;
	wire [4-1:0] node24689;
	wire [4-1:0] node24693;
	wire [4-1:0] node24694;
	wire [4-1:0] node24698;
	wire [4-1:0] node24699;
	wire [4-1:0] node24700;
	wire [4-1:0] node24701;
	wire [4-1:0] node24702;
	wire [4-1:0] node24705;
	wire [4-1:0] node24708;
	wire [4-1:0] node24709;
	wire [4-1:0] node24712;
	wire [4-1:0] node24715;
	wire [4-1:0] node24716;
	wire [4-1:0] node24717;
	wire [4-1:0] node24721;
	wire [4-1:0] node24722;
	wire [4-1:0] node24725;
	wire [4-1:0] node24728;
	wire [4-1:0] node24729;
	wire [4-1:0] node24730;
	wire [4-1:0] node24731;
	wire [4-1:0] node24734;
	wire [4-1:0] node24737;
	wire [4-1:0] node24738;
	wire [4-1:0] node24741;
	wire [4-1:0] node24744;
	wire [4-1:0] node24745;
	wire [4-1:0] node24746;
	wire [4-1:0] node24750;
	wire [4-1:0] node24751;
	wire [4-1:0] node24754;
	wire [4-1:0] node24757;
	wire [4-1:0] node24758;
	wire [4-1:0] node24759;
	wire [4-1:0] node24760;
	wire [4-1:0] node24761;
	wire [4-1:0] node24762;
	wire [4-1:0] node24765;
	wire [4-1:0] node24768;
	wire [4-1:0] node24769;
	wire [4-1:0] node24772;
	wire [4-1:0] node24775;
	wire [4-1:0] node24776;
	wire [4-1:0] node24777;
	wire [4-1:0] node24780;
	wire [4-1:0] node24783;
	wire [4-1:0] node24784;
	wire [4-1:0] node24787;
	wire [4-1:0] node24790;
	wire [4-1:0] node24791;
	wire [4-1:0] node24792;
	wire [4-1:0] node24793;
	wire [4-1:0] node24796;
	wire [4-1:0] node24799;
	wire [4-1:0] node24800;
	wire [4-1:0] node24803;
	wire [4-1:0] node24806;
	wire [4-1:0] node24807;
	wire [4-1:0] node24810;
	wire [4-1:0] node24813;
	wire [4-1:0] node24814;
	wire [4-1:0] node24815;
	wire [4-1:0] node24816;
	wire [4-1:0] node24817;
	wire [4-1:0] node24820;
	wire [4-1:0] node24823;
	wire [4-1:0] node24824;
	wire [4-1:0] node24828;
	wire [4-1:0] node24829;
	wire [4-1:0] node24830;
	wire [4-1:0] node24833;
	wire [4-1:0] node24836;
	wire [4-1:0] node24838;
	wire [4-1:0] node24841;
	wire [4-1:0] node24842;
	wire [4-1:0] node24843;
	wire [4-1:0] node24844;
	wire [4-1:0] node24847;
	wire [4-1:0] node24850;
	wire [4-1:0] node24851;
	wire [4-1:0] node24854;
	wire [4-1:0] node24857;
	wire [4-1:0] node24858;
	wire [4-1:0] node24861;
	wire [4-1:0] node24864;
	wire [4-1:0] node24865;
	wire [4-1:0] node24866;
	wire [4-1:0] node24867;
	wire [4-1:0] node24868;
	wire [4-1:0] node24869;
	wire [4-1:0] node24870;
	wire [4-1:0] node24873;
	wire [4-1:0] node24876;
	wire [4-1:0] node24877;
	wire [4-1:0] node24880;
	wire [4-1:0] node24883;
	wire [4-1:0] node24884;
	wire [4-1:0] node24885;
	wire [4-1:0] node24888;
	wire [4-1:0] node24891;
	wire [4-1:0] node24892;
	wire [4-1:0] node24896;
	wire [4-1:0] node24897;
	wire [4-1:0] node24898;
	wire [4-1:0] node24899;
	wire [4-1:0] node24903;
	wire [4-1:0] node24904;
	wire [4-1:0] node24908;
	wire [4-1:0] node24909;
	wire [4-1:0] node24910;
	wire [4-1:0] node24914;
	wire [4-1:0] node24915;
	wire [4-1:0] node24919;
	wire [4-1:0] node24920;
	wire [4-1:0] node24921;
	wire [4-1:0] node24922;
	wire [4-1:0] node24923;
	wire [4-1:0] node24926;
	wire [4-1:0] node24929;
	wire [4-1:0] node24930;
	wire [4-1:0] node24933;
	wire [4-1:0] node24936;
	wire [4-1:0] node24937;
	wire [4-1:0] node24938;
	wire [4-1:0] node24941;
	wire [4-1:0] node24944;
	wire [4-1:0] node24945;
	wire [4-1:0] node24948;
	wire [4-1:0] node24951;
	wire [4-1:0] node24952;
	wire [4-1:0] node24953;
	wire [4-1:0] node24954;
	wire [4-1:0] node24957;
	wire [4-1:0] node24960;
	wire [4-1:0] node24961;
	wire [4-1:0] node24964;
	wire [4-1:0] node24967;
	wire [4-1:0] node24968;
	wire [4-1:0] node24971;
	wire [4-1:0] node24974;
	wire [4-1:0] node24975;
	wire [4-1:0] node24976;
	wire [4-1:0] node24977;
	wire [4-1:0] node24978;
	wire [4-1:0] node24979;
	wire [4-1:0] node24982;
	wire [4-1:0] node24985;
	wire [4-1:0] node24986;
	wire [4-1:0] node24989;
	wire [4-1:0] node24992;
	wire [4-1:0] node24993;
	wire [4-1:0] node24994;
	wire [4-1:0] node24997;
	wire [4-1:0] node25000;
	wire [4-1:0] node25001;
	wire [4-1:0] node25004;
	wire [4-1:0] node25007;
	wire [4-1:0] node25008;
	wire [4-1:0] node25009;
	wire [4-1:0] node25010;
	wire [4-1:0] node25014;
	wire [4-1:0] node25015;
	wire [4-1:0] node25019;
	wire [4-1:0] node25020;
	wire [4-1:0] node25021;
	wire [4-1:0] node25025;
	wire [4-1:0] node25026;
	wire [4-1:0] node25030;
	wire [4-1:0] node25031;
	wire [4-1:0] node25032;
	wire [4-1:0] node25033;
	wire [4-1:0] node25034;
	wire [4-1:0] node25038;
	wire [4-1:0] node25039;
	wire [4-1:0] node25042;
	wire [4-1:0] node25045;
	wire [4-1:0] node25046;
	wire [4-1:0] node25047;
	wire [4-1:0] node25050;
	wire [4-1:0] node25053;
	wire [4-1:0] node25054;
	wire [4-1:0] node25057;
	wire [4-1:0] node25060;
	wire [4-1:0] node25061;
	wire [4-1:0] node25062;
	wire [4-1:0] node25063;
	wire [4-1:0] node25067;
	wire [4-1:0] node25068;
	wire [4-1:0] node25072;
	wire [4-1:0] node25073;
	wire [4-1:0] node25074;
	wire [4-1:0] node25078;
	wire [4-1:0] node25079;
	wire [4-1:0] node25083;
	wire [4-1:0] node25084;
	wire [4-1:0] node25085;
	wire [4-1:0] node25086;
	wire [4-1:0] node25087;
	wire [4-1:0] node25088;
	wire [4-1:0] node25089;
	wire [4-1:0] node25090;
	wire [4-1:0] node25091;
	wire [4-1:0] node25092;
	wire [4-1:0] node25093;
	wire [4-1:0] node25096;
	wire [4-1:0] node25099;
	wire [4-1:0] node25100;
	wire [4-1:0] node25104;
	wire [4-1:0] node25105;
	wire [4-1:0] node25106;
	wire [4-1:0] node25109;
	wire [4-1:0] node25112;
	wire [4-1:0] node25113;
	wire [4-1:0] node25116;
	wire [4-1:0] node25119;
	wire [4-1:0] node25120;
	wire [4-1:0] node25121;
	wire [4-1:0] node25122;
	wire [4-1:0] node25125;
	wire [4-1:0] node25128;
	wire [4-1:0] node25129;
	wire [4-1:0] node25132;
	wire [4-1:0] node25135;
	wire [4-1:0] node25136;
	wire [4-1:0] node25137;
	wire [4-1:0] node25140;
	wire [4-1:0] node25143;
	wire [4-1:0] node25144;
	wire [4-1:0] node25147;
	wire [4-1:0] node25150;
	wire [4-1:0] node25151;
	wire [4-1:0] node25152;
	wire [4-1:0] node25153;
	wire [4-1:0] node25154;
	wire [4-1:0] node25157;
	wire [4-1:0] node25160;
	wire [4-1:0] node25161;
	wire [4-1:0] node25164;
	wire [4-1:0] node25167;
	wire [4-1:0] node25168;
	wire [4-1:0] node25169;
	wire [4-1:0] node25173;
	wire [4-1:0] node25174;
	wire [4-1:0] node25177;
	wire [4-1:0] node25180;
	wire [4-1:0] node25181;
	wire [4-1:0] node25182;
	wire [4-1:0] node25183;
	wire [4-1:0] node25186;
	wire [4-1:0] node25189;
	wire [4-1:0] node25190;
	wire [4-1:0] node25193;
	wire [4-1:0] node25196;
	wire [4-1:0] node25197;
	wire [4-1:0] node25198;
	wire [4-1:0] node25201;
	wire [4-1:0] node25204;
	wire [4-1:0] node25205;
	wire [4-1:0] node25208;
	wire [4-1:0] node25211;
	wire [4-1:0] node25212;
	wire [4-1:0] node25213;
	wire [4-1:0] node25214;
	wire [4-1:0] node25215;
	wire [4-1:0] node25216;
	wire [4-1:0] node25219;
	wire [4-1:0] node25222;
	wire [4-1:0] node25224;
	wire [4-1:0] node25227;
	wire [4-1:0] node25228;
	wire [4-1:0] node25229;
	wire [4-1:0] node25232;
	wire [4-1:0] node25235;
	wire [4-1:0] node25236;
	wire [4-1:0] node25239;
	wire [4-1:0] node25242;
	wire [4-1:0] node25243;
	wire [4-1:0] node25244;
	wire [4-1:0] node25245;
	wire [4-1:0] node25248;
	wire [4-1:0] node25251;
	wire [4-1:0] node25252;
	wire [4-1:0] node25255;
	wire [4-1:0] node25258;
	wire [4-1:0] node25259;
	wire [4-1:0] node25260;
	wire [4-1:0] node25263;
	wire [4-1:0] node25266;
	wire [4-1:0] node25267;
	wire [4-1:0] node25270;
	wire [4-1:0] node25273;
	wire [4-1:0] node25274;
	wire [4-1:0] node25275;
	wire [4-1:0] node25276;
	wire [4-1:0] node25277;
	wire [4-1:0] node25280;
	wire [4-1:0] node25283;
	wire [4-1:0] node25284;
	wire [4-1:0] node25288;
	wire [4-1:0] node25289;
	wire [4-1:0] node25290;
	wire [4-1:0] node25293;
	wire [4-1:0] node25296;
	wire [4-1:0] node25297;
	wire [4-1:0] node25300;
	wire [4-1:0] node25303;
	wire [4-1:0] node25304;
	wire [4-1:0] node25305;
	wire [4-1:0] node25306;
	wire [4-1:0] node25309;
	wire [4-1:0] node25312;
	wire [4-1:0] node25313;
	wire [4-1:0] node25316;
	wire [4-1:0] node25319;
	wire [4-1:0] node25320;
	wire [4-1:0] node25323;
	wire [4-1:0] node25326;
	wire [4-1:0] node25327;
	wire [4-1:0] node25328;
	wire [4-1:0] node25329;
	wire [4-1:0] node25330;
	wire [4-1:0] node25331;
	wire [4-1:0] node25332;
	wire [4-1:0] node25335;
	wire [4-1:0] node25338;
	wire [4-1:0] node25339;
	wire [4-1:0] node25342;
	wire [4-1:0] node25345;
	wire [4-1:0] node25346;
	wire [4-1:0] node25348;
	wire [4-1:0] node25351;
	wire [4-1:0] node25352;
	wire [4-1:0] node25355;
	wire [4-1:0] node25358;
	wire [4-1:0] node25359;
	wire [4-1:0] node25360;
	wire [4-1:0] node25361;
	wire [4-1:0] node25364;
	wire [4-1:0] node25367;
	wire [4-1:0] node25368;
	wire [4-1:0] node25371;
	wire [4-1:0] node25374;
	wire [4-1:0] node25375;
	wire [4-1:0] node25376;
	wire [4-1:0] node25379;
	wire [4-1:0] node25382;
	wire [4-1:0] node25383;
	wire [4-1:0] node25386;
	wire [4-1:0] node25389;
	wire [4-1:0] node25390;
	wire [4-1:0] node25391;
	wire [4-1:0] node25392;
	wire [4-1:0] node25394;
	wire [4-1:0] node25397;
	wire [4-1:0] node25398;
	wire [4-1:0] node25401;
	wire [4-1:0] node25404;
	wire [4-1:0] node25405;
	wire [4-1:0] node25406;
	wire [4-1:0] node25409;
	wire [4-1:0] node25412;
	wire [4-1:0] node25413;
	wire [4-1:0] node25416;
	wire [4-1:0] node25419;
	wire [4-1:0] node25420;
	wire [4-1:0] node25421;
	wire [4-1:0] node25422;
	wire [4-1:0] node25426;
	wire [4-1:0] node25427;
	wire [4-1:0] node25431;
	wire [4-1:0] node25433;
	wire [4-1:0] node25434;
	wire [4-1:0] node25438;
	wire [4-1:0] node25439;
	wire [4-1:0] node25440;
	wire [4-1:0] node25441;
	wire [4-1:0] node25442;
	wire [4-1:0] node25443;
	wire [4-1:0] node25446;
	wire [4-1:0] node25449;
	wire [4-1:0] node25450;
	wire [4-1:0] node25453;
	wire [4-1:0] node25456;
	wire [4-1:0] node25457;
	wire [4-1:0] node25458;
	wire [4-1:0] node25461;
	wire [4-1:0] node25464;
	wire [4-1:0] node25465;
	wire [4-1:0] node25468;
	wire [4-1:0] node25471;
	wire [4-1:0] node25472;
	wire [4-1:0] node25473;
	wire [4-1:0] node25474;
	wire [4-1:0] node25477;
	wire [4-1:0] node25480;
	wire [4-1:0] node25481;
	wire [4-1:0] node25484;
	wire [4-1:0] node25487;
	wire [4-1:0] node25488;
	wire [4-1:0] node25489;
	wire [4-1:0] node25492;
	wire [4-1:0] node25495;
	wire [4-1:0] node25496;
	wire [4-1:0] node25499;
	wire [4-1:0] node25502;
	wire [4-1:0] node25503;
	wire [4-1:0] node25504;
	wire [4-1:0] node25505;
	wire [4-1:0] node25506;
	wire [4-1:0] node25510;
	wire [4-1:0] node25511;
	wire [4-1:0] node25514;
	wire [4-1:0] node25517;
	wire [4-1:0] node25518;
	wire [4-1:0] node25519;
	wire [4-1:0] node25522;
	wire [4-1:0] node25525;
	wire [4-1:0] node25526;
	wire [4-1:0] node25529;
	wire [4-1:0] node25532;
	wire [4-1:0] node25533;
	wire [4-1:0] node25534;
	wire [4-1:0] node25535;
	wire [4-1:0] node25539;
	wire [4-1:0] node25540;
	wire [4-1:0] node25543;
	wire [4-1:0] node25546;
	wire [4-1:0] node25547;
	wire [4-1:0] node25548;
	wire [4-1:0] node25551;
	wire [4-1:0] node25554;
	wire [4-1:0] node25555;
	wire [4-1:0] node25558;
	wire [4-1:0] node25561;
	wire [4-1:0] node25562;
	wire [4-1:0] node25563;
	wire [4-1:0] node25564;
	wire [4-1:0] node25565;
	wire [4-1:0] node25566;
	wire [4-1:0] node25567;
	wire [4-1:0] node25571;
	wire [4-1:0] node25572;
	wire [4-1:0] node25573;
	wire [4-1:0] node25577;
	wire [4-1:0] node25578;
	wire [4-1:0] node25582;
	wire [4-1:0] node25583;
	wire [4-1:0] node25584;
	wire [4-1:0] node25585;
	wire [4-1:0] node25589;
	wire [4-1:0] node25590;
	wire [4-1:0] node25594;
	wire [4-1:0] node25595;
	wire [4-1:0] node25596;
	wire [4-1:0] node25600;
	wire [4-1:0] node25601;
	wire [4-1:0] node25605;
	wire [4-1:0] node25606;
	wire [4-1:0] node25607;
	wire [4-1:0] node25608;
	wire [4-1:0] node25609;
	wire [4-1:0] node25612;
	wire [4-1:0] node25615;
	wire [4-1:0] node25616;
	wire [4-1:0] node25619;
	wire [4-1:0] node25622;
	wire [4-1:0] node25623;
	wire [4-1:0] node25626;
	wire [4-1:0] node25629;
	wire [4-1:0] node25630;
	wire [4-1:0] node25631;
	wire [4-1:0] node25632;
	wire [4-1:0] node25636;
	wire [4-1:0] node25637;
	wire [4-1:0] node25641;
	wire [4-1:0] node25642;
	wire [4-1:0] node25643;
	wire [4-1:0] node25647;
	wire [4-1:0] node25648;
	wire [4-1:0] node25652;
	wire [4-1:0] node25653;
	wire [4-1:0] node25654;
	wire [4-1:0] node25655;
	wire [4-1:0] node25656;
	wire [4-1:0] node25657;
	wire [4-1:0] node25660;
	wire [4-1:0] node25663;
	wire [4-1:0] node25664;
	wire [4-1:0] node25667;
	wire [4-1:0] node25670;
	wire [4-1:0] node25671;
	wire [4-1:0] node25673;
	wire [4-1:0] node25676;
	wire [4-1:0] node25677;
	wire [4-1:0] node25680;
	wire [4-1:0] node25683;
	wire [4-1:0] node25684;
	wire [4-1:0] node25685;
	wire [4-1:0] node25686;
	wire [4-1:0] node25690;
	wire [4-1:0] node25691;
	wire [4-1:0] node25695;
	wire [4-1:0] node25696;
	wire [4-1:0] node25697;
	wire [4-1:0] node25701;
	wire [4-1:0] node25702;
	wire [4-1:0] node25706;
	wire [4-1:0] node25707;
	wire [4-1:0] node25708;
	wire [4-1:0] node25709;
	wire [4-1:0] node25710;
	wire [4-1:0] node25713;
	wire [4-1:0] node25716;
	wire [4-1:0] node25717;
	wire [4-1:0] node25720;
	wire [4-1:0] node25723;
	wire [4-1:0] node25724;
	wire [4-1:0] node25725;
	wire [4-1:0] node25728;
	wire [4-1:0] node25731;
	wire [4-1:0] node25732;
	wire [4-1:0] node25735;
	wire [4-1:0] node25738;
	wire [4-1:0] node25739;
	wire [4-1:0] node25740;
	wire [4-1:0] node25741;
	wire [4-1:0] node25745;
	wire [4-1:0] node25746;
	wire [4-1:0] node25750;
	wire [4-1:0] node25751;
	wire [4-1:0] node25752;
	wire [4-1:0] node25756;
	wire [4-1:0] node25757;
	wire [4-1:0] node25761;
	wire [4-1:0] node25762;
	wire [4-1:0] node25763;
	wire [4-1:0] node25764;
	wire [4-1:0] node25765;
	wire [4-1:0] node25766;
	wire [4-1:0] node25767;
	wire [4-1:0] node25770;
	wire [4-1:0] node25773;
	wire [4-1:0] node25775;
	wire [4-1:0] node25778;
	wire [4-1:0] node25779;
	wire [4-1:0] node25780;
	wire [4-1:0] node25783;
	wire [4-1:0] node25786;
	wire [4-1:0] node25787;
	wire [4-1:0] node25790;
	wire [4-1:0] node25793;
	wire [4-1:0] node25794;
	wire [4-1:0] node25795;
	wire [4-1:0] node25796;
	wire [4-1:0] node25799;
	wire [4-1:0] node25802;
	wire [4-1:0] node25803;
	wire [4-1:0] node25806;
	wire [4-1:0] node25809;
	wire [4-1:0] node25810;
	wire [4-1:0] node25811;
	wire [4-1:0] node25814;
	wire [4-1:0] node25817;
	wire [4-1:0] node25818;
	wire [4-1:0] node25821;
	wire [4-1:0] node25824;
	wire [4-1:0] node25825;
	wire [4-1:0] node25826;
	wire [4-1:0] node25827;
	wire [4-1:0] node25828;
	wire [4-1:0] node25831;
	wire [4-1:0] node25834;
	wire [4-1:0] node25835;
	wire [4-1:0] node25838;
	wire [4-1:0] node25841;
	wire [4-1:0] node25842;
	wire [4-1:0] node25845;
	wire [4-1:0] node25848;
	wire [4-1:0] node25849;
	wire [4-1:0] node25852;
	wire [4-1:0] node25855;
	wire [4-1:0] node25856;
	wire [4-1:0] node25857;
	wire [4-1:0] node25858;
	wire [4-1:0] node25859;
	wire [4-1:0] node25860;
	wire [4-1:0] node25863;
	wire [4-1:0] node25866;
	wire [4-1:0] node25867;
	wire [4-1:0] node25871;
	wire [4-1:0] node25872;
	wire [4-1:0] node25875;
	wire [4-1:0] node25878;
	wire [4-1:0] node25879;
	wire [4-1:0] node25882;
	wire [4-1:0] node25885;
	wire [4-1:0] node25886;
	wire [4-1:0] node25887;
	wire [4-1:0] node25888;
	wire [4-1:0] node25891;
	wire [4-1:0] node25894;
	wire [4-1:0] node25895;
	wire [4-1:0] node25896;
	wire [4-1:0] node25899;
	wire [4-1:0] node25902;
	wire [4-1:0] node25903;
	wire [4-1:0] node25906;
	wire [4-1:0] node25909;
	wire [4-1:0] node25910;
	wire [4-1:0] node25913;
	wire [4-1:0] node25916;
	wire [4-1:0] node25917;
	wire [4-1:0] node25918;
	wire [4-1:0] node25919;
	wire [4-1:0] node25920;
	wire [4-1:0] node25921;
	wire [4-1:0] node25922;
	wire [4-1:0] node25923;
	wire [4-1:0] node25924;
	wire [4-1:0] node25927;
	wire [4-1:0] node25930;
	wire [4-1:0] node25931;
	wire [4-1:0] node25935;
	wire [4-1:0] node25936;
	wire [4-1:0] node25937;
	wire [4-1:0] node25940;
	wire [4-1:0] node25943;
	wire [4-1:0] node25944;
	wire [4-1:0] node25948;
	wire [4-1:0] node25949;
	wire [4-1:0] node25950;
	wire [4-1:0] node25951;
	wire [4-1:0] node25954;
	wire [4-1:0] node25957;
	wire [4-1:0] node25958;
	wire [4-1:0] node25961;
	wire [4-1:0] node25964;
	wire [4-1:0] node25965;
	wire [4-1:0] node25966;
	wire [4-1:0] node25969;
	wire [4-1:0] node25972;
	wire [4-1:0] node25973;
	wire [4-1:0] node25976;
	wire [4-1:0] node25979;
	wire [4-1:0] node25980;
	wire [4-1:0] node25981;
	wire [4-1:0] node25982;
	wire [4-1:0] node25983;
	wire [4-1:0] node25986;
	wire [4-1:0] node25989;
	wire [4-1:0] node25990;
	wire [4-1:0] node25993;
	wire [4-1:0] node25996;
	wire [4-1:0] node25997;
	wire [4-1:0] node25998;
	wire [4-1:0] node26001;
	wire [4-1:0] node26004;
	wire [4-1:0] node26005;
	wire [4-1:0] node26008;
	wire [4-1:0] node26011;
	wire [4-1:0] node26012;
	wire [4-1:0] node26013;
	wire [4-1:0] node26014;
	wire [4-1:0] node26018;
	wire [4-1:0] node26019;
	wire [4-1:0] node26022;
	wire [4-1:0] node26025;
	wire [4-1:0] node26026;
	wire [4-1:0] node26027;
	wire [4-1:0] node26030;
	wire [4-1:0] node26033;
	wire [4-1:0] node26034;
	wire [4-1:0] node26037;
	wire [4-1:0] node26040;
	wire [4-1:0] node26041;
	wire [4-1:0] node26042;
	wire [4-1:0] node26043;
	wire [4-1:0] node26044;
	wire [4-1:0] node26045;
	wire [4-1:0] node26048;
	wire [4-1:0] node26051;
	wire [4-1:0] node26052;
	wire [4-1:0] node26055;
	wire [4-1:0] node26058;
	wire [4-1:0] node26059;
	wire [4-1:0] node26060;
	wire [4-1:0] node26063;
	wire [4-1:0] node26066;
	wire [4-1:0] node26067;
	wire [4-1:0] node26070;
	wire [4-1:0] node26073;
	wire [4-1:0] node26074;
	wire [4-1:0] node26075;
	wire [4-1:0] node26076;
	wire [4-1:0] node26079;
	wire [4-1:0] node26082;
	wire [4-1:0] node26084;
	wire [4-1:0] node26087;
	wire [4-1:0] node26088;
	wire [4-1:0] node26089;
	wire [4-1:0] node26092;
	wire [4-1:0] node26095;
	wire [4-1:0] node26096;
	wire [4-1:0] node26100;
	wire [4-1:0] node26101;
	wire [4-1:0] node26102;
	wire [4-1:0] node26103;
	wire [4-1:0] node26104;
	wire [4-1:0] node26107;
	wire [4-1:0] node26110;
	wire [4-1:0] node26111;
	wire [4-1:0] node26114;
	wire [4-1:0] node26117;
	wire [4-1:0] node26118;
	wire [4-1:0] node26120;
	wire [4-1:0] node26123;
	wire [4-1:0] node26125;
	wire [4-1:0] node26128;
	wire [4-1:0] node26129;
	wire [4-1:0] node26130;
	wire [4-1:0] node26131;
	wire [4-1:0] node26134;
	wire [4-1:0] node26137;
	wire [4-1:0] node26138;
	wire [4-1:0] node26141;
	wire [4-1:0] node26144;
	wire [4-1:0] node26145;
	wire [4-1:0] node26146;
	wire [4-1:0] node26149;
	wire [4-1:0] node26152;
	wire [4-1:0] node26153;
	wire [4-1:0] node26156;
	wire [4-1:0] node26159;
	wire [4-1:0] node26160;
	wire [4-1:0] node26161;
	wire [4-1:0] node26162;
	wire [4-1:0] node26163;
	wire [4-1:0] node26164;
	wire [4-1:0] node26165;
	wire [4-1:0] node26168;
	wire [4-1:0] node26171;
	wire [4-1:0] node26172;
	wire [4-1:0] node26175;
	wire [4-1:0] node26178;
	wire [4-1:0] node26179;
	wire [4-1:0] node26182;
	wire [4-1:0] node26185;
	wire [4-1:0] node26186;
	wire [4-1:0] node26187;
	wire [4-1:0] node26188;
	wire [4-1:0] node26191;
	wire [4-1:0] node26194;
	wire [4-1:0] node26195;
	wire [4-1:0] node26198;
	wire [4-1:0] node26201;
	wire [4-1:0] node26202;
	wire [4-1:0] node26203;
	wire [4-1:0] node26206;
	wire [4-1:0] node26209;
	wire [4-1:0] node26210;
	wire [4-1:0] node26213;
	wire [4-1:0] node26216;
	wire [4-1:0] node26217;
	wire [4-1:0] node26218;
	wire [4-1:0] node26219;
	wire [4-1:0] node26220;
	wire [4-1:0] node26223;
	wire [4-1:0] node26226;
	wire [4-1:0] node26227;
	wire [4-1:0] node26230;
	wire [4-1:0] node26233;
	wire [4-1:0] node26234;
	wire [4-1:0] node26235;
	wire [4-1:0] node26239;
	wire [4-1:0] node26240;
	wire [4-1:0] node26243;
	wire [4-1:0] node26246;
	wire [4-1:0] node26247;
	wire [4-1:0] node26248;
	wire [4-1:0] node26249;
	wire [4-1:0] node26252;
	wire [4-1:0] node26255;
	wire [4-1:0] node26256;
	wire [4-1:0] node26259;
	wire [4-1:0] node26262;
	wire [4-1:0] node26263;
	wire [4-1:0] node26264;
	wire [4-1:0] node26267;
	wire [4-1:0] node26270;
	wire [4-1:0] node26271;
	wire [4-1:0] node26274;
	wire [4-1:0] node26277;
	wire [4-1:0] node26278;
	wire [4-1:0] node26279;
	wire [4-1:0] node26280;
	wire [4-1:0] node26281;
	wire [4-1:0] node26282;
	wire [4-1:0] node26285;
	wire [4-1:0] node26288;
	wire [4-1:0] node26289;
	wire [4-1:0] node26293;
	wire [4-1:0] node26294;
	wire [4-1:0] node26296;
	wire [4-1:0] node26299;
	wire [4-1:0] node26300;
	wire [4-1:0] node26303;
	wire [4-1:0] node26306;
	wire [4-1:0] node26307;
	wire [4-1:0] node26308;
	wire [4-1:0] node26309;
	wire [4-1:0] node26312;
	wire [4-1:0] node26315;
	wire [4-1:0] node26317;
	wire [4-1:0] node26320;
	wire [4-1:0] node26321;
	wire [4-1:0] node26323;
	wire [4-1:0] node26326;
	wire [4-1:0] node26327;
	wire [4-1:0] node26330;
	wire [4-1:0] node26333;
	wire [4-1:0] node26334;
	wire [4-1:0] node26335;
	wire [4-1:0] node26336;
	wire [4-1:0] node26337;
	wire [4-1:0] node26340;
	wire [4-1:0] node26343;
	wire [4-1:0] node26344;
	wire [4-1:0] node26347;
	wire [4-1:0] node26350;
	wire [4-1:0] node26351;
	wire [4-1:0] node26353;
	wire [4-1:0] node26356;
	wire [4-1:0] node26357;
	wire [4-1:0] node26360;
	wire [4-1:0] node26363;
	wire [4-1:0] node26364;
	wire [4-1:0] node26365;
	wire [4-1:0] node26366;
	wire [4-1:0] node26369;
	wire [4-1:0] node26372;
	wire [4-1:0] node26373;
	wire [4-1:0] node26376;
	wire [4-1:0] node26379;
	wire [4-1:0] node26380;
	wire [4-1:0] node26381;
	wire [4-1:0] node26384;
	wire [4-1:0] node26387;
	wire [4-1:0] node26388;
	wire [4-1:0] node26391;
	wire [4-1:0] node26394;
	wire [4-1:0] node26395;
	wire [4-1:0] node26396;
	wire [4-1:0] node26397;
	wire [4-1:0] node26398;
	wire [4-1:0] node26399;
	wire [4-1:0] node26400;
	wire [4-1:0] node26402;
	wire [4-1:0] node26405;
	wire [4-1:0] node26407;
	wire [4-1:0] node26410;
	wire [4-1:0] node26411;
	wire [4-1:0] node26413;
	wire [4-1:0] node26416;
	wire [4-1:0] node26418;
	wire [4-1:0] node26421;
	wire [4-1:0] node26422;
	wire [4-1:0] node26423;
	wire [4-1:0] node26424;
	wire [4-1:0] node26428;
	wire [4-1:0] node26429;
	wire [4-1:0] node26432;
	wire [4-1:0] node26435;
	wire [4-1:0] node26436;
	wire [4-1:0] node26438;
	wire [4-1:0] node26441;
	wire [4-1:0] node26442;
	wire [4-1:0] node26445;
	wire [4-1:0] node26448;
	wire [4-1:0] node26449;
	wire [4-1:0] node26450;
	wire [4-1:0] node26452;
	wire [4-1:0] node26455;
	wire [4-1:0] node26457;
	wire [4-1:0] node26460;
	wire [4-1:0] node26461;
	wire [4-1:0] node26463;
	wire [4-1:0] node26466;
	wire [4-1:0] node26468;
	wire [4-1:0] node26471;
	wire [4-1:0] node26472;
	wire [4-1:0] node26473;
	wire [4-1:0] node26474;
	wire [4-1:0] node26475;
	wire [4-1:0] node26476;
	wire [4-1:0] node26479;
	wire [4-1:0] node26482;
	wire [4-1:0] node26483;
	wire [4-1:0] node26486;
	wire [4-1:0] node26489;
	wire [4-1:0] node26490;
	wire [4-1:0] node26491;
	wire [4-1:0] node26494;
	wire [4-1:0] node26497;
	wire [4-1:0] node26498;
	wire [4-1:0] node26501;
	wire [4-1:0] node26504;
	wire [4-1:0] node26505;
	wire [4-1:0] node26506;
	wire [4-1:0] node26507;
	wire [4-1:0] node26510;
	wire [4-1:0] node26513;
	wire [4-1:0] node26514;
	wire [4-1:0] node26517;
	wire [4-1:0] node26520;
	wire [4-1:0] node26521;
	wire [4-1:0] node26522;
	wire [4-1:0] node26525;
	wire [4-1:0] node26528;
	wire [4-1:0] node26529;
	wire [4-1:0] node26532;
	wire [4-1:0] node26535;
	wire [4-1:0] node26536;
	wire [4-1:0] node26537;
	wire [4-1:0] node26538;
	wire [4-1:0] node26541;
	wire [4-1:0] node26544;
	wire [4-1:0] node26545;
	wire [4-1:0] node26548;
	wire [4-1:0] node26551;
	wire [4-1:0] node26552;
	wire [4-1:0] node26553;
	wire [4-1:0] node26556;
	wire [4-1:0] node26559;
	wire [4-1:0] node26560;
	wire [4-1:0] node26563;
	wire [4-1:0] node26566;
	wire [4-1:0] node26567;
	wire [4-1:0] node26568;
	wire [4-1:0] node26569;
	wire [4-1:0] node26570;
	wire [4-1:0] node26571;
	wire [4-1:0] node26572;
	wire [4-1:0] node26575;
	wire [4-1:0] node26578;
	wire [4-1:0] node26579;
	wire [4-1:0] node26582;
	wire [4-1:0] node26585;
	wire [4-1:0] node26586;
	wire [4-1:0] node26587;
	wire [4-1:0] node26590;
	wire [4-1:0] node26593;
	wire [4-1:0] node26594;
	wire [4-1:0] node26597;
	wire [4-1:0] node26600;
	wire [4-1:0] node26601;
	wire [4-1:0] node26602;
	wire [4-1:0] node26603;
	wire [4-1:0] node26607;
	wire [4-1:0] node26608;
	wire [4-1:0] node26612;
	wire [4-1:0] node26613;
	wire [4-1:0] node26614;
	wire [4-1:0] node26618;
	wire [4-1:0] node26619;
	wire [4-1:0] node26623;
	wire [4-1:0] node26624;
	wire [4-1:0] node26625;
	wire [4-1:0] node26626;
	wire [4-1:0] node26627;
	wire [4-1:0] node26631;
	wire [4-1:0] node26632;
	wire [4-1:0] node26636;
	wire [4-1:0] node26637;
	wire [4-1:0] node26638;
	wire [4-1:0] node26642;
	wire [4-1:0] node26643;
	wire [4-1:0] node26647;
	wire [4-1:0] node26648;
	wire [4-1:0] node26649;
	wire [4-1:0] node26651;
	wire [4-1:0] node26655;
	wire [4-1:0] node26656;
	wire [4-1:0] node26657;
	wire [4-1:0] node26661;
	wire [4-1:0] node26662;
	wire [4-1:0] node26666;
	wire [4-1:0] node26667;
	wire [4-1:0] node26668;
	wire [4-1:0] node26669;
	wire [4-1:0] node26670;
	wire [4-1:0] node26671;
	wire [4-1:0] node26674;
	wire [4-1:0] node26677;
	wire [4-1:0] node26678;
	wire [4-1:0] node26681;
	wire [4-1:0] node26684;
	wire [4-1:0] node26685;
	wire [4-1:0] node26686;
	wire [4-1:0] node26689;
	wire [4-1:0] node26692;
	wire [4-1:0] node26693;
	wire [4-1:0] node26696;
	wire [4-1:0] node26699;
	wire [4-1:0] node26700;
	wire [4-1:0] node26701;
	wire [4-1:0] node26702;
	wire [4-1:0] node26706;
	wire [4-1:0] node26707;
	wire [4-1:0] node26711;
	wire [4-1:0] node26712;
	wire [4-1:0] node26713;
	wire [4-1:0] node26717;
	wire [4-1:0] node26718;
	wire [4-1:0] node26722;
	wire [4-1:0] node26723;
	wire [4-1:0] node26724;
	wire [4-1:0] node26725;
	wire [4-1:0] node26726;
	wire [4-1:0] node26729;
	wire [4-1:0] node26732;
	wire [4-1:0] node26733;
	wire [4-1:0] node26736;
	wire [4-1:0] node26739;
	wire [4-1:0] node26740;
	wire [4-1:0] node26743;
	wire [4-1:0] node26746;
	wire [4-1:0] node26747;
	wire [4-1:0] node26748;
	wire [4-1:0] node26749;
	wire [4-1:0] node26752;
	wire [4-1:0] node26755;
	wire [4-1:0] node26757;
	wire [4-1:0] node26760;
	wire [4-1:0] node26761;
	wire [4-1:0] node26762;
	wire [4-1:0] node26765;
	wire [4-1:0] node26768;
	wire [4-1:0] node26769;
	wire [4-1:0] node26772;
	wire [4-1:0] node26775;
	wire [4-1:0] node26776;
	wire [4-1:0] node26777;
	wire [4-1:0] node26778;
	wire [4-1:0] node26779;
	wire [4-1:0] node26780;
	wire [4-1:0] node26781;
	wire [4-1:0] node26782;
	wire [4-1:0] node26783;
	wire [4-1:0] node26784;
	wire [4-1:0] node26787;
	wire [4-1:0] node26790;
	wire [4-1:0] node26791;
	wire [4-1:0] node26794;
	wire [4-1:0] node26797;
	wire [4-1:0] node26798;
	wire [4-1:0] node26799;
	wire [4-1:0] node26802;
	wire [4-1:0] node26805;
	wire [4-1:0] node26807;
	wire [4-1:0] node26810;
	wire [4-1:0] node26811;
	wire [4-1:0] node26812;
	wire [4-1:0] node26813;
	wire [4-1:0] node26816;
	wire [4-1:0] node26819;
	wire [4-1:0] node26820;
	wire [4-1:0] node26823;
	wire [4-1:0] node26826;
	wire [4-1:0] node26827;
	wire [4-1:0] node26828;
	wire [4-1:0] node26831;
	wire [4-1:0] node26834;
	wire [4-1:0] node26835;
	wire [4-1:0] node26838;
	wire [4-1:0] node26841;
	wire [4-1:0] node26842;
	wire [4-1:0] node26843;
	wire [4-1:0] node26844;
	wire [4-1:0] node26845;
	wire [4-1:0] node26848;
	wire [4-1:0] node26851;
	wire [4-1:0] node26852;
	wire [4-1:0] node26855;
	wire [4-1:0] node26858;
	wire [4-1:0] node26859;
	wire [4-1:0] node26860;
	wire [4-1:0] node26863;
	wire [4-1:0] node26866;
	wire [4-1:0] node26867;
	wire [4-1:0] node26870;
	wire [4-1:0] node26873;
	wire [4-1:0] node26874;
	wire [4-1:0] node26875;
	wire [4-1:0] node26876;
	wire [4-1:0] node26879;
	wire [4-1:0] node26882;
	wire [4-1:0] node26883;
	wire [4-1:0] node26887;
	wire [4-1:0] node26888;
	wire [4-1:0] node26889;
	wire [4-1:0] node26892;
	wire [4-1:0] node26895;
	wire [4-1:0] node26896;
	wire [4-1:0] node26899;
	wire [4-1:0] node26902;
	wire [4-1:0] node26903;
	wire [4-1:0] node26904;
	wire [4-1:0] node26905;
	wire [4-1:0] node26906;
	wire [4-1:0] node26907;
	wire [4-1:0] node26910;
	wire [4-1:0] node26913;
	wire [4-1:0] node26914;
	wire [4-1:0] node26917;
	wire [4-1:0] node26920;
	wire [4-1:0] node26921;
	wire [4-1:0] node26922;
	wire [4-1:0] node26925;
	wire [4-1:0] node26928;
	wire [4-1:0] node26929;
	wire [4-1:0] node26932;
	wire [4-1:0] node26935;
	wire [4-1:0] node26936;
	wire [4-1:0] node26937;
	wire [4-1:0] node26938;
	wire [4-1:0] node26941;
	wire [4-1:0] node26944;
	wire [4-1:0] node26945;
	wire [4-1:0] node26948;
	wire [4-1:0] node26951;
	wire [4-1:0] node26952;
	wire [4-1:0] node26955;
	wire [4-1:0] node26958;
	wire [4-1:0] node26959;
	wire [4-1:0] node26960;
	wire [4-1:0] node26961;
	wire [4-1:0] node26963;
	wire [4-1:0] node26966;
	wire [4-1:0] node26967;
	wire [4-1:0] node26970;
	wire [4-1:0] node26973;
	wire [4-1:0] node26974;
	wire [4-1:0] node26977;
	wire [4-1:0] node26980;
	wire [4-1:0] node26981;
	wire [4-1:0] node26982;
	wire [4-1:0] node26983;
	wire [4-1:0] node26986;
	wire [4-1:0] node26989;
	wire [4-1:0] node26990;
	wire [4-1:0] node26994;
	wire [4-1:0] node26995;
	wire [4-1:0] node26996;
	wire [4-1:0] node26999;
	wire [4-1:0] node27002;
	wire [4-1:0] node27003;
	wire [4-1:0] node27006;
	wire [4-1:0] node27009;
	wire [4-1:0] node27010;
	wire [4-1:0] node27011;
	wire [4-1:0] node27012;
	wire [4-1:0] node27013;
	wire [4-1:0] node27014;
	wire [4-1:0] node27015;
	wire [4-1:0] node27018;
	wire [4-1:0] node27021;
	wire [4-1:0] node27022;
	wire [4-1:0] node27026;
	wire [4-1:0] node27027;
	wire [4-1:0] node27028;
	wire [4-1:0] node27031;
	wire [4-1:0] node27034;
	wire [4-1:0] node27035;
	wire [4-1:0] node27038;
	wire [4-1:0] node27041;
	wire [4-1:0] node27042;
	wire [4-1:0] node27043;
	wire [4-1:0] node27044;
	wire [4-1:0] node27047;
	wire [4-1:0] node27050;
	wire [4-1:0] node27051;
	wire [4-1:0] node27054;
	wire [4-1:0] node27057;
	wire [4-1:0] node27058;
	wire [4-1:0] node27060;
	wire [4-1:0] node27063;
	wire [4-1:0] node27064;
	wire [4-1:0] node27067;
	wire [4-1:0] node27070;
	wire [4-1:0] node27071;
	wire [4-1:0] node27072;
	wire [4-1:0] node27073;
	wire [4-1:0] node27074;
	wire [4-1:0] node27077;
	wire [4-1:0] node27080;
	wire [4-1:0] node27081;
	wire [4-1:0] node27085;
	wire [4-1:0] node27086;
	wire [4-1:0] node27087;
	wire [4-1:0] node27090;
	wire [4-1:0] node27093;
	wire [4-1:0] node27094;
	wire [4-1:0] node27098;
	wire [4-1:0] node27099;
	wire [4-1:0] node27100;
	wire [4-1:0] node27101;
	wire [4-1:0] node27104;
	wire [4-1:0] node27107;
	wire [4-1:0] node27108;
	wire [4-1:0] node27111;
	wire [4-1:0] node27114;
	wire [4-1:0] node27115;
	wire [4-1:0] node27116;
	wire [4-1:0] node27119;
	wire [4-1:0] node27122;
	wire [4-1:0] node27123;
	wire [4-1:0] node27126;
	wire [4-1:0] node27129;
	wire [4-1:0] node27130;
	wire [4-1:0] node27131;
	wire [4-1:0] node27132;
	wire [4-1:0] node27133;
	wire [4-1:0] node27134;
	wire [4-1:0] node27137;
	wire [4-1:0] node27140;
	wire [4-1:0] node27141;
	wire [4-1:0] node27144;
	wire [4-1:0] node27147;
	wire [4-1:0] node27148;
	wire [4-1:0] node27149;
	wire [4-1:0] node27152;
	wire [4-1:0] node27155;
	wire [4-1:0] node27156;
	wire [4-1:0] node27159;
	wire [4-1:0] node27162;
	wire [4-1:0] node27163;
	wire [4-1:0] node27164;
	wire [4-1:0] node27165;
	wire [4-1:0] node27168;
	wire [4-1:0] node27171;
	wire [4-1:0] node27173;
	wire [4-1:0] node27176;
	wire [4-1:0] node27177;
	wire [4-1:0] node27180;
	wire [4-1:0] node27183;
	wire [4-1:0] node27184;
	wire [4-1:0] node27185;
	wire [4-1:0] node27186;
	wire [4-1:0] node27187;
	wire [4-1:0] node27190;
	wire [4-1:0] node27193;
	wire [4-1:0] node27194;
	wire [4-1:0] node27197;
	wire [4-1:0] node27200;
	wire [4-1:0] node27201;
	wire [4-1:0] node27202;
	wire [4-1:0] node27205;
	wire [4-1:0] node27208;
	wire [4-1:0] node27209;
	wire [4-1:0] node27212;
	wire [4-1:0] node27215;
	wire [4-1:0] node27216;
	wire [4-1:0] node27217;
	wire [4-1:0] node27218;
	wire [4-1:0] node27221;
	wire [4-1:0] node27224;
	wire [4-1:0] node27225;
	wire [4-1:0] node27228;
	wire [4-1:0] node27231;
	wire [4-1:0] node27232;
	wire [4-1:0] node27233;
	wire [4-1:0] node27236;
	wire [4-1:0] node27239;
	wire [4-1:0] node27240;
	wire [4-1:0] node27244;
	wire [4-1:0] node27245;
	wire [4-1:0] node27246;
	wire [4-1:0] node27247;
	wire [4-1:0] node27248;
	wire [4-1:0] node27249;
	wire [4-1:0] node27250;
	wire [4-1:0] node27251;
	wire [4-1:0] node27254;
	wire [4-1:0] node27257;
	wire [4-1:0] node27258;
	wire [4-1:0] node27261;
	wire [4-1:0] node27264;
	wire [4-1:0] node27265;
	wire [4-1:0] node27266;
	wire [4-1:0] node27269;
	wire [4-1:0] node27272;
	wire [4-1:0] node27273;
	wire [4-1:0] node27277;
	wire [4-1:0] node27278;
	wire [4-1:0] node27279;
	wire [4-1:0] node27280;
	wire [4-1:0] node27284;
	wire [4-1:0] node27287;
	wire [4-1:0] node27288;
	wire [4-1:0] node27289;
	wire [4-1:0] node27293;
	wire [4-1:0] node27294;
	wire [4-1:0] node27298;
	wire [4-1:0] node27299;
	wire [4-1:0] node27300;
	wire [4-1:0] node27301;
	wire [4-1:0] node27302;
	wire [4-1:0] node27306;
	wire [4-1:0] node27307;
	wire [4-1:0] node27311;
	wire [4-1:0] node27312;
	wire [4-1:0] node27313;
	wire [4-1:0] node27317;
	wire [4-1:0] node27318;
	wire [4-1:0] node27322;
	wire [4-1:0] node27323;
	wire [4-1:0] node27324;
	wire [4-1:0] node27325;
	wire [4-1:0] node27329;
	wire [4-1:0] node27330;
	wire [4-1:0] node27334;
	wire [4-1:0] node27335;
	wire [4-1:0] node27336;
	wire [4-1:0] node27340;
	wire [4-1:0] node27341;
	wire [4-1:0] node27345;
	wire [4-1:0] node27346;
	wire [4-1:0] node27347;
	wire [4-1:0] node27348;
	wire [4-1:0] node27349;
	wire [4-1:0] node27350;
	wire [4-1:0] node27353;
	wire [4-1:0] node27356;
	wire [4-1:0] node27357;
	wire [4-1:0] node27360;
	wire [4-1:0] node27363;
	wire [4-1:0] node27364;
	wire [4-1:0] node27365;
	wire [4-1:0] node27368;
	wire [4-1:0] node27371;
	wire [4-1:0] node27372;
	wire [4-1:0] node27376;
	wire [4-1:0] node27377;
	wire [4-1:0] node27378;
	wire [4-1:0] node27379;
	wire [4-1:0] node27383;
	wire [4-1:0] node27384;
	wire [4-1:0] node27388;
	wire [4-1:0] node27389;
	wire [4-1:0] node27390;
	wire [4-1:0] node27394;
	wire [4-1:0] node27395;
	wire [4-1:0] node27399;
	wire [4-1:0] node27400;
	wire [4-1:0] node27401;
	wire [4-1:0] node27402;
	wire [4-1:0] node27403;
	wire [4-1:0] node27407;
	wire [4-1:0] node27408;
	wire [4-1:0] node27412;
	wire [4-1:0] node27414;
	wire [4-1:0] node27415;
	wire [4-1:0] node27419;
	wire [4-1:0] node27420;
	wire [4-1:0] node27421;
	wire [4-1:0] node27422;
	wire [4-1:0] node27426;
	wire [4-1:0] node27427;
	wire [4-1:0] node27431;
	wire [4-1:0] node27432;
	wire [4-1:0] node27433;
	wire [4-1:0] node27437;
	wire [4-1:0] node27438;
	wire [4-1:0] node27442;
	wire [4-1:0] node27443;
	wire [4-1:0] node27444;
	wire [4-1:0] node27445;
	wire [4-1:0] node27446;
	wire [4-1:0] node27447;
	wire [4-1:0] node27448;
	wire [4-1:0] node27451;
	wire [4-1:0] node27454;
	wire [4-1:0] node27455;
	wire [4-1:0] node27458;
	wire [4-1:0] node27461;
	wire [4-1:0] node27462;
	wire [4-1:0] node27463;
	wire [4-1:0] node27466;
	wire [4-1:0] node27469;
	wire [4-1:0] node27470;
	wire [4-1:0] node27473;
	wire [4-1:0] node27476;
	wire [4-1:0] node27477;
	wire [4-1:0] node27478;
	wire [4-1:0] node27479;
	wire [4-1:0] node27482;
	wire [4-1:0] node27485;
	wire [4-1:0] node27486;
	wire [4-1:0] node27489;
	wire [4-1:0] node27492;
	wire [4-1:0] node27493;
	wire [4-1:0] node27495;
	wire [4-1:0] node27498;
	wire [4-1:0] node27500;
	wire [4-1:0] node27503;
	wire [4-1:0] node27504;
	wire [4-1:0] node27505;
	wire [4-1:0] node27506;
	wire [4-1:0] node27507;
	wire [4-1:0] node27510;
	wire [4-1:0] node27513;
	wire [4-1:0] node27514;
	wire [4-1:0] node27517;
	wire [4-1:0] node27520;
	wire [4-1:0] node27521;
	wire [4-1:0] node27522;
	wire [4-1:0] node27525;
	wire [4-1:0] node27528;
	wire [4-1:0] node27529;
	wire [4-1:0] node27532;
	wire [4-1:0] node27535;
	wire [4-1:0] node27536;
	wire [4-1:0] node27537;
	wire [4-1:0] node27538;
	wire [4-1:0] node27541;
	wire [4-1:0] node27544;
	wire [4-1:0] node27545;
	wire [4-1:0] node27548;
	wire [4-1:0] node27551;
	wire [4-1:0] node27552;
	wire [4-1:0] node27553;
	wire [4-1:0] node27556;
	wire [4-1:0] node27559;
	wire [4-1:0] node27560;
	wire [4-1:0] node27563;
	wire [4-1:0] node27566;
	wire [4-1:0] node27567;
	wire [4-1:0] node27568;
	wire [4-1:0] node27569;
	wire [4-1:0] node27570;
	wire [4-1:0] node27571;
	wire [4-1:0] node27575;
	wire [4-1:0] node27576;
	wire [4-1:0] node27579;
	wire [4-1:0] node27582;
	wire [4-1:0] node27583;
	wire [4-1:0] node27584;
	wire [4-1:0] node27587;
	wire [4-1:0] node27590;
	wire [4-1:0] node27591;
	wire [4-1:0] node27595;
	wire [4-1:0] node27596;
	wire [4-1:0] node27597;
	wire [4-1:0] node27598;
	wire [4-1:0] node27602;
	wire [4-1:0] node27604;
	wire [4-1:0] node27607;
	wire [4-1:0] node27608;
	wire [4-1:0] node27609;
	wire [4-1:0] node27612;
	wire [4-1:0] node27615;
	wire [4-1:0] node27616;
	wire [4-1:0] node27619;
	wire [4-1:0] node27622;
	wire [4-1:0] node27623;
	wire [4-1:0] node27624;
	wire [4-1:0] node27625;
	wire [4-1:0] node27626;
	wire [4-1:0] node27630;
	wire [4-1:0] node27631;
	wire [4-1:0] node27635;
	wire [4-1:0] node27636;
	wire [4-1:0] node27637;
	wire [4-1:0] node27641;
	wire [4-1:0] node27642;
	wire [4-1:0] node27646;
	wire [4-1:0] node27647;
	wire [4-1:0] node27648;
	wire [4-1:0] node27649;
	wire [4-1:0] node27653;
	wire [4-1:0] node27654;
	wire [4-1:0] node27658;
	wire [4-1:0] node27659;
	wire [4-1:0] node27660;
	wire [4-1:0] node27664;
	wire [4-1:0] node27665;
	wire [4-1:0] node27669;
	wire [4-1:0] node27670;
	wire [4-1:0] node27671;
	wire [4-1:0] node27672;
	wire [4-1:0] node27673;
	wire [4-1:0] node27674;
	wire [4-1:0] node27675;
	wire [4-1:0] node27676;
	wire [4-1:0] node27677;
	wire [4-1:0] node27680;
	wire [4-1:0] node27683;
	wire [4-1:0] node27684;
	wire [4-1:0] node27687;
	wire [4-1:0] node27690;
	wire [4-1:0] node27691;
	wire [4-1:0] node27692;
	wire [4-1:0] node27695;
	wire [4-1:0] node27698;
	wire [4-1:0] node27700;
	wire [4-1:0] node27703;
	wire [4-1:0] node27704;
	wire [4-1:0] node27705;
	wire [4-1:0] node27706;
	wire [4-1:0] node27709;
	wire [4-1:0] node27712;
	wire [4-1:0] node27714;
	wire [4-1:0] node27717;
	wire [4-1:0] node27718;
	wire [4-1:0] node27719;
	wire [4-1:0] node27722;
	wire [4-1:0] node27725;
	wire [4-1:0] node27726;
	wire [4-1:0] node27729;
	wire [4-1:0] node27732;
	wire [4-1:0] node27733;
	wire [4-1:0] node27734;
	wire [4-1:0] node27735;
	wire [4-1:0] node27736;
	wire [4-1:0] node27739;
	wire [4-1:0] node27742;
	wire [4-1:0] node27743;
	wire [4-1:0] node27746;
	wire [4-1:0] node27749;
	wire [4-1:0] node27750;
	wire [4-1:0] node27751;
	wire [4-1:0] node27755;
	wire [4-1:0] node27756;
	wire [4-1:0] node27759;
	wire [4-1:0] node27762;
	wire [4-1:0] node27763;
	wire [4-1:0] node27764;
	wire [4-1:0] node27765;
	wire [4-1:0] node27768;
	wire [4-1:0] node27771;
	wire [4-1:0] node27772;
	wire [4-1:0] node27775;
	wire [4-1:0] node27778;
	wire [4-1:0] node27779;
	wire [4-1:0] node27780;
	wire [4-1:0] node27784;
	wire [4-1:0] node27785;
	wire [4-1:0] node27789;
	wire [4-1:0] node27790;
	wire [4-1:0] node27791;
	wire [4-1:0] node27792;
	wire [4-1:0] node27793;
	wire [4-1:0] node27794;
	wire [4-1:0] node27797;
	wire [4-1:0] node27800;
	wire [4-1:0] node27802;
	wire [4-1:0] node27805;
	wire [4-1:0] node27806;
	wire [4-1:0] node27807;
	wire [4-1:0] node27810;
	wire [4-1:0] node27813;
	wire [4-1:0] node27814;
	wire [4-1:0] node27817;
	wire [4-1:0] node27820;
	wire [4-1:0] node27821;
	wire [4-1:0] node27822;
	wire [4-1:0] node27824;
	wire [4-1:0] node27827;
	wire [4-1:0] node27829;
	wire [4-1:0] node27832;
	wire [4-1:0] node27833;
	wire [4-1:0] node27834;
	wire [4-1:0] node27837;
	wire [4-1:0] node27840;
	wire [4-1:0] node27841;
	wire [4-1:0] node27844;
	wire [4-1:0] node27847;
	wire [4-1:0] node27848;
	wire [4-1:0] node27849;
	wire [4-1:0] node27850;
	wire [4-1:0] node27851;
	wire [4-1:0] node27854;
	wire [4-1:0] node27857;
	wire [4-1:0] node27858;
	wire [4-1:0] node27861;
	wire [4-1:0] node27864;
	wire [4-1:0] node27865;
	wire [4-1:0] node27866;
	wire [4-1:0] node27869;
	wire [4-1:0] node27872;
	wire [4-1:0] node27873;
	wire [4-1:0] node27876;
	wire [4-1:0] node27879;
	wire [4-1:0] node27880;
	wire [4-1:0] node27881;
	wire [4-1:0] node27882;
	wire [4-1:0] node27885;
	wire [4-1:0] node27888;
	wire [4-1:0] node27889;
	wire [4-1:0] node27892;
	wire [4-1:0] node27895;
	wire [4-1:0] node27896;
	wire [4-1:0] node27897;
	wire [4-1:0] node27900;
	wire [4-1:0] node27903;
	wire [4-1:0] node27904;
	wire [4-1:0] node27908;
	wire [4-1:0] node27909;
	wire [4-1:0] node27910;
	wire [4-1:0] node27911;
	wire [4-1:0] node27912;
	wire [4-1:0] node27913;
	wire [4-1:0] node27914;
	wire [4-1:0] node27917;
	wire [4-1:0] node27920;
	wire [4-1:0] node27921;
	wire [4-1:0] node27924;
	wire [4-1:0] node27927;
	wire [4-1:0] node27928;
	wire [4-1:0] node27929;
	wire [4-1:0] node27932;
	wire [4-1:0] node27935;
	wire [4-1:0] node27936;
	wire [4-1:0] node27940;
	wire [4-1:0] node27941;
	wire [4-1:0] node27942;
	wire [4-1:0] node27943;
	wire [4-1:0] node27946;
	wire [4-1:0] node27949;
	wire [4-1:0] node27950;
	wire [4-1:0] node27953;
	wire [4-1:0] node27956;
	wire [4-1:0] node27957;
	wire [4-1:0] node27958;
	wire [4-1:0] node27961;
	wire [4-1:0] node27964;
	wire [4-1:0] node27965;
	wire [4-1:0] node27968;
	wire [4-1:0] node27971;
	wire [4-1:0] node27972;
	wire [4-1:0] node27973;
	wire [4-1:0] node27974;
	wire [4-1:0] node27977;
	wire [4-1:0] node27980;
	wire [4-1:0] node27981;
	wire [4-1:0] node27982;
	wire [4-1:0] node27985;
	wire [4-1:0] node27988;
	wire [4-1:0] node27989;
	wire [4-1:0] node27992;
	wire [4-1:0] node27995;
	wire [4-1:0] node27996;
	wire [4-1:0] node27997;
	wire [4-1:0] node27998;
	wire [4-1:0] node28001;
	wire [4-1:0] node28004;
	wire [4-1:0] node28005;
	wire [4-1:0] node28009;
	wire [4-1:0] node28010;
	wire [4-1:0] node28011;
	wire [4-1:0] node28014;
	wire [4-1:0] node28017;
	wire [4-1:0] node28018;
	wire [4-1:0] node28021;
	wire [4-1:0] node28024;
	wire [4-1:0] node28025;
	wire [4-1:0] node28026;
	wire [4-1:0] node28027;
	wire [4-1:0] node28028;
	wire [4-1:0] node28029;
	wire [4-1:0] node28032;
	wire [4-1:0] node28035;
	wire [4-1:0] node28037;
	wire [4-1:0] node28040;
	wire [4-1:0] node28041;
	wire [4-1:0] node28042;
	wire [4-1:0] node28045;
	wire [4-1:0] node28048;
	wire [4-1:0] node28049;
	wire [4-1:0] node28052;
	wire [4-1:0] node28055;
	wire [4-1:0] node28056;
	wire [4-1:0] node28057;
	wire [4-1:0] node28058;
	wire [4-1:0] node28061;
	wire [4-1:0] node28064;
	wire [4-1:0] node28065;
	wire [4-1:0] node28068;
	wire [4-1:0] node28071;
	wire [4-1:0] node28072;
	wire [4-1:0] node28073;
	wire [4-1:0] node28076;
	wire [4-1:0] node28079;
	wire [4-1:0] node28080;
	wire [4-1:0] node28083;
	wire [4-1:0] node28086;
	wire [4-1:0] node28087;
	wire [4-1:0] node28088;
	wire [4-1:0] node28089;
	wire [4-1:0] node28090;
	wire [4-1:0] node28093;
	wire [4-1:0] node28096;
	wire [4-1:0] node28097;
	wire [4-1:0] node28100;
	wire [4-1:0] node28103;
	wire [4-1:0] node28104;
	wire [4-1:0] node28105;
	wire [4-1:0] node28108;
	wire [4-1:0] node28111;
	wire [4-1:0] node28113;
	wire [4-1:0] node28116;
	wire [4-1:0] node28117;
	wire [4-1:0] node28118;
	wire [4-1:0] node28119;
	wire [4-1:0] node28122;
	wire [4-1:0] node28125;
	wire [4-1:0] node28126;
	wire [4-1:0] node28129;
	wire [4-1:0] node28132;
	wire [4-1:0] node28133;
	wire [4-1:0] node28134;
	wire [4-1:0] node28137;
	wire [4-1:0] node28140;
	wire [4-1:0] node28142;
	wire [4-1:0] node28145;
	wire [4-1:0] node28146;
	wire [4-1:0] node28147;
	wire [4-1:0] node28148;
	wire [4-1:0] node28149;
	wire [4-1:0] node28150;
	wire [4-1:0] node28151;
	wire [4-1:0] node28154;
	wire [4-1:0] node28157;
	wire [4-1:0] node28158;
	wire [4-1:0] node28159;
	wire [4-1:0] node28162;
	wire [4-1:0] node28165;
	wire [4-1:0] node28166;
	wire [4-1:0] node28169;
	wire [4-1:0] node28172;
	wire [4-1:0] node28173;
	wire [4-1:0] node28174;
	wire [4-1:0] node28176;
	wire [4-1:0] node28179;
	wire [4-1:0] node28180;
	wire [4-1:0] node28183;
	wire [4-1:0] node28186;
	wire [4-1:0] node28187;
	wire [4-1:0] node28188;
	wire [4-1:0] node28191;
	wire [4-1:0] node28194;
	wire [4-1:0] node28196;
	wire [4-1:0] node28199;
	wire [4-1:0] node28200;
	wire [4-1:0] node28201;
	wire [4-1:0] node28202;
	wire [4-1:0] node28203;
	wire [4-1:0] node28206;
	wire [4-1:0] node28209;
	wire [4-1:0] node28210;
	wire [4-1:0] node28214;
	wire [4-1:0] node28215;
	wire [4-1:0] node28216;
	wire [4-1:0] node28219;
	wire [4-1:0] node28222;
	wire [4-1:0] node28223;
	wire [4-1:0] node28226;
	wire [4-1:0] node28229;
	wire [4-1:0] node28230;
	wire [4-1:0] node28231;
	wire [4-1:0] node28233;
	wire [4-1:0] node28236;
	wire [4-1:0] node28238;
	wire [4-1:0] node28241;
	wire [4-1:0] node28242;
	wire [4-1:0] node28244;
	wire [4-1:0] node28247;
	wire [4-1:0] node28249;
	wire [4-1:0] node28252;
	wire [4-1:0] node28253;
	wire [4-1:0] node28254;
	wire [4-1:0] node28255;
	wire [4-1:0] node28256;
	wire [4-1:0] node28257;
	wire [4-1:0] node28260;
	wire [4-1:0] node28263;
	wire [4-1:0] node28264;
	wire [4-1:0] node28267;
	wire [4-1:0] node28270;
	wire [4-1:0] node28271;
	wire [4-1:0] node28272;
	wire [4-1:0] node28275;
	wire [4-1:0] node28278;
	wire [4-1:0] node28279;
	wire [4-1:0] node28282;
	wire [4-1:0] node28285;
	wire [4-1:0] node28286;
	wire [4-1:0] node28288;
	wire [4-1:0] node28289;
	wire [4-1:0] node28293;
	wire [4-1:0] node28294;
	wire [4-1:0] node28295;
	wire [4-1:0] node28299;
	wire [4-1:0] node28300;
	wire [4-1:0] node28304;
	wire [4-1:0] node28305;
	wire [4-1:0] node28306;
	wire [4-1:0] node28307;
	wire [4-1:0] node28311;
	wire [4-1:0] node28312;
	wire [4-1:0] node28316;
	wire [4-1:0] node28317;
	wire [4-1:0] node28318;
	wire [4-1:0] node28322;
	wire [4-1:0] node28323;
	wire [4-1:0] node28327;
	wire [4-1:0] node28328;
	wire [4-1:0] node28329;
	wire [4-1:0] node28330;
	wire [4-1:0] node28331;
	wire [4-1:0] node28332;
	wire [4-1:0] node28333;
	wire [4-1:0] node28336;
	wire [4-1:0] node28339;
	wire [4-1:0] node28340;
	wire [4-1:0] node28343;
	wire [4-1:0] node28346;
	wire [4-1:0] node28347;
	wire [4-1:0] node28348;
	wire [4-1:0] node28351;
	wire [4-1:0] node28354;
	wire [4-1:0] node28355;
	wire [4-1:0] node28358;
	wire [4-1:0] node28361;
	wire [4-1:0] node28362;
	wire [4-1:0] node28363;
	wire [4-1:0] node28365;
	wire [4-1:0] node28368;
	wire [4-1:0] node28369;
	wire [4-1:0] node28372;
	wire [4-1:0] node28375;
	wire [4-1:0] node28376;
	wire [4-1:0] node28377;
	wire [4-1:0] node28380;
	wire [4-1:0] node28383;
	wire [4-1:0] node28384;
	wire [4-1:0] node28388;
	wire [4-1:0] node28389;
	wire [4-1:0] node28390;
	wire [4-1:0] node28391;
	wire [4-1:0] node28392;
	wire [4-1:0] node28396;
	wire [4-1:0] node28397;
	wire [4-1:0] node28401;
	wire [4-1:0] node28402;
	wire [4-1:0] node28403;
	wire [4-1:0] node28407;
	wire [4-1:0] node28408;
	wire [4-1:0] node28412;
	wire [4-1:0] node28413;
	wire [4-1:0] node28414;
	wire [4-1:0] node28415;
	wire [4-1:0] node28418;
	wire [4-1:0] node28421;
	wire [4-1:0] node28422;
	wire [4-1:0] node28425;
	wire [4-1:0] node28428;
	wire [4-1:0] node28429;
	wire [4-1:0] node28432;
	wire [4-1:0] node28435;
	wire [4-1:0] node28436;
	wire [4-1:0] node28437;
	wire [4-1:0] node28438;
	wire [4-1:0] node28439;
	wire [4-1:0] node28440;
	wire [4-1:0] node28443;
	wire [4-1:0] node28446;
	wire [4-1:0] node28447;
	wire [4-1:0] node28450;
	wire [4-1:0] node28453;
	wire [4-1:0] node28454;
	wire [4-1:0] node28455;
	wire [4-1:0] node28459;
	wire [4-1:0] node28460;
	wire [4-1:0] node28463;
	wire [4-1:0] node28466;
	wire [4-1:0] node28467;
	wire [4-1:0] node28468;
	wire [4-1:0] node28469;
	wire [4-1:0] node28473;
	wire [4-1:0] node28474;
	wire [4-1:0] node28478;
	wire [4-1:0] node28479;
	wire [4-1:0] node28480;
	wire [4-1:0] node28484;
	wire [4-1:0] node28485;
	wire [4-1:0] node28489;
	wire [4-1:0] node28490;
	wire [4-1:0] node28491;
	wire [4-1:0] node28492;
	wire [4-1:0] node28493;
	wire [4-1:0] node28496;
	wire [4-1:0] node28499;
	wire [4-1:0] node28500;
	wire [4-1:0] node28503;
	wire [4-1:0] node28506;
	wire [4-1:0] node28507;
	wire [4-1:0] node28508;
	wire [4-1:0] node28511;
	wire [4-1:0] node28514;
	wire [4-1:0] node28515;
	wire [4-1:0] node28518;
	wire [4-1:0] node28521;
	wire [4-1:0] node28522;
	wire [4-1:0] node28523;
	wire [4-1:0] node28526;
	wire [4-1:0] node28529;
	wire [4-1:0] node28530;
	wire [4-1:0] node28533;
	wire [4-1:0] node28536;
	wire [4-1:0] node28537;
	wire [4-1:0] node28538;
	wire [4-1:0] node28539;
	wire [4-1:0] node28540;
	wire [4-1:0] node28541;
	wire [4-1:0] node28542;
	wire [4-1:0] node28543;
	wire [4-1:0] node28544;
	wire [4-1:0] node28545;
	wire [4-1:0] node28546;
	wire [4-1:0] node28547;
	wire [4-1:0] node28548;
	wire [4-1:0] node28549;
	wire [4-1:0] node28552;
	wire [4-1:0] node28555;
	wire [4-1:0] node28556;
	wire [4-1:0] node28559;
	wire [4-1:0] node28562;
	wire [4-1:0] node28563;
	wire [4-1:0] node28564;
	wire [4-1:0] node28567;
	wire [4-1:0] node28570;
	wire [4-1:0] node28571;
	wire [4-1:0] node28574;
	wire [4-1:0] node28577;
	wire [4-1:0] node28578;
	wire [4-1:0] node28579;
	wire [4-1:0] node28581;
	wire [4-1:0] node28584;
	wire [4-1:0] node28586;
	wire [4-1:0] node28589;
	wire [4-1:0] node28590;
	wire [4-1:0] node28592;
	wire [4-1:0] node28595;
	wire [4-1:0] node28597;
	wire [4-1:0] node28600;
	wire [4-1:0] node28601;
	wire [4-1:0] node28602;
	wire [4-1:0] node28603;
	wire [4-1:0] node28604;
	wire [4-1:0] node28607;
	wire [4-1:0] node28610;
	wire [4-1:0] node28612;
	wire [4-1:0] node28615;
	wire [4-1:0] node28616;
	wire [4-1:0] node28617;
	wire [4-1:0] node28620;
	wire [4-1:0] node28623;
	wire [4-1:0] node28624;
	wire [4-1:0] node28627;
	wire [4-1:0] node28630;
	wire [4-1:0] node28631;
	wire [4-1:0] node28632;
	wire [4-1:0] node28634;
	wire [4-1:0] node28637;
	wire [4-1:0] node28639;
	wire [4-1:0] node28642;
	wire [4-1:0] node28643;
	wire [4-1:0] node28645;
	wire [4-1:0] node28648;
	wire [4-1:0] node28650;
	wire [4-1:0] node28653;
	wire [4-1:0] node28654;
	wire [4-1:0] node28655;
	wire [4-1:0] node28656;
	wire [4-1:0] node28657;
	wire [4-1:0] node28658;
	wire [4-1:0] node28661;
	wire [4-1:0] node28664;
	wire [4-1:0] node28665;
	wire [4-1:0] node28668;
	wire [4-1:0] node28671;
	wire [4-1:0] node28672;
	wire [4-1:0] node28673;
	wire [4-1:0] node28676;
	wire [4-1:0] node28679;
	wire [4-1:0] node28680;
	wire [4-1:0] node28683;
	wire [4-1:0] node28686;
	wire [4-1:0] node28687;
	wire [4-1:0] node28688;
	wire [4-1:0] node28690;
	wire [4-1:0] node28693;
	wire [4-1:0] node28694;
	wire [4-1:0] node28697;
	wire [4-1:0] node28700;
	wire [4-1:0] node28701;
	wire [4-1:0] node28702;
	wire [4-1:0] node28705;
	wire [4-1:0] node28708;
	wire [4-1:0] node28709;
	wire [4-1:0] node28712;
	wire [4-1:0] node28715;
	wire [4-1:0] node28716;
	wire [4-1:0] node28717;
	wire [4-1:0] node28718;
	wire [4-1:0] node28719;
	wire [4-1:0] node28722;
	wire [4-1:0] node28725;
	wire [4-1:0] node28726;
	wire [4-1:0] node28729;
	wire [4-1:0] node28732;
	wire [4-1:0] node28733;
	wire [4-1:0] node28734;
	wire [4-1:0] node28737;
	wire [4-1:0] node28740;
	wire [4-1:0] node28741;
	wire [4-1:0] node28744;
	wire [4-1:0] node28747;
	wire [4-1:0] node28748;
	wire [4-1:0] node28749;
	wire [4-1:0] node28750;
	wire [4-1:0] node28753;
	wire [4-1:0] node28756;
	wire [4-1:0] node28757;
	wire [4-1:0] node28760;
	wire [4-1:0] node28763;
	wire [4-1:0] node28764;
	wire [4-1:0] node28765;
	wire [4-1:0] node28768;
	wire [4-1:0] node28771;
	wire [4-1:0] node28772;
	wire [4-1:0] node28775;
	wire [4-1:0] node28778;
	wire [4-1:0] node28779;
	wire [4-1:0] node28780;
	wire [4-1:0] node28781;
	wire [4-1:0] node28782;
	wire [4-1:0] node28783;
	wire [4-1:0] node28784;
	wire [4-1:0] node28787;
	wire [4-1:0] node28790;
	wire [4-1:0] node28792;
	wire [4-1:0] node28795;
	wire [4-1:0] node28796;
	wire [4-1:0] node28797;
	wire [4-1:0] node28800;
	wire [4-1:0] node28803;
	wire [4-1:0] node28804;
	wire [4-1:0] node28807;
	wire [4-1:0] node28810;
	wire [4-1:0] node28811;
	wire [4-1:0] node28812;
	wire [4-1:0] node28813;
	wire [4-1:0] node28816;
	wire [4-1:0] node28819;
	wire [4-1:0] node28820;
	wire [4-1:0] node28823;
	wire [4-1:0] node28826;
	wire [4-1:0] node28827;
	wire [4-1:0] node28828;
	wire [4-1:0] node28831;
	wire [4-1:0] node28834;
	wire [4-1:0] node28835;
	wire [4-1:0] node28839;
	wire [4-1:0] node28840;
	wire [4-1:0] node28841;
	wire [4-1:0] node28842;
	wire [4-1:0] node28844;
	wire [4-1:0] node28847;
	wire [4-1:0] node28849;
	wire [4-1:0] node28852;
	wire [4-1:0] node28853;
	wire [4-1:0] node28855;
	wire [4-1:0] node28858;
	wire [4-1:0] node28861;
	wire [4-1:0] node28862;
	wire [4-1:0] node28863;
	wire [4-1:0] node28864;
	wire [4-1:0] node28867;
	wire [4-1:0] node28870;
	wire [4-1:0] node28871;
	wire [4-1:0] node28874;
	wire [4-1:0] node28877;
	wire [4-1:0] node28878;
	wire [4-1:0] node28879;
	wire [4-1:0] node28882;
	wire [4-1:0] node28885;
	wire [4-1:0] node28886;
	wire [4-1:0] node28889;
	wire [4-1:0] node28892;
	wire [4-1:0] node28893;
	wire [4-1:0] node28894;
	wire [4-1:0] node28895;
	wire [4-1:0] node28896;
	wire [4-1:0] node28897;
	wire [4-1:0] node28900;
	wire [4-1:0] node28903;
	wire [4-1:0] node28904;
	wire [4-1:0] node28907;
	wire [4-1:0] node28910;
	wire [4-1:0] node28911;
	wire [4-1:0] node28912;
	wire [4-1:0] node28915;
	wire [4-1:0] node28918;
	wire [4-1:0] node28919;
	wire [4-1:0] node28922;
	wire [4-1:0] node28925;
	wire [4-1:0] node28926;
	wire [4-1:0] node28927;
	wire [4-1:0] node28928;
	wire [4-1:0] node28931;
	wire [4-1:0] node28934;
	wire [4-1:0] node28935;
	wire [4-1:0] node28939;
	wire [4-1:0] node28940;
	wire [4-1:0] node28941;
	wire [4-1:0] node28945;
	wire [4-1:0] node28946;
	wire [4-1:0] node28950;
	wire [4-1:0] node28951;
	wire [4-1:0] node28952;
	wire [4-1:0] node28953;
	wire [4-1:0] node28954;
	wire [4-1:0] node28957;
	wire [4-1:0] node28960;
	wire [4-1:0] node28961;
	wire [4-1:0] node28964;
	wire [4-1:0] node28967;
	wire [4-1:0] node28968;
	wire [4-1:0] node28969;
	wire [4-1:0] node28972;
	wire [4-1:0] node28975;
	wire [4-1:0] node28976;
	wire [4-1:0] node28979;
	wire [4-1:0] node28982;
	wire [4-1:0] node28983;
	wire [4-1:0] node28984;
	wire [4-1:0] node28985;
	wire [4-1:0] node28988;
	wire [4-1:0] node28991;
	wire [4-1:0] node28992;
	wire [4-1:0] node28996;
	wire [4-1:0] node28997;
	wire [4-1:0] node28998;
	wire [4-1:0] node29001;
	wire [4-1:0] node29004;
	wire [4-1:0] node29005;
	wire [4-1:0] node29009;
	wire [4-1:0] node29010;
	wire [4-1:0] node29011;
	wire [4-1:0] node29012;
	wire [4-1:0] node29013;
	wire [4-1:0] node29014;
	wire [4-1:0] node29016;
	wire [4-1:0] node29019;
	wire [4-1:0] node29021;
	wire [4-1:0] node29024;
	wire [4-1:0] node29025;
	wire [4-1:0] node29027;
	wire [4-1:0] node29030;
	wire [4-1:0] node29032;
	wire [4-1:0] node29035;
	wire [4-1:0] node29036;
	wire [4-1:0] node29037;
	wire [4-1:0] node29038;
	wire [4-1:0] node29039;
	wire [4-1:0] node29042;
	wire [4-1:0] node29045;
	wire [4-1:0] node29046;
	wire [4-1:0] node29050;
	wire [4-1:0] node29051;
	wire [4-1:0] node29052;
	wire [4-1:0] node29055;
	wire [4-1:0] node29058;
	wire [4-1:0] node29060;
	wire [4-1:0] node29063;
	wire [4-1:0] node29064;
	wire [4-1:0] node29065;
	wire [4-1:0] node29067;
	wire [4-1:0] node29070;
	wire [4-1:0] node29072;
	wire [4-1:0] node29075;
	wire [4-1:0] node29076;
	wire [4-1:0] node29078;
	wire [4-1:0] node29081;
	wire [4-1:0] node29083;
	wire [4-1:0] node29086;
	wire [4-1:0] node29087;
	wire [4-1:0] node29088;
	wire [4-1:0] node29089;
	wire [4-1:0] node29091;
	wire [4-1:0] node29094;
	wire [4-1:0] node29096;
	wire [4-1:0] node29099;
	wire [4-1:0] node29100;
	wire [4-1:0] node29102;
	wire [4-1:0] node29105;
	wire [4-1:0] node29107;
	wire [4-1:0] node29110;
	wire [4-1:0] node29111;
	wire [4-1:0] node29112;
	wire [4-1:0] node29113;
	wire [4-1:0] node29115;
	wire [4-1:0] node29118;
	wire [4-1:0] node29120;
	wire [4-1:0] node29123;
	wire [4-1:0] node29124;
	wire [4-1:0] node29126;
	wire [4-1:0] node29129;
	wire [4-1:0] node29131;
	wire [4-1:0] node29134;
	wire [4-1:0] node29135;
	wire [4-1:0] node29136;
	wire [4-1:0] node29137;
	wire [4-1:0] node29140;
	wire [4-1:0] node29143;
	wire [4-1:0] node29144;
	wire [4-1:0] node29147;
	wire [4-1:0] node29150;
	wire [4-1:0] node29151;
	wire [4-1:0] node29152;
	wire [4-1:0] node29156;
	wire [4-1:0] node29157;
	wire [4-1:0] node29160;
	wire [4-1:0] node29163;
	wire [4-1:0] node29164;
	wire [4-1:0] node29165;
	wire [4-1:0] node29166;
	wire [4-1:0] node29167;
	wire [4-1:0] node29169;
	wire [4-1:0] node29172;
	wire [4-1:0] node29174;
	wire [4-1:0] node29177;
	wire [4-1:0] node29178;
	wire [4-1:0] node29180;
	wire [4-1:0] node29183;
	wire [4-1:0] node29185;
	wire [4-1:0] node29188;
	wire [4-1:0] node29189;
	wire [4-1:0] node29190;
	wire [4-1:0] node29191;
	wire [4-1:0] node29192;
	wire [4-1:0] node29195;
	wire [4-1:0] node29198;
	wire [4-1:0] node29200;
	wire [4-1:0] node29203;
	wire [4-1:0] node29204;
	wire [4-1:0] node29205;
	wire [4-1:0] node29208;
	wire [4-1:0] node29211;
	wire [4-1:0] node29213;
	wire [4-1:0] node29216;
	wire [4-1:0] node29217;
	wire [4-1:0] node29218;
	wire [4-1:0] node29220;
	wire [4-1:0] node29223;
	wire [4-1:0] node29225;
	wire [4-1:0] node29228;
	wire [4-1:0] node29229;
	wire [4-1:0] node29231;
	wire [4-1:0] node29234;
	wire [4-1:0] node29236;
	wire [4-1:0] node29239;
	wire [4-1:0] node29240;
	wire [4-1:0] node29241;
	wire [4-1:0] node29242;
	wire [4-1:0] node29244;
	wire [4-1:0] node29247;
	wire [4-1:0] node29249;
	wire [4-1:0] node29252;
	wire [4-1:0] node29253;
	wire [4-1:0] node29255;
	wire [4-1:0] node29258;
	wire [4-1:0] node29260;
	wire [4-1:0] node29263;
	wire [4-1:0] node29264;
	wire [4-1:0] node29265;
	wire [4-1:0] node29266;
	wire [4-1:0] node29269;
	wire [4-1:0] node29272;
	wire [4-1:0] node29273;
	wire [4-1:0] node29274;
	wire [4-1:0] node29278;
	wire [4-1:0] node29279;
	wire [4-1:0] node29282;
	wire [4-1:0] node29285;
	wire [4-1:0] node29286;
	wire [4-1:0] node29287;
	wire [4-1:0] node29289;
	wire [4-1:0] node29292;
	wire [4-1:0] node29294;
	wire [4-1:0] node29297;
	wire [4-1:0] node29298;
	wire [4-1:0] node29300;
	wire [4-1:0] node29303;
	wire [4-1:0] node29305;
	wire [4-1:0] node29308;
	wire [4-1:0] node29309;
	wire [4-1:0] node29310;
	wire [4-1:0] node29311;
	wire [4-1:0] node29312;
	wire [4-1:0] node29313;
	wire [4-1:0] node29314;
	wire [4-1:0] node29315;
	wire [4-1:0] node29317;
	wire [4-1:0] node29320;
	wire [4-1:0] node29321;
	wire [4-1:0] node29324;
	wire [4-1:0] node29327;
	wire [4-1:0] node29328;
	wire [4-1:0] node29329;
	wire [4-1:0] node29332;
	wire [4-1:0] node29335;
	wire [4-1:0] node29336;
	wire [4-1:0] node29339;
	wire [4-1:0] node29342;
	wire [4-1:0] node29343;
	wire [4-1:0] node29344;
	wire [4-1:0] node29347;
	wire [4-1:0] node29350;
	wire [4-1:0] node29351;
	wire [4-1:0] node29352;
	wire [4-1:0] node29355;
	wire [4-1:0] node29358;
	wire [4-1:0] node29359;
	wire [4-1:0] node29362;
	wire [4-1:0] node29365;
	wire [4-1:0] node29366;
	wire [4-1:0] node29367;
	wire [4-1:0] node29368;
	wire [4-1:0] node29369;
	wire [4-1:0] node29372;
	wire [4-1:0] node29375;
	wire [4-1:0] node29376;
	wire [4-1:0] node29379;
	wire [4-1:0] node29382;
	wire [4-1:0] node29383;
	wire [4-1:0] node29384;
	wire [4-1:0] node29387;
	wire [4-1:0] node29390;
	wire [4-1:0] node29391;
	wire [4-1:0] node29394;
	wire [4-1:0] node29397;
	wire [4-1:0] node29398;
	wire [4-1:0] node29399;
	wire [4-1:0] node29400;
	wire [4-1:0] node29403;
	wire [4-1:0] node29406;
	wire [4-1:0] node29407;
	wire [4-1:0] node29410;
	wire [4-1:0] node29413;
	wire [4-1:0] node29414;
	wire [4-1:0] node29415;
	wire [4-1:0] node29418;
	wire [4-1:0] node29421;
	wire [4-1:0] node29422;
	wire [4-1:0] node29425;
	wire [4-1:0] node29428;
	wire [4-1:0] node29429;
	wire [4-1:0] node29430;
	wire [4-1:0] node29431;
	wire [4-1:0] node29432;
	wire [4-1:0] node29433;
	wire [4-1:0] node29436;
	wire [4-1:0] node29439;
	wire [4-1:0] node29440;
	wire [4-1:0] node29443;
	wire [4-1:0] node29446;
	wire [4-1:0] node29447;
	wire [4-1:0] node29448;
	wire [4-1:0] node29451;
	wire [4-1:0] node29454;
	wire [4-1:0] node29455;
	wire [4-1:0] node29458;
	wire [4-1:0] node29461;
	wire [4-1:0] node29462;
	wire [4-1:0] node29463;
	wire [4-1:0] node29464;
	wire [4-1:0] node29467;
	wire [4-1:0] node29470;
	wire [4-1:0] node29471;
	wire [4-1:0] node29474;
	wire [4-1:0] node29477;
	wire [4-1:0] node29478;
	wire [4-1:0] node29479;
	wire [4-1:0] node29482;
	wire [4-1:0] node29485;
	wire [4-1:0] node29486;
	wire [4-1:0] node29489;
	wire [4-1:0] node29492;
	wire [4-1:0] node29493;
	wire [4-1:0] node29494;
	wire [4-1:0] node29495;
	wire [4-1:0] node29496;
	wire [4-1:0] node29499;
	wire [4-1:0] node29502;
	wire [4-1:0] node29504;
	wire [4-1:0] node29507;
	wire [4-1:0] node29508;
	wire [4-1:0] node29510;
	wire [4-1:0] node29513;
	wire [4-1:0] node29514;
	wire [4-1:0] node29517;
	wire [4-1:0] node29520;
	wire [4-1:0] node29521;
	wire [4-1:0] node29522;
	wire [4-1:0] node29523;
	wire [4-1:0] node29526;
	wire [4-1:0] node29529;
	wire [4-1:0] node29530;
	wire [4-1:0] node29533;
	wire [4-1:0] node29536;
	wire [4-1:0] node29537;
	wire [4-1:0] node29538;
	wire [4-1:0] node29541;
	wire [4-1:0] node29544;
	wire [4-1:0] node29546;
	wire [4-1:0] node29549;
	wire [4-1:0] node29550;
	wire [4-1:0] node29551;
	wire [4-1:0] node29552;
	wire [4-1:0] node29553;
	wire [4-1:0] node29554;
	wire [4-1:0] node29555;
	wire [4-1:0] node29558;
	wire [4-1:0] node29561;
	wire [4-1:0] node29562;
	wire [4-1:0] node29565;
	wire [4-1:0] node29568;
	wire [4-1:0] node29569;
	wire [4-1:0] node29571;
	wire [4-1:0] node29574;
	wire [4-1:0] node29576;
	wire [4-1:0] node29579;
	wire [4-1:0] node29580;
	wire [4-1:0] node29582;
	wire [4-1:0] node29583;
	wire [4-1:0] node29586;
	wire [4-1:0] node29589;
	wire [4-1:0] node29590;
	wire [4-1:0] node29591;
	wire [4-1:0] node29595;
	wire [4-1:0] node29596;
	wire [4-1:0] node29599;
	wire [4-1:0] node29602;
	wire [4-1:0] node29603;
	wire [4-1:0] node29604;
	wire [4-1:0] node29605;
	wire [4-1:0] node29606;
	wire [4-1:0] node29610;
	wire [4-1:0] node29611;
	wire [4-1:0] node29614;
	wire [4-1:0] node29617;
	wire [4-1:0] node29618;
	wire [4-1:0] node29619;
	wire [4-1:0] node29622;
	wire [4-1:0] node29625;
	wire [4-1:0] node29626;
	wire [4-1:0] node29629;
	wire [4-1:0] node29632;
	wire [4-1:0] node29633;
	wire [4-1:0] node29634;
	wire [4-1:0] node29636;
	wire [4-1:0] node29639;
	wire [4-1:0] node29640;
	wire [4-1:0] node29643;
	wire [4-1:0] node29646;
	wire [4-1:0] node29647;
	wire [4-1:0] node29648;
	wire [4-1:0] node29651;
	wire [4-1:0] node29654;
	wire [4-1:0] node29656;
	wire [4-1:0] node29659;
	wire [4-1:0] node29660;
	wire [4-1:0] node29661;
	wire [4-1:0] node29662;
	wire [4-1:0] node29663;
	wire [4-1:0] node29665;
	wire [4-1:0] node29668;
	wire [4-1:0] node29670;
	wire [4-1:0] node29673;
	wire [4-1:0] node29674;
	wire [4-1:0] node29676;
	wire [4-1:0] node29679;
	wire [4-1:0] node29681;
	wire [4-1:0] node29684;
	wire [4-1:0] node29685;
	wire [4-1:0] node29686;
	wire [4-1:0] node29688;
	wire [4-1:0] node29691;
	wire [4-1:0] node29693;
	wire [4-1:0] node29696;
	wire [4-1:0] node29697;
	wire [4-1:0] node29699;
	wire [4-1:0] node29702;
	wire [4-1:0] node29704;
	wire [4-1:0] node29707;
	wire [4-1:0] node29708;
	wire [4-1:0] node29709;
	wire [4-1:0] node29710;
	wire [4-1:0] node29711;
	wire [4-1:0] node29714;
	wire [4-1:0] node29717;
	wire [4-1:0] node29719;
	wire [4-1:0] node29722;
	wire [4-1:0] node29724;
	wire [4-1:0] node29725;
	wire [4-1:0] node29728;
	wire [4-1:0] node29731;
	wire [4-1:0] node29732;
	wire [4-1:0] node29733;
	wire [4-1:0] node29734;
	wire [4-1:0] node29737;
	wire [4-1:0] node29740;
	wire [4-1:0] node29742;
	wire [4-1:0] node29745;
	wire [4-1:0] node29746;
	wire [4-1:0] node29747;
	wire [4-1:0] node29750;
	wire [4-1:0] node29753;
	wire [4-1:0] node29754;
	wire [4-1:0] node29757;
	wire [4-1:0] node29760;
	wire [4-1:0] node29761;
	wire [4-1:0] node29762;
	wire [4-1:0] node29763;
	wire [4-1:0] node29764;
	wire [4-1:0] node29765;
	wire [4-1:0] node29766;
	wire [4-1:0] node29767;
	wire [4-1:0] node29771;
	wire [4-1:0] node29772;
	wire [4-1:0] node29775;
	wire [4-1:0] node29778;
	wire [4-1:0] node29779;
	wire [4-1:0] node29782;
	wire [4-1:0] node29785;
	wire [4-1:0] node29786;
	wire [4-1:0] node29787;
	wire [4-1:0] node29788;
	wire [4-1:0] node29791;
	wire [4-1:0] node29794;
	wire [4-1:0] node29795;
	wire [4-1:0] node29798;
	wire [4-1:0] node29801;
	wire [4-1:0] node29802;
	wire [4-1:0] node29803;
	wire [4-1:0] node29806;
	wire [4-1:0] node29809;
	wire [4-1:0] node29811;
	wire [4-1:0] node29814;
	wire [4-1:0] node29815;
	wire [4-1:0] node29816;
	wire [4-1:0] node29817;
	wire [4-1:0] node29818;
	wire [4-1:0] node29821;
	wire [4-1:0] node29824;
	wire [4-1:0] node29825;
	wire [4-1:0] node29828;
	wire [4-1:0] node29831;
	wire [4-1:0] node29832;
	wire [4-1:0] node29833;
	wire [4-1:0] node29836;
	wire [4-1:0] node29839;
	wire [4-1:0] node29840;
	wire [4-1:0] node29843;
	wire [4-1:0] node29846;
	wire [4-1:0] node29847;
	wire [4-1:0] node29848;
	wire [4-1:0] node29849;
	wire [4-1:0] node29853;
	wire [4-1:0] node29854;
	wire [4-1:0] node29858;
	wire [4-1:0] node29859;
	wire [4-1:0] node29860;
	wire [4-1:0] node29863;
	wire [4-1:0] node29866;
	wire [4-1:0] node29867;
	wire [4-1:0] node29870;
	wire [4-1:0] node29873;
	wire [4-1:0] node29874;
	wire [4-1:0] node29875;
	wire [4-1:0] node29876;
	wire [4-1:0] node29877;
	wire [4-1:0] node29878;
	wire [4-1:0] node29881;
	wire [4-1:0] node29884;
	wire [4-1:0] node29885;
	wire [4-1:0] node29888;
	wire [4-1:0] node29891;
	wire [4-1:0] node29892;
	wire [4-1:0] node29893;
	wire [4-1:0] node29896;
	wire [4-1:0] node29899;
	wire [4-1:0] node29900;
	wire [4-1:0] node29903;
	wire [4-1:0] node29906;
	wire [4-1:0] node29907;
	wire [4-1:0] node29908;
	wire [4-1:0] node29909;
	wire [4-1:0] node29912;
	wire [4-1:0] node29915;
	wire [4-1:0] node29916;
	wire [4-1:0] node29919;
	wire [4-1:0] node29922;
	wire [4-1:0] node29923;
	wire [4-1:0] node29924;
	wire [4-1:0] node29927;
	wire [4-1:0] node29930;
	wire [4-1:0] node29931;
	wire [4-1:0] node29934;
	wire [4-1:0] node29937;
	wire [4-1:0] node29938;
	wire [4-1:0] node29939;
	wire [4-1:0] node29940;
	wire [4-1:0] node29942;
	wire [4-1:0] node29945;
	wire [4-1:0] node29946;
	wire [4-1:0] node29949;
	wire [4-1:0] node29952;
	wire [4-1:0] node29953;
	wire [4-1:0] node29954;
	wire [4-1:0] node29957;
	wire [4-1:0] node29960;
	wire [4-1:0] node29961;
	wire [4-1:0] node29964;
	wire [4-1:0] node29967;
	wire [4-1:0] node29968;
	wire [4-1:0] node29969;
	wire [4-1:0] node29970;
	wire [4-1:0] node29973;
	wire [4-1:0] node29976;
	wire [4-1:0] node29977;
	wire [4-1:0] node29980;
	wire [4-1:0] node29983;
	wire [4-1:0] node29984;
	wire [4-1:0] node29986;
	wire [4-1:0] node29989;
	wire [4-1:0] node29990;
	wire [4-1:0] node29993;
	wire [4-1:0] node29996;
	wire [4-1:0] node29997;
	wire [4-1:0] node29998;
	wire [4-1:0] node29999;
	wire [4-1:0] node30000;
	wire [4-1:0] node30001;
	wire [4-1:0] node30002;
	wire [4-1:0] node30005;
	wire [4-1:0] node30008;
	wire [4-1:0] node30009;
	wire [4-1:0] node30013;
	wire [4-1:0] node30014;
	wire [4-1:0] node30015;
	wire [4-1:0] node30018;
	wire [4-1:0] node30021;
	wire [4-1:0] node30022;
	wire [4-1:0] node30025;
	wire [4-1:0] node30028;
	wire [4-1:0] node30029;
	wire [4-1:0] node30030;
	wire [4-1:0] node30031;
	wire [4-1:0] node30034;
	wire [4-1:0] node30037;
	wire [4-1:0] node30038;
	wire [4-1:0] node30041;
	wire [4-1:0] node30044;
	wire [4-1:0] node30045;
	wire [4-1:0] node30046;
	wire [4-1:0] node30049;
	wire [4-1:0] node30052;
	wire [4-1:0] node30053;
	wire [4-1:0] node30056;
	wire [4-1:0] node30059;
	wire [4-1:0] node30060;
	wire [4-1:0] node30061;
	wire [4-1:0] node30062;
	wire [4-1:0] node30063;
	wire [4-1:0] node30066;
	wire [4-1:0] node30069;
	wire [4-1:0] node30070;
	wire [4-1:0] node30073;
	wire [4-1:0] node30076;
	wire [4-1:0] node30077;
	wire [4-1:0] node30078;
	wire [4-1:0] node30081;
	wire [4-1:0] node30084;
	wire [4-1:0] node30085;
	wire [4-1:0] node30088;
	wire [4-1:0] node30091;
	wire [4-1:0] node30092;
	wire [4-1:0] node30093;
	wire [4-1:0] node30094;
	wire [4-1:0] node30097;
	wire [4-1:0] node30100;
	wire [4-1:0] node30101;
	wire [4-1:0] node30105;
	wire [4-1:0] node30106;
	wire [4-1:0] node30107;
	wire [4-1:0] node30110;
	wire [4-1:0] node30113;
	wire [4-1:0] node30114;
	wire [4-1:0] node30117;
	wire [4-1:0] node30120;
	wire [4-1:0] node30121;
	wire [4-1:0] node30122;
	wire [4-1:0] node30123;
	wire [4-1:0] node30124;
	wire [4-1:0] node30125;
	wire [4-1:0] node30128;
	wire [4-1:0] node30131;
	wire [4-1:0] node30132;
	wire [4-1:0] node30135;
	wire [4-1:0] node30138;
	wire [4-1:0] node30139;
	wire [4-1:0] node30140;
	wire [4-1:0] node30143;
	wire [4-1:0] node30146;
	wire [4-1:0] node30148;
	wire [4-1:0] node30151;
	wire [4-1:0] node30152;
	wire [4-1:0] node30153;
	wire [4-1:0] node30154;
	wire [4-1:0] node30157;
	wire [4-1:0] node30161;
	wire [4-1:0] node30162;
	wire [4-1:0] node30164;
	wire [4-1:0] node30167;
	wire [4-1:0] node30168;
	wire [4-1:0] node30171;
	wire [4-1:0] node30174;
	wire [4-1:0] node30175;
	wire [4-1:0] node30176;
	wire [4-1:0] node30177;
	wire [4-1:0] node30178;
	wire [4-1:0] node30181;
	wire [4-1:0] node30184;
	wire [4-1:0] node30185;
	wire [4-1:0] node30188;
	wire [4-1:0] node30191;
	wire [4-1:0] node30192;
	wire [4-1:0] node30193;
	wire [4-1:0] node30197;
	wire [4-1:0] node30198;
	wire [4-1:0] node30201;
	wire [4-1:0] node30204;
	wire [4-1:0] node30205;
	wire [4-1:0] node30206;
	wire [4-1:0] node30209;
	wire [4-1:0] node30212;
	wire [4-1:0] node30213;
	wire [4-1:0] node30214;
	wire [4-1:0] node30217;
	wire [4-1:0] node30220;
	wire [4-1:0] node30221;
	wire [4-1:0] node30224;
	wire [4-1:0] node30227;
	wire [4-1:0] node30228;
	wire [4-1:0] node30229;
	wire [4-1:0] node30230;
	wire [4-1:0] node30231;
	wire [4-1:0] node30232;
	wire [4-1:0] node30233;
	wire [4-1:0] node30234;
	wire [4-1:0] node30235;
	wire [4-1:0] node30238;
	wire [4-1:0] node30241;
	wire [4-1:0] node30242;
	wire [4-1:0] node30243;
	wire [4-1:0] node30246;
	wire [4-1:0] node30249;
	wire [4-1:0] node30250;
	wire [4-1:0] node30253;
	wire [4-1:0] node30256;
	wire [4-1:0] node30257;
	wire [4-1:0] node30258;
	wire [4-1:0] node30261;
	wire [4-1:0] node30264;
	wire [4-1:0] node30265;
	wire [4-1:0] node30266;
	wire [4-1:0] node30269;
	wire [4-1:0] node30272;
	wire [4-1:0] node30273;
	wire [4-1:0] node30276;
	wire [4-1:0] node30279;
	wire [4-1:0] node30280;
	wire [4-1:0] node30281;
	wire [4-1:0] node30282;
	wire [4-1:0] node30285;
	wire [4-1:0] node30288;
	wire [4-1:0] node30289;
	wire [4-1:0] node30290;
	wire [4-1:0] node30293;
	wire [4-1:0] node30296;
	wire [4-1:0] node30299;
	wire [4-1:0] node30300;
	wire [4-1:0] node30301;
	wire [4-1:0] node30304;
	wire [4-1:0] node30307;
	wire [4-1:0] node30308;
	wire [4-1:0] node30309;
	wire [4-1:0] node30312;
	wire [4-1:0] node30315;
	wire [4-1:0] node30317;
	wire [4-1:0] node30320;
	wire [4-1:0] node30321;
	wire [4-1:0] node30322;
	wire [4-1:0] node30323;
	wire [4-1:0] node30324;
	wire [4-1:0] node30325;
	wire [4-1:0] node30328;
	wire [4-1:0] node30331;
	wire [4-1:0] node30332;
	wire [4-1:0] node30335;
	wire [4-1:0] node30338;
	wire [4-1:0] node30339;
	wire [4-1:0] node30340;
	wire [4-1:0] node30343;
	wire [4-1:0] node30346;
	wire [4-1:0] node30347;
	wire [4-1:0] node30350;
	wire [4-1:0] node30353;
	wire [4-1:0] node30354;
	wire [4-1:0] node30355;
	wire [4-1:0] node30357;
	wire [4-1:0] node30360;
	wire [4-1:0] node30361;
	wire [4-1:0] node30364;
	wire [4-1:0] node30367;
	wire [4-1:0] node30368;
	wire [4-1:0] node30369;
	wire [4-1:0] node30372;
	wire [4-1:0] node30375;
	wire [4-1:0] node30376;
	wire [4-1:0] node30379;
	wire [4-1:0] node30382;
	wire [4-1:0] node30383;
	wire [4-1:0] node30384;
	wire [4-1:0] node30385;
	wire [4-1:0] node30386;
	wire [4-1:0] node30389;
	wire [4-1:0] node30392;
	wire [4-1:0] node30394;
	wire [4-1:0] node30397;
	wire [4-1:0] node30398;
	wire [4-1:0] node30399;
	wire [4-1:0] node30402;
	wire [4-1:0] node30405;
	wire [4-1:0] node30406;
	wire [4-1:0] node30409;
	wire [4-1:0] node30412;
	wire [4-1:0] node30413;
	wire [4-1:0] node30414;
	wire [4-1:0] node30416;
	wire [4-1:0] node30419;
	wire [4-1:0] node30420;
	wire [4-1:0] node30424;
	wire [4-1:0] node30425;
	wire [4-1:0] node30426;
	wire [4-1:0] node30429;
	wire [4-1:0] node30432;
	wire [4-1:0] node30433;
	wire [4-1:0] node30436;
	wire [4-1:0] node30439;
	wire [4-1:0] node30440;
	wire [4-1:0] node30441;
	wire [4-1:0] node30442;
	wire [4-1:0] node30443;
	wire [4-1:0] node30444;
	wire [4-1:0] node30445;
	wire [4-1:0] node30448;
	wire [4-1:0] node30451;
	wire [4-1:0] node30452;
	wire [4-1:0] node30455;
	wire [4-1:0] node30458;
	wire [4-1:0] node30459;
	wire [4-1:0] node30462;
	wire [4-1:0] node30465;
	wire [4-1:0] node30466;
	wire [4-1:0] node30467;
	wire [4-1:0] node30468;
	wire [4-1:0] node30471;
	wire [4-1:0] node30474;
	wire [4-1:0] node30475;
	wire [4-1:0] node30478;
	wire [4-1:0] node30481;
	wire [4-1:0] node30482;
	wire [4-1:0] node30485;
	wire [4-1:0] node30488;
	wire [4-1:0] node30489;
	wire [4-1:0] node30490;
	wire [4-1:0] node30491;
	wire [4-1:0] node30492;
	wire [4-1:0] node30495;
	wire [4-1:0] node30498;
	wire [4-1:0] node30499;
	wire [4-1:0] node30502;
	wire [4-1:0] node30505;
	wire [4-1:0] node30506;
	wire [4-1:0] node30509;
	wire [4-1:0] node30512;
	wire [4-1:0] node30513;
	wire [4-1:0] node30514;
	wire [4-1:0] node30515;
	wire [4-1:0] node30518;
	wire [4-1:0] node30521;
	wire [4-1:0] node30523;
	wire [4-1:0] node30526;
	wire [4-1:0] node30527;
	wire [4-1:0] node30528;
	wire [4-1:0] node30532;
	wire [4-1:0] node30534;
	wire [4-1:0] node30537;
	wire [4-1:0] node30538;
	wire [4-1:0] node30539;
	wire [4-1:0] node30540;
	wire [4-1:0] node30541;
	wire [4-1:0] node30542;
	wire [4-1:0] node30545;
	wire [4-1:0] node30548;
	wire [4-1:0] node30549;
	wire [4-1:0] node30552;
	wire [4-1:0] node30555;
	wire [4-1:0] node30556;
	wire [4-1:0] node30557;
	wire [4-1:0] node30560;
	wire [4-1:0] node30563;
	wire [4-1:0] node30564;
	wire [4-1:0] node30567;
	wire [4-1:0] node30570;
	wire [4-1:0] node30571;
	wire [4-1:0] node30572;
	wire [4-1:0] node30573;
	wire [4-1:0] node30576;
	wire [4-1:0] node30579;
	wire [4-1:0] node30580;
	wire [4-1:0] node30583;
	wire [4-1:0] node30586;
	wire [4-1:0] node30587;
	wire [4-1:0] node30588;
	wire [4-1:0] node30591;
	wire [4-1:0] node30594;
	wire [4-1:0] node30595;
	wire [4-1:0] node30598;
	wire [4-1:0] node30601;
	wire [4-1:0] node30602;
	wire [4-1:0] node30603;
	wire [4-1:0] node30604;
	wire [4-1:0] node30605;
	wire [4-1:0] node30608;
	wire [4-1:0] node30611;
	wire [4-1:0] node30612;
	wire [4-1:0] node30615;
	wire [4-1:0] node30618;
	wire [4-1:0] node30619;
	wire [4-1:0] node30620;
	wire [4-1:0] node30623;
	wire [4-1:0] node30626;
	wire [4-1:0] node30627;
	wire [4-1:0] node30630;
	wire [4-1:0] node30633;
	wire [4-1:0] node30634;
	wire [4-1:0] node30635;
	wire [4-1:0] node30636;
	wire [4-1:0] node30639;
	wire [4-1:0] node30642;
	wire [4-1:0] node30643;
	wire [4-1:0] node30646;
	wire [4-1:0] node30649;
	wire [4-1:0] node30650;
	wire [4-1:0] node30651;
	wire [4-1:0] node30655;
	wire [4-1:0] node30656;
	wire [4-1:0] node30659;
	wire [4-1:0] node30662;
	wire [4-1:0] node30663;
	wire [4-1:0] node30664;
	wire [4-1:0] node30665;
	wire [4-1:0] node30666;
	wire [4-1:0] node30667;
	wire [4-1:0] node30668;
	wire [4-1:0] node30671;
	wire [4-1:0] node30674;
	wire [4-1:0] node30675;
	wire [4-1:0] node30676;
	wire [4-1:0] node30679;
	wire [4-1:0] node30682;
	wire [4-1:0] node30683;
	wire [4-1:0] node30686;
	wire [4-1:0] node30689;
	wire [4-1:0] node30690;
	wire [4-1:0] node30691;
	wire [4-1:0] node30692;
	wire [4-1:0] node30695;
	wire [4-1:0] node30698;
	wire [4-1:0] node30699;
	wire [4-1:0] node30702;
	wire [4-1:0] node30705;
	wire [4-1:0] node30706;
	wire [4-1:0] node30707;
	wire [4-1:0] node30711;
	wire [4-1:0] node30712;
	wire [4-1:0] node30715;
	wire [4-1:0] node30718;
	wire [4-1:0] node30719;
	wire [4-1:0] node30720;
	wire [4-1:0] node30721;
	wire [4-1:0] node30722;
	wire [4-1:0] node30725;
	wire [4-1:0] node30728;
	wire [4-1:0] node30729;
	wire [4-1:0] node30732;
	wire [4-1:0] node30735;
	wire [4-1:0] node30736;
	wire [4-1:0] node30737;
	wire [4-1:0] node30740;
	wire [4-1:0] node30743;
	wire [4-1:0] node30744;
	wire [4-1:0] node30747;
	wire [4-1:0] node30750;
	wire [4-1:0] node30751;
	wire [4-1:0] node30752;
	wire [4-1:0] node30753;
	wire [4-1:0] node30756;
	wire [4-1:0] node30759;
	wire [4-1:0] node30760;
	wire [4-1:0] node30763;
	wire [4-1:0] node30766;
	wire [4-1:0] node30767;
	wire [4-1:0] node30768;
	wire [4-1:0] node30771;
	wire [4-1:0] node30774;
	wire [4-1:0] node30775;
	wire [4-1:0] node30778;
	wire [4-1:0] node30781;
	wire [4-1:0] node30782;
	wire [4-1:0] node30783;
	wire [4-1:0] node30784;
	wire [4-1:0] node30785;
	wire [4-1:0] node30786;
	wire [4-1:0] node30789;
	wire [4-1:0] node30792;
	wire [4-1:0] node30793;
	wire [4-1:0] node30796;
	wire [4-1:0] node30799;
	wire [4-1:0] node30800;
	wire [4-1:0] node30802;
	wire [4-1:0] node30805;
	wire [4-1:0] node30806;
	wire [4-1:0] node30809;
	wire [4-1:0] node30812;
	wire [4-1:0] node30813;
	wire [4-1:0] node30814;
	wire [4-1:0] node30815;
	wire [4-1:0] node30818;
	wire [4-1:0] node30821;
	wire [4-1:0] node30822;
	wire [4-1:0] node30825;
	wire [4-1:0] node30828;
	wire [4-1:0] node30829;
	wire [4-1:0] node30830;
	wire [4-1:0] node30833;
	wire [4-1:0] node30836;
	wire [4-1:0] node30837;
	wire [4-1:0] node30840;
	wire [4-1:0] node30843;
	wire [4-1:0] node30844;
	wire [4-1:0] node30845;
	wire [4-1:0] node30846;
	wire [4-1:0] node30847;
	wire [4-1:0] node30850;
	wire [4-1:0] node30853;
	wire [4-1:0] node30854;
	wire [4-1:0] node30857;
	wire [4-1:0] node30860;
	wire [4-1:0] node30861;
	wire [4-1:0] node30862;
	wire [4-1:0] node30865;
	wire [4-1:0] node30868;
	wire [4-1:0] node30869;
	wire [4-1:0] node30872;
	wire [4-1:0] node30875;
	wire [4-1:0] node30876;
	wire [4-1:0] node30877;
	wire [4-1:0] node30879;
	wire [4-1:0] node30882;
	wire [4-1:0] node30884;
	wire [4-1:0] node30887;
	wire [4-1:0] node30888;
	wire [4-1:0] node30890;
	wire [4-1:0] node30893;
	wire [4-1:0] node30895;
	wire [4-1:0] node30898;
	wire [4-1:0] node30899;
	wire [4-1:0] node30900;
	wire [4-1:0] node30901;
	wire [4-1:0] node30902;
	wire [4-1:0] node30903;
	wire [4-1:0] node30906;
	wire [4-1:0] node30909;
	wire [4-1:0] node30910;
	wire [4-1:0] node30913;
	wire [4-1:0] node30916;
	wire [4-1:0] node30917;
	wire [4-1:0] node30918;
	wire [4-1:0] node30921;
	wire [4-1:0] node30924;
	wire [4-1:0] node30925;
	wire [4-1:0] node30926;
	wire [4-1:0] node30929;
	wire [4-1:0] node30932;
	wire [4-1:0] node30933;
	wire [4-1:0] node30936;
	wire [4-1:0] node30939;
	wire [4-1:0] node30940;
	wire [4-1:0] node30941;
	wire [4-1:0] node30942;
	wire [4-1:0] node30943;
	wire [4-1:0] node30946;
	wire [4-1:0] node30949;
	wire [4-1:0] node30950;
	wire [4-1:0] node30954;
	wire [4-1:0] node30955;
	wire [4-1:0] node30956;
	wire [4-1:0] node30959;
	wire [4-1:0] node30962;
	wire [4-1:0] node30963;
	wire [4-1:0] node30966;
	wire [4-1:0] node30969;
	wire [4-1:0] node30970;
	wire [4-1:0] node30971;
	wire [4-1:0] node30974;
	wire [4-1:0] node30977;
	wire [4-1:0] node30978;
	wire [4-1:0] node30979;
	wire [4-1:0] node30982;
	wire [4-1:0] node30985;
	wire [4-1:0] node30986;
	wire [4-1:0] node30989;
	wire [4-1:0] node30992;
	wire [4-1:0] node30993;
	wire [4-1:0] node30994;
	wire [4-1:0] node30995;
	wire [4-1:0] node30996;
	wire [4-1:0] node30997;
	wire [4-1:0] node31000;
	wire [4-1:0] node31003;
	wire [4-1:0] node31004;
	wire [4-1:0] node31007;
	wire [4-1:0] node31010;
	wire [4-1:0] node31011;
	wire [4-1:0] node31014;
	wire [4-1:0] node31017;
	wire [4-1:0] node31018;
	wire [4-1:0] node31019;
	wire [4-1:0] node31020;
	wire [4-1:0] node31023;
	wire [4-1:0] node31026;
	wire [4-1:0] node31027;
	wire [4-1:0] node31030;
	wire [4-1:0] node31033;
	wire [4-1:0] node31034;
	wire [4-1:0] node31037;
	wire [4-1:0] node31040;
	wire [4-1:0] node31041;
	wire [4-1:0] node31042;
	wire [4-1:0] node31043;
	wire [4-1:0] node31046;
	wire [4-1:0] node31049;
	wire [4-1:0] node31050;
	wire [4-1:0] node31051;
	wire [4-1:0] node31054;
	wire [4-1:0] node31057;
	wire [4-1:0] node31058;
	wire [4-1:0] node31061;
	wire [4-1:0] node31064;
	wire [4-1:0] node31065;
	wire [4-1:0] node31066;
	wire [4-1:0] node31069;
	wire [4-1:0] node31072;
	wire [4-1:0] node31073;
	wire [4-1:0] node31076;
	wire [4-1:0] node31079;
	wire [4-1:0] node31080;
	wire [4-1:0] node31081;
	wire [4-1:0] node31082;
	wire [4-1:0] node31083;
	wire [4-1:0] node31084;
	wire [4-1:0] node31085;
	wire [4-1:0] node31086;
	wire [4-1:0] node31087;
	wire [4-1:0] node31091;
	wire [4-1:0] node31092;
	wire [4-1:0] node31096;
	wire [4-1:0] node31097;
	wire [4-1:0] node31098;
	wire [4-1:0] node31101;
	wire [4-1:0] node31104;
	wire [4-1:0] node31105;
	wire [4-1:0] node31108;
	wire [4-1:0] node31111;
	wire [4-1:0] node31112;
	wire [4-1:0] node31113;
	wire [4-1:0] node31114;
	wire [4-1:0] node31117;
	wire [4-1:0] node31120;
	wire [4-1:0] node31121;
	wire [4-1:0] node31124;
	wire [4-1:0] node31127;
	wire [4-1:0] node31128;
	wire [4-1:0] node31129;
	wire [4-1:0] node31132;
	wire [4-1:0] node31135;
	wire [4-1:0] node31136;
	wire [4-1:0] node31139;
	wire [4-1:0] node31142;
	wire [4-1:0] node31143;
	wire [4-1:0] node31144;
	wire [4-1:0] node31145;
	wire [4-1:0] node31146;
	wire [4-1:0] node31149;
	wire [4-1:0] node31152;
	wire [4-1:0] node31153;
	wire [4-1:0] node31157;
	wire [4-1:0] node31158;
	wire [4-1:0] node31159;
	wire [4-1:0] node31162;
	wire [4-1:0] node31165;
	wire [4-1:0] node31166;
	wire [4-1:0] node31169;
	wire [4-1:0] node31172;
	wire [4-1:0] node31173;
	wire [4-1:0] node31174;
	wire [4-1:0] node31175;
	wire [4-1:0] node31178;
	wire [4-1:0] node31181;
	wire [4-1:0] node31182;
	wire [4-1:0] node31185;
	wire [4-1:0] node31188;
	wire [4-1:0] node31189;
	wire [4-1:0] node31190;
	wire [4-1:0] node31193;
	wire [4-1:0] node31196;
	wire [4-1:0] node31197;
	wire [4-1:0] node31200;
	wire [4-1:0] node31203;
	wire [4-1:0] node31204;
	wire [4-1:0] node31205;
	wire [4-1:0] node31206;
	wire [4-1:0] node31207;
	wire [4-1:0] node31208;
	wire [4-1:0] node31211;
	wire [4-1:0] node31214;
	wire [4-1:0] node31215;
	wire [4-1:0] node31218;
	wire [4-1:0] node31221;
	wire [4-1:0] node31222;
	wire [4-1:0] node31223;
	wire [4-1:0] node31226;
	wire [4-1:0] node31229;
	wire [4-1:0] node31230;
	wire [4-1:0] node31233;
	wire [4-1:0] node31236;
	wire [4-1:0] node31237;
	wire [4-1:0] node31238;
	wire [4-1:0] node31241;
	wire [4-1:0] node31244;
	wire [4-1:0] node31245;
	wire [4-1:0] node31247;
	wire [4-1:0] node31250;
	wire [4-1:0] node31251;
	wire [4-1:0] node31254;
	wire [4-1:0] node31257;
	wire [4-1:0] node31258;
	wire [4-1:0] node31259;
	wire [4-1:0] node31260;
	wire [4-1:0] node31261;
	wire [4-1:0] node31264;
	wire [4-1:0] node31267;
	wire [4-1:0] node31268;
	wire [4-1:0] node31271;
	wire [4-1:0] node31274;
	wire [4-1:0] node31275;
	wire [4-1:0] node31276;
	wire [4-1:0] node31279;
	wire [4-1:0] node31282;
	wire [4-1:0] node31283;
	wire [4-1:0] node31286;
	wire [4-1:0] node31289;
	wire [4-1:0] node31290;
	wire [4-1:0] node31291;
	wire [4-1:0] node31294;
	wire [4-1:0] node31297;
	wire [4-1:0] node31298;
	wire [4-1:0] node31299;
	wire [4-1:0] node31302;
	wire [4-1:0] node31305;
	wire [4-1:0] node31306;
	wire [4-1:0] node31309;
	wire [4-1:0] node31312;
	wire [4-1:0] node31313;
	wire [4-1:0] node31314;
	wire [4-1:0] node31315;
	wire [4-1:0] node31316;
	wire [4-1:0] node31317;
	wire [4-1:0] node31318;
	wire [4-1:0] node31321;
	wire [4-1:0] node31324;
	wire [4-1:0] node31325;
	wire [4-1:0] node31328;
	wire [4-1:0] node31331;
	wire [4-1:0] node31332;
	wire [4-1:0] node31335;
	wire [4-1:0] node31338;
	wire [4-1:0] node31339;
	wire [4-1:0] node31340;
	wire [4-1:0] node31341;
	wire [4-1:0] node31345;
	wire [4-1:0] node31346;
	wire [4-1:0] node31349;
	wire [4-1:0] node31352;
	wire [4-1:0] node31353;
	wire [4-1:0] node31355;
	wire [4-1:0] node31358;
	wire [4-1:0] node31359;
	wire [4-1:0] node31362;
	wire [4-1:0] node31365;
	wire [4-1:0] node31366;
	wire [4-1:0] node31367;
	wire [4-1:0] node31368;
	wire [4-1:0] node31369;
	wire [4-1:0] node31373;
	wire [4-1:0] node31374;
	wire [4-1:0] node31378;
	wire [4-1:0] node31379;
	wire [4-1:0] node31380;
	wire [4-1:0] node31384;
	wire [4-1:0] node31385;
	wire [4-1:0] node31389;
	wire [4-1:0] node31390;
	wire [4-1:0] node31391;
	wire [4-1:0] node31392;
	wire [4-1:0] node31396;
	wire [4-1:0] node31398;
	wire [4-1:0] node31401;
	wire [4-1:0] node31402;
	wire [4-1:0] node31405;
	wire [4-1:0] node31407;
	wire [4-1:0] node31410;
	wire [4-1:0] node31411;
	wire [4-1:0] node31412;
	wire [4-1:0] node31413;
	wire [4-1:0] node31414;
	wire [4-1:0] node31415;
	wire [4-1:0] node31419;
	wire [4-1:0] node31420;
	wire [4-1:0] node31424;
	wire [4-1:0] node31425;
	wire [4-1:0] node31426;
	wire [4-1:0] node31430;
	wire [4-1:0] node31431;
	wire [4-1:0] node31435;
	wire [4-1:0] node31436;
	wire [4-1:0] node31437;
	wire [4-1:0] node31439;
	wire [4-1:0] node31442;
	wire [4-1:0] node31443;
	wire [4-1:0] node31446;
	wire [4-1:0] node31449;
	wire [4-1:0] node31450;
	wire [4-1:0] node31451;
	wire [4-1:0] node31454;
	wire [4-1:0] node31457;
	wire [4-1:0] node31458;
	wire [4-1:0] node31461;
	wire [4-1:0] node31464;
	wire [4-1:0] node31465;
	wire [4-1:0] node31466;
	wire [4-1:0] node31467;
	wire [4-1:0] node31468;
	wire [4-1:0] node31472;
	wire [4-1:0] node31473;
	wire [4-1:0] node31477;
	wire [4-1:0] node31478;
	wire [4-1:0] node31479;
	wire [4-1:0] node31483;
	wire [4-1:0] node31484;
	wire [4-1:0] node31488;
	wire [4-1:0] node31489;
	wire [4-1:0] node31490;
	wire [4-1:0] node31491;
	wire [4-1:0] node31494;
	wire [4-1:0] node31497;
	wire [4-1:0] node31499;
	wire [4-1:0] node31502;
	wire [4-1:0] node31503;
	wire [4-1:0] node31506;
	wire [4-1:0] node31507;
	wire [4-1:0] node31510;
	wire [4-1:0] node31513;
	wire [4-1:0] node31514;
	wire [4-1:0] node31515;
	wire [4-1:0] node31516;
	wire [4-1:0] node31517;
	wire [4-1:0] node31518;
	wire [4-1:0] node31519;
	wire [4-1:0] node31520;
	wire [4-1:0] node31523;
	wire [4-1:0] node31526;
	wire [4-1:0] node31527;
	wire [4-1:0] node31530;
	wire [4-1:0] node31533;
	wire [4-1:0] node31534;
	wire [4-1:0] node31535;
	wire [4-1:0] node31538;
	wire [4-1:0] node31541;
	wire [4-1:0] node31542;
	wire [4-1:0] node31545;
	wire [4-1:0] node31548;
	wire [4-1:0] node31549;
	wire [4-1:0] node31550;
	wire [4-1:0] node31551;
	wire [4-1:0] node31554;
	wire [4-1:0] node31557;
	wire [4-1:0] node31558;
	wire [4-1:0] node31561;
	wire [4-1:0] node31564;
	wire [4-1:0] node31565;
	wire [4-1:0] node31566;
	wire [4-1:0] node31569;
	wire [4-1:0] node31572;
	wire [4-1:0] node31573;
	wire [4-1:0] node31576;
	wire [4-1:0] node31579;
	wire [4-1:0] node31580;
	wire [4-1:0] node31581;
	wire [4-1:0] node31582;
	wire [4-1:0] node31583;
	wire [4-1:0] node31586;
	wire [4-1:0] node31589;
	wire [4-1:0] node31590;
	wire [4-1:0] node31593;
	wire [4-1:0] node31596;
	wire [4-1:0] node31597;
	wire [4-1:0] node31598;
	wire [4-1:0] node31601;
	wire [4-1:0] node31604;
	wire [4-1:0] node31605;
	wire [4-1:0] node31608;
	wire [4-1:0] node31611;
	wire [4-1:0] node31612;
	wire [4-1:0] node31613;
	wire [4-1:0] node31614;
	wire [4-1:0] node31617;
	wire [4-1:0] node31620;
	wire [4-1:0] node31621;
	wire [4-1:0] node31624;
	wire [4-1:0] node31627;
	wire [4-1:0] node31628;
	wire [4-1:0] node31631;
	wire [4-1:0] node31634;
	wire [4-1:0] node31635;
	wire [4-1:0] node31636;
	wire [4-1:0] node31637;
	wire [4-1:0] node31638;
	wire [4-1:0] node31639;
	wire [4-1:0] node31642;
	wire [4-1:0] node31645;
	wire [4-1:0] node31646;
	wire [4-1:0] node31649;
	wire [4-1:0] node31652;
	wire [4-1:0] node31653;
	wire [4-1:0] node31654;
	wire [4-1:0] node31657;
	wire [4-1:0] node31660;
	wire [4-1:0] node31661;
	wire [4-1:0] node31664;
	wire [4-1:0] node31667;
	wire [4-1:0] node31668;
	wire [4-1:0] node31669;
	wire [4-1:0] node31670;
	wire [4-1:0] node31674;
	wire [4-1:0] node31675;
	wire [4-1:0] node31678;
	wire [4-1:0] node31681;
	wire [4-1:0] node31682;
	wire [4-1:0] node31683;
	wire [4-1:0] node31686;
	wire [4-1:0] node31689;
	wire [4-1:0] node31690;
	wire [4-1:0] node31693;
	wire [4-1:0] node31696;
	wire [4-1:0] node31697;
	wire [4-1:0] node31698;
	wire [4-1:0] node31699;
	wire [4-1:0] node31700;
	wire [4-1:0] node31703;
	wire [4-1:0] node31706;
	wire [4-1:0] node31707;
	wire [4-1:0] node31710;
	wire [4-1:0] node31713;
	wire [4-1:0] node31714;
	wire [4-1:0] node31717;
	wire [4-1:0] node31720;
	wire [4-1:0] node31721;
	wire [4-1:0] node31722;
	wire [4-1:0] node31723;
	wire [4-1:0] node31726;
	wire [4-1:0] node31729;
	wire [4-1:0] node31730;
	wire [4-1:0] node31733;
	wire [4-1:0] node31736;
	wire [4-1:0] node31737;
	wire [4-1:0] node31738;
	wire [4-1:0] node31741;
	wire [4-1:0] node31744;
	wire [4-1:0] node31746;
	wire [4-1:0] node31749;
	wire [4-1:0] node31750;
	wire [4-1:0] node31751;
	wire [4-1:0] node31752;
	wire [4-1:0] node31753;
	wire [4-1:0] node31754;
	wire [4-1:0] node31755;
	wire [4-1:0] node31758;
	wire [4-1:0] node31761;
	wire [4-1:0] node31762;
	wire [4-1:0] node31765;
	wire [4-1:0] node31768;
	wire [4-1:0] node31769;
	wire [4-1:0] node31770;
	wire [4-1:0] node31773;
	wire [4-1:0] node31777;
	wire [4-1:0] node31778;
	wire [4-1:0] node31779;
	wire [4-1:0] node31780;
	wire [4-1:0] node31783;
	wire [4-1:0] node31786;
	wire [4-1:0] node31787;
	wire [4-1:0] node31790;
	wire [4-1:0] node31793;
	wire [4-1:0] node31794;
	wire [4-1:0] node31795;
	wire [4-1:0] node31798;
	wire [4-1:0] node31801;
	wire [4-1:0] node31802;
	wire [4-1:0] node31805;
	wire [4-1:0] node31808;
	wire [4-1:0] node31809;
	wire [4-1:0] node31810;
	wire [4-1:0] node31811;
	wire [4-1:0] node31812;
	wire [4-1:0] node31815;
	wire [4-1:0] node31818;
	wire [4-1:0] node31819;
	wire [4-1:0] node31822;
	wire [4-1:0] node31825;
	wire [4-1:0] node31826;
	wire [4-1:0] node31827;
	wire [4-1:0] node31830;
	wire [4-1:0] node31833;
	wire [4-1:0] node31834;
	wire [4-1:0] node31837;
	wire [4-1:0] node31840;
	wire [4-1:0] node31841;
	wire [4-1:0] node31842;
	wire [4-1:0] node31843;
	wire [4-1:0] node31846;
	wire [4-1:0] node31849;
	wire [4-1:0] node31850;
	wire [4-1:0] node31853;
	wire [4-1:0] node31856;
	wire [4-1:0] node31857;
	wire [4-1:0] node31858;
	wire [4-1:0] node31861;
	wire [4-1:0] node31864;
	wire [4-1:0] node31865;
	wire [4-1:0] node31868;
	wire [4-1:0] node31871;
	wire [4-1:0] node31872;
	wire [4-1:0] node31873;
	wire [4-1:0] node31874;
	wire [4-1:0] node31875;
	wire [4-1:0] node31876;
	wire [4-1:0] node31879;
	wire [4-1:0] node31882;
	wire [4-1:0] node31883;
	wire [4-1:0] node31886;
	wire [4-1:0] node31889;
	wire [4-1:0] node31890;
	wire [4-1:0] node31891;
	wire [4-1:0] node31894;
	wire [4-1:0] node31897;
	wire [4-1:0] node31898;
	wire [4-1:0] node31901;
	wire [4-1:0] node31904;
	wire [4-1:0] node31905;
	wire [4-1:0] node31906;
	wire [4-1:0] node31907;
	wire [4-1:0] node31910;
	wire [4-1:0] node31913;
	wire [4-1:0] node31914;
	wire [4-1:0] node31917;
	wire [4-1:0] node31920;
	wire [4-1:0] node31921;
	wire [4-1:0] node31922;
	wire [4-1:0] node31925;
	wire [4-1:0] node31928;
	wire [4-1:0] node31929;
	wire [4-1:0] node31932;
	wire [4-1:0] node31935;
	wire [4-1:0] node31936;
	wire [4-1:0] node31937;
	wire [4-1:0] node31938;
	wire [4-1:0] node31939;
	wire [4-1:0] node31942;
	wire [4-1:0] node31945;
	wire [4-1:0] node31946;
	wire [4-1:0] node31949;
	wire [4-1:0] node31952;
	wire [4-1:0] node31953;
	wire [4-1:0] node31954;
	wire [4-1:0] node31957;
	wire [4-1:0] node31960;
	wire [4-1:0] node31962;
	wire [4-1:0] node31965;
	wire [4-1:0] node31966;
	wire [4-1:0] node31967;
	wire [4-1:0] node31968;
	wire [4-1:0] node31971;
	wire [4-1:0] node31974;
	wire [4-1:0] node31975;
	wire [4-1:0] node31978;
	wire [4-1:0] node31981;
	wire [4-1:0] node31982;
	wire [4-1:0] node31983;
	wire [4-1:0] node31986;
	wire [4-1:0] node31989;
	wire [4-1:0] node31990;
	wire [4-1:0] node31993;
	wire [4-1:0] node31996;
	wire [4-1:0] node31997;
	wire [4-1:0] node31998;
	wire [4-1:0] node31999;
	wire [4-1:0] node32000;
	wire [4-1:0] node32001;
	wire [4-1:0] node32002;
	wire [4-1:0] node32003;
	wire [4-1:0] node32004;
	wire [4-1:0] node32005;
	wire [4-1:0] node32006;
	wire [4-1:0] node32009;
	wire [4-1:0] node32012;
	wire [4-1:0] node32014;
	wire [4-1:0] node32017;
	wire [4-1:0] node32018;
	wire [4-1:0] node32019;
	wire [4-1:0] node32023;
	wire [4-1:0] node32024;
	wire [4-1:0] node32028;
	wire [4-1:0] node32029;
	wire [4-1:0] node32030;
	wire [4-1:0] node32032;
	wire [4-1:0] node32035;
	wire [4-1:0] node32037;
	wire [4-1:0] node32040;
	wire [4-1:0] node32041;
	wire [4-1:0] node32043;
	wire [4-1:0] node32046;
	wire [4-1:0] node32048;
	wire [4-1:0] node32051;
	wire [4-1:0] node32052;
	wire [4-1:0] node32053;
	wire [4-1:0] node32054;
	wire [4-1:0] node32055;
	wire [4-1:0] node32058;
	wire [4-1:0] node32061;
	wire [4-1:0] node32062;
	wire [4-1:0] node32065;
	wire [4-1:0] node32068;
	wire [4-1:0] node32069;
	wire [4-1:0] node32070;
	wire [4-1:0] node32073;
	wire [4-1:0] node32076;
	wire [4-1:0] node32077;
	wire [4-1:0] node32081;
	wire [4-1:0] node32082;
	wire [4-1:0] node32083;
	wire [4-1:0] node32085;
	wire [4-1:0] node32088;
	wire [4-1:0] node32089;
	wire [4-1:0] node32092;
	wire [4-1:0] node32095;
	wire [4-1:0] node32096;
	wire [4-1:0] node32097;
	wire [4-1:0] node32100;
	wire [4-1:0] node32103;
	wire [4-1:0] node32104;
	wire [4-1:0] node32107;
	wire [4-1:0] node32110;
	wire [4-1:0] node32111;
	wire [4-1:0] node32112;
	wire [4-1:0] node32113;
	wire [4-1:0] node32114;
	wire [4-1:0] node32115;
	wire [4-1:0] node32118;
	wire [4-1:0] node32121;
	wire [4-1:0] node32122;
	wire [4-1:0] node32125;
	wire [4-1:0] node32128;
	wire [4-1:0] node32129;
	wire [4-1:0] node32130;
	wire [4-1:0] node32133;
	wire [4-1:0] node32136;
	wire [4-1:0] node32137;
	wire [4-1:0] node32140;
	wire [4-1:0] node32143;
	wire [4-1:0] node32144;
	wire [4-1:0] node32145;
	wire [4-1:0] node32147;
	wire [4-1:0] node32150;
	wire [4-1:0] node32152;
	wire [4-1:0] node32155;
	wire [4-1:0] node32156;
	wire [4-1:0] node32158;
	wire [4-1:0] node32161;
	wire [4-1:0] node32163;
	wire [4-1:0] node32166;
	wire [4-1:0] node32167;
	wire [4-1:0] node32168;
	wire [4-1:0] node32169;
	wire [4-1:0] node32170;
	wire [4-1:0] node32173;
	wire [4-1:0] node32176;
	wire [4-1:0] node32177;
	wire [4-1:0] node32180;
	wire [4-1:0] node32183;
	wire [4-1:0] node32184;
	wire [4-1:0] node32185;
	wire [4-1:0] node32188;
	wire [4-1:0] node32191;
	wire [4-1:0] node32192;
	wire [4-1:0] node32195;
	wire [4-1:0] node32198;
	wire [4-1:0] node32199;
	wire [4-1:0] node32200;
	wire [4-1:0] node32202;
	wire [4-1:0] node32205;
	wire [4-1:0] node32206;
	wire [4-1:0] node32209;
	wire [4-1:0] node32212;
	wire [4-1:0] node32213;
	wire [4-1:0] node32214;
	wire [4-1:0] node32217;
	wire [4-1:0] node32220;
	wire [4-1:0] node32221;
	wire [4-1:0] node32224;
	wire [4-1:0] node32227;
	wire [4-1:0] node32228;
	wire [4-1:0] node32229;
	wire [4-1:0] node32230;
	wire [4-1:0] node32231;
	wire [4-1:0] node32232;
	wire [4-1:0] node32233;
	wire [4-1:0] node32236;
	wire [4-1:0] node32239;
	wire [4-1:0] node32240;
	wire [4-1:0] node32243;
	wire [4-1:0] node32246;
	wire [4-1:0] node32247;
	wire [4-1:0] node32248;
	wire [4-1:0] node32251;
	wire [4-1:0] node32254;
	wire [4-1:0] node32255;
	wire [4-1:0] node32258;
	wire [4-1:0] node32261;
	wire [4-1:0] node32262;
	wire [4-1:0] node32263;
	wire [4-1:0] node32265;
	wire [4-1:0] node32268;
	wire [4-1:0] node32270;
	wire [4-1:0] node32273;
	wire [4-1:0] node32274;
	wire [4-1:0] node32276;
	wire [4-1:0] node32280;
	wire [4-1:0] node32281;
	wire [4-1:0] node32282;
	wire [4-1:0] node32283;
	wire [4-1:0] node32284;
	wire [4-1:0] node32287;
	wire [4-1:0] node32290;
	wire [4-1:0] node32291;
	wire [4-1:0] node32294;
	wire [4-1:0] node32297;
	wire [4-1:0] node32298;
	wire [4-1:0] node32300;
	wire [4-1:0] node32303;
	wire [4-1:0] node32304;
	wire [4-1:0] node32307;
	wire [4-1:0] node32310;
	wire [4-1:0] node32311;
	wire [4-1:0] node32312;
	wire [4-1:0] node32314;
	wire [4-1:0] node32317;
	wire [4-1:0] node32319;
	wire [4-1:0] node32322;
	wire [4-1:0] node32323;
	wire [4-1:0] node32325;
	wire [4-1:0] node32328;
	wire [4-1:0] node32330;
	wire [4-1:0] node32333;
	wire [4-1:0] node32334;
	wire [4-1:0] node32335;
	wire [4-1:0] node32336;
	wire [4-1:0] node32337;
	wire [4-1:0] node32338;
	wire [4-1:0] node32341;
	wire [4-1:0] node32344;
	wire [4-1:0] node32345;
	wire [4-1:0] node32348;
	wire [4-1:0] node32351;
	wire [4-1:0] node32352;
	wire [4-1:0] node32355;
	wire [4-1:0] node32356;
	wire [4-1:0] node32359;
	wire [4-1:0] node32362;
	wire [4-1:0] node32363;
	wire [4-1:0] node32364;
	wire [4-1:0] node32365;
	wire [4-1:0] node32369;
	wire [4-1:0] node32370;
	wire [4-1:0] node32373;
	wire [4-1:0] node32376;
	wire [4-1:0] node32377;
	wire [4-1:0] node32378;
	wire [4-1:0] node32381;
	wire [4-1:0] node32384;
	wire [4-1:0] node32385;
	wire [4-1:0] node32388;
	wire [4-1:0] node32391;
	wire [4-1:0] node32392;
	wire [4-1:0] node32393;
	wire [4-1:0] node32394;
	wire [4-1:0] node32395;
	wire [4-1:0] node32398;
	wire [4-1:0] node32401;
	wire [4-1:0] node32402;
	wire [4-1:0] node32405;
	wire [4-1:0] node32408;
	wire [4-1:0] node32409;
	wire [4-1:0] node32411;
	wire [4-1:0] node32414;
	wire [4-1:0] node32415;
	wire [4-1:0] node32418;
	wire [4-1:0] node32421;
	wire [4-1:0] node32422;
	wire [4-1:0] node32423;
	wire [4-1:0] node32424;
	wire [4-1:0] node32427;
	wire [4-1:0] node32430;
	wire [4-1:0] node32431;
	wire [4-1:0] node32435;
	wire [4-1:0] node32436;
	wire [4-1:0] node32437;
	wire [4-1:0] node32440;
	wire [4-1:0] node32443;
	wire [4-1:0] node32444;
	wire [4-1:0] node32447;
	wire [4-1:0] node32450;
	wire [4-1:0] node32451;
	wire [4-1:0] node32452;
	wire [4-1:0] node32453;
	wire [4-1:0] node32454;
	wire [4-1:0] node32455;
	wire [4-1:0] node32456;
	wire [4-1:0] node32457;
	wire [4-1:0] node32460;
	wire [4-1:0] node32463;
	wire [4-1:0] node32464;
	wire [4-1:0] node32467;
	wire [4-1:0] node32470;
	wire [4-1:0] node32471;
	wire [4-1:0] node32472;
	wire [4-1:0] node32475;
	wire [4-1:0] node32478;
	wire [4-1:0] node32479;
	wire [4-1:0] node32483;
	wire [4-1:0] node32484;
	wire [4-1:0] node32485;
	wire [4-1:0] node32487;
	wire [4-1:0] node32490;
	wire [4-1:0] node32492;
	wire [4-1:0] node32495;
	wire [4-1:0] node32496;
	wire [4-1:0] node32498;
	wire [4-1:0] node32501;
	wire [4-1:0] node32503;
	wire [4-1:0] node32506;
	wire [4-1:0] node32507;
	wire [4-1:0] node32508;
	wire [4-1:0] node32509;
	wire [4-1:0] node32510;
	wire [4-1:0] node32513;
	wire [4-1:0] node32516;
	wire [4-1:0] node32517;
	wire [4-1:0] node32520;
	wire [4-1:0] node32523;
	wire [4-1:0] node32524;
	wire [4-1:0] node32525;
	wire [4-1:0] node32528;
	wire [4-1:0] node32531;
	wire [4-1:0] node32532;
	wire [4-1:0] node32535;
	wire [4-1:0] node32538;
	wire [4-1:0] node32539;
	wire [4-1:0] node32540;
	wire [4-1:0] node32543;
	wire [4-1:0] node32546;
	wire [4-1:0] node32547;
	wire [4-1:0] node32549;
	wire [4-1:0] node32552;
	wire [4-1:0] node32553;
	wire [4-1:0] node32556;
	wire [4-1:0] node32559;
	wire [4-1:0] node32560;
	wire [4-1:0] node32561;
	wire [4-1:0] node32562;
	wire [4-1:0] node32563;
	wire [4-1:0] node32564;
	wire [4-1:0] node32567;
	wire [4-1:0] node32570;
	wire [4-1:0] node32571;
	wire [4-1:0] node32574;
	wire [4-1:0] node32577;
	wire [4-1:0] node32578;
	wire [4-1:0] node32579;
	wire [4-1:0] node32582;
	wire [4-1:0] node32585;
	wire [4-1:0] node32586;
	wire [4-1:0] node32590;
	wire [4-1:0] node32591;
	wire [4-1:0] node32592;
	wire [4-1:0] node32595;
	wire [4-1:0] node32598;
	wire [4-1:0] node32599;
	wire [4-1:0] node32600;
	wire [4-1:0] node32603;
	wire [4-1:0] node32606;
	wire [4-1:0] node32607;
	wire [4-1:0] node32610;
	wire [4-1:0] node32613;
	wire [4-1:0] node32614;
	wire [4-1:0] node32615;
	wire [4-1:0] node32616;
	wire [4-1:0] node32617;
	wire [4-1:0] node32620;
	wire [4-1:0] node32623;
	wire [4-1:0] node32624;
	wire [4-1:0] node32627;
	wire [4-1:0] node32630;
	wire [4-1:0] node32631;
	wire [4-1:0] node32633;
	wire [4-1:0] node32636;
	wire [4-1:0] node32637;
	wire [4-1:0] node32640;
	wire [4-1:0] node32643;
	wire [4-1:0] node32644;
	wire [4-1:0] node32645;
	wire [4-1:0] node32647;
	wire [4-1:0] node32650;
	wire [4-1:0] node32652;
	wire [4-1:0] node32655;
	wire [4-1:0] node32656;
	wire [4-1:0] node32658;
	wire [4-1:0] node32661;
	wire [4-1:0] node32663;
	wire [4-1:0] node32666;
	wire [4-1:0] node32667;
	wire [4-1:0] node32668;
	wire [4-1:0] node32669;
	wire [4-1:0] node32670;
	wire [4-1:0] node32671;
	wire [4-1:0] node32672;
	wire [4-1:0] node32675;
	wire [4-1:0] node32678;
	wire [4-1:0] node32679;
	wire [4-1:0] node32682;
	wire [4-1:0] node32685;
	wire [4-1:0] node32686;
	wire [4-1:0] node32687;
	wire [4-1:0] node32690;
	wire [4-1:0] node32693;
	wire [4-1:0] node32694;
	wire [4-1:0] node32697;
	wire [4-1:0] node32700;
	wire [4-1:0] node32701;
	wire [4-1:0] node32702;
	wire [4-1:0] node32704;
	wire [4-1:0] node32707;
	wire [4-1:0] node32709;
	wire [4-1:0] node32712;
	wire [4-1:0] node32713;
	wire [4-1:0] node32715;
	wire [4-1:0] node32718;
	wire [4-1:0] node32720;
	wire [4-1:0] node32723;
	wire [4-1:0] node32724;
	wire [4-1:0] node32725;
	wire [4-1:0] node32726;
	wire [4-1:0] node32727;
	wire [4-1:0] node32730;
	wire [4-1:0] node32733;
	wire [4-1:0] node32734;
	wire [4-1:0] node32737;
	wire [4-1:0] node32740;
	wire [4-1:0] node32741;
	wire [4-1:0] node32743;
	wire [4-1:0] node32746;
	wire [4-1:0] node32747;
	wire [4-1:0] node32750;
	wire [4-1:0] node32753;
	wire [4-1:0] node32754;
	wire [4-1:0] node32755;
	wire [4-1:0] node32758;
	wire [4-1:0] node32761;
	wire [4-1:0] node32762;
	wire [4-1:0] node32763;
	wire [4-1:0] node32766;
	wire [4-1:0] node32769;
	wire [4-1:0] node32770;
	wire [4-1:0] node32773;
	wire [4-1:0] node32776;
	wire [4-1:0] node32777;
	wire [4-1:0] node32778;
	wire [4-1:0] node32779;
	wire [4-1:0] node32780;
	wire [4-1:0] node32781;
	wire [4-1:0] node32784;
	wire [4-1:0] node32787;
	wire [4-1:0] node32789;
	wire [4-1:0] node32792;
	wire [4-1:0] node32793;
	wire [4-1:0] node32794;
	wire [4-1:0] node32797;
	wire [4-1:0] node32800;
	wire [4-1:0] node32801;
	wire [4-1:0] node32804;
	wire [4-1:0] node32807;
	wire [4-1:0] node32808;
	wire [4-1:0] node32809;
	wire [4-1:0] node32811;
	wire [4-1:0] node32814;
	wire [4-1:0] node32816;
	wire [4-1:0] node32819;
	wire [4-1:0] node32820;
	wire [4-1:0] node32822;
	wire [4-1:0] node32825;
	wire [4-1:0] node32827;
	wire [4-1:0] node32830;
	wire [4-1:0] node32831;
	wire [4-1:0] node32832;
	wire [4-1:0] node32833;
	wire [4-1:0] node32834;
	wire [4-1:0] node32838;
	wire [4-1:0] node32839;
	wire [4-1:0] node32842;
	wire [4-1:0] node32845;
	wire [4-1:0] node32846;
	wire [4-1:0] node32847;
	wire [4-1:0] node32851;
	wire [4-1:0] node32852;
	wire [4-1:0] node32856;
	wire [4-1:0] node32857;
	wire [4-1:0] node32858;
	wire [4-1:0] node32860;
	wire [4-1:0] node32863;
	wire [4-1:0] node32865;
	wire [4-1:0] node32868;
	wire [4-1:0] node32869;
	wire [4-1:0] node32871;
	wire [4-1:0] node32874;
	wire [4-1:0] node32876;
	wire [4-1:0] node32879;
	wire [4-1:0] node32880;
	wire [4-1:0] node32881;
	wire [4-1:0] node32882;
	wire [4-1:0] node32883;
	wire [4-1:0] node32884;
	wire [4-1:0] node32885;
	wire [4-1:0] node32886;
	wire [4-1:0] node32887;
	wire [4-1:0] node32890;
	wire [4-1:0] node32893;
	wire [4-1:0] node32894;
	wire [4-1:0] node32897;
	wire [4-1:0] node32900;
	wire [4-1:0] node32901;
	wire [4-1:0] node32902;
	wire [4-1:0] node32905;
	wire [4-1:0] node32908;
	wire [4-1:0] node32909;
	wire [4-1:0] node32912;
	wire [4-1:0] node32915;
	wire [4-1:0] node32916;
	wire [4-1:0] node32917;
	wire [4-1:0] node32918;
	wire [4-1:0] node32921;
	wire [4-1:0] node32924;
	wire [4-1:0] node32925;
	wire [4-1:0] node32928;
	wire [4-1:0] node32931;
	wire [4-1:0] node32932;
	wire [4-1:0] node32933;
	wire [4-1:0] node32936;
	wire [4-1:0] node32939;
	wire [4-1:0] node32940;
	wire [4-1:0] node32943;
	wire [4-1:0] node32946;
	wire [4-1:0] node32947;
	wire [4-1:0] node32948;
	wire [4-1:0] node32949;
	wire [4-1:0] node32950;
	wire [4-1:0] node32953;
	wire [4-1:0] node32956;
	wire [4-1:0] node32957;
	wire [4-1:0] node32961;
	wire [4-1:0] node32962;
	wire [4-1:0] node32963;
	wire [4-1:0] node32966;
	wire [4-1:0] node32969;
	wire [4-1:0] node32970;
	wire [4-1:0] node32973;
	wire [4-1:0] node32976;
	wire [4-1:0] node32977;
	wire [4-1:0] node32978;
	wire [4-1:0] node32979;
	wire [4-1:0] node32982;
	wire [4-1:0] node32985;
	wire [4-1:0] node32986;
	wire [4-1:0] node32989;
	wire [4-1:0] node32992;
	wire [4-1:0] node32993;
	wire [4-1:0] node32996;
	wire [4-1:0] node32999;
	wire [4-1:0] node33000;
	wire [4-1:0] node33001;
	wire [4-1:0] node33002;
	wire [4-1:0] node33003;
	wire [4-1:0] node33004;
	wire [4-1:0] node33007;
	wire [4-1:0] node33010;
	wire [4-1:0] node33011;
	wire [4-1:0] node33014;
	wire [4-1:0] node33017;
	wire [4-1:0] node33018;
	wire [4-1:0] node33019;
	wire [4-1:0] node33022;
	wire [4-1:0] node33025;
	wire [4-1:0] node33026;
	wire [4-1:0] node33029;
	wire [4-1:0] node33032;
	wire [4-1:0] node33033;
	wire [4-1:0] node33034;
	wire [4-1:0] node33035;
	wire [4-1:0] node33038;
	wire [4-1:0] node33041;
	wire [4-1:0] node33042;
	wire [4-1:0] node33045;
	wire [4-1:0] node33048;
	wire [4-1:0] node33049;
	wire [4-1:0] node33050;
	wire [4-1:0] node33053;
	wire [4-1:0] node33056;
	wire [4-1:0] node33057;
	wire [4-1:0] node33060;
	wire [4-1:0] node33063;
	wire [4-1:0] node33064;
	wire [4-1:0] node33065;
	wire [4-1:0] node33066;
	wire [4-1:0] node33067;
	wire [4-1:0] node33070;
	wire [4-1:0] node33073;
	wire [4-1:0] node33074;
	wire [4-1:0] node33077;
	wire [4-1:0] node33080;
	wire [4-1:0] node33081;
	wire [4-1:0] node33082;
	wire [4-1:0] node33085;
	wire [4-1:0] node33088;
	wire [4-1:0] node33089;
	wire [4-1:0] node33092;
	wire [4-1:0] node33095;
	wire [4-1:0] node33096;
	wire [4-1:0] node33097;
	wire [4-1:0] node33099;
	wire [4-1:0] node33102;
	wire [4-1:0] node33103;
	wire [4-1:0] node33106;
	wire [4-1:0] node33109;
	wire [4-1:0] node33110;
	wire [4-1:0] node33111;
	wire [4-1:0] node33114;
	wire [4-1:0] node33117;
	wire [4-1:0] node33119;
	wire [4-1:0] node33122;
	wire [4-1:0] node33123;
	wire [4-1:0] node33124;
	wire [4-1:0] node33125;
	wire [4-1:0] node33126;
	wire [4-1:0] node33127;
	wire [4-1:0] node33128;
	wire [4-1:0] node33131;
	wire [4-1:0] node33134;
	wire [4-1:0] node33136;
	wire [4-1:0] node33139;
	wire [4-1:0] node33140;
	wire [4-1:0] node33141;
	wire [4-1:0] node33144;
	wire [4-1:0] node33147;
	wire [4-1:0] node33148;
	wire [4-1:0] node33151;
	wire [4-1:0] node33154;
	wire [4-1:0] node33155;
	wire [4-1:0] node33156;
	wire [4-1:0] node33157;
	wire [4-1:0] node33160;
	wire [4-1:0] node33163;
	wire [4-1:0] node33164;
	wire [4-1:0] node33167;
	wire [4-1:0] node33170;
	wire [4-1:0] node33171;
	wire [4-1:0] node33172;
	wire [4-1:0] node33175;
	wire [4-1:0] node33178;
	wire [4-1:0] node33179;
	wire [4-1:0] node33182;
	wire [4-1:0] node33185;
	wire [4-1:0] node33186;
	wire [4-1:0] node33187;
	wire [4-1:0] node33188;
	wire [4-1:0] node33189;
	wire [4-1:0] node33192;
	wire [4-1:0] node33195;
	wire [4-1:0] node33196;
	wire [4-1:0] node33199;
	wire [4-1:0] node33202;
	wire [4-1:0] node33203;
	wire [4-1:0] node33204;
	wire [4-1:0] node33208;
	wire [4-1:0] node33209;
	wire [4-1:0] node33212;
	wire [4-1:0] node33215;
	wire [4-1:0] node33216;
	wire [4-1:0] node33217;
	wire [4-1:0] node33218;
	wire [4-1:0] node33221;
	wire [4-1:0] node33224;
	wire [4-1:0] node33225;
	wire [4-1:0] node33228;
	wire [4-1:0] node33231;
	wire [4-1:0] node33232;
	wire [4-1:0] node33233;
	wire [4-1:0] node33237;
	wire [4-1:0] node33238;
	wire [4-1:0] node33241;
	wire [4-1:0] node33244;
	wire [4-1:0] node33245;
	wire [4-1:0] node33246;
	wire [4-1:0] node33247;
	wire [4-1:0] node33248;
	wire [4-1:0] node33249;
	wire [4-1:0] node33253;
	wire [4-1:0] node33254;
	wire [4-1:0] node33257;
	wire [4-1:0] node33260;
	wire [4-1:0] node33261;
	wire [4-1:0] node33262;
	wire [4-1:0] node33265;
	wire [4-1:0] node33268;
	wire [4-1:0] node33269;
	wire [4-1:0] node33273;
	wire [4-1:0] node33274;
	wire [4-1:0] node33275;
	wire [4-1:0] node33276;
	wire [4-1:0] node33280;
	wire [4-1:0] node33281;
	wire [4-1:0] node33284;
	wire [4-1:0] node33287;
	wire [4-1:0] node33288;
	wire [4-1:0] node33289;
	wire [4-1:0] node33292;
	wire [4-1:0] node33295;
	wire [4-1:0] node33296;
	wire [4-1:0] node33299;
	wire [4-1:0] node33302;
	wire [4-1:0] node33303;
	wire [4-1:0] node33304;
	wire [4-1:0] node33305;
	wire [4-1:0] node33306;
	wire [4-1:0] node33310;
	wire [4-1:0] node33311;
	wire [4-1:0] node33314;
	wire [4-1:0] node33317;
	wire [4-1:0] node33318;
	wire [4-1:0] node33320;
	wire [4-1:0] node33323;
	wire [4-1:0] node33324;
	wire [4-1:0] node33327;
	wire [4-1:0] node33330;
	wire [4-1:0] node33331;
	wire [4-1:0] node33332;
	wire [4-1:0] node33333;
	wire [4-1:0] node33337;
	wire [4-1:0] node33338;
	wire [4-1:0] node33342;
	wire [4-1:0] node33343;
	wire [4-1:0] node33344;
	wire [4-1:0] node33348;
	wire [4-1:0] node33349;
	wire [4-1:0] node33353;
	wire [4-1:0] node33354;
	wire [4-1:0] node33355;
	wire [4-1:0] node33356;
	wire [4-1:0] node33357;
	wire [4-1:0] node33358;
	wire [4-1:0] node33359;
	wire [4-1:0] node33360;
	wire [4-1:0] node33363;
	wire [4-1:0] node33366;
	wire [4-1:0] node33367;
	wire [4-1:0] node33370;
	wire [4-1:0] node33373;
	wire [4-1:0] node33374;
	wire [4-1:0] node33376;
	wire [4-1:0] node33379;
	wire [4-1:0] node33381;
	wire [4-1:0] node33384;
	wire [4-1:0] node33385;
	wire [4-1:0] node33386;
	wire [4-1:0] node33388;
	wire [4-1:0] node33391;
	wire [4-1:0] node33393;
	wire [4-1:0] node33396;
	wire [4-1:0] node33397;
	wire [4-1:0] node33399;
	wire [4-1:0] node33402;
	wire [4-1:0] node33404;
	wire [4-1:0] node33407;
	wire [4-1:0] node33408;
	wire [4-1:0] node33409;
	wire [4-1:0] node33410;
	wire [4-1:0] node33411;
	wire [4-1:0] node33414;
	wire [4-1:0] node33417;
	wire [4-1:0] node33418;
	wire [4-1:0] node33421;
	wire [4-1:0] node33424;
	wire [4-1:0] node33425;
	wire [4-1:0] node33426;
	wire [4-1:0] node33429;
	wire [4-1:0] node33432;
	wire [4-1:0] node33433;
	wire [4-1:0] node33436;
	wire [4-1:0] node33439;
	wire [4-1:0] node33440;
	wire [4-1:0] node33441;
	wire [4-1:0] node33442;
	wire [4-1:0] node33445;
	wire [4-1:0] node33448;
	wire [4-1:0] node33449;
	wire [4-1:0] node33452;
	wire [4-1:0] node33455;
	wire [4-1:0] node33456;
	wire [4-1:0] node33457;
	wire [4-1:0] node33460;
	wire [4-1:0] node33463;
	wire [4-1:0] node33464;
	wire [4-1:0] node33467;
	wire [4-1:0] node33470;
	wire [4-1:0] node33471;
	wire [4-1:0] node33472;
	wire [4-1:0] node33473;
	wire [4-1:0] node33474;
	wire [4-1:0] node33476;
	wire [4-1:0] node33479;
	wire [4-1:0] node33481;
	wire [4-1:0] node33484;
	wire [4-1:0] node33485;
	wire [4-1:0] node33486;
	wire [4-1:0] node33490;
	wire [4-1:0] node33491;
	wire [4-1:0] node33494;
	wire [4-1:0] node33497;
	wire [4-1:0] node33498;
	wire [4-1:0] node33499;
	wire [4-1:0] node33500;
	wire [4-1:0] node33503;
	wire [4-1:0] node33506;
	wire [4-1:0] node33507;
	wire [4-1:0] node33510;
	wire [4-1:0] node33513;
	wire [4-1:0] node33514;
	wire [4-1:0] node33515;
	wire [4-1:0] node33518;
	wire [4-1:0] node33521;
	wire [4-1:0] node33522;
	wire [4-1:0] node33525;
	wire [4-1:0] node33528;
	wire [4-1:0] node33529;
	wire [4-1:0] node33530;
	wire [4-1:0] node33531;
	wire [4-1:0] node33532;
	wire [4-1:0] node33535;
	wire [4-1:0] node33538;
	wire [4-1:0] node33539;
	wire [4-1:0] node33542;
	wire [4-1:0] node33545;
	wire [4-1:0] node33546;
	wire [4-1:0] node33547;
	wire [4-1:0] node33550;
	wire [4-1:0] node33553;
	wire [4-1:0] node33554;
	wire [4-1:0] node33557;
	wire [4-1:0] node33560;
	wire [4-1:0] node33561;
	wire [4-1:0] node33562;
	wire [4-1:0] node33563;
	wire [4-1:0] node33566;
	wire [4-1:0] node33569;
	wire [4-1:0] node33570;
	wire [4-1:0] node33573;
	wire [4-1:0] node33576;
	wire [4-1:0] node33577;
	wire [4-1:0] node33578;
	wire [4-1:0] node33581;
	wire [4-1:0] node33584;
	wire [4-1:0] node33585;
	wire [4-1:0] node33588;
	wire [4-1:0] node33591;
	wire [4-1:0] node33592;
	wire [4-1:0] node33593;
	wire [4-1:0] node33594;
	wire [4-1:0] node33595;
	wire [4-1:0] node33596;
	wire [4-1:0] node33597;
	wire [4-1:0] node33600;
	wire [4-1:0] node33603;
	wire [4-1:0] node33605;
	wire [4-1:0] node33608;
	wire [4-1:0] node33609;
	wire [4-1:0] node33610;
	wire [4-1:0] node33613;
	wire [4-1:0] node33616;
	wire [4-1:0] node33617;
	wire [4-1:0] node33620;
	wire [4-1:0] node33623;
	wire [4-1:0] node33624;
	wire [4-1:0] node33625;
	wire [4-1:0] node33626;
	wire [4-1:0] node33629;
	wire [4-1:0] node33632;
	wire [4-1:0] node33633;
	wire [4-1:0] node33636;
	wire [4-1:0] node33639;
	wire [4-1:0] node33640;
	wire [4-1:0] node33641;
	wire [4-1:0] node33644;
	wire [4-1:0] node33647;
	wire [4-1:0] node33648;
	wire [4-1:0] node33652;
	wire [4-1:0] node33653;
	wire [4-1:0] node33654;
	wire [4-1:0] node33655;
	wire [4-1:0] node33656;
	wire [4-1:0] node33659;
	wire [4-1:0] node33662;
	wire [4-1:0] node33663;
	wire [4-1:0] node33667;
	wire [4-1:0] node33668;
	wire [4-1:0] node33669;
	wire [4-1:0] node33673;
	wire [4-1:0] node33674;
	wire [4-1:0] node33677;
	wire [4-1:0] node33680;
	wire [4-1:0] node33681;
	wire [4-1:0] node33682;
	wire [4-1:0] node33683;
	wire [4-1:0] node33686;
	wire [4-1:0] node33689;
	wire [4-1:0] node33690;
	wire [4-1:0] node33693;
	wire [4-1:0] node33696;
	wire [4-1:0] node33697;
	wire [4-1:0] node33698;
	wire [4-1:0] node33701;
	wire [4-1:0] node33704;
	wire [4-1:0] node33705;
	wire [4-1:0] node33708;
	wire [4-1:0] node33711;
	wire [4-1:0] node33712;
	wire [4-1:0] node33713;
	wire [4-1:0] node33714;
	wire [4-1:0] node33715;
	wire [4-1:0] node33716;
	wire [4-1:0] node33719;
	wire [4-1:0] node33722;
	wire [4-1:0] node33724;
	wire [4-1:0] node33727;
	wire [4-1:0] node33728;
	wire [4-1:0] node33729;
	wire [4-1:0] node33732;
	wire [4-1:0] node33735;
	wire [4-1:0] node33736;
	wire [4-1:0] node33739;
	wire [4-1:0] node33742;
	wire [4-1:0] node33743;
	wire [4-1:0] node33744;
	wire [4-1:0] node33745;
	wire [4-1:0] node33748;
	wire [4-1:0] node33751;
	wire [4-1:0] node33753;
	wire [4-1:0] node33756;
	wire [4-1:0] node33757;
	wire [4-1:0] node33758;
	wire [4-1:0] node33761;
	wire [4-1:0] node33764;
	wire [4-1:0] node33766;
	wire [4-1:0] node33769;
	wire [4-1:0] node33770;
	wire [4-1:0] node33771;
	wire [4-1:0] node33772;
	wire [4-1:0] node33773;
	wire [4-1:0] node33776;
	wire [4-1:0] node33779;
	wire [4-1:0] node33780;
	wire [4-1:0] node33783;
	wire [4-1:0] node33786;
	wire [4-1:0] node33787;
	wire [4-1:0] node33788;
	wire [4-1:0] node33792;
	wire [4-1:0] node33793;
	wire [4-1:0] node33796;
	wire [4-1:0] node33799;
	wire [4-1:0] node33800;
	wire [4-1:0] node33801;
	wire [4-1:0] node33802;
	wire [4-1:0] node33805;
	wire [4-1:0] node33808;
	wire [4-1:0] node33809;
	wire [4-1:0] node33812;
	wire [4-1:0] node33815;
	wire [4-1:0] node33816;
	wire [4-1:0] node33819;
	wire [4-1:0] node33822;
	wire [4-1:0] node33823;
	wire [4-1:0] node33824;
	wire [4-1:0] node33825;
	wire [4-1:0] node33826;
	wire [4-1:0] node33827;
	wire [4-1:0] node33828;
	wire [4-1:0] node33829;
	wire [4-1:0] node33830;
	wire [4-1:0] node33831;
	wire [4-1:0] node33834;
	wire [4-1:0] node33837;
	wire [4-1:0] node33838;
	wire [4-1:0] node33841;
	wire [4-1:0] node33844;
	wire [4-1:0] node33845;
	wire [4-1:0] node33846;
	wire [4-1:0] node33849;
	wire [4-1:0] node33852;
	wire [4-1:0] node33853;
	wire [4-1:0] node33857;
	wire [4-1:0] node33858;
	wire [4-1:0] node33859;
	wire [4-1:0] node33860;
	wire [4-1:0] node33863;
	wire [4-1:0] node33866;
	wire [4-1:0] node33867;
	wire [4-1:0] node33870;
	wire [4-1:0] node33873;
	wire [4-1:0] node33874;
	wire [4-1:0] node33875;
	wire [4-1:0] node33878;
	wire [4-1:0] node33881;
	wire [4-1:0] node33882;
	wire [4-1:0] node33885;
	wire [4-1:0] node33888;
	wire [4-1:0] node33889;
	wire [4-1:0] node33890;
	wire [4-1:0] node33891;
	wire [4-1:0] node33892;
	wire [4-1:0] node33895;
	wire [4-1:0] node33898;
	wire [4-1:0] node33899;
	wire [4-1:0] node33902;
	wire [4-1:0] node33905;
	wire [4-1:0] node33906;
	wire [4-1:0] node33907;
	wire [4-1:0] node33910;
	wire [4-1:0] node33913;
	wire [4-1:0] node33914;
	wire [4-1:0] node33917;
	wire [4-1:0] node33920;
	wire [4-1:0] node33921;
	wire [4-1:0] node33922;
	wire [4-1:0] node33923;
	wire [4-1:0] node33926;
	wire [4-1:0] node33929;
	wire [4-1:0] node33930;
	wire [4-1:0] node33934;
	wire [4-1:0] node33935;
	wire [4-1:0] node33936;
	wire [4-1:0] node33940;
	wire [4-1:0] node33942;
	wire [4-1:0] node33945;
	wire [4-1:0] node33946;
	wire [4-1:0] node33947;
	wire [4-1:0] node33948;
	wire [4-1:0] node33949;
	wire [4-1:0] node33950;
	wire [4-1:0] node33953;
	wire [4-1:0] node33956;
	wire [4-1:0] node33957;
	wire [4-1:0] node33960;
	wire [4-1:0] node33963;
	wire [4-1:0] node33964;
	wire [4-1:0] node33965;
	wire [4-1:0] node33968;
	wire [4-1:0] node33971;
	wire [4-1:0] node33972;
	wire [4-1:0] node33975;
	wire [4-1:0] node33978;
	wire [4-1:0] node33979;
	wire [4-1:0] node33980;
	wire [4-1:0] node33981;
	wire [4-1:0] node33985;
	wire [4-1:0] node33986;
	wire [4-1:0] node33989;
	wire [4-1:0] node33992;
	wire [4-1:0] node33993;
	wire [4-1:0] node33994;
	wire [4-1:0] node33997;
	wire [4-1:0] node34000;
	wire [4-1:0] node34001;
	wire [4-1:0] node34004;
	wire [4-1:0] node34007;
	wire [4-1:0] node34008;
	wire [4-1:0] node34009;
	wire [4-1:0] node34010;
	wire [4-1:0] node34013;
	wire [4-1:0] node34016;
	wire [4-1:0] node34017;
	wire [4-1:0] node34018;
	wire [4-1:0] node34021;
	wire [4-1:0] node34024;
	wire [4-1:0] node34025;
	wire [4-1:0] node34028;
	wire [4-1:0] node34031;
	wire [4-1:0] node34032;
	wire [4-1:0] node34033;
	wire [4-1:0] node34036;
	wire [4-1:0] node34039;
	wire [4-1:0] node34040;
	wire [4-1:0] node34041;
	wire [4-1:0] node34044;
	wire [4-1:0] node34047;
	wire [4-1:0] node34048;
	wire [4-1:0] node34051;
	wire [4-1:0] node34054;
	wire [4-1:0] node34055;
	wire [4-1:0] node34056;
	wire [4-1:0] node34057;
	wire [4-1:0] node34058;
	wire [4-1:0] node34059;
	wire [4-1:0] node34061;
	wire [4-1:0] node34064;
	wire [4-1:0] node34065;
	wire [4-1:0] node34068;
	wire [4-1:0] node34071;
	wire [4-1:0] node34072;
	wire [4-1:0] node34074;
	wire [4-1:0] node34077;
	wire [4-1:0] node34078;
	wire [4-1:0] node34081;
	wire [4-1:0] node34084;
	wire [4-1:0] node34085;
	wire [4-1:0] node34086;
	wire [4-1:0] node34087;
	wire [4-1:0] node34090;
	wire [4-1:0] node34093;
	wire [4-1:0] node34094;
	wire [4-1:0] node34097;
	wire [4-1:0] node34100;
	wire [4-1:0] node34101;
	wire [4-1:0] node34102;
	wire [4-1:0] node34105;
	wire [4-1:0] node34108;
	wire [4-1:0] node34109;
	wire [4-1:0] node34112;
	wire [4-1:0] node34115;
	wire [4-1:0] node34116;
	wire [4-1:0] node34117;
	wire [4-1:0] node34118;
	wire [4-1:0] node34119;
	wire [4-1:0] node34122;
	wire [4-1:0] node34125;
	wire [4-1:0] node34126;
	wire [4-1:0] node34130;
	wire [4-1:0] node34131;
	wire [4-1:0] node34134;
	wire [4-1:0] node34135;
	wire [4-1:0] node34138;
	wire [4-1:0] node34141;
	wire [4-1:0] node34142;
	wire [4-1:0] node34143;
	wire [4-1:0] node34144;
	wire [4-1:0] node34147;
	wire [4-1:0] node34150;
	wire [4-1:0] node34152;
	wire [4-1:0] node34155;
	wire [4-1:0] node34156;
	wire [4-1:0] node34159;
	wire [4-1:0] node34162;
	wire [4-1:0] node34163;
	wire [4-1:0] node34164;
	wire [4-1:0] node34165;
	wire [4-1:0] node34166;
	wire [4-1:0] node34167;
	wire [4-1:0] node34170;
	wire [4-1:0] node34173;
	wire [4-1:0] node34175;
	wire [4-1:0] node34178;
	wire [4-1:0] node34179;
	wire [4-1:0] node34181;
	wire [4-1:0] node34184;
	wire [4-1:0] node34186;
	wire [4-1:0] node34189;
	wire [4-1:0] node34190;
	wire [4-1:0] node34191;
	wire [4-1:0] node34192;
	wire [4-1:0] node34195;
	wire [4-1:0] node34198;
	wire [4-1:0] node34199;
	wire [4-1:0] node34202;
	wire [4-1:0] node34205;
	wire [4-1:0] node34206;
	wire [4-1:0] node34209;
	wire [4-1:0] node34212;
	wire [4-1:0] node34213;
	wire [4-1:0] node34214;
	wire [4-1:0] node34215;
	wire [4-1:0] node34216;
	wire [4-1:0] node34220;
	wire [4-1:0] node34221;
	wire [4-1:0] node34224;
	wire [4-1:0] node34227;
	wire [4-1:0] node34228;
	wire [4-1:0] node34229;
	wire [4-1:0] node34232;
	wire [4-1:0] node34235;
	wire [4-1:0] node34237;
	wire [4-1:0] node34240;
	wire [4-1:0] node34241;
	wire [4-1:0] node34242;
	wire [4-1:0] node34243;
	wire [4-1:0] node34247;
	wire [4-1:0] node34248;
	wire [4-1:0] node34252;
	wire [4-1:0] node34253;
	wire [4-1:0] node34254;
	wire [4-1:0] node34258;
	wire [4-1:0] node34259;
	wire [4-1:0] node34263;
	wire [4-1:0] node34264;
	wire [4-1:0] node34265;
	wire [4-1:0] node34266;
	wire [4-1:0] node34267;
	wire [4-1:0] node34268;
	wire [4-1:0] node34269;
	wire [4-1:0] node34270;
	wire [4-1:0] node34273;
	wire [4-1:0] node34276;
	wire [4-1:0] node34277;
	wire [4-1:0] node34280;
	wire [4-1:0] node34283;
	wire [4-1:0] node34284;
	wire [4-1:0] node34285;
	wire [4-1:0] node34288;
	wire [4-1:0] node34291;
	wire [4-1:0] node34294;
	wire [4-1:0] node34295;
	wire [4-1:0] node34296;
	wire [4-1:0] node34297;
	wire [4-1:0] node34300;
	wire [4-1:0] node34303;
	wire [4-1:0] node34305;
	wire [4-1:0] node34308;
	wire [4-1:0] node34309;
	wire [4-1:0] node34311;
	wire [4-1:0] node34314;
	wire [4-1:0] node34315;
	wire [4-1:0] node34318;
	wire [4-1:0] node34321;
	wire [4-1:0] node34322;
	wire [4-1:0] node34323;
	wire [4-1:0] node34324;
	wire [4-1:0] node34325;
	wire [4-1:0] node34328;
	wire [4-1:0] node34331;
	wire [4-1:0] node34332;
	wire [4-1:0] node34335;
	wire [4-1:0] node34338;
	wire [4-1:0] node34339;
	wire [4-1:0] node34340;
	wire [4-1:0] node34343;
	wire [4-1:0] node34346;
	wire [4-1:0] node34347;
	wire [4-1:0] node34350;
	wire [4-1:0] node34353;
	wire [4-1:0] node34354;
	wire [4-1:0] node34355;
	wire [4-1:0] node34356;
	wire [4-1:0] node34360;
	wire [4-1:0] node34361;
	wire [4-1:0] node34365;
	wire [4-1:0] node34366;
	wire [4-1:0] node34367;
	wire [4-1:0] node34371;
	wire [4-1:0] node34372;
	wire [4-1:0] node34376;
	wire [4-1:0] node34377;
	wire [4-1:0] node34378;
	wire [4-1:0] node34379;
	wire [4-1:0] node34380;
	wire [4-1:0] node34382;
	wire [4-1:0] node34385;
	wire [4-1:0] node34386;
	wire [4-1:0] node34389;
	wire [4-1:0] node34392;
	wire [4-1:0] node34393;
	wire [4-1:0] node34394;
	wire [4-1:0] node34397;
	wire [4-1:0] node34400;
	wire [4-1:0] node34401;
	wire [4-1:0] node34404;
	wire [4-1:0] node34407;
	wire [4-1:0] node34408;
	wire [4-1:0] node34409;
	wire [4-1:0] node34411;
	wire [4-1:0] node34414;
	wire [4-1:0] node34415;
	wire [4-1:0] node34418;
	wire [4-1:0] node34421;
	wire [4-1:0] node34422;
	wire [4-1:0] node34423;
	wire [4-1:0] node34426;
	wire [4-1:0] node34429;
	wire [4-1:0] node34430;
	wire [4-1:0] node34433;
	wire [4-1:0] node34436;
	wire [4-1:0] node34437;
	wire [4-1:0] node34438;
	wire [4-1:0] node34439;
	wire [4-1:0] node34440;
	wire [4-1:0] node34443;
	wire [4-1:0] node34446;
	wire [4-1:0] node34447;
	wire [4-1:0] node34450;
	wire [4-1:0] node34453;
	wire [4-1:0] node34454;
	wire [4-1:0] node34455;
	wire [4-1:0] node34458;
	wire [4-1:0] node34461;
	wire [4-1:0] node34463;
	wire [4-1:0] node34466;
	wire [4-1:0] node34467;
	wire [4-1:0] node34468;
	wire [4-1:0] node34469;
	wire [4-1:0] node34473;
	wire [4-1:0] node34474;
	wire [4-1:0] node34478;
	wire [4-1:0] node34479;
	wire [4-1:0] node34480;
	wire [4-1:0] node34484;
	wire [4-1:0] node34485;
	wire [4-1:0] node34489;
	wire [4-1:0] node34490;
	wire [4-1:0] node34491;
	wire [4-1:0] node34492;
	wire [4-1:0] node34493;
	wire [4-1:0] node34494;
	wire [4-1:0] node34495;
	wire [4-1:0] node34498;
	wire [4-1:0] node34501;
	wire [4-1:0] node34502;
	wire [4-1:0] node34505;
	wire [4-1:0] node34508;
	wire [4-1:0] node34509;
	wire [4-1:0] node34510;
	wire [4-1:0] node34513;
	wire [4-1:0] node34516;
	wire [4-1:0] node34517;
	wire [4-1:0] node34520;
	wire [4-1:0] node34523;
	wire [4-1:0] node34524;
	wire [4-1:0] node34525;
	wire [4-1:0] node34526;
	wire [4-1:0] node34529;
	wire [4-1:0] node34532;
	wire [4-1:0] node34533;
	wire [4-1:0] node34537;
	wire [4-1:0] node34538;
	wire [4-1:0] node34539;
	wire [4-1:0] node34542;
	wire [4-1:0] node34545;
	wire [4-1:0] node34546;
	wire [4-1:0] node34549;
	wire [4-1:0] node34552;
	wire [4-1:0] node34553;
	wire [4-1:0] node34554;
	wire [4-1:0] node34555;
	wire [4-1:0] node34556;
	wire [4-1:0] node34559;
	wire [4-1:0] node34562;
	wire [4-1:0] node34563;
	wire [4-1:0] node34566;
	wire [4-1:0] node34569;
	wire [4-1:0] node34570;
	wire [4-1:0] node34571;
	wire [4-1:0] node34574;
	wire [4-1:0] node34577;
	wire [4-1:0] node34578;
	wire [4-1:0] node34581;
	wire [4-1:0] node34584;
	wire [4-1:0] node34585;
	wire [4-1:0] node34586;
	wire [4-1:0] node34587;
	wire [4-1:0] node34590;
	wire [4-1:0] node34593;
	wire [4-1:0] node34594;
	wire [4-1:0] node34597;
	wire [4-1:0] node34600;
	wire [4-1:0] node34601;
	wire [4-1:0] node34602;
	wire [4-1:0] node34606;
	wire [4-1:0] node34608;
	wire [4-1:0] node34611;
	wire [4-1:0] node34612;
	wire [4-1:0] node34613;
	wire [4-1:0] node34614;
	wire [4-1:0] node34615;
	wire [4-1:0] node34616;
	wire [4-1:0] node34620;
	wire [4-1:0] node34621;
	wire [4-1:0] node34625;
	wire [4-1:0] node34626;
	wire [4-1:0] node34627;
	wire [4-1:0] node34631;
	wire [4-1:0] node34632;
	wire [4-1:0] node34636;
	wire [4-1:0] node34637;
	wire [4-1:0] node34638;
	wire [4-1:0] node34639;
	wire [4-1:0] node34643;
	wire [4-1:0] node34644;
	wire [4-1:0] node34648;
	wire [4-1:0] node34649;
	wire [4-1:0] node34650;
	wire [4-1:0] node34654;
	wire [4-1:0] node34655;
	wire [4-1:0] node34659;
	wire [4-1:0] node34660;
	wire [4-1:0] node34661;
	wire [4-1:0] node34662;
	wire [4-1:0] node34663;
	wire [4-1:0] node34666;
	wire [4-1:0] node34669;
	wire [4-1:0] node34671;
	wire [4-1:0] node34674;
	wire [4-1:0] node34675;
	wire [4-1:0] node34678;
	wire [4-1:0] node34681;
	wire [4-1:0] node34682;
	wire [4-1:0] node34683;
	wire [4-1:0] node34684;
	wire [4-1:0] node34687;
	wire [4-1:0] node34690;
	wire [4-1:0] node34691;
	wire [4-1:0] node34694;
	wire [4-1:0] node34697;
	wire [4-1:0] node34698;
	wire [4-1:0] node34699;
	wire [4-1:0] node34702;
	wire [4-1:0] node34705;
	wire [4-1:0] node34706;
	wire [4-1:0] node34709;
	wire [4-1:0] node34712;
	wire [4-1:0] node34713;
	wire [4-1:0] node34714;
	wire [4-1:0] node34715;
	wire [4-1:0] node34716;
	wire [4-1:0] node34717;
	wire [4-1:0] node34718;
	wire [4-1:0] node34719;
	wire [4-1:0] node34720;
	wire [4-1:0] node34723;
	wire [4-1:0] node34726;
	wire [4-1:0] node34727;
	wire [4-1:0] node34730;
	wire [4-1:0] node34733;
	wire [4-1:0] node34734;
	wire [4-1:0] node34735;
	wire [4-1:0] node34738;
	wire [4-1:0] node34741;
	wire [4-1:0] node34742;
	wire [4-1:0] node34745;
	wire [4-1:0] node34748;
	wire [4-1:0] node34749;
	wire [4-1:0] node34750;
	wire [4-1:0] node34751;
	wire [4-1:0] node34754;
	wire [4-1:0] node34757;
	wire [4-1:0] node34759;
	wire [4-1:0] node34762;
	wire [4-1:0] node34763;
	wire [4-1:0] node34764;
	wire [4-1:0] node34767;
	wire [4-1:0] node34770;
	wire [4-1:0] node34772;
	wire [4-1:0] node34775;
	wire [4-1:0] node34776;
	wire [4-1:0] node34777;
	wire [4-1:0] node34778;
	wire [4-1:0] node34779;
	wire [4-1:0] node34782;
	wire [4-1:0] node34785;
	wire [4-1:0] node34786;
	wire [4-1:0] node34789;
	wire [4-1:0] node34792;
	wire [4-1:0] node34793;
	wire [4-1:0] node34794;
	wire [4-1:0] node34797;
	wire [4-1:0] node34800;
	wire [4-1:0] node34801;
	wire [4-1:0] node34804;
	wire [4-1:0] node34807;
	wire [4-1:0] node34808;
	wire [4-1:0] node34809;
	wire [4-1:0] node34811;
	wire [4-1:0] node34814;
	wire [4-1:0] node34815;
	wire [4-1:0] node34818;
	wire [4-1:0] node34821;
	wire [4-1:0] node34822;
	wire [4-1:0] node34823;
	wire [4-1:0] node34826;
	wire [4-1:0] node34829;
	wire [4-1:0] node34830;
	wire [4-1:0] node34833;
	wire [4-1:0] node34836;
	wire [4-1:0] node34837;
	wire [4-1:0] node34838;
	wire [4-1:0] node34839;
	wire [4-1:0] node34840;
	wire [4-1:0] node34841;
	wire [4-1:0] node34844;
	wire [4-1:0] node34847;
	wire [4-1:0] node34848;
	wire [4-1:0] node34851;
	wire [4-1:0] node34854;
	wire [4-1:0] node34855;
	wire [4-1:0] node34856;
	wire [4-1:0] node34860;
	wire [4-1:0] node34861;
	wire [4-1:0] node34864;
	wire [4-1:0] node34867;
	wire [4-1:0] node34868;
	wire [4-1:0] node34869;
	wire [4-1:0] node34870;
	wire [4-1:0] node34873;
	wire [4-1:0] node34876;
	wire [4-1:0] node34877;
	wire [4-1:0] node34880;
	wire [4-1:0] node34883;
	wire [4-1:0] node34884;
	wire [4-1:0] node34885;
	wire [4-1:0] node34888;
	wire [4-1:0] node34891;
	wire [4-1:0] node34892;
	wire [4-1:0] node34895;
	wire [4-1:0] node34898;
	wire [4-1:0] node34899;
	wire [4-1:0] node34900;
	wire [4-1:0] node34901;
	wire [4-1:0] node34902;
	wire [4-1:0] node34905;
	wire [4-1:0] node34908;
	wire [4-1:0] node34909;
	wire [4-1:0] node34912;
	wire [4-1:0] node34915;
	wire [4-1:0] node34916;
	wire [4-1:0] node34917;
	wire [4-1:0] node34921;
	wire [4-1:0] node34922;
	wire [4-1:0] node34925;
	wire [4-1:0] node34928;
	wire [4-1:0] node34929;
	wire [4-1:0] node34930;
	wire [4-1:0] node34933;
	wire [4-1:0] node34936;
	wire [4-1:0] node34937;
	wire [4-1:0] node34938;
	wire [4-1:0] node34941;
	wire [4-1:0] node34944;
	wire [4-1:0] node34945;
	wire [4-1:0] node34948;
	wire [4-1:0] node34951;
	wire [4-1:0] node34952;
	wire [4-1:0] node34953;
	wire [4-1:0] node34954;
	wire [4-1:0] node34955;
	wire [4-1:0] node34956;
	wire [4-1:0] node34957;
	wire [4-1:0] node34960;
	wire [4-1:0] node34963;
	wire [4-1:0] node34964;
	wire [4-1:0] node34967;
	wire [4-1:0] node34970;
	wire [4-1:0] node34971;
	wire [4-1:0] node34972;
	wire [4-1:0] node34975;
	wire [4-1:0] node34978;
	wire [4-1:0] node34980;
	wire [4-1:0] node34983;
	wire [4-1:0] node34984;
	wire [4-1:0] node34985;
	wire [4-1:0] node34986;
	wire [4-1:0] node34990;
	wire [4-1:0] node34991;
	wire [4-1:0] node34995;
	wire [4-1:0] node34996;
	wire [4-1:0] node34997;
	wire [4-1:0] node35001;
	wire [4-1:0] node35002;
	wire [4-1:0] node35006;
	wire [4-1:0] node35007;
	wire [4-1:0] node35008;
	wire [4-1:0] node35009;
	wire [4-1:0] node35010;
	wire [4-1:0] node35013;
	wire [4-1:0] node35016;
	wire [4-1:0] node35017;
	wire [4-1:0] node35020;
	wire [4-1:0] node35023;
	wire [4-1:0] node35024;
	wire [4-1:0] node35025;
	wire [4-1:0] node35029;
	wire [4-1:0] node35030;
	wire [4-1:0] node35033;
	wire [4-1:0] node35036;
	wire [4-1:0] node35037;
	wire [4-1:0] node35038;
	wire [4-1:0] node35039;
	wire [4-1:0] node35042;
	wire [4-1:0] node35045;
	wire [4-1:0] node35046;
	wire [4-1:0] node35049;
	wire [4-1:0] node35052;
	wire [4-1:0] node35053;
	wire [4-1:0] node35054;
	wire [4-1:0] node35057;
	wire [4-1:0] node35060;
	wire [4-1:0] node35062;
	wire [4-1:0] node35065;
	wire [4-1:0] node35066;
	wire [4-1:0] node35067;
	wire [4-1:0] node35068;
	wire [4-1:0] node35069;
	wire [4-1:0] node35070;
	wire [4-1:0] node35073;
	wire [4-1:0] node35076;
	wire [4-1:0] node35077;
	wire [4-1:0] node35080;
	wire [4-1:0] node35083;
	wire [4-1:0] node35084;
	wire [4-1:0] node35085;
	wire [4-1:0] node35088;
	wire [4-1:0] node35091;
	wire [4-1:0] node35092;
	wire [4-1:0] node35095;
	wire [4-1:0] node35098;
	wire [4-1:0] node35099;
	wire [4-1:0] node35100;
	wire [4-1:0] node35101;
	wire [4-1:0] node35105;
	wire [4-1:0] node35106;
	wire [4-1:0] node35110;
	wire [4-1:0] node35111;
	wire [4-1:0] node35112;
	wire [4-1:0] node35116;
	wire [4-1:0] node35117;
	wire [4-1:0] node35121;
	wire [4-1:0] node35122;
	wire [4-1:0] node35123;
	wire [4-1:0] node35124;
	wire [4-1:0] node35126;
	wire [4-1:0] node35129;
	wire [4-1:0] node35130;
	wire [4-1:0] node35133;
	wire [4-1:0] node35136;
	wire [4-1:0] node35137;
	wire [4-1:0] node35138;
	wire [4-1:0] node35141;
	wire [4-1:0] node35144;
	wire [4-1:0] node35145;
	wire [4-1:0] node35149;
	wire [4-1:0] node35150;
	wire [4-1:0] node35151;
	wire [4-1:0] node35152;
	wire [4-1:0] node35155;
	wire [4-1:0] node35158;
	wire [4-1:0] node35159;
	wire [4-1:0] node35162;
	wire [4-1:0] node35165;
	wire [4-1:0] node35166;
	wire [4-1:0] node35167;
	wire [4-1:0] node35170;
	wire [4-1:0] node35173;
	wire [4-1:0] node35174;
	wire [4-1:0] node35177;
	wire [4-1:0] node35180;
	wire [4-1:0] node35181;
	wire [4-1:0] node35182;
	wire [4-1:0] node35183;
	wire [4-1:0] node35184;
	wire [4-1:0] node35185;
	wire [4-1:0] node35186;
	wire [4-1:0] node35187;
	wire [4-1:0] node35190;
	wire [4-1:0] node35193;
	wire [4-1:0] node35194;
	wire [4-1:0] node35197;
	wire [4-1:0] node35200;
	wire [4-1:0] node35201;
	wire [4-1:0] node35202;
	wire [4-1:0] node35206;
	wire [4-1:0] node35207;
	wire [4-1:0] node35210;
	wire [4-1:0] node35213;
	wire [4-1:0] node35214;
	wire [4-1:0] node35215;
	wire [4-1:0] node35216;
	wire [4-1:0] node35220;
	wire [4-1:0] node35221;
	wire [4-1:0] node35224;
	wire [4-1:0] node35227;
	wire [4-1:0] node35228;
	wire [4-1:0] node35229;
	wire [4-1:0] node35232;
	wire [4-1:0] node35235;
	wire [4-1:0] node35236;
	wire [4-1:0] node35240;
	wire [4-1:0] node35241;
	wire [4-1:0] node35242;
	wire [4-1:0] node35243;
	wire [4-1:0] node35244;
	wire [4-1:0] node35247;
	wire [4-1:0] node35250;
	wire [4-1:0] node35251;
	wire [4-1:0] node35254;
	wire [4-1:0] node35257;
	wire [4-1:0] node35258;
	wire [4-1:0] node35259;
	wire [4-1:0] node35262;
	wire [4-1:0] node35265;
	wire [4-1:0] node35267;
	wire [4-1:0] node35270;
	wire [4-1:0] node35271;
	wire [4-1:0] node35272;
	wire [4-1:0] node35273;
	wire [4-1:0] node35277;
	wire [4-1:0] node35278;
	wire [4-1:0] node35282;
	wire [4-1:0] node35283;
	wire [4-1:0] node35284;
	wire [4-1:0] node35288;
	wire [4-1:0] node35289;
	wire [4-1:0] node35293;
	wire [4-1:0] node35294;
	wire [4-1:0] node35295;
	wire [4-1:0] node35296;
	wire [4-1:0] node35297;
	wire [4-1:0] node35298;
	wire [4-1:0] node35301;
	wire [4-1:0] node35304;
	wire [4-1:0] node35305;
	wire [4-1:0] node35308;
	wire [4-1:0] node35311;
	wire [4-1:0] node35312;
	wire [4-1:0] node35313;
	wire [4-1:0] node35316;
	wire [4-1:0] node35319;
	wire [4-1:0] node35321;
	wire [4-1:0] node35324;
	wire [4-1:0] node35325;
	wire [4-1:0] node35326;
	wire [4-1:0] node35327;
	wire [4-1:0] node35331;
	wire [4-1:0] node35332;
	wire [4-1:0] node35336;
	wire [4-1:0] node35337;
	wire [4-1:0] node35338;
	wire [4-1:0] node35342;
	wire [4-1:0] node35343;
	wire [4-1:0] node35347;
	wire [4-1:0] node35348;
	wire [4-1:0] node35349;
	wire [4-1:0] node35350;
	wire [4-1:0] node35351;
	wire [4-1:0] node35354;
	wire [4-1:0] node35357;
	wire [4-1:0] node35358;
	wire [4-1:0] node35361;
	wire [4-1:0] node35364;
	wire [4-1:0] node35365;
	wire [4-1:0] node35366;
	wire [4-1:0] node35370;
	wire [4-1:0] node35371;
	wire [4-1:0] node35374;
	wire [4-1:0] node35377;
	wire [4-1:0] node35378;
	wire [4-1:0] node35379;
	wire [4-1:0] node35380;
	wire [4-1:0] node35383;
	wire [4-1:0] node35386;
	wire [4-1:0] node35387;
	wire [4-1:0] node35390;
	wire [4-1:0] node35393;
	wire [4-1:0] node35394;
	wire [4-1:0] node35395;
	wire [4-1:0] node35398;
	wire [4-1:0] node35401;
	wire [4-1:0] node35402;
	wire [4-1:0] node35405;
	wire [4-1:0] node35408;
	wire [4-1:0] node35409;
	wire [4-1:0] node35410;
	wire [4-1:0] node35411;
	wire [4-1:0] node35412;
	wire [4-1:0] node35413;
	wire [4-1:0] node35414;
	wire [4-1:0] node35417;
	wire [4-1:0] node35420;
	wire [4-1:0] node35421;
	wire [4-1:0] node35424;
	wire [4-1:0] node35427;
	wire [4-1:0] node35428;
	wire [4-1:0] node35429;
	wire [4-1:0] node35432;
	wire [4-1:0] node35435;
	wire [4-1:0] node35436;
	wire [4-1:0] node35439;
	wire [4-1:0] node35442;
	wire [4-1:0] node35443;
	wire [4-1:0] node35444;
	wire [4-1:0] node35445;
	wire [4-1:0] node35448;
	wire [4-1:0] node35451;
	wire [4-1:0] node35452;
	wire [4-1:0] node35455;
	wire [4-1:0] node35458;
	wire [4-1:0] node35459;
	wire [4-1:0] node35460;
	wire [4-1:0] node35463;
	wire [4-1:0] node35466;
	wire [4-1:0] node35467;
	wire [4-1:0] node35470;
	wire [4-1:0] node35473;
	wire [4-1:0] node35474;
	wire [4-1:0] node35475;
	wire [4-1:0] node35476;
	wire [4-1:0] node35477;
	wire [4-1:0] node35480;
	wire [4-1:0] node35483;
	wire [4-1:0] node35484;
	wire [4-1:0] node35487;
	wire [4-1:0] node35490;
	wire [4-1:0] node35491;
	wire [4-1:0] node35492;
	wire [4-1:0] node35495;
	wire [4-1:0] node35498;
	wire [4-1:0] node35499;
	wire [4-1:0] node35503;
	wire [4-1:0] node35504;
	wire [4-1:0] node35505;
	wire [4-1:0] node35507;
	wire [4-1:0] node35510;
	wire [4-1:0] node35511;
	wire [4-1:0] node35514;
	wire [4-1:0] node35517;
	wire [4-1:0] node35518;
	wire [4-1:0] node35519;
	wire [4-1:0] node35522;
	wire [4-1:0] node35525;
	wire [4-1:0] node35526;
	wire [4-1:0] node35529;
	wire [4-1:0] node35532;
	wire [4-1:0] node35533;
	wire [4-1:0] node35534;
	wire [4-1:0] node35535;
	wire [4-1:0] node35536;
	wire [4-1:0] node35537;
	wire [4-1:0] node35540;
	wire [4-1:0] node35543;
	wire [4-1:0] node35544;
	wire [4-1:0] node35547;
	wire [4-1:0] node35550;
	wire [4-1:0] node35551;
	wire [4-1:0] node35552;
	wire [4-1:0] node35556;
	wire [4-1:0] node35557;
	wire [4-1:0] node35560;
	wire [4-1:0] node35563;
	wire [4-1:0] node35564;
	wire [4-1:0] node35565;
	wire [4-1:0] node35566;
	wire [4-1:0] node35569;
	wire [4-1:0] node35572;
	wire [4-1:0] node35573;
	wire [4-1:0] node35576;
	wire [4-1:0] node35579;
	wire [4-1:0] node35580;
	wire [4-1:0] node35581;
	wire [4-1:0] node35584;
	wire [4-1:0] node35587;
	wire [4-1:0] node35588;
	wire [4-1:0] node35591;
	wire [4-1:0] node35594;
	wire [4-1:0] node35595;
	wire [4-1:0] node35596;
	wire [4-1:0] node35597;
	wire [4-1:0] node35598;
	wire [4-1:0] node35601;
	wire [4-1:0] node35604;
	wire [4-1:0] node35605;
	wire [4-1:0] node35608;
	wire [4-1:0] node35611;
	wire [4-1:0] node35612;
	wire [4-1:0] node35613;
	wire [4-1:0] node35616;
	wire [4-1:0] node35619;
	wire [4-1:0] node35620;
	wire [4-1:0] node35623;
	wire [4-1:0] node35626;
	wire [4-1:0] node35627;
	wire [4-1:0] node35628;
	wire [4-1:0] node35629;
	wire [4-1:0] node35632;
	wire [4-1:0] node35635;
	wire [4-1:0] node35636;
	wire [4-1:0] node35639;
	wire [4-1:0] node35642;
	wire [4-1:0] node35643;
	wire [4-1:0] node35644;
	wire [4-1:0] node35647;
	wire [4-1:0] node35650;
	wire [4-1:0] node35651;
	wire [4-1:0] node35654;
	wire [4-1:0] node35657;
	wire [4-1:0] node35658;
	wire [4-1:0] node35659;
	wire [4-1:0] node35660;
	wire [4-1:0] node35661;
	wire [4-1:0] node35662;
	wire [4-1:0] node35663;
	wire [4-1:0] node35664;
	wire [4-1:0] node35665;
	wire [4-1:0] node35666;
	wire [4-1:0] node35667;
	wire [4-1:0] node35668;
	wire [4-1:0] node35672;
	wire [4-1:0] node35673;
	wire [4-1:0] node35677;
	wire [4-1:0] node35678;
	wire [4-1:0] node35679;
	wire [4-1:0] node35683;
	wire [4-1:0] node35684;
	wire [4-1:0] node35688;
	wire [4-1:0] node35689;
	wire [4-1:0] node35690;
	wire [4-1:0] node35691;
	wire [4-1:0] node35694;
	wire [4-1:0] node35697;
	wire [4-1:0] node35698;
	wire [4-1:0] node35701;
	wire [4-1:0] node35704;
	wire [4-1:0] node35705;
	wire [4-1:0] node35706;
	wire [4-1:0] node35709;
	wire [4-1:0] node35712;
	wire [4-1:0] node35713;
	wire [4-1:0] node35716;
	wire [4-1:0] node35719;
	wire [4-1:0] node35720;
	wire [4-1:0] node35721;
	wire [4-1:0] node35722;
	wire [4-1:0] node35723;
	wire [4-1:0] node35726;
	wire [4-1:0] node35729;
	wire [4-1:0] node35730;
	wire [4-1:0] node35733;
	wire [4-1:0] node35736;
	wire [4-1:0] node35737;
	wire [4-1:0] node35740;
	wire [4-1:0] node35743;
	wire [4-1:0] node35744;
	wire [4-1:0] node35745;
	wire [4-1:0] node35746;
	wire [4-1:0] node35749;
	wire [4-1:0] node35752;
	wire [4-1:0] node35754;
	wire [4-1:0] node35757;
	wire [4-1:0] node35758;
	wire [4-1:0] node35759;
	wire [4-1:0] node35763;
	wire [4-1:0] node35764;
	wire [4-1:0] node35767;
	wire [4-1:0] node35770;
	wire [4-1:0] node35771;
	wire [4-1:0] node35772;
	wire [4-1:0] node35773;
	wire [4-1:0] node35774;
	wire [4-1:0] node35775;
	wire [4-1:0] node35779;
	wire [4-1:0] node35780;
	wire [4-1:0] node35784;
	wire [4-1:0] node35785;
	wire [4-1:0] node35786;
	wire [4-1:0] node35790;
	wire [4-1:0] node35791;
	wire [4-1:0] node35795;
	wire [4-1:0] node35796;
	wire [4-1:0] node35797;
	wire [4-1:0] node35798;
	wire [4-1:0] node35801;
	wire [4-1:0] node35804;
	wire [4-1:0] node35806;
	wire [4-1:0] node35809;
	wire [4-1:0] node35810;
	wire [4-1:0] node35811;
	wire [4-1:0] node35815;
	wire [4-1:0] node35816;
	wire [4-1:0] node35820;
	wire [4-1:0] node35821;
	wire [4-1:0] node35822;
	wire [4-1:0] node35823;
	wire [4-1:0] node35824;
	wire [4-1:0] node35828;
	wire [4-1:0] node35829;
	wire [4-1:0] node35833;
	wire [4-1:0] node35834;
	wire [4-1:0] node35835;
	wire [4-1:0] node35839;
	wire [4-1:0] node35840;
	wire [4-1:0] node35844;
	wire [4-1:0] node35845;
	wire [4-1:0] node35846;
	wire [4-1:0] node35847;
	wire [4-1:0] node35850;
	wire [4-1:0] node35853;
	wire [4-1:0] node35854;
	wire [4-1:0] node35858;
	wire [4-1:0] node35859;
	wire [4-1:0] node35860;
	wire [4-1:0] node35863;
	wire [4-1:0] node35866;
	wire [4-1:0] node35867;
	wire [4-1:0] node35870;
	wire [4-1:0] node35873;
	wire [4-1:0] node35874;
	wire [4-1:0] node35875;
	wire [4-1:0] node35876;
	wire [4-1:0] node35877;
	wire [4-1:0] node35878;
	wire [4-1:0] node35879;
	wire [4-1:0] node35882;
	wire [4-1:0] node35885;
	wire [4-1:0] node35887;
	wire [4-1:0] node35890;
	wire [4-1:0] node35891;
	wire [4-1:0] node35892;
	wire [4-1:0] node35896;
	wire [4-1:0] node35897;
	wire [4-1:0] node35900;
	wire [4-1:0] node35903;
	wire [4-1:0] node35904;
	wire [4-1:0] node35905;
	wire [4-1:0] node35908;
	wire [4-1:0] node35911;
	wire [4-1:0] node35912;
	wire [4-1:0] node35914;
	wire [4-1:0] node35917;
	wire [4-1:0] node35918;
	wire [4-1:0] node35921;
	wire [4-1:0] node35924;
	wire [4-1:0] node35925;
	wire [4-1:0] node35926;
	wire [4-1:0] node35927;
	wire [4-1:0] node35928;
	wire [4-1:0] node35931;
	wire [4-1:0] node35934;
	wire [4-1:0] node35935;
	wire [4-1:0] node35938;
	wire [4-1:0] node35941;
	wire [4-1:0] node35942;
	wire [4-1:0] node35943;
	wire [4-1:0] node35946;
	wire [4-1:0] node35949;
	wire [4-1:0] node35950;
	wire [4-1:0] node35954;
	wire [4-1:0] node35955;
	wire [4-1:0] node35956;
	wire [4-1:0] node35958;
	wire [4-1:0] node35961;
	wire [4-1:0] node35963;
	wire [4-1:0] node35966;
	wire [4-1:0] node35967;
	wire [4-1:0] node35969;
	wire [4-1:0] node35972;
	wire [4-1:0] node35974;
	wire [4-1:0] node35977;
	wire [4-1:0] node35978;
	wire [4-1:0] node35979;
	wire [4-1:0] node35980;
	wire [4-1:0] node35981;
	wire [4-1:0] node35982;
	wire [4-1:0] node35985;
	wire [4-1:0] node35988;
	wire [4-1:0] node35990;
	wire [4-1:0] node35993;
	wire [4-1:0] node35994;
	wire [4-1:0] node35995;
	wire [4-1:0] node35998;
	wire [4-1:0] node36001;
	wire [4-1:0] node36002;
	wire [4-1:0] node36005;
	wire [4-1:0] node36008;
	wire [4-1:0] node36009;
	wire [4-1:0] node36010;
	wire [4-1:0] node36012;
	wire [4-1:0] node36015;
	wire [4-1:0] node36017;
	wire [4-1:0] node36020;
	wire [4-1:0] node36021;
	wire [4-1:0] node36023;
	wire [4-1:0] node36026;
	wire [4-1:0] node36028;
	wire [4-1:0] node36031;
	wire [4-1:0] node36032;
	wire [4-1:0] node36033;
	wire [4-1:0] node36034;
	wire [4-1:0] node36035;
	wire [4-1:0] node36038;
	wire [4-1:0] node36041;
	wire [4-1:0] node36042;
	wire [4-1:0] node36045;
	wire [4-1:0] node36048;
	wire [4-1:0] node36049;
	wire [4-1:0] node36050;
	wire [4-1:0] node36053;
	wire [4-1:0] node36056;
	wire [4-1:0] node36057;
	wire [4-1:0] node36060;
	wire [4-1:0] node36063;
	wire [4-1:0] node36064;
	wire [4-1:0] node36065;
	wire [4-1:0] node36067;
	wire [4-1:0] node36070;
	wire [4-1:0] node36072;
	wire [4-1:0] node36075;
	wire [4-1:0] node36076;
	wire [4-1:0] node36078;
	wire [4-1:0] node36081;
	wire [4-1:0] node36083;
	wire [4-1:0] node36086;
	wire [4-1:0] node36087;
	wire [4-1:0] node36088;
	wire [4-1:0] node36089;
	wire [4-1:0] node36090;
	wire [4-1:0] node36091;
	wire [4-1:0] node36092;
	wire [4-1:0] node36093;
	wire [4-1:0] node36096;
	wire [4-1:0] node36099;
	wire [4-1:0] node36100;
	wire [4-1:0] node36103;
	wire [4-1:0] node36106;
	wire [4-1:0] node36107;
	wire [4-1:0] node36108;
	wire [4-1:0] node36111;
	wire [4-1:0] node36114;
	wire [4-1:0] node36115;
	wire [4-1:0] node36119;
	wire [4-1:0] node36120;
	wire [4-1:0] node36121;
	wire [4-1:0] node36123;
	wire [4-1:0] node36126;
	wire [4-1:0] node36128;
	wire [4-1:0] node36131;
	wire [4-1:0] node36132;
	wire [4-1:0] node36134;
	wire [4-1:0] node36137;
	wire [4-1:0] node36139;
	wire [4-1:0] node36142;
	wire [4-1:0] node36143;
	wire [4-1:0] node36144;
	wire [4-1:0] node36145;
	wire [4-1:0] node36146;
	wire [4-1:0] node36149;
	wire [4-1:0] node36152;
	wire [4-1:0] node36153;
	wire [4-1:0] node36156;
	wire [4-1:0] node36159;
	wire [4-1:0] node36160;
	wire [4-1:0] node36161;
	wire [4-1:0] node36164;
	wire [4-1:0] node36167;
	wire [4-1:0] node36168;
	wire [4-1:0] node36171;
	wire [4-1:0] node36174;
	wire [4-1:0] node36175;
	wire [4-1:0] node36176;
	wire [4-1:0] node36177;
	wire [4-1:0] node36180;
	wire [4-1:0] node36183;
	wire [4-1:0] node36184;
	wire [4-1:0] node36187;
	wire [4-1:0] node36190;
	wire [4-1:0] node36191;
	wire [4-1:0] node36192;
	wire [4-1:0] node36195;
	wire [4-1:0] node36198;
	wire [4-1:0] node36199;
	wire [4-1:0] node36202;
	wire [4-1:0] node36205;
	wire [4-1:0] node36206;
	wire [4-1:0] node36207;
	wire [4-1:0] node36208;
	wire [4-1:0] node36209;
	wire [4-1:0] node36210;
	wire [4-1:0] node36213;
	wire [4-1:0] node36216;
	wire [4-1:0] node36217;
	wire [4-1:0] node36220;
	wire [4-1:0] node36223;
	wire [4-1:0] node36224;
	wire [4-1:0] node36225;
	wire [4-1:0] node36228;
	wire [4-1:0] node36231;
	wire [4-1:0] node36232;
	wire [4-1:0] node36235;
	wire [4-1:0] node36238;
	wire [4-1:0] node36239;
	wire [4-1:0] node36240;
	wire [4-1:0] node36243;
	wire [4-1:0] node36246;
	wire [4-1:0] node36247;
	wire [4-1:0] node36248;
	wire [4-1:0] node36251;
	wire [4-1:0] node36254;
	wire [4-1:0] node36255;
	wire [4-1:0] node36258;
	wire [4-1:0] node36261;
	wire [4-1:0] node36262;
	wire [4-1:0] node36263;
	wire [4-1:0] node36264;
	wire [4-1:0] node36265;
	wire [4-1:0] node36268;
	wire [4-1:0] node36271;
	wire [4-1:0] node36272;
	wire [4-1:0] node36276;
	wire [4-1:0] node36277;
	wire [4-1:0] node36279;
	wire [4-1:0] node36282;
	wire [4-1:0] node36283;
	wire [4-1:0] node36286;
	wire [4-1:0] node36289;
	wire [4-1:0] node36290;
	wire [4-1:0] node36291;
	wire [4-1:0] node36293;
	wire [4-1:0] node36296;
	wire [4-1:0] node36298;
	wire [4-1:0] node36301;
	wire [4-1:0] node36302;
	wire [4-1:0] node36304;
	wire [4-1:0] node36307;
	wire [4-1:0] node36309;
	wire [4-1:0] node36312;
	wire [4-1:0] node36313;
	wire [4-1:0] node36314;
	wire [4-1:0] node36315;
	wire [4-1:0] node36316;
	wire [4-1:0] node36317;
	wire [4-1:0] node36318;
	wire [4-1:0] node36321;
	wire [4-1:0] node36324;
	wire [4-1:0] node36325;
	wire [4-1:0] node36328;
	wire [4-1:0] node36331;
	wire [4-1:0] node36332;
	wire [4-1:0] node36333;
	wire [4-1:0] node36336;
	wire [4-1:0] node36339;
	wire [4-1:0] node36340;
	wire [4-1:0] node36343;
	wire [4-1:0] node36346;
	wire [4-1:0] node36347;
	wire [4-1:0] node36348;
	wire [4-1:0] node36349;
	wire [4-1:0] node36352;
	wire [4-1:0] node36355;
	wire [4-1:0] node36356;
	wire [4-1:0] node36360;
	wire [4-1:0] node36361;
	wire [4-1:0] node36362;
	wire [4-1:0] node36365;
	wire [4-1:0] node36368;
	wire [4-1:0] node36369;
	wire [4-1:0] node36372;
	wire [4-1:0] node36375;
	wire [4-1:0] node36376;
	wire [4-1:0] node36377;
	wire [4-1:0] node36378;
	wire [4-1:0] node36379;
	wire [4-1:0] node36382;
	wire [4-1:0] node36385;
	wire [4-1:0] node36386;
	wire [4-1:0] node36389;
	wire [4-1:0] node36392;
	wire [4-1:0] node36393;
	wire [4-1:0] node36394;
	wire [4-1:0] node36397;
	wire [4-1:0] node36400;
	wire [4-1:0] node36401;
	wire [4-1:0] node36404;
	wire [4-1:0] node36407;
	wire [4-1:0] node36408;
	wire [4-1:0] node36409;
	wire [4-1:0] node36410;
	wire [4-1:0] node36413;
	wire [4-1:0] node36416;
	wire [4-1:0] node36418;
	wire [4-1:0] node36421;
	wire [4-1:0] node36422;
	wire [4-1:0] node36423;
	wire [4-1:0] node36427;
	wire [4-1:0] node36428;
	wire [4-1:0] node36431;
	wire [4-1:0] node36434;
	wire [4-1:0] node36435;
	wire [4-1:0] node36436;
	wire [4-1:0] node36437;
	wire [4-1:0] node36438;
	wire [4-1:0] node36439;
	wire [4-1:0] node36443;
	wire [4-1:0] node36444;
	wire [4-1:0] node36448;
	wire [4-1:0] node36449;
	wire [4-1:0] node36450;
	wire [4-1:0] node36454;
	wire [4-1:0] node36455;
	wire [4-1:0] node36459;
	wire [4-1:0] node36460;
	wire [4-1:0] node36461;
	wire [4-1:0] node36462;
	wire [4-1:0] node36465;
	wire [4-1:0] node36468;
	wire [4-1:0] node36469;
	wire [4-1:0] node36472;
	wire [4-1:0] node36475;
	wire [4-1:0] node36476;
	wire [4-1:0] node36477;
	wire [4-1:0] node36480;
	wire [4-1:0] node36483;
	wire [4-1:0] node36484;
	wire [4-1:0] node36487;
	wire [4-1:0] node36490;
	wire [4-1:0] node36491;
	wire [4-1:0] node36492;
	wire [4-1:0] node36493;
	wire [4-1:0] node36494;
	wire [4-1:0] node36498;
	wire [4-1:0] node36499;
	wire [4-1:0] node36503;
	wire [4-1:0] node36504;
	wire [4-1:0] node36505;
	wire [4-1:0] node36509;
	wire [4-1:0] node36510;
	wire [4-1:0] node36514;
	wire [4-1:0] node36515;
	wire [4-1:0] node36516;
	wire [4-1:0] node36517;
	wire [4-1:0] node36520;
	wire [4-1:0] node36523;
	wire [4-1:0] node36524;
	wire [4-1:0] node36527;
	wire [4-1:0] node36530;
	wire [4-1:0] node36531;
	wire [4-1:0] node36532;
	wire [4-1:0] node36535;
	wire [4-1:0] node36538;
	wire [4-1:0] node36539;
	wire [4-1:0] node36542;
	wire [4-1:0] node36545;
	wire [4-1:0] node36546;
	wire [4-1:0] node36547;
	wire [4-1:0] node36548;
	wire [4-1:0] node36549;
	wire [4-1:0] node36550;
	wire [4-1:0] node36551;
	wire [4-1:0] node36552;
	wire [4-1:0] node36553;
	wire [4-1:0] node36557;
	wire [4-1:0] node36558;
	wire [4-1:0] node36561;
	wire [4-1:0] node36564;
	wire [4-1:0] node36565;
	wire [4-1:0] node36566;
	wire [4-1:0] node36569;
	wire [4-1:0] node36572;
	wire [4-1:0] node36574;
	wire [4-1:0] node36577;
	wire [4-1:0] node36578;
	wire [4-1:0] node36579;
	wire [4-1:0] node36581;
	wire [4-1:0] node36584;
	wire [4-1:0] node36586;
	wire [4-1:0] node36589;
	wire [4-1:0] node36590;
	wire [4-1:0] node36592;
	wire [4-1:0] node36595;
	wire [4-1:0] node36597;
	wire [4-1:0] node36600;
	wire [4-1:0] node36601;
	wire [4-1:0] node36602;
	wire [4-1:0] node36603;
	wire [4-1:0] node36604;
	wire [4-1:0] node36607;
	wire [4-1:0] node36610;
	wire [4-1:0] node36611;
	wire [4-1:0] node36614;
	wire [4-1:0] node36617;
	wire [4-1:0] node36618;
	wire [4-1:0] node36620;
	wire [4-1:0] node36623;
	wire [4-1:0] node36624;
	wire [4-1:0] node36627;
	wire [4-1:0] node36630;
	wire [4-1:0] node36631;
	wire [4-1:0] node36632;
	wire [4-1:0] node36634;
	wire [4-1:0] node36637;
	wire [4-1:0] node36639;
	wire [4-1:0] node36642;
	wire [4-1:0] node36643;
	wire [4-1:0] node36645;
	wire [4-1:0] node36648;
	wire [4-1:0] node36650;
	wire [4-1:0] node36653;
	wire [4-1:0] node36654;
	wire [4-1:0] node36655;
	wire [4-1:0] node36656;
	wire [4-1:0] node36657;
	wire [4-1:0] node36658;
	wire [4-1:0] node36661;
	wire [4-1:0] node36664;
	wire [4-1:0] node36665;
	wire [4-1:0] node36668;
	wire [4-1:0] node36671;
	wire [4-1:0] node36672;
	wire [4-1:0] node36674;
	wire [4-1:0] node36677;
	wire [4-1:0] node36679;
	wire [4-1:0] node36682;
	wire [4-1:0] node36683;
	wire [4-1:0] node36684;
	wire [4-1:0] node36685;
	wire [4-1:0] node36688;
	wire [4-1:0] node36691;
	wire [4-1:0] node36692;
	wire [4-1:0] node36695;
	wire [4-1:0] node36698;
	wire [4-1:0] node36699;
	wire [4-1:0] node36700;
	wire [4-1:0] node36703;
	wire [4-1:0] node36706;
	wire [4-1:0] node36707;
	wire [4-1:0] node36711;
	wire [4-1:0] node36712;
	wire [4-1:0] node36713;
	wire [4-1:0] node36714;
	wire [4-1:0] node36715;
	wire [4-1:0] node36718;
	wire [4-1:0] node36721;
	wire [4-1:0] node36722;
	wire [4-1:0] node36725;
	wire [4-1:0] node36728;
	wire [4-1:0] node36729;
	wire [4-1:0] node36730;
	wire [4-1:0] node36733;
	wire [4-1:0] node36736;
	wire [4-1:0] node36737;
	wire [4-1:0] node36740;
	wire [4-1:0] node36743;
	wire [4-1:0] node36744;
	wire [4-1:0] node36745;
	wire [4-1:0] node36748;
	wire [4-1:0] node36751;
	wire [4-1:0] node36752;
	wire [4-1:0] node36753;
	wire [4-1:0] node36756;
	wire [4-1:0] node36759;
	wire [4-1:0] node36760;
	wire [4-1:0] node36763;
	wire [4-1:0] node36766;
	wire [4-1:0] node36767;
	wire [4-1:0] node36768;
	wire [4-1:0] node36769;
	wire [4-1:0] node36770;
	wire [4-1:0] node36771;
	wire [4-1:0] node36772;
	wire [4-1:0] node36775;
	wire [4-1:0] node36778;
	wire [4-1:0] node36780;
	wire [4-1:0] node36783;
	wire [4-1:0] node36784;
	wire [4-1:0] node36785;
	wire [4-1:0] node36788;
	wire [4-1:0] node36791;
	wire [4-1:0] node36792;
	wire [4-1:0] node36795;
	wire [4-1:0] node36798;
	wire [4-1:0] node36799;
	wire [4-1:0] node36800;
	wire [4-1:0] node36802;
	wire [4-1:0] node36805;
	wire [4-1:0] node36807;
	wire [4-1:0] node36810;
	wire [4-1:0] node36811;
	wire [4-1:0] node36813;
	wire [4-1:0] node36816;
	wire [4-1:0] node36818;
	wire [4-1:0] node36821;
	wire [4-1:0] node36822;
	wire [4-1:0] node36823;
	wire [4-1:0] node36824;
	wire [4-1:0] node36825;
	wire [4-1:0] node36828;
	wire [4-1:0] node36831;
	wire [4-1:0] node36832;
	wire [4-1:0] node36835;
	wire [4-1:0] node36838;
	wire [4-1:0] node36839;
	wire [4-1:0] node36841;
	wire [4-1:0] node36844;
	wire [4-1:0] node36845;
	wire [4-1:0] node36848;
	wire [4-1:0] node36851;
	wire [4-1:0] node36852;
	wire [4-1:0] node36853;
	wire [4-1:0] node36854;
	wire [4-1:0] node36857;
	wire [4-1:0] node36860;
	wire [4-1:0] node36861;
	wire [4-1:0] node36864;
	wire [4-1:0] node36867;
	wire [4-1:0] node36868;
	wire [4-1:0] node36871;
	wire [4-1:0] node36874;
	wire [4-1:0] node36875;
	wire [4-1:0] node36876;
	wire [4-1:0] node36877;
	wire [4-1:0] node36878;
	wire [4-1:0] node36879;
	wire [4-1:0] node36883;
	wire [4-1:0] node36884;
	wire [4-1:0] node36887;
	wire [4-1:0] node36890;
	wire [4-1:0] node36891;
	wire [4-1:0] node36892;
	wire [4-1:0] node36896;
	wire [4-1:0] node36897;
	wire [4-1:0] node36901;
	wire [4-1:0] node36902;
	wire [4-1:0] node36903;
	wire [4-1:0] node36904;
	wire [4-1:0] node36908;
	wire [4-1:0] node36909;
	wire [4-1:0] node36913;
	wire [4-1:0] node36914;
	wire [4-1:0] node36915;
	wire [4-1:0] node36919;
	wire [4-1:0] node36920;
	wire [4-1:0] node36924;
	wire [4-1:0] node36925;
	wire [4-1:0] node36926;
	wire [4-1:0] node36927;
	wire [4-1:0] node36928;
	wire [4-1:0] node36932;
	wire [4-1:0] node36933;
	wire [4-1:0] node36937;
	wire [4-1:0] node36938;
	wire [4-1:0] node36940;
	wire [4-1:0] node36943;
	wire [4-1:0] node36945;
	wire [4-1:0] node36948;
	wire [4-1:0] node36949;
	wire [4-1:0] node36950;
	wire [4-1:0] node36951;
	wire [4-1:0] node36954;
	wire [4-1:0] node36957;
	wire [4-1:0] node36958;
	wire [4-1:0] node36961;
	wire [4-1:0] node36964;
	wire [4-1:0] node36965;
	wire [4-1:0] node36966;
	wire [4-1:0] node36969;
	wire [4-1:0] node36972;
	wire [4-1:0] node36973;
	wire [4-1:0] node36976;
	wire [4-1:0] node36979;
	wire [4-1:0] node36980;
	wire [4-1:0] node36981;
	wire [4-1:0] node36982;
	wire [4-1:0] node36983;
	wire [4-1:0] node36984;
	wire [4-1:0] node36985;
	wire [4-1:0] node36986;
	wire [4-1:0] node36989;
	wire [4-1:0] node36992;
	wire [4-1:0] node36993;
	wire [4-1:0] node36996;
	wire [4-1:0] node36999;
	wire [4-1:0] node37000;
	wire [4-1:0] node37001;
	wire [4-1:0] node37004;
	wire [4-1:0] node37007;
	wire [4-1:0] node37008;
	wire [4-1:0] node37011;
	wire [4-1:0] node37014;
	wire [4-1:0] node37015;
	wire [4-1:0] node37016;
	wire [4-1:0] node37020;
	wire [4-1:0] node37021;
	wire [4-1:0] node37023;
	wire [4-1:0] node37026;
	wire [4-1:0] node37028;
	wire [4-1:0] node37031;
	wire [4-1:0] node37032;
	wire [4-1:0] node37033;
	wire [4-1:0] node37034;
	wire [4-1:0] node37035;
	wire [4-1:0] node37038;
	wire [4-1:0] node37041;
	wire [4-1:0] node37042;
	wire [4-1:0] node37045;
	wire [4-1:0] node37048;
	wire [4-1:0] node37049;
	wire [4-1:0] node37050;
	wire [4-1:0] node37053;
	wire [4-1:0] node37056;
	wire [4-1:0] node37057;
	wire [4-1:0] node37060;
	wire [4-1:0] node37063;
	wire [4-1:0] node37064;
	wire [4-1:0] node37065;
	wire [4-1:0] node37066;
	wire [4-1:0] node37069;
	wire [4-1:0] node37072;
	wire [4-1:0] node37074;
	wire [4-1:0] node37077;
	wire [4-1:0] node37078;
	wire [4-1:0] node37079;
	wire [4-1:0] node37082;
	wire [4-1:0] node37085;
	wire [4-1:0] node37086;
	wire [4-1:0] node37089;
	wire [4-1:0] node37092;
	wire [4-1:0] node37093;
	wire [4-1:0] node37094;
	wire [4-1:0] node37095;
	wire [4-1:0] node37096;
	wire [4-1:0] node37097;
	wire [4-1:0] node37100;
	wire [4-1:0] node37103;
	wire [4-1:0] node37104;
	wire [4-1:0] node37107;
	wire [4-1:0] node37110;
	wire [4-1:0] node37111;
	wire [4-1:0] node37112;
	wire [4-1:0] node37115;
	wire [4-1:0] node37118;
	wire [4-1:0] node37119;
	wire [4-1:0] node37122;
	wire [4-1:0] node37125;
	wire [4-1:0] node37126;
	wire [4-1:0] node37127;
	wire [4-1:0] node37128;
	wire [4-1:0] node37131;
	wire [4-1:0] node37134;
	wire [4-1:0] node37135;
	wire [4-1:0] node37138;
	wire [4-1:0] node37141;
	wire [4-1:0] node37142;
	wire [4-1:0] node37143;
	wire [4-1:0] node37146;
	wire [4-1:0] node37149;
	wire [4-1:0] node37150;
	wire [4-1:0] node37153;
	wire [4-1:0] node37156;
	wire [4-1:0] node37157;
	wire [4-1:0] node37158;
	wire [4-1:0] node37159;
	wire [4-1:0] node37161;
	wire [4-1:0] node37164;
	wire [4-1:0] node37165;
	wire [4-1:0] node37168;
	wire [4-1:0] node37171;
	wire [4-1:0] node37172;
	wire [4-1:0] node37173;
	wire [4-1:0] node37176;
	wire [4-1:0] node37179;
	wire [4-1:0] node37180;
	wire [4-1:0] node37183;
	wire [4-1:0] node37186;
	wire [4-1:0] node37187;
	wire [4-1:0] node37188;
	wire [4-1:0] node37189;
	wire [4-1:0] node37192;
	wire [4-1:0] node37195;
	wire [4-1:0] node37196;
	wire [4-1:0] node37199;
	wire [4-1:0] node37202;
	wire [4-1:0] node37203;
	wire [4-1:0] node37206;
	wire [4-1:0] node37209;
	wire [4-1:0] node37210;
	wire [4-1:0] node37211;
	wire [4-1:0] node37212;
	wire [4-1:0] node37213;
	wire [4-1:0] node37214;
	wire [4-1:0] node37215;
	wire [4-1:0] node37218;
	wire [4-1:0] node37221;
	wire [4-1:0] node37222;
	wire [4-1:0] node37226;
	wire [4-1:0] node37227;
	wire [4-1:0] node37228;
	wire [4-1:0] node37231;
	wire [4-1:0] node37234;
	wire [4-1:0] node37235;
	wire [4-1:0] node37238;
	wire [4-1:0] node37241;
	wire [4-1:0] node37242;
	wire [4-1:0] node37243;
	wire [4-1:0] node37244;
	wire [4-1:0] node37247;
	wire [4-1:0] node37250;
	wire [4-1:0] node37251;
	wire [4-1:0] node37255;
	wire [4-1:0] node37256;
	wire [4-1:0] node37257;
	wire [4-1:0] node37260;
	wire [4-1:0] node37263;
	wire [4-1:0] node37264;
	wire [4-1:0] node37267;
	wire [4-1:0] node37270;
	wire [4-1:0] node37271;
	wire [4-1:0] node37272;
	wire [4-1:0] node37273;
	wire [4-1:0] node37274;
	wire [4-1:0] node37277;
	wire [4-1:0] node37280;
	wire [4-1:0] node37281;
	wire [4-1:0] node37285;
	wire [4-1:0] node37286;
	wire [4-1:0] node37287;
	wire [4-1:0] node37290;
	wire [4-1:0] node37293;
	wire [4-1:0] node37295;
	wire [4-1:0] node37298;
	wire [4-1:0] node37299;
	wire [4-1:0] node37300;
	wire [4-1:0] node37301;
	wire [4-1:0] node37304;
	wire [4-1:0] node37307;
	wire [4-1:0] node37308;
	wire [4-1:0] node37311;
	wire [4-1:0] node37314;
	wire [4-1:0] node37315;
	wire [4-1:0] node37316;
	wire [4-1:0] node37319;
	wire [4-1:0] node37322;
	wire [4-1:0] node37323;
	wire [4-1:0] node37326;
	wire [4-1:0] node37329;
	wire [4-1:0] node37330;
	wire [4-1:0] node37331;
	wire [4-1:0] node37332;
	wire [4-1:0] node37333;
	wire [4-1:0] node37334;
	wire [4-1:0] node37337;
	wire [4-1:0] node37340;
	wire [4-1:0] node37341;
	wire [4-1:0] node37345;
	wire [4-1:0] node37346;
	wire [4-1:0] node37347;
	wire [4-1:0] node37351;
	wire [4-1:0] node37352;
	wire [4-1:0] node37355;
	wire [4-1:0] node37358;
	wire [4-1:0] node37359;
	wire [4-1:0] node37360;
	wire [4-1:0] node37361;
	wire [4-1:0] node37364;
	wire [4-1:0] node37367;
	wire [4-1:0] node37368;
	wire [4-1:0] node37371;
	wire [4-1:0] node37374;
	wire [4-1:0] node37375;
	wire [4-1:0] node37376;
	wire [4-1:0] node37379;
	wire [4-1:0] node37382;
	wire [4-1:0] node37383;
	wire [4-1:0] node37386;
	wire [4-1:0] node37389;
	wire [4-1:0] node37390;
	wire [4-1:0] node37391;
	wire [4-1:0] node37392;
	wire [4-1:0] node37393;
	wire [4-1:0] node37396;
	wire [4-1:0] node37399;
	wire [4-1:0] node37400;
	wire [4-1:0] node37403;
	wire [4-1:0] node37406;
	wire [4-1:0] node37407;
	wire [4-1:0] node37408;
	wire [4-1:0] node37411;
	wire [4-1:0] node37414;
	wire [4-1:0] node37415;
	wire [4-1:0] node37418;
	wire [4-1:0] node37421;
	wire [4-1:0] node37422;
	wire [4-1:0] node37423;
	wire [4-1:0] node37426;
	wire [4-1:0] node37429;
	wire [4-1:0] node37430;
	wire [4-1:0] node37433;
	wire [4-1:0] node37436;
	wire [4-1:0] node37437;
	wire [4-1:0] node37438;
	wire [4-1:0] node37439;
	wire [4-1:0] node37440;
	wire [4-1:0] node37441;
	wire [4-1:0] node37442;
	wire [4-1:0] node37443;
	wire [4-1:0] node37444;
	wire [4-1:0] node37445;
	wire [4-1:0] node37448;
	wire [4-1:0] node37451;
	wire [4-1:0] node37452;
	wire [4-1:0] node37455;
	wire [4-1:0] node37458;
	wire [4-1:0] node37459;
	wire [4-1:0] node37462;
	wire [4-1:0] node37465;
	wire [4-1:0] node37466;
	wire [4-1:0] node37467;
	wire [4-1:0] node37468;
	wire [4-1:0] node37471;
	wire [4-1:0] node37474;
	wire [4-1:0] node37475;
	wire [4-1:0] node37478;
	wire [4-1:0] node37481;
	wire [4-1:0] node37482;
	wire [4-1:0] node37483;
	wire [4-1:0] node37486;
	wire [4-1:0] node37489;
	wire [4-1:0] node37491;
	wire [4-1:0] node37494;
	wire [4-1:0] node37495;
	wire [4-1:0] node37496;
	wire [4-1:0] node37497;
	wire [4-1:0] node37498;
	wire [4-1:0] node37501;
	wire [4-1:0] node37504;
	wire [4-1:0] node37505;
	wire [4-1:0] node37508;
	wire [4-1:0] node37511;
	wire [4-1:0] node37512;
	wire [4-1:0] node37515;
	wire [4-1:0] node37518;
	wire [4-1:0] node37519;
	wire [4-1:0] node37520;
	wire [4-1:0] node37521;
	wire [4-1:0] node37524;
	wire [4-1:0] node37527;
	wire [4-1:0] node37528;
	wire [4-1:0] node37532;
	wire [4-1:0] node37533;
	wire [4-1:0] node37535;
	wire [4-1:0] node37538;
	wire [4-1:0] node37539;
	wire [4-1:0] node37542;
	wire [4-1:0] node37545;
	wire [4-1:0] node37546;
	wire [4-1:0] node37547;
	wire [4-1:0] node37548;
	wire [4-1:0] node37549;
	wire [4-1:0] node37550;
	wire [4-1:0] node37554;
	wire [4-1:0] node37555;
	wire [4-1:0] node37558;
	wire [4-1:0] node37561;
	wire [4-1:0] node37562;
	wire [4-1:0] node37563;
	wire [4-1:0] node37566;
	wire [4-1:0] node37569;
	wire [4-1:0] node37570;
	wire [4-1:0] node37573;
	wire [4-1:0] node37576;
	wire [4-1:0] node37577;
	wire [4-1:0] node37578;
	wire [4-1:0] node37579;
	wire [4-1:0] node37582;
	wire [4-1:0] node37585;
	wire [4-1:0] node37586;
	wire [4-1:0] node37589;
	wire [4-1:0] node37592;
	wire [4-1:0] node37593;
	wire [4-1:0] node37594;
	wire [4-1:0] node37597;
	wire [4-1:0] node37600;
	wire [4-1:0] node37601;
	wire [4-1:0] node37604;
	wire [4-1:0] node37607;
	wire [4-1:0] node37608;
	wire [4-1:0] node37609;
	wire [4-1:0] node37610;
	wire [4-1:0] node37611;
	wire [4-1:0] node37614;
	wire [4-1:0] node37617;
	wire [4-1:0] node37618;
	wire [4-1:0] node37621;
	wire [4-1:0] node37624;
	wire [4-1:0] node37625;
	wire [4-1:0] node37626;
	wire [4-1:0] node37629;
	wire [4-1:0] node37632;
	wire [4-1:0] node37633;
	wire [4-1:0] node37636;
	wire [4-1:0] node37639;
	wire [4-1:0] node37640;
	wire [4-1:0] node37641;
	wire [4-1:0] node37642;
	wire [4-1:0] node37645;
	wire [4-1:0] node37648;
	wire [4-1:0] node37649;
	wire [4-1:0] node37652;
	wire [4-1:0] node37655;
	wire [4-1:0] node37656;
	wire [4-1:0] node37657;
	wire [4-1:0] node37660;
	wire [4-1:0] node37663;
	wire [4-1:0] node37664;
	wire [4-1:0] node37668;
	wire [4-1:0] node37669;
	wire [4-1:0] node37670;
	wire [4-1:0] node37671;
	wire [4-1:0] node37672;
	wire [4-1:0] node37673;
	wire [4-1:0] node37674;
	wire [4-1:0] node37677;
	wire [4-1:0] node37680;
	wire [4-1:0] node37681;
	wire [4-1:0] node37685;
	wire [4-1:0] node37686;
	wire [4-1:0] node37687;
	wire [4-1:0] node37690;
	wire [4-1:0] node37693;
	wire [4-1:0] node37695;
	wire [4-1:0] node37698;
	wire [4-1:0] node37699;
	wire [4-1:0] node37700;
	wire [4-1:0] node37701;
	wire [4-1:0] node37704;
	wire [4-1:0] node37707;
	wire [4-1:0] node37708;
	wire [4-1:0] node37711;
	wire [4-1:0] node37714;
	wire [4-1:0] node37715;
	wire [4-1:0] node37716;
	wire [4-1:0] node37719;
	wire [4-1:0] node37722;
	wire [4-1:0] node37723;
	wire [4-1:0] node37726;
	wire [4-1:0] node37729;
	wire [4-1:0] node37730;
	wire [4-1:0] node37731;
	wire [4-1:0] node37732;
	wire [4-1:0] node37733;
	wire [4-1:0] node37736;
	wire [4-1:0] node37739;
	wire [4-1:0] node37740;
	wire [4-1:0] node37743;
	wire [4-1:0] node37746;
	wire [4-1:0] node37747;
	wire [4-1:0] node37748;
	wire [4-1:0] node37751;
	wire [4-1:0] node37754;
	wire [4-1:0] node37755;
	wire [4-1:0] node37759;
	wire [4-1:0] node37760;
	wire [4-1:0] node37761;
	wire [4-1:0] node37762;
	wire [4-1:0] node37766;
	wire [4-1:0] node37767;
	wire [4-1:0] node37770;
	wire [4-1:0] node37773;
	wire [4-1:0] node37774;
	wire [4-1:0] node37777;
	wire [4-1:0] node37780;
	wire [4-1:0] node37781;
	wire [4-1:0] node37782;
	wire [4-1:0] node37783;
	wire [4-1:0] node37784;
	wire [4-1:0] node37785;
	wire [4-1:0] node37788;
	wire [4-1:0] node37791;
	wire [4-1:0] node37792;
	wire [4-1:0] node37795;
	wire [4-1:0] node37798;
	wire [4-1:0] node37799;
	wire [4-1:0] node37800;
	wire [4-1:0] node37804;
	wire [4-1:0] node37805;
	wire [4-1:0] node37808;
	wire [4-1:0] node37811;
	wire [4-1:0] node37812;
	wire [4-1:0] node37813;
	wire [4-1:0] node37814;
	wire [4-1:0] node37818;
	wire [4-1:0] node37819;
	wire [4-1:0] node37823;
	wire [4-1:0] node37824;
	wire [4-1:0] node37825;
	wire [4-1:0] node37829;
	wire [4-1:0] node37830;
	wire [4-1:0] node37834;
	wire [4-1:0] node37835;
	wire [4-1:0] node37836;
	wire [4-1:0] node37837;
	wire [4-1:0] node37838;
	wire [4-1:0] node37841;
	wire [4-1:0] node37844;
	wire [4-1:0] node37845;
	wire [4-1:0] node37848;
	wire [4-1:0] node37851;
	wire [4-1:0] node37852;
	wire [4-1:0] node37853;
	wire [4-1:0] node37856;
	wire [4-1:0] node37859;
	wire [4-1:0] node37860;
	wire [4-1:0] node37863;
	wire [4-1:0] node37866;
	wire [4-1:0] node37867;
	wire [4-1:0] node37868;
	wire [4-1:0] node37869;
	wire [4-1:0] node37873;
	wire [4-1:0] node37874;
	wire [4-1:0] node37878;
	wire [4-1:0] node37879;
	wire [4-1:0] node37880;
	wire [4-1:0] node37884;
	wire [4-1:0] node37885;
	wire [4-1:0] node37889;
	wire [4-1:0] node37890;
	wire [4-1:0] node37891;
	wire [4-1:0] node37892;
	wire [4-1:0] node37893;
	wire [4-1:0] node37894;
	wire [4-1:0] node37895;
	wire [4-1:0] node37896;
	wire [4-1:0] node37899;
	wire [4-1:0] node37902;
	wire [4-1:0] node37903;
	wire [4-1:0] node37907;
	wire [4-1:0] node37908;
	wire [4-1:0] node37911;
	wire [4-1:0] node37912;
	wire [4-1:0] node37915;
	wire [4-1:0] node37918;
	wire [4-1:0] node37919;
	wire [4-1:0] node37920;
	wire [4-1:0] node37921;
	wire [4-1:0] node37924;
	wire [4-1:0] node37927;
	wire [4-1:0] node37928;
	wire [4-1:0] node37931;
	wire [4-1:0] node37934;
	wire [4-1:0] node37935;
	wire [4-1:0] node37936;
	wire [4-1:0] node37939;
	wire [4-1:0] node37942;
	wire [4-1:0] node37943;
	wire [4-1:0] node37947;
	wire [4-1:0] node37948;
	wire [4-1:0] node37949;
	wire [4-1:0] node37950;
	wire [4-1:0] node37951;
	wire [4-1:0] node37954;
	wire [4-1:0] node37957;
	wire [4-1:0] node37958;
	wire [4-1:0] node37961;
	wire [4-1:0] node37964;
	wire [4-1:0] node37965;
	wire [4-1:0] node37966;
	wire [4-1:0] node37970;
	wire [4-1:0] node37971;
	wire [4-1:0] node37975;
	wire [4-1:0] node37976;
	wire [4-1:0] node37977;
	wire [4-1:0] node37978;
	wire [4-1:0] node37982;
	wire [4-1:0] node37983;
	wire [4-1:0] node37987;
	wire [4-1:0] node37988;
	wire [4-1:0] node37989;
	wire [4-1:0] node37993;
	wire [4-1:0] node37994;
	wire [4-1:0] node37998;
	wire [4-1:0] node37999;
	wire [4-1:0] node38000;
	wire [4-1:0] node38001;
	wire [4-1:0] node38002;
	wire [4-1:0] node38003;
	wire [4-1:0] node38006;
	wire [4-1:0] node38009;
	wire [4-1:0] node38011;
	wire [4-1:0] node38014;
	wire [4-1:0] node38015;
	wire [4-1:0] node38016;
	wire [4-1:0] node38019;
	wire [4-1:0] node38022;
	wire [4-1:0] node38024;
	wire [4-1:0] node38027;
	wire [4-1:0] node38028;
	wire [4-1:0] node38029;
	wire [4-1:0] node38030;
	wire [4-1:0] node38034;
	wire [4-1:0] node38035;
	wire [4-1:0] node38039;
	wire [4-1:0] node38040;
	wire [4-1:0] node38041;
	wire [4-1:0] node38045;
	wire [4-1:0] node38046;
	wire [4-1:0] node38050;
	wire [4-1:0] node38051;
	wire [4-1:0] node38052;
	wire [4-1:0] node38053;
	wire [4-1:0] node38054;
	wire [4-1:0] node38057;
	wire [4-1:0] node38060;
	wire [4-1:0] node38061;
	wire [4-1:0] node38064;
	wire [4-1:0] node38067;
	wire [4-1:0] node38068;
	wire [4-1:0] node38069;
	wire [4-1:0] node38072;
	wire [4-1:0] node38075;
	wire [4-1:0] node38076;
	wire [4-1:0] node38079;
	wire [4-1:0] node38082;
	wire [4-1:0] node38083;
	wire [4-1:0] node38084;
	wire [4-1:0] node38085;
	wire [4-1:0] node38088;
	wire [4-1:0] node38091;
	wire [4-1:0] node38092;
	wire [4-1:0] node38095;
	wire [4-1:0] node38098;
	wire [4-1:0] node38099;
	wire [4-1:0] node38100;
	wire [4-1:0] node38103;
	wire [4-1:0] node38106;
	wire [4-1:0] node38107;
	wire [4-1:0] node38110;
	wire [4-1:0] node38113;
	wire [4-1:0] node38114;
	wire [4-1:0] node38115;
	wire [4-1:0] node38116;
	wire [4-1:0] node38117;
	wire [4-1:0] node38118;
	wire [4-1:0] node38119;
	wire [4-1:0] node38122;
	wire [4-1:0] node38125;
	wire [4-1:0] node38126;
	wire [4-1:0] node38129;
	wire [4-1:0] node38132;
	wire [4-1:0] node38133;
	wire [4-1:0] node38134;
	wire [4-1:0] node38137;
	wire [4-1:0] node38140;
	wire [4-1:0] node38141;
	wire [4-1:0] node38145;
	wire [4-1:0] node38146;
	wire [4-1:0] node38147;
	wire [4-1:0] node38148;
	wire [4-1:0] node38152;
	wire [4-1:0] node38153;
	wire [4-1:0] node38157;
	wire [4-1:0] node38158;
	wire [4-1:0] node38159;
	wire [4-1:0] node38163;
	wire [4-1:0] node38164;
	wire [4-1:0] node38168;
	wire [4-1:0] node38169;
	wire [4-1:0] node38170;
	wire [4-1:0] node38171;
	wire [4-1:0] node38172;
	wire [4-1:0] node38176;
	wire [4-1:0] node38177;
	wire [4-1:0] node38181;
	wire [4-1:0] node38182;
	wire [4-1:0] node38183;
	wire [4-1:0] node38186;
	wire [4-1:0] node38189;
	wire [4-1:0] node38190;
	wire [4-1:0] node38193;
	wire [4-1:0] node38196;
	wire [4-1:0] node38197;
	wire [4-1:0] node38198;
	wire [4-1:0] node38199;
	wire [4-1:0] node38203;
	wire [4-1:0] node38204;
	wire [4-1:0] node38208;
	wire [4-1:0] node38209;
	wire [4-1:0] node38210;
	wire [4-1:0] node38214;
	wire [4-1:0] node38216;
	wire [4-1:0] node38219;
	wire [4-1:0] node38220;
	wire [4-1:0] node38221;
	wire [4-1:0] node38222;
	wire [4-1:0] node38223;
	wire [4-1:0] node38224;
	wire [4-1:0] node38227;
	wire [4-1:0] node38230;
	wire [4-1:0] node38231;
	wire [4-1:0] node38234;
	wire [4-1:0] node38237;
	wire [4-1:0] node38238;
	wire [4-1:0] node38239;
	wire [4-1:0] node38242;
	wire [4-1:0] node38245;
	wire [4-1:0] node38246;
	wire [4-1:0] node38250;
	wire [4-1:0] node38251;
	wire [4-1:0] node38252;
	wire [4-1:0] node38253;
	wire [4-1:0] node38256;
	wire [4-1:0] node38259;
	wire [4-1:0] node38260;
	wire [4-1:0] node38263;
	wire [4-1:0] node38266;
	wire [4-1:0] node38267;
	wire [4-1:0] node38270;
	wire [4-1:0] node38273;
	wire [4-1:0] node38274;
	wire [4-1:0] node38275;
	wire [4-1:0] node38276;
	wire [4-1:0] node38277;
	wire [4-1:0] node38280;
	wire [4-1:0] node38283;
	wire [4-1:0] node38284;
	wire [4-1:0] node38288;
	wire [4-1:0] node38289;
	wire [4-1:0] node38290;
	wire [4-1:0] node38293;
	wire [4-1:0] node38296;
	wire [4-1:0] node38297;
	wire [4-1:0] node38300;
	wire [4-1:0] node38303;
	wire [4-1:0] node38304;
	wire [4-1:0] node38305;
	wire [4-1:0] node38306;
	wire [4-1:0] node38310;
	wire [4-1:0] node38311;
	wire [4-1:0] node38315;
	wire [4-1:0] node38316;
	wire [4-1:0] node38317;
	wire [4-1:0] node38321;
	wire [4-1:0] node38322;
	wire [4-1:0] node38326;
	wire [4-1:0] node38327;
	wire [4-1:0] node38328;
	wire [4-1:0] node38329;
	wire [4-1:0] node38330;
	wire [4-1:0] node38331;
	wire [4-1:0] node38332;
	wire [4-1:0] node38333;
	wire [4-1:0] node38334;
	wire [4-1:0] node38337;
	wire [4-1:0] node38340;
	wire [4-1:0] node38341;
	wire [4-1:0] node38344;
	wire [4-1:0] node38347;
	wire [4-1:0] node38348;
	wire [4-1:0] node38349;
	wire [4-1:0] node38353;
	wire [4-1:0] node38354;
	wire [4-1:0] node38357;
	wire [4-1:0] node38360;
	wire [4-1:0] node38361;
	wire [4-1:0] node38362;
	wire [4-1:0] node38363;
	wire [4-1:0] node38366;
	wire [4-1:0] node38369;
	wire [4-1:0] node38370;
	wire [4-1:0] node38373;
	wire [4-1:0] node38376;
	wire [4-1:0] node38377;
	wire [4-1:0] node38380;
	wire [4-1:0] node38383;
	wire [4-1:0] node38384;
	wire [4-1:0] node38385;
	wire [4-1:0] node38386;
	wire [4-1:0] node38387;
	wire [4-1:0] node38390;
	wire [4-1:0] node38393;
	wire [4-1:0] node38395;
	wire [4-1:0] node38398;
	wire [4-1:0] node38399;
	wire [4-1:0] node38400;
	wire [4-1:0] node38404;
	wire [4-1:0] node38405;
	wire [4-1:0] node38408;
	wire [4-1:0] node38411;
	wire [4-1:0] node38412;
	wire [4-1:0] node38413;
	wire [4-1:0] node38414;
	wire [4-1:0] node38417;
	wire [4-1:0] node38420;
	wire [4-1:0] node38421;
	wire [4-1:0] node38424;
	wire [4-1:0] node38427;
	wire [4-1:0] node38428;
	wire [4-1:0] node38431;
	wire [4-1:0] node38434;
	wire [4-1:0] node38435;
	wire [4-1:0] node38436;
	wire [4-1:0] node38437;
	wire [4-1:0] node38438;
	wire [4-1:0] node38439;
	wire [4-1:0] node38442;
	wire [4-1:0] node38445;
	wire [4-1:0] node38446;
	wire [4-1:0] node38449;
	wire [4-1:0] node38452;
	wire [4-1:0] node38453;
	wire [4-1:0] node38454;
	wire [4-1:0] node38457;
	wire [4-1:0] node38460;
	wire [4-1:0] node38461;
	wire [4-1:0] node38464;
	wire [4-1:0] node38467;
	wire [4-1:0] node38468;
	wire [4-1:0] node38469;
	wire [4-1:0] node38470;
	wire [4-1:0] node38474;
	wire [4-1:0] node38475;
	wire [4-1:0] node38479;
	wire [4-1:0] node38480;
	wire [4-1:0] node38481;
	wire [4-1:0] node38485;
	wire [4-1:0] node38486;
	wire [4-1:0] node38490;
	wire [4-1:0] node38491;
	wire [4-1:0] node38492;
	wire [4-1:0] node38493;
	wire [4-1:0] node38494;
	wire [4-1:0] node38497;
	wire [4-1:0] node38500;
	wire [4-1:0] node38502;
	wire [4-1:0] node38505;
	wire [4-1:0] node38506;
	wire [4-1:0] node38507;
	wire [4-1:0] node38510;
	wire [4-1:0] node38513;
	wire [4-1:0] node38514;
	wire [4-1:0] node38517;
	wire [4-1:0] node38520;
	wire [4-1:0] node38521;
	wire [4-1:0] node38522;
	wire [4-1:0] node38523;
	wire [4-1:0] node38526;
	wire [4-1:0] node38529;
	wire [4-1:0] node38530;
	wire [4-1:0] node38534;
	wire [4-1:0] node38535;
	wire [4-1:0] node38536;
	wire [4-1:0] node38539;
	wire [4-1:0] node38542;
	wire [4-1:0] node38543;
	wire [4-1:0] node38546;
	wire [4-1:0] node38549;
	wire [4-1:0] node38550;
	wire [4-1:0] node38551;
	wire [4-1:0] node38552;
	wire [4-1:0] node38553;
	wire [4-1:0] node38554;
	wire [4-1:0] node38556;
	wire [4-1:0] node38559;
	wire [4-1:0] node38560;
	wire [4-1:0] node38563;
	wire [4-1:0] node38566;
	wire [4-1:0] node38567;
	wire [4-1:0] node38568;
	wire [4-1:0] node38571;
	wire [4-1:0] node38574;
	wire [4-1:0] node38575;
	wire [4-1:0] node38579;
	wire [4-1:0] node38580;
	wire [4-1:0] node38581;
	wire [4-1:0] node38582;
	wire [4-1:0] node38586;
	wire [4-1:0] node38587;
	wire [4-1:0] node38591;
	wire [4-1:0] node38592;
	wire [4-1:0] node38593;
	wire [4-1:0] node38597;
	wire [4-1:0] node38598;
	wire [4-1:0] node38602;
	wire [4-1:0] node38603;
	wire [4-1:0] node38604;
	wire [4-1:0] node38605;
	wire [4-1:0] node38606;
	wire [4-1:0] node38609;
	wire [4-1:0] node38612;
	wire [4-1:0] node38613;
	wire [4-1:0] node38616;
	wire [4-1:0] node38619;
	wire [4-1:0] node38620;
	wire [4-1:0] node38622;
	wire [4-1:0] node38625;
	wire [4-1:0] node38626;
	wire [4-1:0] node38630;
	wire [4-1:0] node38631;
	wire [4-1:0] node38632;
	wire [4-1:0] node38633;
	wire [4-1:0] node38636;
	wire [4-1:0] node38639;
	wire [4-1:0] node38640;
	wire [4-1:0] node38643;
	wire [4-1:0] node38646;
	wire [4-1:0] node38647;
	wire [4-1:0] node38648;
	wire [4-1:0] node38651;
	wire [4-1:0] node38654;
	wire [4-1:0] node38655;
	wire [4-1:0] node38658;
	wire [4-1:0] node38661;
	wire [4-1:0] node38662;
	wire [4-1:0] node38663;
	wire [4-1:0] node38664;
	wire [4-1:0] node38665;
	wire [4-1:0] node38667;
	wire [4-1:0] node38670;
	wire [4-1:0] node38671;
	wire [4-1:0] node38674;
	wire [4-1:0] node38677;
	wire [4-1:0] node38678;
	wire [4-1:0] node38679;
	wire [4-1:0] node38682;
	wire [4-1:0] node38685;
	wire [4-1:0] node38686;
	wire [4-1:0] node38690;
	wire [4-1:0] node38691;
	wire [4-1:0] node38692;
	wire [4-1:0] node38693;
	wire [4-1:0] node38696;
	wire [4-1:0] node38699;
	wire [4-1:0] node38700;
	wire [4-1:0] node38703;
	wire [4-1:0] node38706;
	wire [4-1:0] node38707;
	wire [4-1:0] node38708;
	wire [4-1:0] node38711;
	wire [4-1:0] node38714;
	wire [4-1:0] node38715;
	wire [4-1:0] node38718;
	wire [4-1:0] node38721;
	wire [4-1:0] node38722;
	wire [4-1:0] node38723;
	wire [4-1:0] node38724;
	wire [4-1:0] node38725;
	wire [4-1:0] node38728;
	wire [4-1:0] node38731;
	wire [4-1:0] node38732;
	wire [4-1:0] node38735;
	wire [4-1:0] node38738;
	wire [4-1:0] node38739;
	wire [4-1:0] node38740;
	wire [4-1:0] node38744;
	wire [4-1:0] node38745;
	wire [4-1:0] node38749;
	wire [4-1:0] node38750;
	wire [4-1:0] node38751;
	wire [4-1:0] node38752;
	wire [4-1:0] node38755;
	wire [4-1:0] node38758;
	wire [4-1:0] node38759;
	wire [4-1:0] node38762;
	wire [4-1:0] node38765;
	wire [4-1:0] node38766;
	wire [4-1:0] node38769;
	wire [4-1:0] node38772;
	wire [4-1:0] node38773;
	wire [4-1:0] node38774;
	wire [4-1:0] node38775;
	wire [4-1:0] node38776;
	wire [4-1:0] node38777;
	wire [4-1:0] node38778;
	wire [4-1:0] node38779;
	wire [4-1:0] node38782;
	wire [4-1:0] node38785;
	wire [4-1:0] node38786;
	wire [4-1:0] node38789;
	wire [4-1:0] node38792;
	wire [4-1:0] node38793;
	wire [4-1:0] node38794;
	wire [4-1:0] node38797;
	wire [4-1:0] node38800;
	wire [4-1:0] node38801;
	wire [4-1:0] node38804;
	wire [4-1:0] node38807;
	wire [4-1:0] node38808;
	wire [4-1:0] node38809;
	wire [4-1:0] node38810;
	wire [4-1:0] node38814;
	wire [4-1:0] node38815;
	wire [4-1:0] node38819;
	wire [4-1:0] node38820;
	wire [4-1:0] node38821;
	wire [4-1:0] node38825;
	wire [4-1:0] node38826;
	wire [4-1:0] node38830;
	wire [4-1:0] node38831;
	wire [4-1:0] node38832;
	wire [4-1:0] node38833;
	wire [4-1:0] node38834;
	wire [4-1:0] node38837;
	wire [4-1:0] node38840;
	wire [4-1:0] node38841;
	wire [4-1:0] node38844;
	wire [4-1:0] node38847;
	wire [4-1:0] node38848;
	wire [4-1:0] node38849;
	wire [4-1:0] node38852;
	wire [4-1:0] node38855;
	wire [4-1:0] node38856;
	wire [4-1:0] node38860;
	wire [4-1:0] node38861;
	wire [4-1:0] node38862;
	wire [4-1:0] node38863;
	wire [4-1:0] node38866;
	wire [4-1:0] node38869;
	wire [4-1:0] node38870;
	wire [4-1:0] node38873;
	wire [4-1:0] node38876;
	wire [4-1:0] node38877;
	wire [4-1:0] node38878;
	wire [4-1:0] node38882;
	wire [4-1:0] node38884;
	wire [4-1:0] node38887;
	wire [4-1:0] node38888;
	wire [4-1:0] node38889;
	wire [4-1:0] node38890;
	wire [4-1:0] node38891;
	wire [4-1:0] node38892;
	wire [4-1:0] node38895;
	wire [4-1:0] node38898;
	wire [4-1:0] node38899;
	wire [4-1:0] node38902;
	wire [4-1:0] node38905;
	wire [4-1:0] node38906;
	wire [4-1:0] node38907;
	wire [4-1:0] node38911;
	wire [4-1:0] node38912;
	wire [4-1:0] node38915;
	wire [4-1:0] node38918;
	wire [4-1:0] node38919;
	wire [4-1:0] node38920;
	wire [4-1:0] node38922;
	wire [4-1:0] node38925;
	wire [4-1:0] node38926;
	wire [4-1:0] node38929;
	wire [4-1:0] node38932;
	wire [4-1:0] node38933;
	wire [4-1:0] node38934;
	wire [4-1:0] node38937;
	wire [4-1:0] node38940;
	wire [4-1:0] node38941;
	wire [4-1:0] node38944;
	wire [4-1:0] node38947;
	wire [4-1:0] node38948;
	wire [4-1:0] node38949;
	wire [4-1:0] node38950;
	wire [4-1:0] node38951;
	wire [4-1:0] node38954;
	wire [4-1:0] node38957;
	wire [4-1:0] node38958;
	wire [4-1:0] node38961;
	wire [4-1:0] node38964;
	wire [4-1:0] node38965;
	wire [4-1:0] node38966;
	wire [4-1:0] node38969;
	wire [4-1:0] node38972;
	wire [4-1:0] node38974;
	wire [4-1:0] node38977;
	wire [4-1:0] node38978;
	wire [4-1:0] node38979;
	wire [4-1:0] node38980;
	wire [4-1:0] node38983;
	wire [4-1:0] node38986;
	wire [4-1:0] node38988;
	wire [4-1:0] node38991;
	wire [4-1:0] node38992;
	wire [4-1:0] node38995;
	wire [4-1:0] node38998;
	wire [4-1:0] node38999;
	wire [4-1:0] node39000;
	wire [4-1:0] node39001;
	wire [4-1:0] node39002;
	wire [4-1:0] node39003;
	wire [4-1:0] node39004;
	wire [4-1:0] node39007;
	wire [4-1:0] node39010;
	wire [4-1:0] node39011;
	wire [4-1:0] node39014;
	wire [4-1:0] node39017;
	wire [4-1:0] node39018;
	wire [4-1:0] node39019;
	wire [4-1:0] node39022;
	wire [4-1:0] node39025;
	wire [4-1:0] node39026;
	wire [4-1:0] node39030;
	wire [4-1:0] node39031;
	wire [4-1:0] node39032;
	wire [4-1:0] node39033;
	wire [4-1:0] node39037;
	wire [4-1:0] node39038;
	wire [4-1:0] node39042;
	wire [4-1:0] node39043;
	wire [4-1:0] node39044;
	wire [4-1:0] node39048;
	wire [4-1:0] node39049;
	wire [4-1:0] node39053;
	wire [4-1:0] node39054;
	wire [4-1:0] node39055;
	wire [4-1:0] node39056;
	wire [4-1:0] node39057;
	wire [4-1:0] node39060;
	wire [4-1:0] node39063;
	wire [4-1:0] node39065;
	wire [4-1:0] node39068;
	wire [4-1:0] node39069;
	wire [4-1:0] node39070;
	wire [4-1:0] node39073;
	wire [4-1:0] node39076;
	wire [4-1:0] node39077;
	wire [4-1:0] node39081;
	wire [4-1:0] node39082;
	wire [4-1:0] node39083;
	wire [4-1:0] node39084;
	wire [4-1:0] node39087;
	wire [4-1:0] node39090;
	wire [4-1:0] node39091;
	wire [4-1:0] node39095;
	wire [4-1:0] node39096;
	wire [4-1:0] node39097;
	wire [4-1:0] node39100;
	wire [4-1:0] node39103;
	wire [4-1:0] node39104;
	wire [4-1:0] node39107;
	wire [4-1:0] node39110;
	wire [4-1:0] node39111;
	wire [4-1:0] node39112;
	wire [4-1:0] node39113;
	wire [4-1:0] node39114;
	wire [4-1:0] node39115;
	wire [4-1:0] node39118;
	wire [4-1:0] node39121;
	wire [4-1:0] node39122;
	wire [4-1:0] node39126;
	wire [4-1:0] node39127;
	wire [4-1:0] node39129;
	wire [4-1:0] node39132;
	wire [4-1:0] node39133;
	wire [4-1:0] node39136;
	wire [4-1:0] node39139;
	wire [4-1:0] node39140;
	wire [4-1:0] node39141;
	wire [4-1:0] node39142;
	wire [4-1:0] node39146;
	wire [4-1:0] node39147;
	wire [4-1:0] node39151;
	wire [4-1:0] node39152;
	wire [4-1:0] node39153;
	wire [4-1:0] node39157;
	wire [4-1:0] node39158;
	wire [4-1:0] node39162;
	wire [4-1:0] node39163;
	wire [4-1:0] node39164;
	wire [4-1:0] node39165;
	wire [4-1:0] node39166;
	wire [4-1:0] node39169;
	wire [4-1:0] node39172;
	wire [4-1:0] node39174;
	wire [4-1:0] node39177;
	wire [4-1:0] node39178;
	wire [4-1:0] node39179;
	wire [4-1:0] node39182;
	wire [4-1:0] node39185;
	wire [4-1:0] node39186;
	wire [4-1:0] node39189;
	wire [4-1:0] node39192;
	wire [4-1:0] node39193;
	wire [4-1:0] node39194;
	wire [4-1:0] node39195;
	wire [4-1:0] node39198;
	wire [4-1:0] node39201;
	wire [4-1:0] node39202;
	wire [4-1:0] node39205;
	wire [4-1:0] node39208;
	wire [4-1:0] node39209;
	wire [4-1:0] node39210;
	wire [4-1:0] node39213;
	wire [4-1:0] node39216;
	wire [4-1:0] node39217;
	wire [4-1:0] node39220;
	wire [4-1:0] node39223;
	wire [4-1:0] node39224;
	wire [4-1:0] node39225;
	wire [4-1:0] node39226;
	wire [4-1:0] node39227;
	wire [4-1:0] node39228;
	wire [4-1:0] node39229;
	wire [4-1:0] node39230;
	wire [4-1:0] node39231;
	wire [4-1:0] node39232;
	wire [4-1:0] node39233;
	wire [4-1:0] node39236;
	wire [4-1:0] node39239;
	wire [4-1:0] node39240;
	wire [4-1:0] node39243;
	wire [4-1:0] node39246;
	wire [4-1:0] node39247;
	wire [4-1:0] node39248;
	wire [4-1:0] node39252;
	wire [4-1:0] node39253;
	wire [4-1:0] node39256;
	wire [4-1:0] node39259;
	wire [4-1:0] node39260;
	wire [4-1:0] node39261;
	wire [4-1:0] node39262;
	wire [4-1:0] node39265;
	wire [4-1:0] node39268;
	wire [4-1:0] node39269;
	wire [4-1:0] node39272;
	wire [4-1:0] node39275;
	wire [4-1:0] node39276;
	wire [4-1:0] node39277;
	wire [4-1:0] node39280;
	wire [4-1:0] node39283;
	wire [4-1:0] node39284;
	wire [4-1:0] node39287;
	wire [4-1:0] node39290;
	wire [4-1:0] node39291;
	wire [4-1:0] node39292;
	wire [4-1:0] node39293;
	wire [4-1:0] node39294;
	wire [4-1:0] node39297;
	wire [4-1:0] node39300;
	wire [4-1:0] node39301;
	wire [4-1:0] node39304;
	wire [4-1:0] node39307;
	wire [4-1:0] node39308;
	wire [4-1:0] node39309;
	wire [4-1:0] node39313;
	wire [4-1:0] node39314;
	wire [4-1:0] node39317;
	wire [4-1:0] node39320;
	wire [4-1:0] node39321;
	wire [4-1:0] node39322;
	wire [4-1:0] node39323;
	wire [4-1:0] node39326;
	wire [4-1:0] node39329;
	wire [4-1:0] node39330;
	wire [4-1:0] node39333;
	wire [4-1:0] node39336;
	wire [4-1:0] node39337;
	wire [4-1:0] node39338;
	wire [4-1:0] node39341;
	wire [4-1:0] node39344;
	wire [4-1:0] node39345;
	wire [4-1:0] node39348;
	wire [4-1:0] node39351;
	wire [4-1:0] node39352;
	wire [4-1:0] node39353;
	wire [4-1:0] node39354;
	wire [4-1:0] node39355;
	wire [4-1:0] node39356;
	wire [4-1:0] node39359;
	wire [4-1:0] node39362;
	wire [4-1:0] node39363;
	wire [4-1:0] node39366;
	wire [4-1:0] node39369;
	wire [4-1:0] node39370;
	wire [4-1:0] node39371;
	wire [4-1:0] node39374;
	wire [4-1:0] node39377;
	wire [4-1:0] node39378;
	wire [4-1:0] node39381;
	wire [4-1:0] node39384;
	wire [4-1:0] node39385;
	wire [4-1:0] node39386;
	wire [4-1:0] node39387;
	wire [4-1:0] node39390;
	wire [4-1:0] node39393;
	wire [4-1:0] node39394;
	wire [4-1:0] node39397;
	wire [4-1:0] node39400;
	wire [4-1:0] node39401;
	wire [4-1:0] node39402;
	wire [4-1:0] node39405;
	wire [4-1:0] node39408;
	wire [4-1:0] node39410;
	wire [4-1:0] node39413;
	wire [4-1:0] node39414;
	wire [4-1:0] node39415;
	wire [4-1:0] node39416;
	wire [4-1:0] node39417;
	wire [4-1:0] node39420;
	wire [4-1:0] node39423;
	wire [4-1:0] node39424;
	wire [4-1:0] node39427;
	wire [4-1:0] node39430;
	wire [4-1:0] node39431;
	wire [4-1:0] node39432;
	wire [4-1:0] node39435;
	wire [4-1:0] node39438;
	wire [4-1:0] node39439;
	wire [4-1:0] node39442;
	wire [4-1:0] node39445;
	wire [4-1:0] node39446;
	wire [4-1:0] node39447;
	wire [4-1:0] node39448;
	wire [4-1:0] node39451;
	wire [4-1:0] node39454;
	wire [4-1:0] node39456;
	wire [4-1:0] node39459;
	wire [4-1:0] node39460;
	wire [4-1:0] node39461;
	wire [4-1:0] node39464;
	wire [4-1:0] node39467;
	wire [4-1:0] node39469;
	wire [4-1:0] node39472;
	wire [4-1:0] node39473;
	wire [4-1:0] node39474;
	wire [4-1:0] node39475;
	wire [4-1:0] node39476;
	wire [4-1:0] node39477;
	wire [4-1:0] node39478;
	wire [4-1:0] node39482;
	wire [4-1:0] node39483;
	wire [4-1:0] node39486;
	wire [4-1:0] node39489;
	wire [4-1:0] node39490;
	wire [4-1:0] node39491;
	wire [4-1:0] node39494;
	wire [4-1:0] node39497;
	wire [4-1:0] node39498;
	wire [4-1:0] node39501;
	wire [4-1:0] node39504;
	wire [4-1:0] node39505;
	wire [4-1:0] node39506;
	wire [4-1:0] node39507;
	wire [4-1:0] node39510;
	wire [4-1:0] node39513;
	wire [4-1:0] node39514;
	wire [4-1:0] node39517;
	wire [4-1:0] node39520;
	wire [4-1:0] node39521;
	wire [4-1:0] node39522;
	wire [4-1:0] node39525;
	wire [4-1:0] node39528;
	wire [4-1:0] node39529;
	wire [4-1:0] node39532;
	wire [4-1:0] node39535;
	wire [4-1:0] node39536;
	wire [4-1:0] node39537;
	wire [4-1:0] node39538;
	wire [4-1:0] node39539;
	wire [4-1:0] node39542;
	wire [4-1:0] node39545;
	wire [4-1:0] node39546;
	wire [4-1:0] node39549;
	wire [4-1:0] node39552;
	wire [4-1:0] node39553;
	wire [4-1:0] node39554;
	wire [4-1:0] node39557;
	wire [4-1:0] node39560;
	wire [4-1:0] node39561;
	wire [4-1:0] node39565;
	wire [4-1:0] node39566;
	wire [4-1:0] node39567;
	wire [4-1:0] node39568;
	wire [4-1:0] node39571;
	wire [4-1:0] node39574;
	wire [4-1:0] node39575;
	wire [4-1:0] node39578;
	wire [4-1:0] node39581;
	wire [4-1:0] node39582;
	wire [4-1:0] node39583;
	wire [4-1:0] node39586;
	wire [4-1:0] node39589;
	wire [4-1:0] node39590;
	wire [4-1:0] node39593;
	wire [4-1:0] node39596;
	wire [4-1:0] node39597;
	wire [4-1:0] node39598;
	wire [4-1:0] node39599;
	wire [4-1:0] node39600;
	wire [4-1:0] node39601;
	wire [4-1:0] node39604;
	wire [4-1:0] node39607;
	wire [4-1:0] node39608;
	wire [4-1:0] node39611;
	wire [4-1:0] node39614;
	wire [4-1:0] node39615;
	wire [4-1:0] node39616;
	wire [4-1:0] node39619;
	wire [4-1:0] node39622;
	wire [4-1:0] node39623;
	wire [4-1:0] node39626;
	wire [4-1:0] node39629;
	wire [4-1:0] node39630;
	wire [4-1:0] node39631;
	wire [4-1:0] node39632;
	wire [4-1:0] node39635;
	wire [4-1:0] node39638;
	wire [4-1:0] node39639;
	wire [4-1:0] node39642;
	wire [4-1:0] node39645;
	wire [4-1:0] node39646;
	wire [4-1:0] node39647;
	wire [4-1:0] node39650;
	wire [4-1:0] node39653;
	wire [4-1:0] node39654;
	wire [4-1:0] node39657;
	wire [4-1:0] node39660;
	wire [4-1:0] node39661;
	wire [4-1:0] node39662;
	wire [4-1:0] node39663;
	wire [4-1:0] node39664;
	wire [4-1:0] node39667;
	wire [4-1:0] node39670;
	wire [4-1:0] node39671;
	wire [4-1:0] node39674;
	wire [4-1:0] node39677;
	wire [4-1:0] node39678;
	wire [4-1:0] node39679;
	wire [4-1:0] node39682;
	wire [4-1:0] node39685;
	wire [4-1:0] node39686;
	wire [4-1:0] node39689;
	wire [4-1:0] node39692;
	wire [4-1:0] node39693;
	wire [4-1:0] node39694;
	wire [4-1:0] node39696;
	wire [4-1:0] node39699;
	wire [4-1:0] node39700;
	wire [4-1:0] node39703;
	wire [4-1:0] node39706;
	wire [4-1:0] node39707;
	wire [4-1:0] node39709;
	wire [4-1:0] node39712;
	wire [4-1:0] node39713;
	wire [4-1:0] node39716;
	wire [4-1:0] node39719;
	wire [4-1:0] node39720;
	wire [4-1:0] node39721;
	wire [4-1:0] node39722;
	wire [4-1:0] node39723;
	wire [4-1:0] node39724;
	wire [4-1:0] node39725;
	wire [4-1:0] node39726;
	wire [4-1:0] node39729;
	wire [4-1:0] node39732;
	wire [4-1:0] node39733;
	wire [4-1:0] node39736;
	wire [4-1:0] node39739;
	wire [4-1:0] node39740;
	wire [4-1:0] node39741;
	wire [4-1:0] node39744;
	wire [4-1:0] node39747;
	wire [4-1:0] node39748;
	wire [4-1:0] node39751;
	wire [4-1:0] node39754;
	wire [4-1:0] node39755;
	wire [4-1:0] node39756;
	wire [4-1:0] node39757;
	wire [4-1:0] node39760;
	wire [4-1:0] node39763;
	wire [4-1:0] node39764;
	wire [4-1:0] node39767;
	wire [4-1:0] node39770;
	wire [4-1:0] node39771;
	wire [4-1:0] node39773;
	wire [4-1:0] node39776;
	wire [4-1:0] node39777;
	wire [4-1:0] node39780;
	wire [4-1:0] node39783;
	wire [4-1:0] node39784;
	wire [4-1:0] node39785;
	wire [4-1:0] node39786;
	wire [4-1:0] node39787;
	wire [4-1:0] node39790;
	wire [4-1:0] node39793;
	wire [4-1:0] node39794;
	wire [4-1:0] node39797;
	wire [4-1:0] node39800;
	wire [4-1:0] node39801;
	wire [4-1:0] node39802;
	wire [4-1:0] node39805;
	wire [4-1:0] node39808;
	wire [4-1:0] node39809;
	wire [4-1:0] node39812;
	wire [4-1:0] node39815;
	wire [4-1:0] node39816;
	wire [4-1:0] node39817;
	wire [4-1:0] node39818;
	wire [4-1:0] node39821;
	wire [4-1:0] node39824;
	wire [4-1:0] node39825;
	wire [4-1:0] node39828;
	wire [4-1:0] node39831;
	wire [4-1:0] node39832;
	wire [4-1:0] node39833;
	wire [4-1:0] node39836;
	wire [4-1:0] node39839;
	wire [4-1:0] node39840;
	wire [4-1:0] node39843;
	wire [4-1:0] node39846;
	wire [4-1:0] node39847;
	wire [4-1:0] node39848;
	wire [4-1:0] node39849;
	wire [4-1:0] node39850;
	wire [4-1:0] node39851;
	wire [4-1:0] node39854;
	wire [4-1:0] node39857;
	wire [4-1:0] node39858;
	wire [4-1:0] node39861;
	wire [4-1:0] node39864;
	wire [4-1:0] node39865;
	wire [4-1:0] node39866;
	wire [4-1:0] node39869;
	wire [4-1:0] node39872;
	wire [4-1:0] node39873;
	wire [4-1:0] node39876;
	wire [4-1:0] node39879;
	wire [4-1:0] node39880;
	wire [4-1:0] node39881;
	wire [4-1:0] node39882;
	wire [4-1:0] node39885;
	wire [4-1:0] node39888;
	wire [4-1:0] node39889;
	wire [4-1:0] node39892;
	wire [4-1:0] node39895;
	wire [4-1:0] node39896;
	wire [4-1:0] node39898;
	wire [4-1:0] node39901;
	wire [4-1:0] node39903;
	wire [4-1:0] node39906;
	wire [4-1:0] node39907;
	wire [4-1:0] node39908;
	wire [4-1:0] node39909;
	wire [4-1:0] node39910;
	wire [4-1:0] node39913;
	wire [4-1:0] node39916;
	wire [4-1:0] node39917;
	wire [4-1:0] node39920;
	wire [4-1:0] node39923;
	wire [4-1:0] node39924;
	wire [4-1:0] node39925;
	wire [4-1:0] node39928;
	wire [4-1:0] node39931;
	wire [4-1:0] node39932;
	wire [4-1:0] node39935;
	wire [4-1:0] node39938;
	wire [4-1:0] node39939;
	wire [4-1:0] node39940;
	wire [4-1:0] node39941;
	wire [4-1:0] node39944;
	wire [4-1:0] node39947;
	wire [4-1:0] node39948;
	wire [4-1:0] node39951;
	wire [4-1:0] node39954;
	wire [4-1:0] node39955;
	wire [4-1:0] node39956;
	wire [4-1:0] node39959;
	wire [4-1:0] node39962;
	wire [4-1:0] node39963;
	wire [4-1:0] node39966;
	wire [4-1:0] node39969;
	wire [4-1:0] node39970;
	wire [4-1:0] node39971;
	wire [4-1:0] node39972;
	wire [4-1:0] node39973;
	wire [4-1:0] node39974;
	wire [4-1:0] node39975;
	wire [4-1:0] node39978;
	wire [4-1:0] node39981;
	wire [4-1:0] node39982;
	wire [4-1:0] node39985;
	wire [4-1:0] node39988;
	wire [4-1:0] node39989;
	wire [4-1:0] node39990;
	wire [4-1:0] node39993;
	wire [4-1:0] node39996;
	wire [4-1:0] node39997;
	wire [4-1:0] node40000;
	wire [4-1:0] node40003;
	wire [4-1:0] node40004;
	wire [4-1:0] node40005;
	wire [4-1:0] node40006;
	wire [4-1:0] node40009;
	wire [4-1:0] node40012;
	wire [4-1:0] node40013;
	wire [4-1:0] node40016;
	wire [4-1:0] node40019;
	wire [4-1:0] node40020;
	wire [4-1:0] node40021;
	wire [4-1:0] node40024;
	wire [4-1:0] node40027;
	wire [4-1:0] node40028;
	wire [4-1:0] node40031;
	wire [4-1:0] node40034;
	wire [4-1:0] node40035;
	wire [4-1:0] node40036;
	wire [4-1:0] node40037;
	wire [4-1:0] node40038;
	wire [4-1:0] node40041;
	wire [4-1:0] node40044;
	wire [4-1:0] node40045;
	wire [4-1:0] node40048;
	wire [4-1:0] node40051;
	wire [4-1:0] node40052;
	wire [4-1:0] node40053;
	wire [4-1:0] node40056;
	wire [4-1:0] node40059;
	wire [4-1:0] node40060;
	wire [4-1:0] node40063;
	wire [4-1:0] node40066;
	wire [4-1:0] node40067;
	wire [4-1:0] node40068;
	wire [4-1:0] node40069;
	wire [4-1:0] node40072;
	wire [4-1:0] node40075;
	wire [4-1:0] node40076;
	wire [4-1:0] node40079;
	wire [4-1:0] node40082;
	wire [4-1:0] node40083;
	wire [4-1:0] node40084;
	wire [4-1:0] node40087;
	wire [4-1:0] node40090;
	wire [4-1:0] node40091;
	wire [4-1:0] node40094;
	wire [4-1:0] node40097;
	wire [4-1:0] node40098;
	wire [4-1:0] node40099;
	wire [4-1:0] node40100;
	wire [4-1:0] node40101;
	wire [4-1:0] node40102;
	wire [4-1:0] node40105;
	wire [4-1:0] node40108;
	wire [4-1:0] node40109;
	wire [4-1:0] node40112;
	wire [4-1:0] node40115;
	wire [4-1:0] node40116;
	wire [4-1:0] node40118;
	wire [4-1:0] node40121;
	wire [4-1:0] node40122;
	wire [4-1:0] node40125;
	wire [4-1:0] node40128;
	wire [4-1:0] node40129;
	wire [4-1:0] node40130;
	wire [4-1:0] node40131;
	wire [4-1:0] node40134;
	wire [4-1:0] node40137;
	wire [4-1:0] node40138;
	wire [4-1:0] node40141;
	wire [4-1:0] node40144;
	wire [4-1:0] node40145;
	wire [4-1:0] node40146;
	wire [4-1:0] node40149;
	wire [4-1:0] node40152;
	wire [4-1:0] node40153;
	wire [4-1:0] node40156;
	wire [4-1:0] node40159;
	wire [4-1:0] node40160;
	wire [4-1:0] node40161;
	wire [4-1:0] node40162;
	wire [4-1:0] node40163;
	wire [4-1:0] node40166;
	wire [4-1:0] node40169;
	wire [4-1:0] node40170;
	wire [4-1:0] node40173;
	wire [4-1:0] node40176;
	wire [4-1:0] node40177;
	wire [4-1:0] node40178;
	wire [4-1:0] node40181;
	wire [4-1:0] node40184;
	wire [4-1:0] node40185;
	wire [4-1:0] node40188;
	wire [4-1:0] node40191;
	wire [4-1:0] node40192;
	wire [4-1:0] node40193;
	wire [4-1:0] node40194;
	wire [4-1:0] node40197;
	wire [4-1:0] node40200;
	wire [4-1:0] node40203;
	wire [4-1:0] node40204;
	wire [4-1:0] node40205;
	wire [4-1:0] node40208;
	wire [4-1:0] node40211;
	wire [4-1:0] node40212;
	wire [4-1:0] node40215;
	wire [4-1:0] node40218;
	wire [4-1:0] node40219;
	wire [4-1:0] node40220;
	wire [4-1:0] node40221;
	wire [4-1:0] node40222;
	wire [4-1:0] node40223;
	wire [4-1:0] node40224;
	wire [4-1:0] node40225;
	wire [4-1:0] node40226;
	wire [4-1:0] node40229;
	wire [4-1:0] node40232;
	wire [4-1:0] node40233;
	wire [4-1:0] node40236;
	wire [4-1:0] node40239;
	wire [4-1:0] node40240;
	wire [4-1:0] node40241;
	wire [4-1:0] node40244;
	wire [4-1:0] node40247;
	wire [4-1:0] node40248;
	wire [4-1:0] node40251;
	wire [4-1:0] node40254;
	wire [4-1:0] node40255;
	wire [4-1:0] node40256;
	wire [4-1:0] node40257;
	wire [4-1:0] node40260;
	wire [4-1:0] node40263;
	wire [4-1:0] node40264;
	wire [4-1:0] node40267;
	wire [4-1:0] node40270;
	wire [4-1:0] node40271;
	wire [4-1:0] node40273;
	wire [4-1:0] node40276;
	wire [4-1:0] node40277;
	wire [4-1:0] node40280;
	wire [4-1:0] node40283;
	wire [4-1:0] node40284;
	wire [4-1:0] node40285;
	wire [4-1:0] node40286;
	wire [4-1:0] node40287;
	wire [4-1:0] node40290;
	wire [4-1:0] node40293;
	wire [4-1:0] node40294;
	wire [4-1:0] node40297;
	wire [4-1:0] node40300;
	wire [4-1:0] node40301;
	wire [4-1:0] node40302;
	wire [4-1:0] node40305;
	wire [4-1:0] node40308;
	wire [4-1:0] node40309;
	wire [4-1:0] node40312;
	wire [4-1:0] node40315;
	wire [4-1:0] node40316;
	wire [4-1:0] node40317;
	wire [4-1:0] node40318;
	wire [4-1:0] node40321;
	wire [4-1:0] node40324;
	wire [4-1:0] node40325;
	wire [4-1:0] node40328;
	wire [4-1:0] node40331;
	wire [4-1:0] node40332;
	wire [4-1:0] node40333;
	wire [4-1:0] node40336;
	wire [4-1:0] node40339;
	wire [4-1:0] node40340;
	wire [4-1:0] node40343;
	wire [4-1:0] node40346;
	wire [4-1:0] node40347;
	wire [4-1:0] node40348;
	wire [4-1:0] node40349;
	wire [4-1:0] node40350;
	wire [4-1:0] node40351;
	wire [4-1:0] node40354;
	wire [4-1:0] node40357;
	wire [4-1:0] node40358;
	wire [4-1:0] node40361;
	wire [4-1:0] node40364;
	wire [4-1:0] node40365;
	wire [4-1:0] node40366;
	wire [4-1:0] node40369;
	wire [4-1:0] node40372;
	wire [4-1:0] node40373;
	wire [4-1:0] node40376;
	wire [4-1:0] node40379;
	wire [4-1:0] node40380;
	wire [4-1:0] node40381;
	wire [4-1:0] node40382;
	wire [4-1:0] node40385;
	wire [4-1:0] node40388;
	wire [4-1:0] node40389;
	wire [4-1:0] node40392;
	wire [4-1:0] node40395;
	wire [4-1:0] node40396;
	wire [4-1:0] node40397;
	wire [4-1:0] node40400;
	wire [4-1:0] node40403;
	wire [4-1:0] node40404;
	wire [4-1:0] node40407;
	wire [4-1:0] node40410;
	wire [4-1:0] node40411;
	wire [4-1:0] node40412;
	wire [4-1:0] node40413;
	wire [4-1:0] node40414;
	wire [4-1:0] node40417;
	wire [4-1:0] node40420;
	wire [4-1:0] node40421;
	wire [4-1:0] node40424;
	wire [4-1:0] node40427;
	wire [4-1:0] node40428;
	wire [4-1:0] node40429;
	wire [4-1:0] node40432;
	wire [4-1:0] node40435;
	wire [4-1:0] node40436;
	wire [4-1:0] node40439;
	wire [4-1:0] node40442;
	wire [4-1:0] node40443;
	wire [4-1:0] node40444;
	wire [4-1:0] node40445;
	wire [4-1:0] node40448;
	wire [4-1:0] node40451;
	wire [4-1:0] node40452;
	wire [4-1:0] node40455;
	wire [4-1:0] node40458;
	wire [4-1:0] node40459;
	wire [4-1:0] node40460;
	wire [4-1:0] node40464;
	wire [4-1:0] node40465;
	wire [4-1:0] node40468;
	wire [4-1:0] node40471;
	wire [4-1:0] node40472;
	wire [4-1:0] node40473;
	wire [4-1:0] node40474;
	wire [4-1:0] node40475;
	wire [4-1:0] node40476;
	wire [4-1:0] node40477;
	wire [4-1:0] node40481;
	wire [4-1:0] node40483;
	wire [4-1:0] node40486;
	wire [4-1:0] node40487;
	wire [4-1:0] node40488;
	wire [4-1:0] node40491;
	wire [4-1:0] node40494;
	wire [4-1:0] node40495;
	wire [4-1:0] node40498;
	wire [4-1:0] node40501;
	wire [4-1:0] node40502;
	wire [4-1:0] node40503;
	wire [4-1:0] node40504;
	wire [4-1:0] node40508;
	wire [4-1:0] node40509;
	wire [4-1:0] node40512;
	wire [4-1:0] node40515;
	wire [4-1:0] node40516;
	wire [4-1:0] node40517;
	wire [4-1:0] node40520;
	wire [4-1:0] node40523;
	wire [4-1:0] node40524;
	wire [4-1:0] node40527;
	wire [4-1:0] node40530;
	wire [4-1:0] node40531;
	wire [4-1:0] node40532;
	wire [4-1:0] node40533;
	wire [4-1:0] node40534;
	wire [4-1:0] node40537;
	wire [4-1:0] node40540;
	wire [4-1:0] node40541;
	wire [4-1:0] node40544;
	wire [4-1:0] node40547;
	wire [4-1:0] node40548;
	wire [4-1:0] node40549;
	wire [4-1:0] node40552;
	wire [4-1:0] node40555;
	wire [4-1:0] node40558;
	wire [4-1:0] node40559;
	wire [4-1:0] node40560;
	wire [4-1:0] node40561;
	wire [4-1:0] node40564;
	wire [4-1:0] node40567;
	wire [4-1:0] node40569;
	wire [4-1:0] node40572;
	wire [4-1:0] node40573;
	wire [4-1:0] node40574;
	wire [4-1:0] node40577;
	wire [4-1:0] node40580;
	wire [4-1:0] node40581;
	wire [4-1:0] node40584;
	wire [4-1:0] node40587;
	wire [4-1:0] node40588;
	wire [4-1:0] node40589;
	wire [4-1:0] node40590;
	wire [4-1:0] node40591;
	wire [4-1:0] node40592;
	wire [4-1:0] node40595;
	wire [4-1:0] node40598;
	wire [4-1:0] node40599;
	wire [4-1:0] node40602;
	wire [4-1:0] node40605;
	wire [4-1:0] node40606;
	wire [4-1:0] node40607;
	wire [4-1:0] node40610;
	wire [4-1:0] node40613;
	wire [4-1:0] node40614;
	wire [4-1:0] node40617;
	wire [4-1:0] node40620;
	wire [4-1:0] node40621;
	wire [4-1:0] node40622;
	wire [4-1:0] node40623;
	wire [4-1:0] node40627;
	wire [4-1:0] node40628;
	wire [4-1:0] node40631;
	wire [4-1:0] node40634;
	wire [4-1:0] node40635;
	wire [4-1:0] node40636;
	wire [4-1:0] node40639;
	wire [4-1:0] node40642;
	wire [4-1:0] node40643;
	wire [4-1:0] node40646;
	wire [4-1:0] node40649;
	wire [4-1:0] node40650;
	wire [4-1:0] node40651;
	wire [4-1:0] node40652;
	wire [4-1:0] node40653;
	wire [4-1:0] node40656;
	wire [4-1:0] node40659;
	wire [4-1:0] node40660;
	wire [4-1:0] node40663;
	wire [4-1:0] node40666;
	wire [4-1:0] node40667;
	wire [4-1:0] node40669;
	wire [4-1:0] node40672;
	wire [4-1:0] node40673;
	wire [4-1:0] node40676;
	wire [4-1:0] node40679;
	wire [4-1:0] node40680;
	wire [4-1:0] node40681;
	wire [4-1:0] node40682;
	wire [4-1:0] node40685;
	wire [4-1:0] node40688;
	wire [4-1:0] node40690;
	wire [4-1:0] node40693;
	wire [4-1:0] node40694;
	wire [4-1:0] node40695;
	wire [4-1:0] node40699;
	wire [4-1:0] node40700;
	wire [4-1:0] node40703;
	wire [4-1:0] node40706;
	wire [4-1:0] node40707;
	wire [4-1:0] node40708;
	wire [4-1:0] node40709;
	wire [4-1:0] node40710;
	wire [4-1:0] node40711;
	wire [4-1:0] node40712;
	wire [4-1:0] node40713;
	wire [4-1:0] node40716;
	wire [4-1:0] node40719;
	wire [4-1:0] node40720;
	wire [4-1:0] node40723;
	wire [4-1:0] node40726;
	wire [4-1:0] node40727;
	wire [4-1:0] node40728;
	wire [4-1:0] node40731;
	wire [4-1:0] node40734;
	wire [4-1:0] node40737;
	wire [4-1:0] node40738;
	wire [4-1:0] node40739;
	wire [4-1:0] node40740;
	wire [4-1:0] node40743;
	wire [4-1:0] node40746;
	wire [4-1:0] node40747;
	wire [4-1:0] node40750;
	wire [4-1:0] node40753;
	wire [4-1:0] node40754;
	wire [4-1:0] node40755;
	wire [4-1:0] node40758;
	wire [4-1:0] node40761;
	wire [4-1:0] node40762;
	wire [4-1:0] node40765;
	wire [4-1:0] node40768;
	wire [4-1:0] node40769;
	wire [4-1:0] node40770;
	wire [4-1:0] node40771;
	wire [4-1:0] node40772;
	wire [4-1:0] node40775;
	wire [4-1:0] node40778;
	wire [4-1:0] node40779;
	wire [4-1:0] node40782;
	wire [4-1:0] node40785;
	wire [4-1:0] node40786;
	wire [4-1:0] node40787;
	wire [4-1:0] node40790;
	wire [4-1:0] node40793;
	wire [4-1:0] node40795;
	wire [4-1:0] node40798;
	wire [4-1:0] node40799;
	wire [4-1:0] node40800;
	wire [4-1:0] node40801;
	wire [4-1:0] node40804;
	wire [4-1:0] node40807;
	wire [4-1:0] node40808;
	wire [4-1:0] node40811;
	wire [4-1:0] node40814;
	wire [4-1:0] node40815;
	wire [4-1:0] node40816;
	wire [4-1:0] node40819;
	wire [4-1:0] node40822;
	wire [4-1:0] node40823;
	wire [4-1:0] node40826;
	wire [4-1:0] node40829;
	wire [4-1:0] node40830;
	wire [4-1:0] node40831;
	wire [4-1:0] node40832;
	wire [4-1:0] node40833;
	wire [4-1:0] node40834;
	wire [4-1:0] node40837;
	wire [4-1:0] node40840;
	wire [4-1:0] node40841;
	wire [4-1:0] node40844;
	wire [4-1:0] node40847;
	wire [4-1:0] node40848;
	wire [4-1:0] node40849;
	wire [4-1:0] node40852;
	wire [4-1:0] node40855;
	wire [4-1:0] node40856;
	wire [4-1:0] node40859;
	wire [4-1:0] node40862;
	wire [4-1:0] node40863;
	wire [4-1:0] node40864;
	wire [4-1:0] node40865;
	wire [4-1:0] node40868;
	wire [4-1:0] node40871;
	wire [4-1:0] node40872;
	wire [4-1:0] node40875;
	wire [4-1:0] node40878;
	wire [4-1:0] node40879;
	wire [4-1:0] node40880;
	wire [4-1:0] node40883;
	wire [4-1:0] node40886;
	wire [4-1:0] node40887;
	wire [4-1:0] node40890;
	wire [4-1:0] node40893;
	wire [4-1:0] node40894;
	wire [4-1:0] node40895;
	wire [4-1:0] node40896;
	wire [4-1:0] node40897;
	wire [4-1:0] node40900;
	wire [4-1:0] node40903;
	wire [4-1:0] node40904;
	wire [4-1:0] node40907;
	wire [4-1:0] node40910;
	wire [4-1:0] node40911;
	wire [4-1:0] node40912;
	wire [4-1:0] node40915;
	wire [4-1:0] node40918;
	wire [4-1:0] node40919;
	wire [4-1:0] node40922;
	wire [4-1:0] node40925;
	wire [4-1:0] node40926;
	wire [4-1:0] node40927;
	wire [4-1:0] node40928;
	wire [4-1:0] node40931;
	wire [4-1:0] node40934;
	wire [4-1:0] node40935;
	wire [4-1:0] node40938;
	wire [4-1:0] node40941;
	wire [4-1:0] node40942;
	wire [4-1:0] node40943;
	wire [4-1:0] node40946;
	wire [4-1:0] node40949;
	wire [4-1:0] node40950;
	wire [4-1:0] node40953;
	wire [4-1:0] node40956;
	wire [4-1:0] node40957;
	wire [4-1:0] node40958;
	wire [4-1:0] node40959;
	wire [4-1:0] node40960;
	wire [4-1:0] node40961;
	wire [4-1:0] node40962;
	wire [4-1:0] node40965;
	wire [4-1:0] node40968;
	wire [4-1:0] node40969;
	wire [4-1:0] node40972;
	wire [4-1:0] node40975;
	wire [4-1:0] node40976;
	wire [4-1:0] node40979;
	wire [4-1:0] node40980;
	wire [4-1:0] node40983;
	wire [4-1:0] node40986;
	wire [4-1:0] node40987;
	wire [4-1:0] node40988;
	wire [4-1:0] node40989;
	wire [4-1:0] node40992;
	wire [4-1:0] node40995;
	wire [4-1:0] node40996;
	wire [4-1:0] node40999;
	wire [4-1:0] node41002;
	wire [4-1:0] node41003;
	wire [4-1:0] node41004;
	wire [4-1:0] node41007;
	wire [4-1:0] node41010;
	wire [4-1:0] node41011;
	wire [4-1:0] node41014;
	wire [4-1:0] node41017;
	wire [4-1:0] node41018;
	wire [4-1:0] node41019;
	wire [4-1:0] node41020;
	wire [4-1:0] node41021;
	wire [4-1:0] node41024;
	wire [4-1:0] node41027;
	wire [4-1:0] node41028;
	wire [4-1:0] node41031;
	wire [4-1:0] node41034;
	wire [4-1:0] node41035;
	wire [4-1:0] node41036;
	wire [4-1:0] node41039;
	wire [4-1:0] node41042;
	wire [4-1:0] node41043;
	wire [4-1:0] node41046;
	wire [4-1:0] node41049;
	wire [4-1:0] node41050;
	wire [4-1:0] node41051;
	wire [4-1:0] node41052;
	wire [4-1:0] node41055;
	wire [4-1:0] node41058;
	wire [4-1:0] node41059;
	wire [4-1:0] node41063;
	wire [4-1:0] node41064;
	wire [4-1:0] node41065;
	wire [4-1:0] node41068;
	wire [4-1:0] node41071;
	wire [4-1:0] node41072;
	wire [4-1:0] node41075;
	wire [4-1:0] node41078;
	wire [4-1:0] node41079;
	wire [4-1:0] node41080;
	wire [4-1:0] node41081;
	wire [4-1:0] node41082;
	wire [4-1:0] node41083;
	wire [4-1:0] node41086;
	wire [4-1:0] node41089;
	wire [4-1:0] node41090;
	wire [4-1:0] node41093;
	wire [4-1:0] node41096;
	wire [4-1:0] node41097;
	wire [4-1:0] node41098;
	wire [4-1:0] node41101;
	wire [4-1:0] node41104;
	wire [4-1:0] node41105;
	wire [4-1:0] node41108;
	wire [4-1:0] node41111;
	wire [4-1:0] node41112;
	wire [4-1:0] node41113;
	wire [4-1:0] node41114;
	wire [4-1:0] node41117;
	wire [4-1:0] node41120;
	wire [4-1:0] node41121;
	wire [4-1:0] node41124;
	wire [4-1:0] node41127;
	wire [4-1:0] node41128;
	wire [4-1:0] node41129;
	wire [4-1:0] node41132;
	wire [4-1:0] node41135;
	wire [4-1:0] node41136;
	wire [4-1:0] node41139;
	wire [4-1:0] node41142;
	wire [4-1:0] node41143;
	wire [4-1:0] node41144;
	wire [4-1:0] node41145;
	wire [4-1:0] node41146;
	wire [4-1:0] node41149;
	wire [4-1:0] node41152;
	wire [4-1:0] node41153;
	wire [4-1:0] node41156;
	wire [4-1:0] node41159;
	wire [4-1:0] node41160;
	wire [4-1:0] node41161;
	wire [4-1:0] node41164;
	wire [4-1:0] node41167;
	wire [4-1:0] node41168;
	wire [4-1:0] node41171;
	wire [4-1:0] node41174;
	wire [4-1:0] node41175;
	wire [4-1:0] node41176;
	wire [4-1:0] node41177;
	wire [4-1:0] node41180;
	wire [4-1:0] node41183;
	wire [4-1:0] node41185;
	wire [4-1:0] node41188;
	wire [4-1:0] node41189;
	wire [4-1:0] node41190;
	wire [4-1:0] node41194;
	wire [4-1:0] node41195;
	wire [4-1:0] node41198;
	wire [4-1:0] node41201;
	wire [4-1:0] node41202;
	wire [4-1:0] node41203;
	wire [4-1:0] node41204;
	wire [4-1:0] node41205;
	wire [4-1:0] node41206;
	wire [4-1:0] node41207;
	wire [4-1:0] node41208;
	wire [4-1:0] node41209;
	wire [4-1:0] node41210;
	wire [4-1:0] node41213;
	wire [4-1:0] node41216;
	wire [4-1:0] node41217;
	wire [4-1:0] node41220;
	wire [4-1:0] node41223;
	wire [4-1:0] node41224;
	wire [4-1:0] node41225;
	wire [4-1:0] node41228;
	wire [4-1:0] node41231;
	wire [4-1:0] node41232;
	wire [4-1:0] node41235;
	wire [4-1:0] node41238;
	wire [4-1:0] node41239;
	wire [4-1:0] node41240;
	wire [4-1:0] node41241;
	wire [4-1:0] node41244;
	wire [4-1:0] node41247;
	wire [4-1:0] node41248;
	wire [4-1:0] node41251;
	wire [4-1:0] node41254;
	wire [4-1:0] node41255;
	wire [4-1:0] node41256;
	wire [4-1:0] node41259;
	wire [4-1:0] node41262;
	wire [4-1:0] node41263;
	wire [4-1:0] node41266;
	wire [4-1:0] node41269;
	wire [4-1:0] node41270;
	wire [4-1:0] node41271;
	wire [4-1:0] node41272;
	wire [4-1:0] node41273;
	wire [4-1:0] node41276;
	wire [4-1:0] node41279;
	wire [4-1:0] node41281;
	wire [4-1:0] node41284;
	wire [4-1:0] node41285;
	wire [4-1:0] node41286;
	wire [4-1:0] node41289;
	wire [4-1:0] node41292;
	wire [4-1:0] node41293;
	wire [4-1:0] node41296;
	wire [4-1:0] node41299;
	wire [4-1:0] node41300;
	wire [4-1:0] node41301;
	wire [4-1:0] node41302;
	wire [4-1:0] node41305;
	wire [4-1:0] node41308;
	wire [4-1:0] node41309;
	wire [4-1:0] node41312;
	wire [4-1:0] node41315;
	wire [4-1:0] node41316;
	wire [4-1:0] node41317;
	wire [4-1:0] node41320;
	wire [4-1:0] node41323;
	wire [4-1:0] node41325;
	wire [4-1:0] node41328;
	wire [4-1:0] node41329;
	wire [4-1:0] node41330;
	wire [4-1:0] node41331;
	wire [4-1:0] node41332;
	wire [4-1:0] node41335;
	wire [4-1:0] node41338;
	wire [4-1:0] node41339;
	wire [4-1:0] node41340;
	wire [4-1:0] node41343;
	wire [4-1:0] node41346;
	wire [4-1:0] node41347;
	wire [4-1:0] node41350;
	wire [4-1:0] node41353;
	wire [4-1:0] node41354;
	wire [4-1:0] node41355;
	wire [4-1:0] node41357;
	wire [4-1:0] node41360;
	wire [4-1:0] node41362;
	wire [4-1:0] node41365;
	wire [4-1:0] node41366;
	wire [4-1:0] node41368;
	wire [4-1:0] node41371;
	wire [4-1:0] node41373;
	wire [4-1:0] node41376;
	wire [4-1:0] node41377;
	wire [4-1:0] node41378;
	wire [4-1:0] node41379;
	wire [4-1:0] node41382;
	wire [4-1:0] node41385;
	wire [4-1:0] node41386;
	wire [4-1:0] node41387;
	wire [4-1:0] node41390;
	wire [4-1:0] node41393;
	wire [4-1:0] node41394;
	wire [4-1:0] node41397;
	wire [4-1:0] node41400;
	wire [4-1:0] node41401;
	wire [4-1:0] node41402;
	wire [4-1:0] node41403;
	wire [4-1:0] node41406;
	wire [4-1:0] node41409;
	wire [4-1:0] node41410;
	wire [4-1:0] node41413;
	wire [4-1:0] node41416;
	wire [4-1:0] node41417;
	wire [4-1:0] node41418;
	wire [4-1:0] node41421;
	wire [4-1:0] node41424;
	wire [4-1:0] node41425;
	wire [4-1:0] node41428;
	wire [4-1:0] node41431;
	wire [4-1:0] node41432;
	wire [4-1:0] node41433;
	wire [4-1:0] node41434;
	wire [4-1:0] node41435;
	wire [4-1:0] node41436;
	wire [4-1:0] node41437;
	wire [4-1:0] node41440;
	wire [4-1:0] node41443;
	wire [4-1:0] node41444;
	wire [4-1:0] node41448;
	wire [4-1:0] node41449;
	wire [4-1:0] node41450;
	wire [4-1:0] node41453;
	wire [4-1:0] node41456;
	wire [4-1:0] node41457;
	wire [4-1:0] node41460;
	wire [4-1:0] node41463;
	wire [4-1:0] node41464;
	wire [4-1:0] node41465;
	wire [4-1:0] node41466;
	wire [4-1:0] node41469;
	wire [4-1:0] node41472;
	wire [4-1:0] node41473;
	wire [4-1:0] node41476;
	wire [4-1:0] node41479;
	wire [4-1:0] node41480;
	wire [4-1:0] node41481;
	wire [4-1:0] node41484;
	wire [4-1:0] node41487;
	wire [4-1:0] node41488;
	wire [4-1:0] node41491;
	wire [4-1:0] node41494;
	wire [4-1:0] node41495;
	wire [4-1:0] node41496;
	wire [4-1:0] node41497;
	wire [4-1:0] node41498;
	wire [4-1:0] node41501;
	wire [4-1:0] node41504;
	wire [4-1:0] node41505;
	wire [4-1:0] node41508;
	wire [4-1:0] node41511;
	wire [4-1:0] node41512;
	wire [4-1:0] node41513;
	wire [4-1:0] node41516;
	wire [4-1:0] node41519;
	wire [4-1:0] node41520;
	wire [4-1:0] node41523;
	wire [4-1:0] node41526;
	wire [4-1:0] node41527;
	wire [4-1:0] node41528;
	wire [4-1:0] node41529;
	wire [4-1:0] node41532;
	wire [4-1:0] node41535;
	wire [4-1:0] node41536;
	wire [4-1:0] node41539;
	wire [4-1:0] node41542;
	wire [4-1:0] node41543;
	wire [4-1:0] node41544;
	wire [4-1:0] node41548;
	wire [4-1:0] node41550;
	wire [4-1:0] node41553;
	wire [4-1:0] node41554;
	wire [4-1:0] node41555;
	wire [4-1:0] node41556;
	wire [4-1:0] node41557;
	wire [4-1:0] node41558;
	wire [4-1:0] node41561;
	wire [4-1:0] node41564;
	wire [4-1:0] node41566;
	wire [4-1:0] node41569;
	wire [4-1:0] node41570;
	wire [4-1:0] node41571;
	wire [4-1:0] node41574;
	wire [4-1:0] node41577;
	wire [4-1:0] node41578;
	wire [4-1:0] node41581;
	wire [4-1:0] node41584;
	wire [4-1:0] node41585;
	wire [4-1:0] node41586;
	wire [4-1:0] node41587;
	wire [4-1:0] node41590;
	wire [4-1:0] node41593;
	wire [4-1:0] node41594;
	wire [4-1:0] node41597;
	wire [4-1:0] node41600;
	wire [4-1:0] node41601;
	wire [4-1:0] node41602;
	wire [4-1:0] node41605;
	wire [4-1:0] node41608;
	wire [4-1:0] node41609;
	wire [4-1:0] node41612;
	wire [4-1:0] node41615;
	wire [4-1:0] node41616;
	wire [4-1:0] node41617;
	wire [4-1:0] node41618;
	wire [4-1:0] node41621;
	wire [4-1:0] node41624;
	wire [4-1:0] node41625;
	wire [4-1:0] node41626;
	wire [4-1:0] node41629;
	wire [4-1:0] node41632;
	wire [4-1:0] node41633;
	wire [4-1:0] node41637;
	wire [4-1:0] node41638;
	wire [4-1:0] node41639;
	wire [4-1:0] node41640;
	wire [4-1:0] node41643;
	wire [4-1:0] node41646;
	wire [4-1:0] node41647;
	wire [4-1:0] node41650;
	wire [4-1:0] node41653;
	wire [4-1:0] node41654;
	wire [4-1:0] node41657;
	wire [4-1:0] node41660;
	wire [4-1:0] node41661;
	wire [4-1:0] node41662;
	wire [4-1:0] node41663;
	wire [4-1:0] node41664;
	wire [4-1:0] node41665;
	wire [4-1:0] node41666;
	wire [4-1:0] node41667;
	wire [4-1:0] node41670;
	wire [4-1:0] node41673;
	wire [4-1:0] node41674;
	wire [4-1:0] node41677;
	wire [4-1:0] node41680;
	wire [4-1:0] node41681;
	wire [4-1:0] node41682;
	wire [4-1:0] node41685;
	wire [4-1:0] node41688;
	wire [4-1:0] node41689;
	wire [4-1:0] node41692;
	wire [4-1:0] node41695;
	wire [4-1:0] node41696;
	wire [4-1:0] node41697;
	wire [4-1:0] node41698;
	wire [4-1:0] node41701;
	wire [4-1:0] node41704;
	wire [4-1:0] node41705;
	wire [4-1:0] node41709;
	wire [4-1:0] node41710;
	wire [4-1:0] node41711;
	wire [4-1:0] node41714;
	wire [4-1:0] node41717;
	wire [4-1:0] node41718;
	wire [4-1:0] node41721;
	wire [4-1:0] node41724;
	wire [4-1:0] node41725;
	wire [4-1:0] node41726;
	wire [4-1:0] node41727;
	wire [4-1:0] node41728;
	wire [4-1:0] node41731;
	wire [4-1:0] node41734;
	wire [4-1:0] node41735;
	wire [4-1:0] node41738;
	wire [4-1:0] node41741;
	wire [4-1:0] node41742;
	wire [4-1:0] node41743;
	wire [4-1:0] node41746;
	wire [4-1:0] node41749;
	wire [4-1:0] node41750;
	wire [4-1:0] node41753;
	wire [4-1:0] node41756;
	wire [4-1:0] node41757;
	wire [4-1:0] node41758;
	wire [4-1:0] node41759;
	wire [4-1:0] node41762;
	wire [4-1:0] node41765;
	wire [4-1:0] node41767;
	wire [4-1:0] node41770;
	wire [4-1:0] node41771;
	wire [4-1:0] node41772;
	wire [4-1:0] node41775;
	wire [4-1:0] node41778;
	wire [4-1:0] node41779;
	wire [4-1:0] node41782;
	wire [4-1:0] node41785;
	wire [4-1:0] node41786;
	wire [4-1:0] node41787;
	wire [4-1:0] node41788;
	wire [4-1:0] node41789;
	wire [4-1:0] node41790;
	wire [4-1:0] node41793;
	wire [4-1:0] node41796;
	wire [4-1:0] node41797;
	wire [4-1:0] node41800;
	wire [4-1:0] node41803;
	wire [4-1:0] node41804;
	wire [4-1:0] node41805;
	wire [4-1:0] node41808;
	wire [4-1:0] node41811;
	wire [4-1:0] node41812;
	wire [4-1:0] node41815;
	wire [4-1:0] node41818;
	wire [4-1:0] node41819;
	wire [4-1:0] node41820;
	wire [4-1:0] node41821;
	wire [4-1:0] node41824;
	wire [4-1:0] node41827;
	wire [4-1:0] node41828;
	wire [4-1:0] node41831;
	wire [4-1:0] node41834;
	wire [4-1:0] node41835;
	wire [4-1:0] node41836;
	wire [4-1:0] node41839;
	wire [4-1:0] node41842;
	wire [4-1:0] node41843;
	wire [4-1:0] node41846;
	wire [4-1:0] node41849;
	wire [4-1:0] node41850;
	wire [4-1:0] node41851;
	wire [4-1:0] node41852;
	wire [4-1:0] node41855;
	wire [4-1:0] node41858;
	wire [4-1:0] node41859;
	wire [4-1:0] node41862;
	wire [4-1:0] node41865;
	wire [4-1:0] node41866;
	wire [4-1:0] node41867;
	wire [4-1:0] node41868;
	wire [4-1:0] node41871;
	wire [4-1:0] node41874;
	wire [4-1:0] node41875;
	wire [4-1:0] node41878;
	wire [4-1:0] node41881;
	wire [4-1:0] node41882;
	wire [4-1:0] node41883;
	wire [4-1:0] node41886;
	wire [4-1:0] node41889;
	wire [4-1:0] node41890;
	wire [4-1:0] node41893;
	wire [4-1:0] node41896;
	wire [4-1:0] node41897;
	wire [4-1:0] node41898;
	wire [4-1:0] node41899;
	wire [4-1:0] node41900;
	wire [4-1:0] node41901;
	wire [4-1:0] node41902;
	wire [4-1:0] node41905;
	wire [4-1:0] node41908;
	wire [4-1:0] node41909;
	wire [4-1:0] node41912;
	wire [4-1:0] node41915;
	wire [4-1:0] node41916;
	wire [4-1:0] node41917;
	wire [4-1:0] node41920;
	wire [4-1:0] node41923;
	wire [4-1:0] node41924;
	wire [4-1:0] node41927;
	wire [4-1:0] node41930;
	wire [4-1:0] node41931;
	wire [4-1:0] node41932;
	wire [4-1:0] node41933;
	wire [4-1:0] node41936;
	wire [4-1:0] node41939;
	wire [4-1:0] node41940;
	wire [4-1:0] node41943;
	wire [4-1:0] node41946;
	wire [4-1:0] node41947;
	wire [4-1:0] node41948;
	wire [4-1:0] node41951;
	wire [4-1:0] node41954;
	wire [4-1:0] node41955;
	wire [4-1:0] node41958;
	wire [4-1:0] node41961;
	wire [4-1:0] node41962;
	wire [4-1:0] node41963;
	wire [4-1:0] node41964;
	wire [4-1:0] node41966;
	wire [4-1:0] node41969;
	wire [4-1:0] node41970;
	wire [4-1:0] node41973;
	wire [4-1:0] node41976;
	wire [4-1:0] node41977;
	wire [4-1:0] node41978;
	wire [4-1:0] node41981;
	wire [4-1:0] node41984;
	wire [4-1:0] node41985;
	wire [4-1:0] node41988;
	wire [4-1:0] node41991;
	wire [4-1:0] node41992;
	wire [4-1:0] node41993;
	wire [4-1:0] node41994;
	wire [4-1:0] node41997;
	wire [4-1:0] node42000;
	wire [4-1:0] node42001;
	wire [4-1:0] node42005;
	wire [4-1:0] node42006;
	wire [4-1:0] node42007;
	wire [4-1:0] node42010;
	wire [4-1:0] node42013;
	wire [4-1:0] node42014;
	wire [4-1:0] node42017;
	wire [4-1:0] node42020;
	wire [4-1:0] node42021;
	wire [4-1:0] node42022;
	wire [4-1:0] node42023;
	wire [4-1:0] node42024;
	wire [4-1:0] node42025;
	wire [4-1:0] node42028;
	wire [4-1:0] node42031;
	wire [4-1:0] node42032;
	wire [4-1:0] node42035;
	wire [4-1:0] node42038;
	wire [4-1:0] node42039;
	wire [4-1:0] node42040;
	wire [4-1:0] node42043;
	wire [4-1:0] node42046;
	wire [4-1:0] node42047;
	wire [4-1:0] node42050;
	wire [4-1:0] node42053;
	wire [4-1:0] node42054;
	wire [4-1:0] node42055;
	wire [4-1:0] node42056;
	wire [4-1:0] node42059;
	wire [4-1:0] node42062;
	wire [4-1:0] node42063;
	wire [4-1:0] node42066;
	wire [4-1:0] node42069;
	wire [4-1:0] node42070;
	wire [4-1:0] node42073;
	wire [4-1:0] node42076;
	wire [4-1:0] node42077;
	wire [4-1:0] node42078;
	wire [4-1:0] node42079;
	wire [4-1:0] node42080;
	wire [4-1:0] node42083;
	wire [4-1:0] node42086;
	wire [4-1:0] node42088;
	wire [4-1:0] node42091;
	wire [4-1:0] node42092;
	wire [4-1:0] node42093;
	wire [4-1:0] node42096;
	wire [4-1:0] node42099;
	wire [4-1:0] node42100;
	wire [4-1:0] node42103;
	wire [4-1:0] node42106;
	wire [4-1:0] node42107;
	wire [4-1:0] node42108;
	wire [4-1:0] node42109;
	wire [4-1:0] node42112;
	wire [4-1:0] node42115;
	wire [4-1:0] node42116;
	wire [4-1:0] node42119;
	wire [4-1:0] node42122;
	wire [4-1:0] node42123;
	wire [4-1:0] node42126;
	wire [4-1:0] node42129;
	wire [4-1:0] node42130;
	wire [4-1:0] node42131;
	wire [4-1:0] node42132;
	wire [4-1:0] node42133;
	wire [4-1:0] node42134;
	wire [4-1:0] node42135;
	wire [4-1:0] node42136;
	wire [4-1:0] node42137;
	wire [4-1:0] node42140;
	wire [4-1:0] node42143;
	wire [4-1:0] node42144;
	wire [4-1:0] node42147;
	wire [4-1:0] node42150;
	wire [4-1:0] node42151;
	wire [4-1:0] node42152;
	wire [4-1:0] node42155;
	wire [4-1:0] node42158;
	wire [4-1:0] node42159;
	wire [4-1:0] node42162;
	wire [4-1:0] node42165;
	wire [4-1:0] node42166;
	wire [4-1:0] node42167;
	wire [4-1:0] node42168;
	wire [4-1:0] node42171;
	wire [4-1:0] node42174;
	wire [4-1:0] node42175;
	wire [4-1:0] node42178;
	wire [4-1:0] node42181;
	wire [4-1:0] node42182;
	wire [4-1:0] node42183;
	wire [4-1:0] node42186;
	wire [4-1:0] node42189;
	wire [4-1:0] node42190;
	wire [4-1:0] node42193;
	wire [4-1:0] node42196;
	wire [4-1:0] node42197;
	wire [4-1:0] node42198;
	wire [4-1:0] node42199;
	wire [4-1:0] node42200;
	wire [4-1:0] node42203;
	wire [4-1:0] node42206;
	wire [4-1:0] node42207;
	wire [4-1:0] node42210;
	wire [4-1:0] node42213;
	wire [4-1:0] node42214;
	wire [4-1:0] node42215;
	wire [4-1:0] node42218;
	wire [4-1:0] node42221;
	wire [4-1:0] node42222;
	wire [4-1:0] node42225;
	wire [4-1:0] node42228;
	wire [4-1:0] node42229;
	wire [4-1:0] node42230;
	wire [4-1:0] node42232;
	wire [4-1:0] node42235;
	wire [4-1:0] node42236;
	wire [4-1:0] node42239;
	wire [4-1:0] node42242;
	wire [4-1:0] node42243;
	wire [4-1:0] node42244;
	wire [4-1:0] node42247;
	wire [4-1:0] node42250;
	wire [4-1:0] node42251;
	wire [4-1:0] node42254;
	wire [4-1:0] node42257;
	wire [4-1:0] node42258;
	wire [4-1:0] node42259;
	wire [4-1:0] node42260;
	wire [4-1:0] node42261;
	wire [4-1:0] node42262;
	wire [4-1:0] node42265;
	wire [4-1:0] node42268;
	wire [4-1:0] node42269;
	wire [4-1:0] node42272;
	wire [4-1:0] node42275;
	wire [4-1:0] node42276;
	wire [4-1:0] node42277;
	wire [4-1:0] node42280;
	wire [4-1:0] node42283;
	wire [4-1:0] node42284;
	wire [4-1:0] node42287;
	wire [4-1:0] node42290;
	wire [4-1:0] node42291;
	wire [4-1:0] node42292;
	wire [4-1:0] node42293;
	wire [4-1:0] node42296;
	wire [4-1:0] node42299;
	wire [4-1:0] node42300;
	wire [4-1:0] node42303;
	wire [4-1:0] node42306;
	wire [4-1:0] node42307;
	wire [4-1:0] node42308;
	wire [4-1:0] node42311;
	wire [4-1:0] node42314;
	wire [4-1:0] node42316;
	wire [4-1:0] node42319;
	wire [4-1:0] node42320;
	wire [4-1:0] node42321;
	wire [4-1:0] node42322;
	wire [4-1:0] node42324;
	wire [4-1:0] node42327;
	wire [4-1:0] node42328;
	wire [4-1:0] node42331;
	wire [4-1:0] node42334;
	wire [4-1:0] node42335;
	wire [4-1:0] node42336;
	wire [4-1:0] node42339;
	wire [4-1:0] node42342;
	wire [4-1:0] node42343;
	wire [4-1:0] node42346;
	wire [4-1:0] node42349;
	wire [4-1:0] node42350;
	wire [4-1:0] node42351;
	wire [4-1:0] node42352;
	wire [4-1:0] node42355;
	wire [4-1:0] node42358;
	wire [4-1:0] node42359;
	wire [4-1:0] node42362;
	wire [4-1:0] node42365;
	wire [4-1:0] node42366;
	wire [4-1:0] node42367;
	wire [4-1:0] node42370;
	wire [4-1:0] node42373;
	wire [4-1:0] node42374;
	wire [4-1:0] node42377;
	wire [4-1:0] node42380;
	wire [4-1:0] node42381;
	wire [4-1:0] node42382;
	wire [4-1:0] node42383;
	wire [4-1:0] node42384;
	wire [4-1:0] node42385;
	wire [4-1:0] node42386;
	wire [4-1:0] node42389;
	wire [4-1:0] node42392;
	wire [4-1:0] node42393;
	wire [4-1:0] node42397;
	wire [4-1:0] node42398;
	wire [4-1:0] node42399;
	wire [4-1:0] node42402;
	wire [4-1:0] node42405;
	wire [4-1:0] node42406;
	wire [4-1:0] node42409;
	wire [4-1:0] node42412;
	wire [4-1:0] node42413;
	wire [4-1:0] node42414;
	wire [4-1:0] node42415;
	wire [4-1:0] node42418;
	wire [4-1:0] node42421;
	wire [4-1:0] node42422;
	wire [4-1:0] node42425;
	wire [4-1:0] node42428;
	wire [4-1:0] node42429;
	wire [4-1:0] node42430;
	wire [4-1:0] node42434;
	wire [4-1:0] node42435;
	wire [4-1:0] node42438;
	wire [4-1:0] node42441;
	wire [4-1:0] node42442;
	wire [4-1:0] node42443;
	wire [4-1:0] node42444;
	wire [4-1:0] node42445;
	wire [4-1:0] node42448;
	wire [4-1:0] node42451;
	wire [4-1:0] node42452;
	wire [4-1:0] node42455;
	wire [4-1:0] node42458;
	wire [4-1:0] node42459;
	wire [4-1:0] node42460;
	wire [4-1:0] node42463;
	wire [4-1:0] node42466;
	wire [4-1:0] node42467;
	wire [4-1:0] node42470;
	wire [4-1:0] node42473;
	wire [4-1:0] node42474;
	wire [4-1:0] node42475;
	wire [4-1:0] node42476;
	wire [4-1:0] node42479;
	wire [4-1:0] node42482;
	wire [4-1:0] node42483;
	wire [4-1:0] node42486;
	wire [4-1:0] node42489;
	wire [4-1:0] node42490;
	wire [4-1:0] node42491;
	wire [4-1:0] node42494;
	wire [4-1:0] node42497;
	wire [4-1:0] node42498;
	wire [4-1:0] node42501;
	wire [4-1:0] node42504;
	wire [4-1:0] node42505;
	wire [4-1:0] node42506;
	wire [4-1:0] node42507;
	wire [4-1:0] node42508;
	wire [4-1:0] node42510;
	wire [4-1:0] node42513;
	wire [4-1:0] node42514;
	wire [4-1:0] node42517;
	wire [4-1:0] node42520;
	wire [4-1:0] node42521;
	wire [4-1:0] node42522;
	wire [4-1:0] node42525;
	wire [4-1:0] node42528;
	wire [4-1:0] node42529;
	wire [4-1:0] node42532;
	wire [4-1:0] node42535;
	wire [4-1:0] node42536;
	wire [4-1:0] node42537;
	wire [4-1:0] node42538;
	wire [4-1:0] node42541;
	wire [4-1:0] node42544;
	wire [4-1:0] node42545;
	wire [4-1:0] node42548;
	wire [4-1:0] node42551;
	wire [4-1:0] node42552;
	wire [4-1:0] node42553;
	wire [4-1:0] node42556;
	wire [4-1:0] node42559;
	wire [4-1:0] node42560;
	wire [4-1:0] node42563;
	wire [4-1:0] node42566;
	wire [4-1:0] node42567;
	wire [4-1:0] node42568;
	wire [4-1:0] node42569;
	wire [4-1:0] node42570;
	wire [4-1:0] node42574;
	wire [4-1:0] node42575;
	wire [4-1:0] node42578;
	wire [4-1:0] node42581;
	wire [4-1:0] node42582;
	wire [4-1:0] node42585;
	wire [4-1:0] node42588;
	wire [4-1:0] node42589;
	wire [4-1:0] node42590;
	wire [4-1:0] node42591;
	wire [4-1:0] node42594;
	wire [4-1:0] node42597;
	wire [4-1:0] node42598;
	wire [4-1:0] node42601;
	wire [4-1:0] node42604;
	wire [4-1:0] node42605;
	wire [4-1:0] node42606;
	wire [4-1:0] node42609;
	wire [4-1:0] node42612;
	wire [4-1:0] node42613;
	wire [4-1:0] node42616;
	wire [4-1:0] node42619;
	wire [4-1:0] node42620;
	wire [4-1:0] node42621;
	wire [4-1:0] node42622;
	wire [4-1:0] node42623;
	wire [4-1:0] node42624;
	wire [4-1:0] node42625;
	wire [4-1:0] node42626;
	wire [4-1:0] node42629;
	wire [4-1:0] node42632;
	wire [4-1:0] node42633;
	wire [4-1:0] node42636;
	wire [4-1:0] node42639;
	wire [4-1:0] node42640;
	wire [4-1:0] node42641;
	wire [4-1:0] node42644;
	wire [4-1:0] node42647;
	wire [4-1:0] node42649;
	wire [4-1:0] node42652;
	wire [4-1:0] node42653;
	wire [4-1:0] node42654;
	wire [4-1:0] node42656;
	wire [4-1:0] node42659;
	wire [4-1:0] node42660;
	wire [4-1:0] node42663;
	wire [4-1:0] node42666;
	wire [4-1:0] node42667;
	wire [4-1:0] node42668;
	wire [4-1:0] node42671;
	wire [4-1:0] node42674;
	wire [4-1:0] node42675;
	wire [4-1:0] node42678;
	wire [4-1:0] node42681;
	wire [4-1:0] node42682;
	wire [4-1:0] node42683;
	wire [4-1:0] node42684;
	wire [4-1:0] node42685;
	wire [4-1:0] node42688;
	wire [4-1:0] node42691;
	wire [4-1:0] node42692;
	wire [4-1:0] node42695;
	wire [4-1:0] node42698;
	wire [4-1:0] node42699;
	wire [4-1:0] node42700;
	wire [4-1:0] node42703;
	wire [4-1:0] node42706;
	wire [4-1:0] node42707;
	wire [4-1:0] node42711;
	wire [4-1:0] node42712;
	wire [4-1:0] node42713;
	wire [4-1:0] node42714;
	wire [4-1:0] node42717;
	wire [4-1:0] node42720;
	wire [4-1:0] node42721;
	wire [4-1:0] node42724;
	wire [4-1:0] node42727;
	wire [4-1:0] node42728;
	wire [4-1:0] node42729;
	wire [4-1:0] node42732;
	wire [4-1:0] node42735;
	wire [4-1:0] node42736;
	wire [4-1:0] node42739;
	wire [4-1:0] node42742;
	wire [4-1:0] node42743;
	wire [4-1:0] node42744;
	wire [4-1:0] node42745;
	wire [4-1:0] node42746;
	wire [4-1:0] node42748;
	wire [4-1:0] node42751;
	wire [4-1:0] node42753;
	wire [4-1:0] node42756;
	wire [4-1:0] node42757;
	wire [4-1:0] node42759;
	wire [4-1:0] node42762;
	wire [4-1:0] node42764;
	wire [4-1:0] node42767;
	wire [4-1:0] node42768;
	wire [4-1:0] node42769;
	wire [4-1:0] node42770;
	wire [4-1:0] node42773;
	wire [4-1:0] node42776;
	wire [4-1:0] node42777;
	wire [4-1:0] node42780;
	wire [4-1:0] node42783;
	wire [4-1:0] node42784;
	wire [4-1:0] node42785;
	wire [4-1:0] node42789;
	wire [4-1:0] node42790;
	wire [4-1:0] node42793;
	wire [4-1:0] node42796;
	wire [4-1:0] node42797;
	wire [4-1:0] node42798;
	wire [4-1:0] node42799;
	wire [4-1:0] node42800;
	wire [4-1:0] node42804;
	wire [4-1:0] node42805;
	wire [4-1:0] node42809;
	wire [4-1:0] node42810;
	wire [4-1:0] node42811;
	wire [4-1:0] node42815;
	wire [4-1:0] node42816;
	wire [4-1:0] node42820;
	wire [4-1:0] node42821;
	wire [4-1:0] node42822;
	wire [4-1:0] node42823;
	wire [4-1:0] node42827;
	wire [4-1:0] node42828;
	wire [4-1:0] node42832;
	wire [4-1:0] node42833;
	wire [4-1:0] node42834;
	wire [4-1:0] node42838;
	wire [4-1:0] node42839;
	wire [4-1:0] node42843;
	wire [4-1:0] node42844;
	wire [4-1:0] node42845;
	wire [4-1:0] node42846;
	wire [4-1:0] node42847;
	wire [4-1:0] node42848;
	wire [4-1:0] node42849;
	wire [4-1:0] node42852;
	wire [4-1:0] node42855;
	wire [4-1:0] node42856;
	wire [4-1:0] node42859;
	wire [4-1:0] node42862;
	wire [4-1:0] node42863;
	wire [4-1:0] node42864;
	wire [4-1:0] node42867;
	wire [4-1:0] node42870;
	wire [4-1:0] node42871;
	wire [4-1:0] node42874;
	wire [4-1:0] node42877;
	wire [4-1:0] node42878;
	wire [4-1:0] node42879;
	wire [4-1:0] node42880;
	wire [4-1:0] node42883;
	wire [4-1:0] node42886;
	wire [4-1:0] node42887;
	wire [4-1:0] node42890;
	wire [4-1:0] node42893;
	wire [4-1:0] node42894;
	wire [4-1:0] node42895;
	wire [4-1:0] node42898;
	wire [4-1:0] node42901;
	wire [4-1:0] node42902;
	wire [4-1:0] node42905;
	wire [4-1:0] node42908;
	wire [4-1:0] node42909;
	wire [4-1:0] node42910;
	wire [4-1:0] node42911;
	wire [4-1:0] node42912;
	wire [4-1:0] node42915;
	wire [4-1:0] node42918;
	wire [4-1:0] node42920;
	wire [4-1:0] node42923;
	wire [4-1:0] node42924;
	wire [4-1:0] node42925;
	wire [4-1:0] node42928;
	wire [4-1:0] node42931;
	wire [4-1:0] node42932;
	wire [4-1:0] node42935;
	wire [4-1:0] node42938;
	wire [4-1:0] node42939;
	wire [4-1:0] node42940;
	wire [4-1:0] node42941;
	wire [4-1:0] node42944;
	wire [4-1:0] node42947;
	wire [4-1:0] node42949;
	wire [4-1:0] node42952;
	wire [4-1:0] node42953;
	wire [4-1:0] node42954;
	wire [4-1:0] node42957;
	wire [4-1:0] node42960;
	wire [4-1:0] node42961;
	wire [4-1:0] node42964;
	wire [4-1:0] node42967;
	wire [4-1:0] node42968;
	wire [4-1:0] node42969;
	wire [4-1:0] node42970;
	wire [4-1:0] node42971;
	wire [4-1:0] node42973;
	wire [4-1:0] node42976;
	wire [4-1:0] node42978;
	wire [4-1:0] node42981;
	wire [4-1:0] node42982;
	wire [4-1:0] node42985;
	wire [4-1:0] node42987;
	wire [4-1:0] node42990;
	wire [4-1:0] node42991;
	wire [4-1:0] node42992;
	wire [4-1:0] node42995;
	wire [4-1:0] node42996;
	wire [4-1:0] node43000;
	wire [4-1:0] node43001;
	wire [4-1:0] node43002;
	wire [4-1:0] node43006;
	wire [4-1:0] node43007;
	wire [4-1:0] node43011;
	wire [4-1:0] node43012;
	wire [4-1:0] node43013;
	wire [4-1:0] node43014;
	wire [4-1:0] node43015;
	wire [4-1:0] node43018;
	wire [4-1:0] node43021;
	wire [4-1:0] node43022;
	wire [4-1:0] node43025;
	wire [4-1:0] node43028;
	wire [4-1:0] node43029;
	wire [4-1:0] node43030;
	wire [4-1:0] node43033;
	wire [4-1:0] node43036;
	wire [4-1:0] node43037;
	wire [4-1:0] node43040;
	wire [4-1:0] node43043;
	wire [4-1:0] node43044;
	wire [4-1:0] node43045;
	wire [4-1:0] node43046;
	wire [4-1:0] node43050;
	wire [4-1:0] node43051;
	wire [4-1:0] node43055;
	wire [4-1:0] node43056;
	wire [4-1:0] node43057;
	wire [4-1:0] node43061;
	wire [4-1:0] node43062;
	wire [4-1:0] node43066;
	wire [4-1:0] node43067;
	wire [4-1:0] node43068;
	wire [4-1:0] node43069;
	wire [4-1:0] node43070;
	wire [4-1:0] node43071;
	wire [4-1:0] node43072;
	wire [4-1:0] node43073;
	wire [4-1:0] node43074;
	wire [4-1:0] node43075;
	wire [4-1:0] node43076;
	wire [4-1:0] node43077;
	wire [4-1:0] node43078;
	wire [4-1:0] node43081;
	wire [4-1:0] node43084;
	wire [4-1:0] node43086;
	wire [4-1:0] node43089;
	wire [4-1:0] node43090;
	wire [4-1:0] node43091;
	wire [4-1:0] node43095;
	wire [4-1:0] node43096;
	wire [4-1:0] node43099;
	wire [4-1:0] node43102;
	wire [4-1:0] node43103;
	wire [4-1:0] node43104;
	wire [4-1:0] node43105;
	wire [4-1:0] node43109;
	wire [4-1:0] node43110;
	wire [4-1:0] node43113;
	wire [4-1:0] node43116;
	wire [4-1:0] node43117;
	wire [4-1:0] node43120;
	wire [4-1:0] node43123;
	wire [4-1:0] node43124;
	wire [4-1:0] node43125;
	wire [4-1:0] node43126;
	wire [4-1:0] node43127;
	wire [4-1:0] node43130;
	wire [4-1:0] node43133;
	wire [4-1:0] node43134;
	wire [4-1:0] node43137;
	wire [4-1:0] node43140;
	wire [4-1:0] node43141;
	wire [4-1:0] node43142;
	wire [4-1:0] node43145;
	wire [4-1:0] node43148;
	wire [4-1:0] node43149;
	wire [4-1:0] node43152;
	wire [4-1:0] node43155;
	wire [4-1:0] node43156;
	wire [4-1:0] node43157;
	wire [4-1:0] node43158;
	wire [4-1:0] node43162;
	wire [4-1:0] node43163;
	wire [4-1:0] node43167;
	wire [4-1:0] node43168;
	wire [4-1:0] node43169;
	wire [4-1:0] node43173;
	wire [4-1:0] node43174;
	wire [4-1:0] node43178;
	wire [4-1:0] node43179;
	wire [4-1:0] node43180;
	wire [4-1:0] node43181;
	wire [4-1:0] node43182;
	wire [4-1:0] node43183;
	wire [4-1:0] node43187;
	wire [4-1:0] node43188;
	wire [4-1:0] node43191;
	wire [4-1:0] node43194;
	wire [4-1:0] node43195;
	wire [4-1:0] node43197;
	wire [4-1:0] node43200;
	wire [4-1:0] node43201;
	wire [4-1:0] node43204;
	wire [4-1:0] node43207;
	wire [4-1:0] node43208;
	wire [4-1:0] node43209;
	wire [4-1:0] node43210;
	wire [4-1:0] node43215;
	wire [4-1:0] node43216;
	wire [4-1:0] node43217;
	wire [4-1:0] node43221;
	wire [4-1:0] node43222;
	wire [4-1:0] node43226;
	wire [4-1:0] node43227;
	wire [4-1:0] node43228;
	wire [4-1:0] node43229;
	wire [4-1:0] node43231;
	wire [4-1:0] node43234;
	wire [4-1:0] node43235;
	wire [4-1:0] node43238;
	wire [4-1:0] node43241;
	wire [4-1:0] node43242;
	wire [4-1:0] node43243;
	wire [4-1:0] node43246;
	wire [4-1:0] node43249;
	wire [4-1:0] node43250;
	wire [4-1:0] node43253;
	wire [4-1:0] node43256;
	wire [4-1:0] node43257;
	wire [4-1:0] node43258;
	wire [4-1:0] node43259;
	wire [4-1:0] node43262;
	wire [4-1:0] node43265;
	wire [4-1:0] node43266;
	wire [4-1:0] node43269;
	wire [4-1:0] node43272;
	wire [4-1:0] node43273;
	wire [4-1:0] node43276;
	wire [4-1:0] node43279;
	wire [4-1:0] node43280;
	wire [4-1:0] node43281;
	wire [4-1:0] node43282;
	wire [4-1:0] node43283;
	wire [4-1:0] node43284;
	wire [4-1:0] node43285;
	wire [4-1:0] node43288;
	wire [4-1:0] node43291;
	wire [4-1:0] node43292;
	wire [4-1:0] node43295;
	wire [4-1:0] node43298;
	wire [4-1:0] node43299;
	wire [4-1:0] node43300;
	wire [4-1:0] node43303;
	wire [4-1:0] node43306;
	wire [4-1:0] node43308;
	wire [4-1:0] node43311;
	wire [4-1:0] node43312;
	wire [4-1:0] node43313;
	wire [4-1:0] node43314;
	wire [4-1:0] node43317;
	wire [4-1:0] node43320;
	wire [4-1:0] node43321;
	wire [4-1:0] node43324;
	wire [4-1:0] node43327;
	wire [4-1:0] node43328;
	wire [4-1:0] node43329;
	wire [4-1:0] node43332;
	wire [4-1:0] node43335;
	wire [4-1:0] node43336;
	wire [4-1:0] node43339;
	wire [4-1:0] node43342;
	wire [4-1:0] node43343;
	wire [4-1:0] node43344;
	wire [4-1:0] node43345;
	wire [4-1:0] node43346;
	wire [4-1:0] node43349;
	wire [4-1:0] node43352;
	wire [4-1:0] node43353;
	wire [4-1:0] node43356;
	wire [4-1:0] node43359;
	wire [4-1:0] node43360;
	wire [4-1:0] node43361;
	wire [4-1:0] node43364;
	wire [4-1:0] node43367;
	wire [4-1:0] node43369;
	wire [4-1:0] node43372;
	wire [4-1:0] node43373;
	wire [4-1:0] node43374;
	wire [4-1:0] node43375;
	wire [4-1:0] node43378;
	wire [4-1:0] node43381;
	wire [4-1:0] node43382;
	wire [4-1:0] node43385;
	wire [4-1:0] node43388;
	wire [4-1:0] node43389;
	wire [4-1:0] node43392;
	wire [4-1:0] node43395;
	wire [4-1:0] node43396;
	wire [4-1:0] node43397;
	wire [4-1:0] node43398;
	wire [4-1:0] node43399;
	wire [4-1:0] node43401;
	wire [4-1:0] node43404;
	wire [4-1:0] node43405;
	wire [4-1:0] node43408;
	wire [4-1:0] node43411;
	wire [4-1:0] node43412;
	wire [4-1:0] node43413;
	wire [4-1:0] node43416;
	wire [4-1:0] node43419;
	wire [4-1:0] node43420;
	wire [4-1:0] node43423;
	wire [4-1:0] node43426;
	wire [4-1:0] node43427;
	wire [4-1:0] node43428;
	wire [4-1:0] node43429;
	wire [4-1:0] node43432;
	wire [4-1:0] node43435;
	wire [4-1:0] node43436;
	wire [4-1:0] node43439;
	wire [4-1:0] node43442;
	wire [4-1:0] node43443;
	wire [4-1:0] node43446;
	wire [4-1:0] node43449;
	wire [4-1:0] node43450;
	wire [4-1:0] node43451;
	wire [4-1:0] node43452;
	wire [4-1:0] node43453;
	wire [4-1:0] node43457;
	wire [4-1:0] node43458;
	wire [4-1:0] node43461;
	wire [4-1:0] node43464;
	wire [4-1:0] node43465;
	wire [4-1:0] node43466;
	wire [4-1:0] node43470;
	wire [4-1:0] node43471;
	wire [4-1:0] node43474;
	wire [4-1:0] node43477;
	wire [4-1:0] node43478;
	wire [4-1:0] node43479;
	wire [4-1:0] node43480;
	wire [4-1:0] node43483;
	wire [4-1:0] node43486;
	wire [4-1:0] node43487;
	wire [4-1:0] node43490;
	wire [4-1:0] node43493;
	wire [4-1:0] node43494;
	wire [4-1:0] node43497;
	wire [4-1:0] node43500;
	wire [4-1:0] node43501;
	wire [4-1:0] node43502;
	wire [4-1:0] node43503;
	wire [4-1:0] node43504;
	wire [4-1:0] node43505;
	wire [4-1:0] node43506;
	wire [4-1:0] node43507;
	wire [4-1:0] node43510;
	wire [4-1:0] node43513;
	wire [4-1:0] node43514;
	wire [4-1:0] node43517;
	wire [4-1:0] node43520;
	wire [4-1:0] node43521;
	wire [4-1:0] node43522;
	wire [4-1:0] node43526;
	wire [4-1:0] node43527;
	wire [4-1:0] node43530;
	wire [4-1:0] node43533;
	wire [4-1:0] node43534;
	wire [4-1:0] node43535;
	wire [4-1:0] node43536;
	wire [4-1:0] node43539;
	wire [4-1:0] node43542;
	wire [4-1:0] node43543;
	wire [4-1:0] node43546;
	wire [4-1:0] node43549;
	wire [4-1:0] node43550;
	wire [4-1:0] node43551;
	wire [4-1:0] node43554;
	wire [4-1:0] node43557;
	wire [4-1:0] node43558;
	wire [4-1:0] node43561;
	wire [4-1:0] node43564;
	wire [4-1:0] node43565;
	wire [4-1:0] node43566;
	wire [4-1:0] node43567;
	wire [4-1:0] node43568;
	wire [4-1:0] node43571;
	wire [4-1:0] node43574;
	wire [4-1:0] node43575;
	wire [4-1:0] node43578;
	wire [4-1:0] node43581;
	wire [4-1:0] node43582;
	wire [4-1:0] node43583;
	wire [4-1:0] node43586;
	wire [4-1:0] node43589;
	wire [4-1:0] node43590;
	wire [4-1:0] node43594;
	wire [4-1:0] node43595;
	wire [4-1:0] node43596;
	wire [4-1:0] node43597;
	wire [4-1:0] node43600;
	wire [4-1:0] node43603;
	wire [4-1:0] node43604;
	wire [4-1:0] node43607;
	wire [4-1:0] node43610;
	wire [4-1:0] node43611;
	wire [4-1:0] node43612;
	wire [4-1:0] node43615;
	wire [4-1:0] node43618;
	wire [4-1:0] node43619;
	wire [4-1:0] node43622;
	wire [4-1:0] node43625;
	wire [4-1:0] node43626;
	wire [4-1:0] node43627;
	wire [4-1:0] node43628;
	wire [4-1:0] node43629;
	wire [4-1:0] node43631;
	wire [4-1:0] node43634;
	wire [4-1:0] node43636;
	wire [4-1:0] node43639;
	wire [4-1:0] node43640;
	wire [4-1:0] node43641;
	wire [4-1:0] node43645;
	wire [4-1:0] node43646;
	wire [4-1:0] node43649;
	wire [4-1:0] node43652;
	wire [4-1:0] node43653;
	wire [4-1:0] node43654;
	wire [4-1:0] node43655;
	wire [4-1:0] node43658;
	wire [4-1:0] node43661;
	wire [4-1:0] node43662;
	wire [4-1:0] node43665;
	wire [4-1:0] node43668;
	wire [4-1:0] node43669;
	wire [4-1:0] node43670;
	wire [4-1:0] node43673;
	wire [4-1:0] node43676;
	wire [4-1:0] node43677;
	wire [4-1:0] node43680;
	wire [4-1:0] node43683;
	wire [4-1:0] node43684;
	wire [4-1:0] node43685;
	wire [4-1:0] node43686;
	wire [4-1:0] node43687;
	wire [4-1:0] node43690;
	wire [4-1:0] node43693;
	wire [4-1:0] node43695;
	wire [4-1:0] node43698;
	wire [4-1:0] node43699;
	wire [4-1:0] node43701;
	wire [4-1:0] node43704;
	wire [4-1:0] node43705;
	wire [4-1:0] node43708;
	wire [4-1:0] node43711;
	wire [4-1:0] node43712;
	wire [4-1:0] node43713;
	wire [4-1:0] node43714;
	wire [4-1:0] node43718;
	wire [4-1:0] node43719;
	wire [4-1:0] node43723;
	wire [4-1:0] node43724;
	wire [4-1:0] node43725;
	wire [4-1:0] node43729;
	wire [4-1:0] node43730;
	wire [4-1:0] node43734;
	wire [4-1:0] node43735;
	wire [4-1:0] node43736;
	wire [4-1:0] node43737;
	wire [4-1:0] node43738;
	wire [4-1:0] node43739;
	wire [4-1:0] node43740;
	wire [4-1:0] node43744;
	wire [4-1:0] node43745;
	wire [4-1:0] node43749;
	wire [4-1:0] node43750;
	wire [4-1:0] node43751;
	wire [4-1:0] node43755;
	wire [4-1:0] node43756;
	wire [4-1:0] node43759;
	wire [4-1:0] node43762;
	wire [4-1:0] node43763;
	wire [4-1:0] node43764;
	wire [4-1:0] node43765;
	wire [4-1:0] node43768;
	wire [4-1:0] node43771;
	wire [4-1:0] node43772;
	wire [4-1:0] node43775;
	wire [4-1:0] node43778;
	wire [4-1:0] node43779;
	wire [4-1:0] node43780;
	wire [4-1:0] node43783;
	wire [4-1:0] node43786;
	wire [4-1:0] node43787;
	wire [4-1:0] node43790;
	wire [4-1:0] node43793;
	wire [4-1:0] node43794;
	wire [4-1:0] node43795;
	wire [4-1:0] node43796;
	wire [4-1:0] node43797;
	wire [4-1:0] node43800;
	wire [4-1:0] node43803;
	wire [4-1:0] node43804;
	wire [4-1:0] node43807;
	wire [4-1:0] node43810;
	wire [4-1:0] node43811;
	wire [4-1:0] node43813;
	wire [4-1:0] node43816;
	wire [4-1:0] node43817;
	wire [4-1:0] node43820;
	wire [4-1:0] node43823;
	wire [4-1:0] node43824;
	wire [4-1:0] node43825;
	wire [4-1:0] node43826;
	wire [4-1:0] node43830;
	wire [4-1:0] node43831;
	wire [4-1:0] node43835;
	wire [4-1:0] node43836;
	wire [4-1:0] node43837;
	wire [4-1:0] node43841;
	wire [4-1:0] node43842;
	wire [4-1:0] node43846;
	wire [4-1:0] node43847;
	wire [4-1:0] node43848;
	wire [4-1:0] node43849;
	wire [4-1:0] node43850;
	wire [4-1:0] node43851;
	wire [4-1:0] node43854;
	wire [4-1:0] node43857;
	wire [4-1:0] node43858;
	wire [4-1:0] node43861;
	wire [4-1:0] node43864;
	wire [4-1:0] node43865;
	wire [4-1:0] node43866;
	wire [4-1:0] node43869;
	wire [4-1:0] node43872;
	wire [4-1:0] node43873;
	wire [4-1:0] node43876;
	wire [4-1:0] node43879;
	wire [4-1:0] node43880;
	wire [4-1:0] node43881;
	wire [4-1:0] node43882;
	wire [4-1:0] node43886;
	wire [4-1:0] node43887;
	wire [4-1:0] node43891;
	wire [4-1:0] node43892;
	wire [4-1:0] node43893;
	wire [4-1:0] node43897;
	wire [4-1:0] node43898;
	wire [4-1:0] node43902;
	wire [4-1:0] node43903;
	wire [4-1:0] node43904;
	wire [4-1:0] node43905;
	wire [4-1:0] node43906;
	wire [4-1:0] node43909;
	wire [4-1:0] node43912;
	wire [4-1:0] node43913;
	wire [4-1:0] node43916;
	wire [4-1:0] node43919;
	wire [4-1:0] node43920;
	wire [4-1:0] node43922;
	wire [4-1:0] node43925;
	wire [4-1:0] node43926;
	wire [4-1:0] node43930;
	wire [4-1:0] node43931;
	wire [4-1:0] node43932;
	wire [4-1:0] node43933;
	wire [4-1:0] node43936;
	wire [4-1:0] node43939;
	wire [4-1:0] node43940;
	wire [4-1:0] node43944;
	wire [4-1:0] node43945;
	wire [4-1:0] node43948;
	wire [4-1:0] node43951;
	wire [4-1:0] node43952;
	wire [4-1:0] node43953;
	wire [4-1:0] node43954;
	wire [4-1:0] node43955;
	wire [4-1:0] node43956;
	wire [4-1:0] node43957;
	wire [4-1:0] node43958;
	wire [4-1:0] node43959;
	wire [4-1:0] node43962;
	wire [4-1:0] node43965;
	wire [4-1:0] node43966;
	wire [4-1:0] node43970;
	wire [4-1:0] node43971;
	wire [4-1:0] node43972;
	wire [4-1:0] node43975;
	wire [4-1:0] node43978;
	wire [4-1:0] node43979;
	wire [4-1:0] node43982;
	wire [4-1:0] node43985;
	wire [4-1:0] node43986;
	wire [4-1:0] node43987;
	wire [4-1:0] node43989;
	wire [4-1:0] node43992;
	wire [4-1:0] node43993;
	wire [4-1:0] node43996;
	wire [4-1:0] node43999;
	wire [4-1:0] node44000;
	wire [4-1:0] node44001;
	wire [4-1:0] node44004;
	wire [4-1:0] node44007;
	wire [4-1:0] node44008;
	wire [4-1:0] node44011;
	wire [4-1:0] node44014;
	wire [4-1:0] node44015;
	wire [4-1:0] node44016;
	wire [4-1:0] node44017;
	wire [4-1:0] node44018;
	wire [4-1:0] node44021;
	wire [4-1:0] node44024;
	wire [4-1:0] node44025;
	wire [4-1:0] node44028;
	wire [4-1:0] node44031;
	wire [4-1:0] node44032;
	wire [4-1:0] node44033;
	wire [4-1:0] node44036;
	wire [4-1:0] node44039;
	wire [4-1:0] node44040;
	wire [4-1:0] node44043;
	wire [4-1:0] node44046;
	wire [4-1:0] node44047;
	wire [4-1:0] node44048;
	wire [4-1:0] node44049;
	wire [4-1:0] node44052;
	wire [4-1:0] node44055;
	wire [4-1:0] node44056;
	wire [4-1:0] node44059;
	wire [4-1:0] node44062;
	wire [4-1:0] node44063;
	wire [4-1:0] node44064;
	wire [4-1:0] node44067;
	wire [4-1:0] node44070;
	wire [4-1:0] node44071;
	wire [4-1:0] node44074;
	wire [4-1:0] node44077;
	wire [4-1:0] node44078;
	wire [4-1:0] node44079;
	wire [4-1:0] node44080;
	wire [4-1:0] node44081;
	wire [4-1:0] node44082;
	wire [4-1:0] node44086;
	wire [4-1:0] node44087;
	wire [4-1:0] node44091;
	wire [4-1:0] node44092;
	wire [4-1:0] node44093;
	wire [4-1:0] node44097;
	wire [4-1:0] node44098;
	wire [4-1:0] node44102;
	wire [4-1:0] node44103;
	wire [4-1:0] node44104;
	wire [4-1:0] node44105;
	wire [4-1:0] node44108;
	wire [4-1:0] node44111;
	wire [4-1:0] node44112;
	wire [4-1:0] node44115;
	wire [4-1:0] node44118;
	wire [4-1:0] node44119;
	wire [4-1:0] node44121;
	wire [4-1:0] node44124;
	wire [4-1:0] node44125;
	wire [4-1:0] node44128;
	wire [4-1:0] node44131;
	wire [4-1:0] node44132;
	wire [4-1:0] node44133;
	wire [4-1:0] node44134;
	wire [4-1:0] node44135;
	wire [4-1:0] node44138;
	wire [4-1:0] node44141;
	wire [4-1:0] node44142;
	wire [4-1:0] node44145;
	wire [4-1:0] node44148;
	wire [4-1:0] node44149;
	wire [4-1:0] node44152;
	wire [4-1:0] node44155;
	wire [4-1:0] node44156;
	wire [4-1:0] node44157;
	wire [4-1:0] node44158;
	wire [4-1:0] node44161;
	wire [4-1:0] node44164;
	wire [4-1:0] node44165;
	wire [4-1:0] node44168;
	wire [4-1:0] node44171;
	wire [4-1:0] node44172;
	wire [4-1:0] node44173;
	wire [4-1:0] node44176;
	wire [4-1:0] node44179;
	wire [4-1:0] node44180;
	wire [4-1:0] node44184;
	wire [4-1:0] node44185;
	wire [4-1:0] node44186;
	wire [4-1:0] node44187;
	wire [4-1:0] node44188;
	wire [4-1:0] node44189;
	wire [4-1:0] node44190;
	wire [4-1:0] node44193;
	wire [4-1:0] node44196;
	wire [4-1:0] node44197;
	wire [4-1:0] node44200;
	wire [4-1:0] node44203;
	wire [4-1:0] node44204;
	wire [4-1:0] node44205;
	wire [4-1:0] node44208;
	wire [4-1:0] node44211;
	wire [4-1:0] node44212;
	wire [4-1:0] node44215;
	wire [4-1:0] node44218;
	wire [4-1:0] node44219;
	wire [4-1:0] node44220;
	wire [4-1:0] node44221;
	wire [4-1:0] node44224;
	wire [4-1:0] node44227;
	wire [4-1:0] node44228;
	wire [4-1:0] node44231;
	wire [4-1:0] node44234;
	wire [4-1:0] node44235;
	wire [4-1:0] node44238;
	wire [4-1:0] node44241;
	wire [4-1:0] node44242;
	wire [4-1:0] node44243;
	wire [4-1:0] node44244;
	wire [4-1:0] node44245;
	wire [4-1:0] node44248;
	wire [4-1:0] node44251;
	wire [4-1:0] node44252;
	wire [4-1:0] node44255;
	wire [4-1:0] node44258;
	wire [4-1:0] node44259;
	wire [4-1:0] node44260;
	wire [4-1:0] node44263;
	wire [4-1:0] node44266;
	wire [4-1:0] node44267;
	wire [4-1:0] node44270;
	wire [4-1:0] node44273;
	wire [4-1:0] node44274;
	wire [4-1:0] node44275;
	wire [4-1:0] node44276;
	wire [4-1:0] node44279;
	wire [4-1:0] node44282;
	wire [4-1:0] node44284;
	wire [4-1:0] node44287;
	wire [4-1:0] node44288;
	wire [4-1:0] node44291;
	wire [4-1:0] node44294;
	wire [4-1:0] node44295;
	wire [4-1:0] node44296;
	wire [4-1:0] node44297;
	wire [4-1:0] node44298;
	wire [4-1:0] node44299;
	wire [4-1:0] node44302;
	wire [4-1:0] node44305;
	wire [4-1:0] node44306;
	wire [4-1:0] node44310;
	wire [4-1:0] node44311;
	wire [4-1:0] node44312;
	wire [4-1:0] node44316;
	wire [4-1:0] node44317;
	wire [4-1:0] node44320;
	wire [4-1:0] node44323;
	wire [4-1:0] node44324;
	wire [4-1:0] node44325;
	wire [4-1:0] node44326;
	wire [4-1:0] node44329;
	wire [4-1:0] node44332;
	wire [4-1:0] node44334;
	wire [4-1:0] node44337;
	wire [4-1:0] node44338;
	wire [4-1:0] node44339;
	wire [4-1:0] node44342;
	wire [4-1:0] node44345;
	wire [4-1:0] node44346;
	wire [4-1:0] node44349;
	wire [4-1:0] node44352;
	wire [4-1:0] node44353;
	wire [4-1:0] node44354;
	wire [4-1:0] node44355;
	wire [4-1:0] node44358;
	wire [4-1:0] node44359;
	wire [4-1:0] node44362;
	wire [4-1:0] node44365;
	wire [4-1:0] node44366;
	wire [4-1:0] node44367;
	wire [4-1:0] node44370;
	wire [4-1:0] node44373;
	wire [4-1:0] node44374;
	wire [4-1:0] node44378;
	wire [4-1:0] node44379;
	wire [4-1:0] node44380;
	wire [4-1:0] node44381;
	wire [4-1:0] node44384;
	wire [4-1:0] node44387;
	wire [4-1:0] node44388;
	wire [4-1:0] node44391;
	wire [4-1:0] node44394;
	wire [4-1:0] node44395;
	wire [4-1:0] node44398;
	wire [4-1:0] node44401;
	wire [4-1:0] node44402;
	wire [4-1:0] node44403;
	wire [4-1:0] node44404;
	wire [4-1:0] node44405;
	wire [4-1:0] node44406;
	wire [4-1:0] node44407;
	wire [4-1:0] node44408;
	wire [4-1:0] node44411;
	wire [4-1:0] node44414;
	wire [4-1:0] node44415;
	wire [4-1:0] node44418;
	wire [4-1:0] node44421;
	wire [4-1:0] node44422;
	wire [4-1:0] node44423;
	wire [4-1:0] node44426;
	wire [4-1:0] node44429;
	wire [4-1:0] node44430;
	wire [4-1:0] node44433;
	wire [4-1:0] node44436;
	wire [4-1:0] node44437;
	wire [4-1:0] node44438;
	wire [4-1:0] node44439;
	wire [4-1:0] node44442;
	wire [4-1:0] node44445;
	wire [4-1:0] node44446;
	wire [4-1:0] node44449;
	wire [4-1:0] node44452;
	wire [4-1:0] node44453;
	wire [4-1:0] node44456;
	wire [4-1:0] node44459;
	wire [4-1:0] node44460;
	wire [4-1:0] node44461;
	wire [4-1:0] node44462;
	wire [4-1:0] node44463;
	wire [4-1:0] node44467;
	wire [4-1:0] node44468;
	wire [4-1:0] node44471;
	wire [4-1:0] node44474;
	wire [4-1:0] node44475;
	wire [4-1:0] node44476;
	wire [4-1:0] node44479;
	wire [4-1:0] node44482;
	wire [4-1:0] node44483;
	wire [4-1:0] node44486;
	wire [4-1:0] node44489;
	wire [4-1:0] node44490;
	wire [4-1:0] node44491;
	wire [4-1:0] node44492;
	wire [4-1:0] node44496;
	wire [4-1:0] node44497;
	wire [4-1:0] node44501;
	wire [4-1:0] node44502;
	wire [4-1:0] node44503;
	wire [4-1:0] node44507;
	wire [4-1:0] node44508;
	wire [4-1:0] node44512;
	wire [4-1:0] node44513;
	wire [4-1:0] node44514;
	wire [4-1:0] node44515;
	wire [4-1:0] node44516;
	wire [4-1:0] node44518;
	wire [4-1:0] node44521;
	wire [4-1:0] node44522;
	wire [4-1:0] node44525;
	wire [4-1:0] node44528;
	wire [4-1:0] node44529;
	wire [4-1:0] node44530;
	wire [4-1:0] node44533;
	wire [4-1:0] node44536;
	wire [4-1:0] node44537;
	wire [4-1:0] node44540;
	wire [4-1:0] node44543;
	wire [4-1:0] node44544;
	wire [4-1:0] node44545;
	wire [4-1:0] node44546;
	wire [4-1:0] node44550;
	wire [4-1:0] node44551;
	wire [4-1:0] node44555;
	wire [4-1:0] node44556;
	wire [4-1:0] node44557;
	wire [4-1:0] node44561;
	wire [4-1:0] node44562;
	wire [4-1:0] node44566;
	wire [4-1:0] node44567;
	wire [4-1:0] node44568;
	wire [4-1:0] node44569;
	wire [4-1:0] node44570;
	wire [4-1:0] node44573;
	wire [4-1:0] node44576;
	wire [4-1:0] node44577;
	wire [4-1:0] node44580;
	wire [4-1:0] node44583;
	wire [4-1:0] node44584;
	wire [4-1:0] node44585;
	wire [4-1:0] node44588;
	wire [4-1:0] node44591;
	wire [4-1:0] node44592;
	wire [4-1:0] node44595;
	wire [4-1:0] node44598;
	wire [4-1:0] node44599;
	wire [4-1:0] node44600;
	wire [4-1:0] node44601;
	wire [4-1:0] node44604;
	wire [4-1:0] node44607;
	wire [4-1:0] node44608;
	wire [4-1:0] node44611;
	wire [4-1:0] node44614;
	wire [4-1:0] node44615;
	wire [4-1:0] node44618;
	wire [4-1:0] node44621;
	wire [4-1:0] node44622;
	wire [4-1:0] node44623;
	wire [4-1:0] node44624;
	wire [4-1:0] node44625;
	wire [4-1:0] node44626;
	wire [4-1:0] node44627;
	wire [4-1:0] node44630;
	wire [4-1:0] node44633;
	wire [4-1:0] node44634;
	wire [4-1:0] node44638;
	wire [4-1:0] node44639;
	wire [4-1:0] node44640;
	wire [4-1:0] node44643;
	wire [4-1:0] node44646;
	wire [4-1:0] node44647;
	wire [4-1:0] node44650;
	wire [4-1:0] node44653;
	wire [4-1:0] node44654;
	wire [4-1:0] node44655;
	wire [4-1:0] node44656;
	wire [4-1:0] node44659;
	wire [4-1:0] node44662;
	wire [4-1:0] node44663;
	wire [4-1:0] node44666;
	wire [4-1:0] node44669;
	wire [4-1:0] node44670;
	wire [4-1:0] node44671;
	wire [4-1:0] node44674;
	wire [4-1:0] node44677;
	wire [4-1:0] node44678;
	wire [4-1:0] node44681;
	wire [4-1:0] node44684;
	wire [4-1:0] node44685;
	wire [4-1:0] node44686;
	wire [4-1:0] node44687;
	wire [4-1:0] node44688;
	wire [4-1:0] node44691;
	wire [4-1:0] node44694;
	wire [4-1:0] node44695;
	wire [4-1:0] node44698;
	wire [4-1:0] node44701;
	wire [4-1:0] node44702;
	wire [4-1:0] node44703;
	wire [4-1:0] node44706;
	wire [4-1:0] node44709;
	wire [4-1:0] node44710;
	wire [4-1:0] node44713;
	wire [4-1:0] node44716;
	wire [4-1:0] node44717;
	wire [4-1:0] node44718;
	wire [4-1:0] node44719;
	wire [4-1:0] node44723;
	wire [4-1:0] node44724;
	wire [4-1:0] node44728;
	wire [4-1:0] node44729;
	wire [4-1:0] node44730;
	wire [4-1:0] node44734;
	wire [4-1:0] node44735;
	wire [4-1:0] node44739;
	wire [4-1:0] node44740;
	wire [4-1:0] node44741;
	wire [4-1:0] node44742;
	wire [4-1:0] node44743;
	wire [4-1:0] node44744;
	wire [4-1:0] node44748;
	wire [4-1:0] node44749;
	wire [4-1:0] node44752;
	wire [4-1:0] node44755;
	wire [4-1:0] node44756;
	wire [4-1:0] node44757;
	wire [4-1:0] node44760;
	wire [4-1:0] node44763;
	wire [4-1:0] node44764;
	wire [4-1:0] node44768;
	wire [4-1:0] node44769;
	wire [4-1:0] node44770;
	wire [4-1:0] node44771;
	wire [4-1:0] node44774;
	wire [4-1:0] node44777;
	wire [4-1:0] node44778;
	wire [4-1:0] node44781;
	wire [4-1:0] node44784;
	wire [4-1:0] node44785;
	wire [4-1:0] node44786;
	wire [4-1:0] node44789;
	wire [4-1:0] node44792;
	wire [4-1:0] node44793;
	wire [4-1:0] node44796;
	wire [4-1:0] node44799;
	wire [4-1:0] node44800;
	wire [4-1:0] node44801;
	wire [4-1:0] node44802;
	wire [4-1:0] node44804;
	wire [4-1:0] node44807;
	wire [4-1:0] node44808;
	wire [4-1:0] node44812;
	wire [4-1:0] node44813;
	wire [4-1:0] node44814;
	wire [4-1:0] node44817;
	wire [4-1:0] node44820;
	wire [4-1:0] node44821;
	wire [4-1:0] node44824;
	wire [4-1:0] node44827;
	wire [4-1:0] node44828;
	wire [4-1:0] node44829;
	wire [4-1:0] node44830;
	wire [4-1:0] node44833;
	wire [4-1:0] node44836;
	wire [4-1:0] node44837;
	wire [4-1:0] node44840;
	wire [4-1:0] node44843;
	wire [4-1:0] node44844;
	wire [4-1:0] node44847;
	wire [4-1:0] node44850;
	wire [4-1:0] node44851;
	wire [4-1:0] node44852;
	wire [4-1:0] node44853;
	wire [4-1:0] node44854;
	wire [4-1:0] node44855;
	wire [4-1:0] node44856;
	wire [4-1:0] node44857;
	wire [4-1:0] node44858;
	wire [4-1:0] node44859;
	wire [4-1:0] node44862;
	wire [4-1:0] node44865;
	wire [4-1:0] node44866;
	wire [4-1:0] node44869;
	wire [4-1:0] node44872;
	wire [4-1:0] node44873;
	wire [4-1:0] node44874;
	wire [4-1:0] node44877;
	wire [4-1:0] node44880;
	wire [4-1:0] node44881;
	wire [4-1:0] node44884;
	wire [4-1:0] node44887;
	wire [4-1:0] node44888;
	wire [4-1:0] node44889;
	wire [4-1:0] node44890;
	wire [4-1:0] node44893;
	wire [4-1:0] node44896;
	wire [4-1:0] node44897;
	wire [4-1:0] node44900;
	wire [4-1:0] node44903;
	wire [4-1:0] node44904;
	wire [4-1:0] node44905;
	wire [4-1:0] node44908;
	wire [4-1:0] node44911;
	wire [4-1:0] node44912;
	wire [4-1:0] node44915;
	wire [4-1:0] node44918;
	wire [4-1:0] node44919;
	wire [4-1:0] node44920;
	wire [4-1:0] node44921;
	wire [4-1:0] node44922;
	wire [4-1:0] node44925;
	wire [4-1:0] node44928;
	wire [4-1:0] node44930;
	wire [4-1:0] node44933;
	wire [4-1:0] node44934;
	wire [4-1:0] node44935;
	wire [4-1:0] node44939;
	wire [4-1:0] node44940;
	wire [4-1:0] node44944;
	wire [4-1:0] node44945;
	wire [4-1:0] node44946;
	wire [4-1:0] node44947;
	wire [4-1:0] node44950;
	wire [4-1:0] node44954;
	wire [4-1:0] node44955;
	wire [4-1:0] node44956;
	wire [4-1:0] node44959;
	wire [4-1:0] node44962;
	wire [4-1:0] node44963;
	wire [4-1:0] node44966;
	wire [4-1:0] node44969;
	wire [4-1:0] node44970;
	wire [4-1:0] node44971;
	wire [4-1:0] node44972;
	wire [4-1:0] node44973;
	wire [4-1:0] node44974;
	wire [4-1:0] node44978;
	wire [4-1:0] node44979;
	wire [4-1:0] node44983;
	wire [4-1:0] node44984;
	wire [4-1:0] node44985;
	wire [4-1:0] node44989;
	wire [4-1:0] node44990;
	wire [4-1:0] node44994;
	wire [4-1:0] node44995;
	wire [4-1:0] node44996;
	wire [4-1:0] node44997;
	wire [4-1:0] node45001;
	wire [4-1:0] node45002;
	wire [4-1:0] node45006;
	wire [4-1:0] node45007;
	wire [4-1:0] node45008;
	wire [4-1:0] node45012;
	wire [4-1:0] node45013;
	wire [4-1:0] node45017;
	wire [4-1:0] node45018;
	wire [4-1:0] node45019;
	wire [4-1:0] node45020;
	wire [4-1:0] node45022;
	wire [4-1:0] node45025;
	wire [4-1:0] node45026;
	wire [4-1:0] node45029;
	wire [4-1:0] node45032;
	wire [4-1:0] node45033;
	wire [4-1:0] node45034;
	wire [4-1:0] node45037;
	wire [4-1:0] node45040;
	wire [4-1:0] node45041;
	wire [4-1:0] node45044;
	wire [4-1:0] node45047;
	wire [4-1:0] node45048;
	wire [4-1:0] node45049;
	wire [4-1:0] node45050;
	wire [4-1:0] node45053;
	wire [4-1:0] node45056;
	wire [4-1:0] node45057;
	wire [4-1:0] node45060;
	wire [4-1:0] node45063;
	wire [4-1:0] node45064;
	wire [4-1:0] node45067;
	wire [4-1:0] node45070;
	wire [4-1:0] node45071;
	wire [4-1:0] node45072;
	wire [4-1:0] node45073;
	wire [4-1:0] node45074;
	wire [4-1:0] node45075;
	wire [4-1:0] node45076;
	wire [4-1:0] node45079;
	wire [4-1:0] node45082;
	wire [4-1:0] node45083;
	wire [4-1:0] node45086;
	wire [4-1:0] node45089;
	wire [4-1:0] node45090;
	wire [4-1:0] node45091;
	wire [4-1:0] node45094;
	wire [4-1:0] node45097;
	wire [4-1:0] node45098;
	wire [4-1:0] node45101;
	wire [4-1:0] node45104;
	wire [4-1:0] node45105;
	wire [4-1:0] node45106;
	wire [4-1:0] node45107;
	wire [4-1:0] node45111;
	wire [4-1:0] node45112;
	wire [4-1:0] node45116;
	wire [4-1:0] node45117;
	wire [4-1:0] node45118;
	wire [4-1:0] node45122;
	wire [4-1:0] node45123;
	wire [4-1:0] node45127;
	wire [4-1:0] node45128;
	wire [4-1:0] node45129;
	wire [4-1:0] node45130;
	wire [4-1:0] node45131;
	wire [4-1:0] node45134;
	wire [4-1:0] node45137;
	wire [4-1:0] node45138;
	wire [4-1:0] node45141;
	wire [4-1:0] node45144;
	wire [4-1:0] node45145;
	wire [4-1:0] node45147;
	wire [4-1:0] node45150;
	wire [4-1:0] node45151;
	wire [4-1:0] node45154;
	wire [4-1:0] node45157;
	wire [4-1:0] node45158;
	wire [4-1:0] node45159;
	wire [4-1:0] node45160;
	wire [4-1:0] node45164;
	wire [4-1:0] node45165;
	wire [4-1:0] node45169;
	wire [4-1:0] node45170;
	wire [4-1:0] node45171;
	wire [4-1:0] node45175;
	wire [4-1:0] node45176;
	wire [4-1:0] node45180;
	wire [4-1:0] node45181;
	wire [4-1:0] node45182;
	wire [4-1:0] node45183;
	wire [4-1:0] node45184;
	wire [4-1:0] node45185;
	wire [4-1:0] node45188;
	wire [4-1:0] node45191;
	wire [4-1:0] node45192;
	wire [4-1:0] node45195;
	wire [4-1:0] node45198;
	wire [4-1:0] node45199;
	wire [4-1:0] node45200;
	wire [4-1:0] node45203;
	wire [4-1:0] node45206;
	wire [4-1:0] node45207;
	wire [4-1:0] node45210;
	wire [4-1:0] node45213;
	wire [4-1:0] node45214;
	wire [4-1:0] node45215;
	wire [4-1:0] node45216;
	wire [4-1:0] node45219;
	wire [4-1:0] node45222;
	wire [4-1:0] node45223;
	wire [4-1:0] node45226;
	wire [4-1:0] node45229;
	wire [4-1:0] node45230;
	wire [4-1:0] node45233;
	wire [4-1:0] node45236;
	wire [4-1:0] node45237;
	wire [4-1:0] node45238;
	wire [4-1:0] node45239;
	wire [4-1:0] node45240;
	wire [4-1:0] node45243;
	wire [4-1:0] node45246;
	wire [4-1:0] node45247;
	wire [4-1:0] node45250;
	wire [4-1:0] node45253;
	wire [4-1:0] node45254;
	wire [4-1:0] node45256;
	wire [4-1:0] node45259;
	wire [4-1:0] node45260;
	wire [4-1:0] node45263;
	wire [4-1:0] node45266;
	wire [4-1:0] node45267;
	wire [4-1:0] node45268;
	wire [4-1:0] node45269;
	wire [4-1:0] node45272;
	wire [4-1:0] node45275;
	wire [4-1:0] node45276;
	wire [4-1:0] node45279;
	wire [4-1:0] node45282;
	wire [4-1:0] node45283;
	wire [4-1:0] node45284;
	wire [4-1:0] node45287;
	wire [4-1:0] node45290;
	wire [4-1:0] node45291;
	wire [4-1:0] node45294;
	wire [4-1:0] node45297;
	wire [4-1:0] node45298;
	wire [4-1:0] node45299;
	wire [4-1:0] node45300;
	wire [4-1:0] node45301;
	wire [4-1:0] node45302;
	wire [4-1:0] node45303;
	wire [4-1:0] node45304;
	wire [4-1:0] node45307;
	wire [4-1:0] node45310;
	wire [4-1:0] node45311;
	wire [4-1:0] node45314;
	wire [4-1:0] node45317;
	wire [4-1:0] node45318;
	wire [4-1:0] node45319;
	wire [4-1:0] node45322;
	wire [4-1:0] node45325;
	wire [4-1:0] node45327;
	wire [4-1:0] node45330;
	wire [4-1:0] node45331;
	wire [4-1:0] node45332;
	wire [4-1:0] node45333;
	wire [4-1:0] node45337;
	wire [4-1:0] node45338;
	wire [4-1:0] node45342;
	wire [4-1:0] node45343;
	wire [4-1:0] node45344;
	wire [4-1:0] node45348;
	wire [4-1:0] node45349;
	wire [4-1:0] node45353;
	wire [4-1:0] node45354;
	wire [4-1:0] node45355;
	wire [4-1:0] node45356;
	wire [4-1:0] node45357;
	wire [4-1:0] node45360;
	wire [4-1:0] node45363;
	wire [4-1:0] node45364;
	wire [4-1:0] node45367;
	wire [4-1:0] node45370;
	wire [4-1:0] node45371;
	wire [4-1:0] node45372;
	wire [4-1:0] node45375;
	wire [4-1:0] node45378;
	wire [4-1:0] node45379;
	wire [4-1:0] node45382;
	wire [4-1:0] node45385;
	wire [4-1:0] node45386;
	wire [4-1:0] node45387;
	wire [4-1:0] node45388;
	wire [4-1:0] node45391;
	wire [4-1:0] node45394;
	wire [4-1:0] node45395;
	wire [4-1:0] node45399;
	wire [4-1:0] node45400;
	wire [4-1:0] node45401;
	wire [4-1:0] node45404;
	wire [4-1:0] node45407;
	wire [4-1:0] node45408;
	wire [4-1:0] node45411;
	wire [4-1:0] node45414;
	wire [4-1:0] node45415;
	wire [4-1:0] node45416;
	wire [4-1:0] node45417;
	wire [4-1:0] node45418;
	wire [4-1:0] node45419;
	wire [4-1:0] node45422;
	wire [4-1:0] node45425;
	wire [4-1:0] node45427;
	wire [4-1:0] node45430;
	wire [4-1:0] node45431;
	wire [4-1:0] node45432;
	wire [4-1:0] node45435;
	wire [4-1:0] node45438;
	wire [4-1:0] node45440;
	wire [4-1:0] node45443;
	wire [4-1:0] node45444;
	wire [4-1:0] node45445;
	wire [4-1:0] node45446;
	wire [4-1:0] node45449;
	wire [4-1:0] node45452;
	wire [4-1:0] node45453;
	wire [4-1:0] node45456;
	wire [4-1:0] node45459;
	wire [4-1:0] node45460;
	wire [4-1:0] node45461;
	wire [4-1:0] node45464;
	wire [4-1:0] node45467;
	wire [4-1:0] node45468;
	wire [4-1:0] node45471;
	wire [4-1:0] node45474;
	wire [4-1:0] node45475;
	wire [4-1:0] node45476;
	wire [4-1:0] node45477;
	wire [4-1:0] node45478;
	wire [4-1:0] node45481;
	wire [4-1:0] node45484;
	wire [4-1:0] node45485;
	wire [4-1:0] node45488;
	wire [4-1:0] node45491;
	wire [4-1:0] node45492;
	wire [4-1:0] node45493;
	wire [4-1:0] node45496;
	wire [4-1:0] node45499;
	wire [4-1:0] node45500;
	wire [4-1:0] node45503;
	wire [4-1:0] node45506;
	wire [4-1:0] node45507;
	wire [4-1:0] node45508;
	wire [4-1:0] node45509;
	wire [4-1:0] node45513;
	wire [4-1:0] node45514;
	wire [4-1:0] node45518;
	wire [4-1:0] node45519;
	wire [4-1:0] node45520;
	wire [4-1:0] node45524;
	wire [4-1:0] node45525;
	wire [4-1:0] node45529;
	wire [4-1:0] node45530;
	wire [4-1:0] node45531;
	wire [4-1:0] node45532;
	wire [4-1:0] node45533;
	wire [4-1:0] node45534;
	wire [4-1:0] node45535;
	wire [4-1:0] node45538;
	wire [4-1:0] node45541;
	wire [4-1:0] node45542;
	wire [4-1:0] node45545;
	wire [4-1:0] node45548;
	wire [4-1:0] node45549;
	wire [4-1:0] node45550;
	wire [4-1:0] node45553;
	wire [4-1:0] node45556;
	wire [4-1:0] node45557;
	wire [4-1:0] node45560;
	wire [4-1:0] node45563;
	wire [4-1:0] node45564;
	wire [4-1:0] node45565;
	wire [4-1:0] node45567;
	wire [4-1:0] node45570;
	wire [4-1:0] node45571;
	wire [4-1:0] node45574;
	wire [4-1:0] node45577;
	wire [4-1:0] node45578;
	wire [4-1:0] node45579;
	wire [4-1:0] node45582;
	wire [4-1:0] node45585;
	wire [4-1:0] node45586;
	wire [4-1:0] node45589;
	wire [4-1:0] node45592;
	wire [4-1:0] node45593;
	wire [4-1:0] node45594;
	wire [4-1:0] node45595;
	wire [4-1:0] node45596;
	wire [4-1:0] node45599;
	wire [4-1:0] node45602;
	wire [4-1:0] node45603;
	wire [4-1:0] node45606;
	wire [4-1:0] node45609;
	wire [4-1:0] node45610;
	wire [4-1:0] node45611;
	wire [4-1:0] node45614;
	wire [4-1:0] node45617;
	wire [4-1:0] node45618;
	wire [4-1:0] node45622;
	wire [4-1:0] node45623;
	wire [4-1:0] node45624;
	wire [4-1:0] node45625;
	wire [4-1:0] node45628;
	wire [4-1:0] node45631;
	wire [4-1:0] node45632;
	wire [4-1:0] node45635;
	wire [4-1:0] node45638;
	wire [4-1:0] node45639;
	wire [4-1:0] node45640;
	wire [4-1:0] node45643;
	wire [4-1:0] node45646;
	wire [4-1:0] node45647;
	wire [4-1:0] node45650;
	wire [4-1:0] node45653;
	wire [4-1:0] node45654;
	wire [4-1:0] node45655;
	wire [4-1:0] node45656;
	wire [4-1:0] node45657;
	wire [4-1:0] node45658;
	wire [4-1:0] node45661;
	wire [4-1:0] node45664;
	wire [4-1:0] node45665;
	wire [4-1:0] node45668;
	wire [4-1:0] node45671;
	wire [4-1:0] node45672;
	wire [4-1:0] node45673;
	wire [4-1:0] node45676;
	wire [4-1:0] node45679;
	wire [4-1:0] node45680;
	wire [4-1:0] node45683;
	wire [4-1:0] node45686;
	wire [4-1:0] node45687;
	wire [4-1:0] node45688;
	wire [4-1:0] node45690;
	wire [4-1:0] node45693;
	wire [4-1:0] node45694;
	wire [4-1:0] node45697;
	wire [4-1:0] node45700;
	wire [4-1:0] node45701;
	wire [4-1:0] node45702;
	wire [4-1:0] node45705;
	wire [4-1:0] node45708;
	wire [4-1:0] node45709;
	wire [4-1:0] node45712;
	wire [4-1:0] node45715;
	wire [4-1:0] node45716;
	wire [4-1:0] node45717;
	wire [4-1:0] node45718;
	wire [4-1:0] node45719;
	wire [4-1:0] node45722;
	wire [4-1:0] node45725;
	wire [4-1:0] node45726;
	wire [4-1:0] node45729;
	wire [4-1:0] node45732;
	wire [4-1:0] node45733;
	wire [4-1:0] node45734;
	wire [4-1:0] node45737;
	wire [4-1:0] node45740;
	wire [4-1:0] node45741;
	wire [4-1:0] node45744;
	wire [4-1:0] node45747;
	wire [4-1:0] node45748;
	wire [4-1:0] node45749;
	wire [4-1:0] node45750;
	wire [4-1:0] node45753;
	wire [4-1:0] node45756;
	wire [4-1:0] node45757;
	wire [4-1:0] node45760;
	wire [4-1:0] node45763;
	wire [4-1:0] node45764;
	wire [4-1:0] node45765;
	wire [4-1:0] node45768;
	wire [4-1:0] node45771;
	wire [4-1:0] node45772;
	wire [4-1:0] node45775;
	wire [4-1:0] node45778;
	wire [4-1:0] node45779;
	wire [4-1:0] node45780;
	wire [4-1:0] node45781;
	wire [4-1:0] node45782;
	wire [4-1:0] node45783;
	wire [4-1:0] node45784;
	wire [4-1:0] node45785;
	wire [4-1:0] node45786;
	wire [4-1:0] node45789;
	wire [4-1:0] node45792;
	wire [4-1:0] node45793;
	wire [4-1:0] node45796;
	wire [4-1:0] node45799;
	wire [4-1:0] node45800;
	wire [4-1:0] node45803;
	wire [4-1:0] node45804;
	wire [4-1:0] node45807;
	wire [4-1:0] node45810;
	wire [4-1:0] node45811;
	wire [4-1:0] node45812;
	wire [4-1:0] node45813;
	wire [4-1:0] node45816;
	wire [4-1:0] node45819;
	wire [4-1:0] node45820;
	wire [4-1:0] node45823;
	wire [4-1:0] node45826;
	wire [4-1:0] node45827;
	wire [4-1:0] node45830;
	wire [4-1:0] node45833;
	wire [4-1:0] node45834;
	wire [4-1:0] node45835;
	wire [4-1:0] node45836;
	wire [4-1:0] node45838;
	wire [4-1:0] node45841;
	wire [4-1:0] node45843;
	wire [4-1:0] node45846;
	wire [4-1:0] node45847;
	wire [4-1:0] node45848;
	wire [4-1:0] node45851;
	wire [4-1:0] node45854;
	wire [4-1:0] node45855;
	wire [4-1:0] node45858;
	wire [4-1:0] node45861;
	wire [4-1:0] node45862;
	wire [4-1:0] node45863;
	wire [4-1:0] node45864;
	wire [4-1:0] node45868;
	wire [4-1:0] node45869;
	wire [4-1:0] node45873;
	wire [4-1:0] node45874;
	wire [4-1:0] node45875;
	wire [4-1:0] node45879;
	wire [4-1:0] node45880;
	wire [4-1:0] node45884;
	wire [4-1:0] node45885;
	wire [4-1:0] node45886;
	wire [4-1:0] node45887;
	wire [4-1:0] node45888;
	wire [4-1:0] node45889;
	wire [4-1:0] node45892;
	wire [4-1:0] node45895;
	wire [4-1:0] node45896;
	wire [4-1:0] node45899;
	wire [4-1:0] node45902;
	wire [4-1:0] node45903;
	wire [4-1:0] node45904;
	wire [4-1:0] node45907;
	wire [4-1:0] node45910;
	wire [4-1:0] node45911;
	wire [4-1:0] node45915;
	wire [4-1:0] node45916;
	wire [4-1:0] node45917;
	wire [4-1:0] node45918;
	wire [4-1:0] node45922;
	wire [4-1:0] node45923;
	wire [4-1:0] node45927;
	wire [4-1:0] node45928;
	wire [4-1:0] node45929;
	wire [4-1:0] node45933;
	wire [4-1:0] node45934;
	wire [4-1:0] node45938;
	wire [4-1:0] node45939;
	wire [4-1:0] node45940;
	wire [4-1:0] node45941;
	wire [4-1:0] node45942;
	wire [4-1:0] node45945;
	wire [4-1:0] node45948;
	wire [4-1:0] node45949;
	wire [4-1:0] node45953;
	wire [4-1:0] node45954;
	wire [4-1:0] node45955;
	wire [4-1:0] node45958;
	wire [4-1:0] node45961;
	wire [4-1:0] node45962;
	wire [4-1:0] node45965;
	wire [4-1:0] node45968;
	wire [4-1:0] node45969;
	wire [4-1:0] node45970;
	wire [4-1:0] node45971;
	wire [4-1:0] node45974;
	wire [4-1:0] node45977;
	wire [4-1:0] node45978;
	wire [4-1:0] node45981;
	wire [4-1:0] node45984;
	wire [4-1:0] node45985;
	wire [4-1:0] node45987;
	wire [4-1:0] node45990;
	wire [4-1:0] node45991;
	wire [4-1:0] node45994;
	wire [4-1:0] node45997;
	wire [4-1:0] node45998;
	wire [4-1:0] node45999;
	wire [4-1:0] node46000;
	wire [4-1:0] node46001;
	wire [4-1:0] node46002;
	wire [4-1:0] node46003;
	wire [4-1:0] node46007;
	wire [4-1:0] node46008;
	wire [4-1:0] node46011;
	wire [4-1:0] node46014;
	wire [4-1:0] node46015;
	wire [4-1:0] node46017;
	wire [4-1:0] node46020;
	wire [4-1:0] node46021;
	wire [4-1:0] node46024;
	wire [4-1:0] node46027;
	wire [4-1:0] node46028;
	wire [4-1:0] node46029;
	wire [4-1:0] node46030;
	wire [4-1:0] node46033;
	wire [4-1:0] node46036;
	wire [4-1:0] node46037;
	wire [4-1:0] node46040;
	wire [4-1:0] node46043;
	wire [4-1:0] node46044;
	wire [4-1:0] node46045;
	wire [4-1:0] node46048;
	wire [4-1:0] node46051;
	wire [4-1:0] node46052;
	wire [4-1:0] node46055;
	wire [4-1:0] node46058;
	wire [4-1:0] node46059;
	wire [4-1:0] node46060;
	wire [4-1:0] node46061;
	wire [4-1:0] node46063;
	wire [4-1:0] node46066;
	wire [4-1:0] node46067;
	wire [4-1:0] node46070;
	wire [4-1:0] node46073;
	wire [4-1:0] node46074;
	wire [4-1:0] node46075;
	wire [4-1:0] node46078;
	wire [4-1:0] node46081;
	wire [4-1:0] node46082;
	wire [4-1:0] node46085;
	wire [4-1:0] node46088;
	wire [4-1:0] node46089;
	wire [4-1:0] node46090;
	wire [4-1:0] node46091;
	wire [4-1:0] node46095;
	wire [4-1:0] node46096;
	wire [4-1:0] node46100;
	wire [4-1:0] node46101;
	wire [4-1:0] node46102;
	wire [4-1:0] node46106;
	wire [4-1:0] node46107;
	wire [4-1:0] node46111;
	wire [4-1:0] node46112;
	wire [4-1:0] node46113;
	wire [4-1:0] node46114;
	wire [4-1:0] node46115;
	wire [4-1:0] node46116;
	wire [4-1:0] node46119;
	wire [4-1:0] node46122;
	wire [4-1:0] node46124;
	wire [4-1:0] node46127;
	wire [4-1:0] node46128;
	wire [4-1:0] node46130;
	wire [4-1:0] node46133;
	wire [4-1:0] node46134;
	wire [4-1:0] node46137;
	wire [4-1:0] node46140;
	wire [4-1:0] node46141;
	wire [4-1:0] node46142;
	wire [4-1:0] node46143;
	wire [4-1:0] node46146;
	wire [4-1:0] node46149;
	wire [4-1:0] node46150;
	wire [4-1:0] node46153;
	wire [4-1:0] node46156;
	wire [4-1:0] node46157;
	wire [4-1:0] node46160;
	wire [4-1:0] node46163;
	wire [4-1:0] node46164;
	wire [4-1:0] node46165;
	wire [4-1:0] node46166;
	wire [4-1:0] node46167;
	wire [4-1:0] node46170;
	wire [4-1:0] node46173;
	wire [4-1:0] node46174;
	wire [4-1:0] node46177;
	wire [4-1:0] node46180;
	wire [4-1:0] node46181;
	wire [4-1:0] node46182;
	wire [4-1:0] node46185;
	wire [4-1:0] node46188;
	wire [4-1:0] node46189;
	wire [4-1:0] node46192;
	wire [4-1:0] node46195;
	wire [4-1:0] node46196;
	wire [4-1:0] node46197;
	wire [4-1:0] node46198;
	wire [4-1:0] node46201;
	wire [4-1:0] node46204;
	wire [4-1:0] node46205;
	wire [4-1:0] node46208;
	wire [4-1:0] node46211;
	wire [4-1:0] node46212;
	wire [4-1:0] node46215;
	wire [4-1:0] node46218;
	wire [4-1:0] node46219;
	wire [4-1:0] node46220;
	wire [4-1:0] node46221;
	wire [4-1:0] node46222;
	wire [4-1:0] node46223;
	wire [4-1:0] node46224;
	wire [4-1:0] node46225;
	wire [4-1:0] node46229;
	wire [4-1:0] node46230;
	wire [4-1:0] node46234;
	wire [4-1:0] node46235;
	wire [4-1:0] node46236;
	wire [4-1:0] node46239;
	wire [4-1:0] node46242;
	wire [4-1:0] node46243;
	wire [4-1:0] node46246;
	wire [4-1:0] node46249;
	wire [4-1:0] node46250;
	wire [4-1:0] node46251;
	wire [4-1:0] node46252;
	wire [4-1:0] node46255;
	wire [4-1:0] node46258;
	wire [4-1:0] node46259;
	wire [4-1:0] node46262;
	wire [4-1:0] node46265;
	wire [4-1:0] node46266;
	wire [4-1:0] node46267;
	wire [4-1:0] node46271;
	wire [4-1:0] node46272;
	wire [4-1:0] node46276;
	wire [4-1:0] node46277;
	wire [4-1:0] node46278;
	wire [4-1:0] node46279;
	wire [4-1:0] node46280;
	wire [4-1:0] node46283;
	wire [4-1:0] node46286;
	wire [4-1:0] node46287;
	wire [4-1:0] node46290;
	wire [4-1:0] node46293;
	wire [4-1:0] node46294;
	wire [4-1:0] node46295;
	wire [4-1:0] node46298;
	wire [4-1:0] node46301;
	wire [4-1:0] node46302;
	wire [4-1:0] node46305;
	wire [4-1:0] node46308;
	wire [4-1:0] node46309;
	wire [4-1:0] node46310;
	wire [4-1:0] node46311;
	wire [4-1:0] node46315;
	wire [4-1:0] node46316;
	wire [4-1:0] node46320;
	wire [4-1:0] node46321;
	wire [4-1:0] node46322;
	wire [4-1:0] node46326;
	wire [4-1:0] node46327;
	wire [4-1:0] node46331;
	wire [4-1:0] node46332;
	wire [4-1:0] node46333;
	wire [4-1:0] node46334;
	wire [4-1:0] node46335;
	wire [4-1:0] node46337;
	wire [4-1:0] node46340;
	wire [4-1:0] node46342;
	wire [4-1:0] node46345;
	wire [4-1:0] node46346;
	wire [4-1:0] node46347;
	wire [4-1:0] node46350;
	wire [4-1:0] node46353;
	wire [4-1:0] node46354;
	wire [4-1:0] node46357;
	wire [4-1:0] node46360;
	wire [4-1:0] node46361;
	wire [4-1:0] node46362;
	wire [4-1:0] node46363;
	wire [4-1:0] node46366;
	wire [4-1:0] node46369;
	wire [4-1:0] node46370;
	wire [4-1:0] node46373;
	wire [4-1:0] node46376;
	wire [4-1:0] node46377;
	wire [4-1:0] node46378;
	wire [4-1:0] node46381;
	wire [4-1:0] node46384;
	wire [4-1:0] node46385;
	wire [4-1:0] node46389;
	wire [4-1:0] node46390;
	wire [4-1:0] node46391;
	wire [4-1:0] node46392;
	wire [4-1:0] node46393;
	wire [4-1:0] node46396;
	wire [4-1:0] node46399;
	wire [4-1:0] node46400;
	wire [4-1:0] node46403;
	wire [4-1:0] node46406;
	wire [4-1:0] node46407;
	wire [4-1:0] node46408;
	wire [4-1:0] node46411;
	wire [4-1:0] node46414;
	wire [4-1:0] node46415;
	wire [4-1:0] node46418;
	wire [4-1:0] node46421;
	wire [4-1:0] node46422;
	wire [4-1:0] node46423;
	wire [4-1:0] node46424;
	wire [4-1:0] node46427;
	wire [4-1:0] node46430;
	wire [4-1:0] node46431;
	wire [4-1:0] node46434;
	wire [4-1:0] node46437;
	wire [4-1:0] node46438;
	wire [4-1:0] node46441;
	wire [4-1:0] node46444;
	wire [4-1:0] node46445;
	wire [4-1:0] node46446;
	wire [4-1:0] node46447;
	wire [4-1:0] node46448;
	wire [4-1:0] node46449;
	wire [4-1:0] node46450;
	wire [4-1:0] node46453;
	wire [4-1:0] node46456;
	wire [4-1:0] node46457;
	wire [4-1:0] node46460;
	wire [4-1:0] node46463;
	wire [4-1:0] node46464;
	wire [4-1:0] node46465;
	wire [4-1:0] node46468;
	wire [4-1:0] node46471;
	wire [4-1:0] node46472;
	wire [4-1:0] node46475;
	wire [4-1:0] node46478;
	wire [4-1:0] node46479;
	wire [4-1:0] node46480;
	wire [4-1:0] node46481;
	wire [4-1:0] node46484;
	wire [4-1:0] node46487;
	wire [4-1:0] node46489;
	wire [4-1:0] node46492;
	wire [4-1:0] node46493;
	wire [4-1:0] node46495;
	wire [4-1:0] node46498;
	wire [4-1:0] node46499;
	wire [4-1:0] node46502;
	wire [4-1:0] node46505;
	wire [4-1:0] node46506;
	wire [4-1:0] node46507;
	wire [4-1:0] node46508;
	wire [4-1:0] node46509;
	wire [4-1:0] node46512;
	wire [4-1:0] node46515;
	wire [4-1:0] node46517;
	wire [4-1:0] node46520;
	wire [4-1:0] node46521;
	wire [4-1:0] node46522;
	wire [4-1:0] node46525;
	wire [4-1:0] node46528;
	wire [4-1:0] node46529;
	wire [4-1:0] node46532;
	wire [4-1:0] node46535;
	wire [4-1:0] node46536;
	wire [4-1:0] node46537;
	wire [4-1:0] node46538;
	wire [4-1:0] node46541;
	wire [4-1:0] node46544;
	wire [4-1:0] node46546;
	wire [4-1:0] node46549;
	wire [4-1:0] node46550;
	wire [4-1:0] node46551;
	wire [4-1:0] node46554;
	wire [4-1:0] node46557;
	wire [4-1:0] node46558;
	wire [4-1:0] node46561;
	wire [4-1:0] node46564;
	wire [4-1:0] node46565;
	wire [4-1:0] node46566;
	wire [4-1:0] node46567;
	wire [4-1:0] node46568;
	wire [4-1:0] node46569;
	wire [4-1:0] node46572;
	wire [4-1:0] node46575;
	wire [4-1:0] node46576;
	wire [4-1:0] node46579;
	wire [4-1:0] node46582;
	wire [4-1:0] node46583;
	wire [4-1:0] node46584;
	wire [4-1:0] node46587;
	wire [4-1:0] node46590;
	wire [4-1:0] node46591;
	wire [4-1:0] node46594;
	wire [4-1:0] node46597;
	wire [4-1:0] node46598;
	wire [4-1:0] node46599;
	wire [4-1:0] node46600;
	wire [4-1:0] node46603;
	wire [4-1:0] node46606;
	wire [4-1:0] node46607;
	wire [4-1:0] node46610;
	wire [4-1:0] node46613;
	wire [4-1:0] node46614;
	wire [4-1:0] node46615;
	wire [4-1:0] node46618;
	wire [4-1:0] node46621;
	wire [4-1:0] node46622;
	wire [4-1:0] node46625;
	wire [4-1:0] node46628;
	wire [4-1:0] node46629;
	wire [4-1:0] node46630;
	wire [4-1:0] node46631;
	wire [4-1:0] node46632;
	wire [4-1:0] node46635;
	wire [4-1:0] node46638;
	wire [4-1:0] node46639;
	wire [4-1:0] node46642;
	wire [4-1:0] node46645;
	wire [4-1:0] node46646;
	wire [4-1:0] node46647;
	wire [4-1:0] node46650;
	wire [4-1:0] node46653;
	wire [4-1:0] node46654;
	wire [4-1:0] node46657;
	wire [4-1:0] node46660;
	wire [4-1:0] node46661;
	wire [4-1:0] node46662;
	wire [4-1:0] node46663;
	wire [4-1:0] node46666;
	wire [4-1:0] node46669;
	wire [4-1:0] node46670;
	wire [4-1:0] node46673;
	wire [4-1:0] node46676;
	wire [4-1:0] node46677;
	wire [4-1:0] node46678;
	wire [4-1:0] node46681;
	wire [4-1:0] node46684;
	wire [4-1:0] node46685;
	wire [4-1:0] node46688;
	wire [4-1:0] node46691;
	wire [4-1:0] node46692;
	wire [4-1:0] node46693;
	wire [4-1:0] node46694;
	wire [4-1:0] node46695;
	wire [4-1:0] node46696;
	wire [4-1:0] node46697;
	wire [4-1:0] node46698;
	wire [4-1:0] node46699;
	wire [4-1:0] node46700;
	wire [4-1:0] node46702;
	wire [4-1:0] node46705;
	wire [4-1:0] node46707;
	wire [4-1:0] node46710;
	wire [4-1:0] node46711;
	wire [4-1:0] node46712;
	wire [4-1:0] node46715;
	wire [4-1:0] node46718;
	wire [4-1:0] node46719;
	wire [4-1:0] node46723;
	wire [4-1:0] node46724;
	wire [4-1:0] node46725;
	wire [4-1:0] node46726;
	wire [4-1:0] node46729;
	wire [4-1:0] node46732;
	wire [4-1:0] node46733;
	wire [4-1:0] node46736;
	wire [4-1:0] node46739;
	wire [4-1:0] node46740;
	wire [4-1:0] node46742;
	wire [4-1:0] node46745;
	wire [4-1:0] node46746;
	wire [4-1:0] node46749;
	wire [4-1:0] node46752;
	wire [4-1:0] node46753;
	wire [4-1:0] node46754;
	wire [4-1:0] node46755;
	wire [4-1:0] node46757;
	wire [4-1:0] node46760;
	wire [4-1:0] node46762;
	wire [4-1:0] node46765;
	wire [4-1:0] node46766;
	wire [4-1:0] node46767;
	wire [4-1:0] node46770;
	wire [4-1:0] node46773;
	wire [4-1:0] node46774;
	wire [4-1:0] node46777;
	wire [4-1:0] node46780;
	wire [4-1:0] node46781;
	wire [4-1:0] node46782;
	wire [4-1:0] node46783;
	wire [4-1:0] node46787;
	wire [4-1:0] node46788;
	wire [4-1:0] node46792;
	wire [4-1:0] node46793;
	wire [4-1:0] node46794;
	wire [4-1:0] node46798;
	wire [4-1:0] node46799;
	wire [4-1:0] node46803;
	wire [4-1:0] node46804;
	wire [4-1:0] node46805;
	wire [4-1:0] node46806;
	wire [4-1:0] node46807;
	wire [4-1:0] node46808;
	wire [4-1:0] node46811;
	wire [4-1:0] node46814;
	wire [4-1:0] node46815;
	wire [4-1:0] node46818;
	wire [4-1:0] node46821;
	wire [4-1:0] node46822;
	wire [4-1:0] node46823;
	wire [4-1:0] node46826;
	wire [4-1:0] node46829;
	wire [4-1:0] node46830;
	wire [4-1:0] node46834;
	wire [4-1:0] node46835;
	wire [4-1:0] node46836;
	wire [4-1:0] node46837;
	wire [4-1:0] node46841;
	wire [4-1:0] node46842;
	wire [4-1:0] node46846;
	wire [4-1:0] node46847;
	wire [4-1:0] node46848;
	wire [4-1:0] node46852;
	wire [4-1:0] node46855;
	wire [4-1:0] node46856;
	wire [4-1:0] node46857;
	wire [4-1:0] node46858;
	wire [4-1:0] node46859;
	wire [4-1:0] node46862;
	wire [4-1:0] node46865;
	wire [4-1:0] node46866;
	wire [4-1:0] node46869;
	wire [4-1:0] node46872;
	wire [4-1:0] node46873;
	wire [4-1:0] node46875;
	wire [4-1:0] node46878;
	wire [4-1:0] node46879;
	wire [4-1:0] node46882;
	wire [4-1:0] node46885;
	wire [4-1:0] node46886;
	wire [4-1:0] node46887;
	wire [4-1:0] node46888;
	wire [4-1:0] node46891;
	wire [4-1:0] node46894;
	wire [4-1:0] node46895;
	wire [4-1:0] node46898;
	wire [4-1:0] node46901;
	wire [4-1:0] node46902;
	wire [4-1:0] node46905;
	wire [4-1:0] node46908;
	wire [4-1:0] node46909;
	wire [4-1:0] node46910;
	wire [4-1:0] node46911;
	wire [4-1:0] node46912;
	wire [4-1:0] node46913;
	wire [4-1:0] node46914;
	wire [4-1:0] node46917;
	wire [4-1:0] node46920;
	wire [4-1:0] node46921;
	wire [4-1:0] node46924;
	wire [4-1:0] node46927;
	wire [4-1:0] node46928;
	wire [4-1:0] node46930;
	wire [4-1:0] node46933;
	wire [4-1:0] node46934;
	wire [4-1:0] node46937;
	wire [4-1:0] node46940;
	wire [4-1:0] node46941;
	wire [4-1:0] node46942;
	wire [4-1:0] node46943;
	wire [4-1:0] node46946;
	wire [4-1:0] node46949;
	wire [4-1:0] node46950;
	wire [4-1:0] node46953;
	wire [4-1:0] node46956;
	wire [4-1:0] node46957;
	wire [4-1:0] node46960;
	wire [4-1:0] node46963;
	wire [4-1:0] node46964;
	wire [4-1:0] node46965;
	wire [4-1:0] node46966;
	wire [4-1:0] node46967;
	wire [4-1:0] node46970;
	wire [4-1:0] node46973;
	wire [4-1:0] node46974;
	wire [4-1:0] node46977;
	wire [4-1:0] node46980;
	wire [4-1:0] node46981;
	wire [4-1:0] node46982;
	wire [4-1:0] node46986;
	wire [4-1:0] node46987;
	wire [4-1:0] node46990;
	wire [4-1:0] node46993;
	wire [4-1:0] node46994;
	wire [4-1:0] node46995;
	wire [4-1:0] node46996;
	wire [4-1:0] node46999;
	wire [4-1:0] node47002;
	wire [4-1:0] node47003;
	wire [4-1:0] node47006;
	wire [4-1:0] node47009;
	wire [4-1:0] node47010;
	wire [4-1:0] node47011;
	wire [4-1:0] node47014;
	wire [4-1:0] node47017;
	wire [4-1:0] node47018;
	wire [4-1:0] node47021;
	wire [4-1:0] node47024;
	wire [4-1:0] node47025;
	wire [4-1:0] node47026;
	wire [4-1:0] node47027;
	wire [4-1:0] node47028;
	wire [4-1:0] node47030;
	wire [4-1:0] node47033;
	wire [4-1:0] node47034;
	wire [4-1:0] node47037;
	wire [4-1:0] node47040;
	wire [4-1:0] node47041;
	wire [4-1:0] node47042;
	wire [4-1:0] node47045;
	wire [4-1:0] node47048;
	wire [4-1:0] node47049;
	wire [4-1:0] node47053;
	wire [4-1:0] node47054;
	wire [4-1:0] node47055;
	wire [4-1:0] node47056;
	wire [4-1:0] node47060;
	wire [4-1:0] node47061;
	wire [4-1:0] node47065;
	wire [4-1:0] node47066;
	wire [4-1:0] node47067;
	wire [4-1:0] node47071;
	wire [4-1:0] node47072;
	wire [4-1:0] node47076;
	wire [4-1:0] node47077;
	wire [4-1:0] node47078;
	wire [4-1:0] node47079;
	wire [4-1:0] node47080;
	wire [4-1:0] node47083;
	wire [4-1:0] node47086;
	wire [4-1:0] node47087;
	wire [4-1:0] node47090;
	wire [4-1:0] node47093;
	wire [4-1:0] node47094;
	wire [4-1:0] node47095;
	wire [4-1:0] node47098;
	wire [4-1:0] node47101;
	wire [4-1:0] node47104;
	wire [4-1:0] node47105;
	wire [4-1:0] node47106;
	wire [4-1:0] node47107;
	wire [4-1:0] node47110;
	wire [4-1:0] node47113;
	wire [4-1:0] node47114;
	wire [4-1:0] node47117;
	wire [4-1:0] node47120;
	wire [4-1:0] node47121;
	wire [4-1:0] node47124;
	wire [4-1:0] node47127;
	wire [4-1:0] node47128;
	wire [4-1:0] node47129;
	wire [4-1:0] node47130;
	wire [4-1:0] node47131;
	wire [4-1:0] node47132;
	wire [4-1:0] node47133;
	wire [4-1:0] node47134;
	wire [4-1:0] node47137;
	wire [4-1:0] node47140;
	wire [4-1:0] node47141;
	wire [4-1:0] node47144;
	wire [4-1:0] node47147;
	wire [4-1:0] node47148;
	wire [4-1:0] node47149;
	wire [4-1:0] node47152;
	wire [4-1:0] node47155;
	wire [4-1:0] node47157;
	wire [4-1:0] node47160;
	wire [4-1:0] node47161;
	wire [4-1:0] node47162;
	wire [4-1:0] node47163;
	wire [4-1:0] node47167;
	wire [4-1:0] node47168;
	wire [4-1:0] node47172;
	wire [4-1:0] node47173;
	wire [4-1:0] node47174;
	wire [4-1:0] node47178;
	wire [4-1:0] node47179;
	wire [4-1:0] node47183;
	wire [4-1:0] node47184;
	wire [4-1:0] node47185;
	wire [4-1:0] node47186;
	wire [4-1:0] node47187;
	wire [4-1:0] node47190;
	wire [4-1:0] node47193;
	wire [4-1:0] node47194;
	wire [4-1:0] node47197;
	wire [4-1:0] node47200;
	wire [4-1:0] node47201;
	wire [4-1:0] node47202;
	wire [4-1:0] node47205;
	wire [4-1:0] node47208;
	wire [4-1:0] node47209;
	wire [4-1:0] node47212;
	wire [4-1:0] node47215;
	wire [4-1:0] node47216;
	wire [4-1:0] node47217;
	wire [4-1:0] node47218;
	wire [4-1:0] node47221;
	wire [4-1:0] node47224;
	wire [4-1:0] node47225;
	wire [4-1:0] node47228;
	wire [4-1:0] node47231;
	wire [4-1:0] node47232;
	wire [4-1:0] node47233;
	wire [4-1:0] node47236;
	wire [4-1:0] node47239;
	wire [4-1:0] node47240;
	wire [4-1:0] node47243;
	wire [4-1:0] node47246;
	wire [4-1:0] node47247;
	wire [4-1:0] node47248;
	wire [4-1:0] node47249;
	wire [4-1:0] node47250;
	wire [4-1:0] node47251;
	wire [4-1:0] node47255;
	wire [4-1:0] node47256;
	wire [4-1:0] node47259;
	wire [4-1:0] node47262;
	wire [4-1:0] node47263;
	wire [4-1:0] node47264;
	wire [4-1:0] node47267;
	wire [4-1:0] node47270;
	wire [4-1:0] node47271;
	wire [4-1:0] node47274;
	wire [4-1:0] node47277;
	wire [4-1:0] node47278;
	wire [4-1:0] node47279;
	wire [4-1:0] node47280;
	wire [4-1:0] node47284;
	wire [4-1:0] node47285;
	wire [4-1:0] node47289;
	wire [4-1:0] node47290;
	wire [4-1:0] node47291;
	wire [4-1:0] node47295;
	wire [4-1:0] node47296;
	wire [4-1:0] node47300;
	wire [4-1:0] node47301;
	wire [4-1:0] node47302;
	wire [4-1:0] node47303;
	wire [4-1:0] node47304;
	wire [4-1:0] node47308;
	wire [4-1:0] node47309;
	wire [4-1:0] node47312;
	wire [4-1:0] node47315;
	wire [4-1:0] node47316;
	wire [4-1:0] node47317;
	wire [4-1:0] node47320;
	wire [4-1:0] node47323;
	wire [4-1:0] node47324;
	wire [4-1:0] node47327;
	wire [4-1:0] node47330;
	wire [4-1:0] node47331;
	wire [4-1:0] node47332;
	wire [4-1:0] node47333;
	wire [4-1:0] node47337;
	wire [4-1:0] node47338;
	wire [4-1:0] node47342;
	wire [4-1:0] node47344;
	wire [4-1:0] node47345;
	wire [4-1:0] node47349;
	wire [4-1:0] node47350;
	wire [4-1:0] node47351;
	wire [4-1:0] node47352;
	wire [4-1:0] node47353;
	wire [4-1:0] node47354;
	wire [4-1:0] node47355;
	wire [4-1:0] node47358;
	wire [4-1:0] node47361;
	wire [4-1:0] node47362;
	wire [4-1:0] node47365;
	wire [4-1:0] node47368;
	wire [4-1:0] node47369;
	wire [4-1:0] node47371;
	wire [4-1:0] node47374;
	wire [4-1:0] node47376;
	wire [4-1:0] node47379;
	wire [4-1:0] node47380;
	wire [4-1:0] node47381;
	wire [4-1:0] node47382;
	wire [4-1:0] node47386;
	wire [4-1:0] node47387;
	wire [4-1:0] node47391;
	wire [4-1:0] node47392;
	wire [4-1:0] node47393;
	wire [4-1:0] node47397;
	wire [4-1:0] node47398;
	wire [4-1:0] node47402;
	wire [4-1:0] node47403;
	wire [4-1:0] node47404;
	wire [4-1:0] node47405;
	wire [4-1:0] node47406;
	wire [4-1:0] node47409;
	wire [4-1:0] node47412;
	wire [4-1:0] node47413;
	wire [4-1:0] node47416;
	wire [4-1:0] node47419;
	wire [4-1:0] node47420;
	wire [4-1:0] node47421;
	wire [4-1:0] node47424;
	wire [4-1:0] node47427;
	wire [4-1:0] node47428;
	wire [4-1:0] node47431;
	wire [4-1:0] node47434;
	wire [4-1:0] node47435;
	wire [4-1:0] node47436;
	wire [4-1:0] node47437;
	wire [4-1:0] node47441;
	wire [4-1:0] node47442;
	wire [4-1:0] node47445;
	wire [4-1:0] node47448;
	wire [4-1:0] node47449;
	wire [4-1:0] node47450;
	wire [4-1:0] node47453;
	wire [4-1:0] node47456;
	wire [4-1:0] node47457;
	wire [4-1:0] node47460;
	wire [4-1:0] node47463;
	wire [4-1:0] node47464;
	wire [4-1:0] node47465;
	wire [4-1:0] node47466;
	wire [4-1:0] node47467;
	wire [4-1:0] node47468;
	wire [4-1:0] node47471;
	wire [4-1:0] node47474;
	wire [4-1:0] node47475;
	wire [4-1:0] node47478;
	wire [4-1:0] node47481;
	wire [4-1:0] node47482;
	wire [4-1:0] node47483;
	wire [4-1:0] node47486;
	wire [4-1:0] node47489;
	wire [4-1:0] node47490;
	wire [4-1:0] node47493;
	wire [4-1:0] node47496;
	wire [4-1:0] node47497;
	wire [4-1:0] node47498;
	wire [4-1:0] node47499;
	wire [4-1:0] node47502;
	wire [4-1:0] node47505;
	wire [4-1:0] node47506;
	wire [4-1:0] node47509;
	wire [4-1:0] node47512;
	wire [4-1:0] node47513;
	wire [4-1:0] node47516;
	wire [4-1:0] node47519;
	wire [4-1:0] node47520;
	wire [4-1:0] node47521;
	wire [4-1:0] node47522;
	wire [4-1:0] node47523;
	wire [4-1:0] node47526;
	wire [4-1:0] node47529;
	wire [4-1:0] node47530;
	wire [4-1:0] node47533;
	wire [4-1:0] node47536;
	wire [4-1:0] node47537;
	wire [4-1:0] node47538;
	wire [4-1:0] node47541;
	wire [4-1:0] node47544;
	wire [4-1:0] node47545;
	wire [4-1:0] node47548;
	wire [4-1:0] node47551;
	wire [4-1:0] node47552;
	wire [4-1:0] node47553;
	wire [4-1:0] node47554;
	wire [4-1:0] node47557;
	wire [4-1:0] node47560;
	wire [4-1:0] node47561;
	wire [4-1:0] node47564;
	wire [4-1:0] node47567;
	wire [4-1:0] node47568;
	wire [4-1:0] node47571;
	wire [4-1:0] node47574;
	wire [4-1:0] node47575;
	wire [4-1:0] node47576;
	wire [4-1:0] node47577;
	wire [4-1:0] node47578;
	wire [4-1:0] node47579;
	wire [4-1:0] node47580;
	wire [4-1:0] node47581;
	wire [4-1:0] node47582;
	wire [4-1:0] node47586;
	wire [4-1:0] node47587;
	wire [4-1:0] node47590;
	wire [4-1:0] node47593;
	wire [4-1:0] node47594;
	wire [4-1:0] node47595;
	wire [4-1:0] node47598;
	wire [4-1:0] node47601;
	wire [4-1:0] node47603;
	wire [4-1:0] node47606;
	wire [4-1:0] node47607;
	wire [4-1:0] node47608;
	wire [4-1:0] node47609;
	wire [4-1:0] node47613;
	wire [4-1:0] node47614;
	wire [4-1:0] node47618;
	wire [4-1:0] node47619;
	wire [4-1:0] node47620;
	wire [4-1:0] node47624;
	wire [4-1:0] node47625;
	wire [4-1:0] node47629;
	wire [4-1:0] node47630;
	wire [4-1:0] node47631;
	wire [4-1:0] node47632;
	wire [4-1:0] node47633;
	wire [4-1:0] node47636;
	wire [4-1:0] node47639;
	wire [4-1:0] node47640;
	wire [4-1:0] node47643;
	wire [4-1:0] node47646;
	wire [4-1:0] node47647;
	wire [4-1:0] node47648;
	wire [4-1:0] node47651;
	wire [4-1:0] node47654;
	wire [4-1:0] node47655;
	wire [4-1:0] node47659;
	wire [4-1:0] node47660;
	wire [4-1:0] node47661;
	wire [4-1:0] node47662;
	wire [4-1:0] node47665;
	wire [4-1:0] node47668;
	wire [4-1:0] node47669;
	wire [4-1:0] node47672;
	wire [4-1:0] node47675;
	wire [4-1:0] node47676;
	wire [4-1:0] node47677;
	wire [4-1:0] node47680;
	wire [4-1:0] node47683;
	wire [4-1:0] node47684;
	wire [4-1:0] node47687;
	wire [4-1:0] node47690;
	wire [4-1:0] node47691;
	wire [4-1:0] node47692;
	wire [4-1:0] node47693;
	wire [4-1:0] node47694;
	wire [4-1:0] node47695;
	wire [4-1:0] node47698;
	wire [4-1:0] node47701;
	wire [4-1:0] node47702;
	wire [4-1:0] node47705;
	wire [4-1:0] node47708;
	wire [4-1:0] node47709;
	wire [4-1:0] node47710;
	wire [4-1:0] node47713;
	wire [4-1:0] node47716;
	wire [4-1:0] node47717;
	wire [4-1:0] node47720;
	wire [4-1:0] node47723;
	wire [4-1:0] node47724;
	wire [4-1:0] node47725;
	wire [4-1:0] node47726;
	wire [4-1:0] node47730;
	wire [4-1:0] node47731;
	wire [4-1:0] node47735;
	wire [4-1:0] node47736;
	wire [4-1:0] node47737;
	wire [4-1:0] node47741;
	wire [4-1:0] node47742;
	wire [4-1:0] node47746;
	wire [4-1:0] node47747;
	wire [4-1:0] node47748;
	wire [4-1:0] node47749;
	wire [4-1:0] node47750;
	wire [4-1:0] node47753;
	wire [4-1:0] node47756;
	wire [4-1:0] node47757;
	wire [4-1:0] node47761;
	wire [4-1:0] node47762;
	wire [4-1:0] node47763;
	wire [4-1:0] node47766;
	wire [4-1:0] node47769;
	wire [4-1:0] node47770;
	wire [4-1:0] node47773;
	wire [4-1:0] node47776;
	wire [4-1:0] node47777;
	wire [4-1:0] node47778;
	wire [4-1:0] node47779;
	wire [4-1:0] node47782;
	wire [4-1:0] node47785;
	wire [4-1:0] node47786;
	wire [4-1:0] node47789;
	wire [4-1:0] node47792;
	wire [4-1:0] node47793;
	wire [4-1:0] node47796;
	wire [4-1:0] node47799;
	wire [4-1:0] node47800;
	wire [4-1:0] node47801;
	wire [4-1:0] node47802;
	wire [4-1:0] node47803;
	wire [4-1:0] node47804;
	wire [4-1:0] node47807;
	wire [4-1:0] node47808;
	wire [4-1:0] node47811;
	wire [4-1:0] node47814;
	wire [4-1:0] node47815;
	wire [4-1:0] node47816;
	wire [4-1:0] node47819;
	wire [4-1:0] node47822;
	wire [4-1:0] node47823;
	wire [4-1:0] node47826;
	wire [4-1:0] node47829;
	wire [4-1:0] node47830;
	wire [4-1:0] node47831;
	wire [4-1:0] node47832;
	wire [4-1:0] node47835;
	wire [4-1:0] node47838;
	wire [4-1:0] node47839;
	wire [4-1:0] node47842;
	wire [4-1:0] node47845;
	wire [4-1:0] node47846;
	wire [4-1:0] node47847;
	wire [4-1:0] node47850;
	wire [4-1:0] node47853;
	wire [4-1:0] node47854;
	wire [4-1:0] node47857;
	wire [4-1:0] node47860;
	wire [4-1:0] node47861;
	wire [4-1:0] node47862;
	wire [4-1:0] node47863;
	wire [4-1:0] node47864;
	wire [4-1:0] node47867;
	wire [4-1:0] node47870;
	wire [4-1:0] node47871;
	wire [4-1:0] node47874;
	wire [4-1:0] node47877;
	wire [4-1:0] node47878;
	wire [4-1:0] node47879;
	wire [4-1:0] node47883;
	wire [4-1:0] node47884;
	wire [4-1:0] node47887;
	wire [4-1:0] node47890;
	wire [4-1:0] node47891;
	wire [4-1:0] node47892;
	wire [4-1:0] node47893;
	wire [4-1:0] node47896;
	wire [4-1:0] node47899;
	wire [4-1:0] node47900;
	wire [4-1:0] node47903;
	wire [4-1:0] node47906;
	wire [4-1:0] node47907;
	wire [4-1:0] node47909;
	wire [4-1:0] node47912;
	wire [4-1:0] node47913;
	wire [4-1:0] node47916;
	wire [4-1:0] node47919;
	wire [4-1:0] node47920;
	wire [4-1:0] node47921;
	wire [4-1:0] node47922;
	wire [4-1:0] node47923;
	wire [4-1:0] node47924;
	wire [4-1:0] node47927;
	wire [4-1:0] node47930;
	wire [4-1:0] node47931;
	wire [4-1:0] node47934;
	wire [4-1:0] node47937;
	wire [4-1:0] node47938;
	wire [4-1:0] node47939;
	wire [4-1:0] node47943;
	wire [4-1:0] node47944;
	wire [4-1:0] node47947;
	wire [4-1:0] node47950;
	wire [4-1:0] node47951;
	wire [4-1:0] node47952;
	wire [4-1:0] node47953;
	wire [4-1:0] node47957;
	wire [4-1:0] node47958;
	wire [4-1:0] node47962;
	wire [4-1:0] node47963;
	wire [4-1:0] node47964;
	wire [4-1:0] node47968;
	wire [4-1:0] node47969;
	wire [4-1:0] node47973;
	wire [4-1:0] node47974;
	wire [4-1:0] node47975;
	wire [4-1:0] node47976;
	wire [4-1:0] node47977;
	wire [4-1:0] node47980;
	wire [4-1:0] node47983;
	wire [4-1:0] node47984;
	wire [4-1:0] node47987;
	wire [4-1:0] node47990;
	wire [4-1:0] node47991;
	wire [4-1:0] node47992;
	wire [4-1:0] node47995;
	wire [4-1:0] node47998;
	wire [4-1:0] node47999;
	wire [4-1:0] node48002;
	wire [4-1:0] node48005;
	wire [4-1:0] node48006;
	wire [4-1:0] node48007;
	wire [4-1:0] node48008;
	wire [4-1:0] node48011;
	wire [4-1:0] node48014;
	wire [4-1:0] node48015;
	wire [4-1:0] node48018;
	wire [4-1:0] node48021;
	wire [4-1:0] node48022;
	wire [4-1:0] node48025;
	wire [4-1:0] node48028;
	wire [4-1:0] node48029;
	wire [4-1:0] node48030;
	wire [4-1:0] node48031;
	wire [4-1:0] node48032;
	wire [4-1:0] node48033;
	wire [4-1:0] node48034;
	wire [4-1:0] node48035;
	wire [4-1:0] node48038;
	wire [4-1:0] node48041;
	wire [4-1:0] node48042;
	wire [4-1:0] node48045;
	wire [4-1:0] node48048;
	wire [4-1:0] node48049;
	wire [4-1:0] node48050;
	wire [4-1:0] node48053;
	wire [4-1:0] node48056;
	wire [4-1:0] node48057;
	wire [4-1:0] node48060;
	wire [4-1:0] node48063;
	wire [4-1:0] node48064;
	wire [4-1:0] node48065;
	wire [4-1:0] node48066;
	wire [4-1:0] node48069;
	wire [4-1:0] node48072;
	wire [4-1:0] node48073;
	wire [4-1:0] node48076;
	wire [4-1:0] node48079;
	wire [4-1:0] node48080;
	wire [4-1:0] node48081;
	wire [4-1:0] node48084;
	wire [4-1:0] node48087;
	wire [4-1:0] node48088;
	wire [4-1:0] node48092;
	wire [4-1:0] node48093;
	wire [4-1:0] node48094;
	wire [4-1:0] node48095;
	wire [4-1:0] node48096;
	wire [4-1:0] node48099;
	wire [4-1:0] node48102;
	wire [4-1:0] node48103;
	wire [4-1:0] node48106;
	wire [4-1:0] node48109;
	wire [4-1:0] node48110;
	wire [4-1:0] node48112;
	wire [4-1:0] node48115;
	wire [4-1:0] node48117;
	wire [4-1:0] node48120;
	wire [4-1:0] node48121;
	wire [4-1:0] node48122;
	wire [4-1:0] node48123;
	wire [4-1:0] node48126;
	wire [4-1:0] node48129;
	wire [4-1:0] node48130;
	wire [4-1:0] node48133;
	wire [4-1:0] node48136;
	wire [4-1:0] node48137;
	wire [4-1:0] node48138;
	wire [4-1:0] node48141;
	wire [4-1:0] node48144;
	wire [4-1:0] node48145;
	wire [4-1:0] node48149;
	wire [4-1:0] node48150;
	wire [4-1:0] node48151;
	wire [4-1:0] node48152;
	wire [4-1:0] node48153;
	wire [4-1:0] node48155;
	wire [4-1:0] node48158;
	wire [4-1:0] node48160;
	wire [4-1:0] node48163;
	wire [4-1:0] node48164;
	wire [4-1:0] node48165;
	wire [4-1:0] node48168;
	wire [4-1:0] node48171;
	wire [4-1:0] node48172;
	wire [4-1:0] node48176;
	wire [4-1:0] node48177;
	wire [4-1:0] node48178;
	wire [4-1:0] node48179;
	wire [4-1:0] node48182;
	wire [4-1:0] node48185;
	wire [4-1:0] node48186;
	wire [4-1:0] node48189;
	wire [4-1:0] node48192;
	wire [4-1:0] node48193;
	wire [4-1:0] node48194;
	wire [4-1:0] node48197;
	wire [4-1:0] node48200;
	wire [4-1:0] node48201;
	wire [4-1:0] node48205;
	wire [4-1:0] node48206;
	wire [4-1:0] node48207;
	wire [4-1:0] node48208;
	wire [4-1:0] node48209;
	wire [4-1:0] node48212;
	wire [4-1:0] node48215;
	wire [4-1:0] node48217;
	wire [4-1:0] node48220;
	wire [4-1:0] node48221;
	wire [4-1:0] node48223;
	wire [4-1:0] node48226;
	wire [4-1:0] node48228;
	wire [4-1:0] node48231;
	wire [4-1:0] node48232;
	wire [4-1:0] node48233;
	wire [4-1:0] node48234;
	wire [4-1:0] node48238;
	wire [4-1:0] node48239;
	wire [4-1:0] node48243;
	wire [4-1:0] node48244;
	wire [4-1:0] node48245;
	wire [4-1:0] node48249;
	wire [4-1:0] node48250;
	wire [4-1:0] node48254;
	wire [4-1:0] node48255;
	wire [4-1:0] node48256;
	wire [4-1:0] node48257;
	wire [4-1:0] node48258;
	wire [4-1:0] node48259;
	wire [4-1:0] node48260;
	wire [4-1:0] node48263;
	wire [4-1:0] node48266;
	wire [4-1:0] node48267;
	wire [4-1:0] node48270;
	wire [4-1:0] node48273;
	wire [4-1:0] node48274;
	wire [4-1:0] node48275;
	wire [4-1:0] node48279;
	wire [4-1:0] node48280;
	wire [4-1:0] node48283;
	wire [4-1:0] node48286;
	wire [4-1:0] node48287;
	wire [4-1:0] node48288;
	wire [4-1:0] node48289;
	wire [4-1:0] node48293;
	wire [4-1:0] node48294;
	wire [4-1:0] node48298;
	wire [4-1:0] node48299;
	wire [4-1:0] node48300;
	wire [4-1:0] node48304;
	wire [4-1:0] node48305;
	wire [4-1:0] node48309;
	wire [4-1:0] node48310;
	wire [4-1:0] node48311;
	wire [4-1:0] node48312;
	wire [4-1:0] node48313;
	wire [4-1:0] node48316;
	wire [4-1:0] node48319;
	wire [4-1:0] node48320;
	wire [4-1:0] node48324;
	wire [4-1:0] node48325;
	wire [4-1:0] node48326;
	wire [4-1:0] node48329;
	wire [4-1:0] node48332;
	wire [4-1:0] node48334;
	wire [4-1:0] node48337;
	wire [4-1:0] node48338;
	wire [4-1:0] node48339;
	wire [4-1:0] node48340;
	wire [4-1:0] node48343;
	wire [4-1:0] node48346;
	wire [4-1:0] node48347;
	wire [4-1:0] node48350;
	wire [4-1:0] node48353;
	wire [4-1:0] node48354;
	wire [4-1:0] node48355;
	wire [4-1:0] node48358;
	wire [4-1:0] node48361;
	wire [4-1:0] node48363;
	wire [4-1:0] node48366;
	wire [4-1:0] node48367;
	wire [4-1:0] node48368;
	wire [4-1:0] node48369;
	wire [4-1:0] node48370;
	wire [4-1:0] node48371;
	wire [4-1:0] node48374;
	wire [4-1:0] node48377;
	wire [4-1:0] node48379;
	wire [4-1:0] node48382;
	wire [4-1:0] node48383;
	wire [4-1:0] node48384;
	wire [4-1:0] node48387;
	wire [4-1:0] node48390;
	wire [4-1:0] node48391;
	wire [4-1:0] node48394;
	wire [4-1:0] node48397;
	wire [4-1:0] node48398;
	wire [4-1:0] node48399;
	wire [4-1:0] node48400;
	wire [4-1:0] node48404;
	wire [4-1:0] node48405;
	wire [4-1:0] node48409;
	wire [4-1:0] node48410;
	wire [4-1:0] node48411;
	wire [4-1:0] node48415;
	wire [4-1:0] node48416;
	wire [4-1:0] node48420;
	wire [4-1:0] node48421;
	wire [4-1:0] node48422;
	wire [4-1:0] node48423;
	wire [4-1:0] node48424;
	wire [4-1:0] node48427;
	wire [4-1:0] node48430;
	wire [4-1:0] node48431;
	wire [4-1:0] node48434;
	wire [4-1:0] node48437;
	wire [4-1:0] node48438;
	wire [4-1:0] node48439;
	wire [4-1:0] node48442;
	wire [4-1:0] node48445;
	wire [4-1:0] node48446;
	wire [4-1:0] node48449;
	wire [4-1:0] node48452;
	wire [4-1:0] node48453;
	wire [4-1:0] node48454;
	wire [4-1:0] node48455;
	wire [4-1:0] node48459;
	wire [4-1:0] node48460;
	wire [4-1:0] node48464;
	wire [4-1:0] node48465;
	wire [4-1:0] node48466;
	wire [4-1:0] node48470;
	wire [4-1:0] node48471;
	wire [4-1:0] node48475;
	wire [4-1:0] node48476;
	wire [4-1:0] node48477;
	wire [4-1:0] node48478;
	wire [4-1:0] node48479;
	wire [4-1:0] node48480;
	wire [4-1:0] node48481;
	wire [4-1:0] node48482;
	wire [4-1:0] node48483;
	wire [4-1:0] node48484;
	wire [4-1:0] node48487;
	wire [4-1:0] node48490;
	wire [4-1:0] node48491;
	wire [4-1:0] node48494;
	wire [4-1:0] node48497;
	wire [4-1:0] node48499;
	wire [4-1:0] node48500;
	wire [4-1:0] node48503;
	wire [4-1:0] node48506;
	wire [4-1:0] node48507;
	wire [4-1:0] node48508;
	wire [4-1:0] node48509;
	wire [4-1:0] node48512;
	wire [4-1:0] node48515;
	wire [4-1:0] node48516;
	wire [4-1:0] node48520;
	wire [4-1:0] node48521;
	wire [4-1:0] node48522;
	wire [4-1:0] node48525;
	wire [4-1:0] node48528;
	wire [4-1:0] node48529;
	wire [4-1:0] node48532;
	wire [4-1:0] node48535;
	wire [4-1:0] node48536;
	wire [4-1:0] node48537;
	wire [4-1:0] node48538;
	wire [4-1:0] node48539;
	wire [4-1:0] node48542;
	wire [4-1:0] node48545;
	wire [4-1:0] node48546;
	wire [4-1:0] node48549;
	wire [4-1:0] node48552;
	wire [4-1:0] node48553;
	wire [4-1:0] node48554;
	wire [4-1:0] node48557;
	wire [4-1:0] node48560;
	wire [4-1:0] node48561;
	wire [4-1:0] node48564;
	wire [4-1:0] node48567;
	wire [4-1:0] node48568;
	wire [4-1:0] node48569;
	wire [4-1:0] node48571;
	wire [4-1:0] node48574;
	wire [4-1:0] node48575;
	wire [4-1:0] node48578;
	wire [4-1:0] node48581;
	wire [4-1:0] node48582;
	wire [4-1:0] node48583;
	wire [4-1:0] node48586;
	wire [4-1:0] node48589;
	wire [4-1:0] node48590;
	wire [4-1:0] node48593;
	wire [4-1:0] node48596;
	wire [4-1:0] node48597;
	wire [4-1:0] node48598;
	wire [4-1:0] node48599;
	wire [4-1:0] node48600;
	wire [4-1:0] node48601;
	wire [4-1:0] node48604;
	wire [4-1:0] node48607;
	wire [4-1:0] node48608;
	wire [4-1:0] node48611;
	wire [4-1:0] node48614;
	wire [4-1:0] node48615;
	wire [4-1:0] node48616;
	wire [4-1:0] node48619;
	wire [4-1:0] node48622;
	wire [4-1:0] node48623;
	wire [4-1:0] node48626;
	wire [4-1:0] node48629;
	wire [4-1:0] node48630;
	wire [4-1:0] node48631;
	wire [4-1:0] node48632;
	wire [4-1:0] node48635;
	wire [4-1:0] node48638;
	wire [4-1:0] node48640;
	wire [4-1:0] node48643;
	wire [4-1:0] node48644;
	wire [4-1:0] node48647;
	wire [4-1:0] node48650;
	wire [4-1:0] node48651;
	wire [4-1:0] node48652;
	wire [4-1:0] node48653;
	wire [4-1:0] node48654;
	wire [4-1:0] node48658;
	wire [4-1:0] node48659;
	wire [4-1:0] node48662;
	wire [4-1:0] node48665;
	wire [4-1:0] node48666;
	wire [4-1:0] node48667;
	wire [4-1:0] node48670;
	wire [4-1:0] node48673;
	wire [4-1:0] node48674;
	wire [4-1:0] node48677;
	wire [4-1:0] node48680;
	wire [4-1:0] node48681;
	wire [4-1:0] node48682;
	wire [4-1:0] node48683;
	wire [4-1:0] node48686;
	wire [4-1:0] node48689;
	wire [4-1:0] node48691;
	wire [4-1:0] node48694;
	wire [4-1:0] node48695;
	wire [4-1:0] node48696;
	wire [4-1:0] node48699;
	wire [4-1:0] node48702;
	wire [4-1:0] node48703;
	wire [4-1:0] node48706;
	wire [4-1:0] node48709;
	wire [4-1:0] node48710;
	wire [4-1:0] node48711;
	wire [4-1:0] node48712;
	wire [4-1:0] node48713;
	wire [4-1:0] node48714;
	wire [4-1:0] node48715;
	wire [4-1:0] node48718;
	wire [4-1:0] node48721;
	wire [4-1:0] node48723;
	wire [4-1:0] node48726;
	wire [4-1:0] node48727;
	wire [4-1:0] node48728;
	wire [4-1:0] node48731;
	wire [4-1:0] node48734;
	wire [4-1:0] node48736;
	wire [4-1:0] node48739;
	wire [4-1:0] node48740;
	wire [4-1:0] node48741;
	wire [4-1:0] node48742;
	wire [4-1:0] node48745;
	wire [4-1:0] node48748;
	wire [4-1:0] node48749;
	wire [4-1:0] node48752;
	wire [4-1:0] node48755;
	wire [4-1:0] node48756;
	wire [4-1:0] node48757;
	wire [4-1:0] node48760;
	wire [4-1:0] node48763;
	wire [4-1:0] node48764;
	wire [4-1:0] node48767;
	wire [4-1:0] node48770;
	wire [4-1:0] node48771;
	wire [4-1:0] node48772;
	wire [4-1:0] node48773;
	wire [4-1:0] node48774;
	wire [4-1:0] node48777;
	wire [4-1:0] node48780;
	wire [4-1:0] node48781;
	wire [4-1:0] node48784;
	wire [4-1:0] node48787;
	wire [4-1:0] node48788;
	wire [4-1:0] node48789;
	wire [4-1:0] node48792;
	wire [4-1:0] node48795;
	wire [4-1:0] node48797;
	wire [4-1:0] node48800;
	wire [4-1:0] node48801;
	wire [4-1:0] node48802;
	wire [4-1:0] node48803;
	wire [4-1:0] node48806;
	wire [4-1:0] node48809;
	wire [4-1:0] node48811;
	wire [4-1:0] node48814;
	wire [4-1:0] node48815;
	wire [4-1:0] node48816;
	wire [4-1:0] node48819;
	wire [4-1:0] node48822;
	wire [4-1:0] node48823;
	wire [4-1:0] node48826;
	wire [4-1:0] node48829;
	wire [4-1:0] node48830;
	wire [4-1:0] node48831;
	wire [4-1:0] node48832;
	wire [4-1:0] node48833;
	wire [4-1:0] node48835;
	wire [4-1:0] node48838;
	wire [4-1:0] node48840;
	wire [4-1:0] node48843;
	wire [4-1:0] node48844;
	wire [4-1:0] node48845;
	wire [4-1:0] node48848;
	wire [4-1:0] node48851;
	wire [4-1:0] node48852;
	wire [4-1:0] node48856;
	wire [4-1:0] node48857;
	wire [4-1:0] node48858;
	wire [4-1:0] node48859;
	wire [4-1:0] node48863;
	wire [4-1:0] node48864;
	wire [4-1:0] node48868;
	wire [4-1:0] node48869;
	wire [4-1:0] node48870;
	wire [4-1:0] node48874;
	wire [4-1:0] node48875;
	wire [4-1:0] node48879;
	wire [4-1:0] node48880;
	wire [4-1:0] node48881;
	wire [4-1:0] node48882;
	wire [4-1:0] node48884;
	wire [4-1:0] node48887;
	wire [4-1:0] node48888;
	wire [4-1:0] node48891;
	wire [4-1:0] node48894;
	wire [4-1:0] node48895;
	wire [4-1:0] node48896;
	wire [4-1:0] node48899;
	wire [4-1:0] node48902;
	wire [4-1:0] node48903;
	wire [4-1:0] node48907;
	wire [4-1:0] node48908;
	wire [4-1:0] node48909;
	wire [4-1:0] node48910;
	wire [4-1:0] node48914;
	wire [4-1:0] node48915;
	wire [4-1:0] node48919;
	wire [4-1:0] node48920;
	wire [4-1:0] node48921;
	wire [4-1:0] node48925;
	wire [4-1:0] node48926;
	wire [4-1:0] node48930;
	wire [4-1:0] node48931;
	wire [4-1:0] node48932;
	wire [4-1:0] node48933;
	wire [4-1:0] node48934;
	wire [4-1:0] node48935;
	wire [4-1:0] node48936;
	wire [4-1:0] node48937;
	wire [4-1:0] node48940;
	wire [4-1:0] node48943;
	wire [4-1:0] node48944;
	wire [4-1:0] node48947;
	wire [4-1:0] node48950;
	wire [4-1:0] node48951;
	wire [4-1:0] node48952;
	wire [4-1:0] node48955;
	wire [4-1:0] node48958;
	wire [4-1:0] node48959;
	wire [4-1:0] node48962;
	wire [4-1:0] node48965;
	wire [4-1:0] node48966;
	wire [4-1:0] node48967;
	wire [4-1:0] node48968;
	wire [4-1:0] node48972;
	wire [4-1:0] node48973;
	wire [4-1:0] node48977;
	wire [4-1:0] node48978;
	wire [4-1:0] node48979;
	wire [4-1:0] node48983;
	wire [4-1:0] node48984;
	wire [4-1:0] node48988;
	wire [4-1:0] node48989;
	wire [4-1:0] node48990;
	wire [4-1:0] node48991;
	wire [4-1:0] node48992;
	wire [4-1:0] node48995;
	wire [4-1:0] node48998;
	wire [4-1:0] node48999;
	wire [4-1:0] node49002;
	wire [4-1:0] node49005;
	wire [4-1:0] node49006;
	wire [4-1:0] node49008;
	wire [4-1:0] node49011;
	wire [4-1:0] node49012;
	wire [4-1:0] node49015;
	wire [4-1:0] node49018;
	wire [4-1:0] node49019;
	wire [4-1:0] node49020;
	wire [4-1:0] node49021;
	wire [4-1:0] node49025;
	wire [4-1:0] node49026;
	wire [4-1:0] node49030;
	wire [4-1:0] node49031;
	wire [4-1:0] node49032;
	wire [4-1:0] node49036;
	wire [4-1:0] node49037;
	wire [4-1:0] node49041;
	wire [4-1:0] node49042;
	wire [4-1:0] node49043;
	wire [4-1:0] node49044;
	wire [4-1:0] node49045;
	wire [4-1:0] node49046;
	wire [4-1:0] node49049;
	wire [4-1:0] node49052;
	wire [4-1:0] node49053;
	wire [4-1:0] node49056;
	wire [4-1:0] node49059;
	wire [4-1:0] node49060;
	wire [4-1:0] node49061;
	wire [4-1:0] node49064;
	wire [4-1:0] node49067;
	wire [4-1:0] node49069;
	wire [4-1:0] node49072;
	wire [4-1:0] node49073;
	wire [4-1:0] node49074;
	wire [4-1:0] node49075;
	wire [4-1:0] node49079;
	wire [4-1:0] node49080;
	wire [4-1:0] node49084;
	wire [4-1:0] node49085;
	wire [4-1:0] node49086;
	wire [4-1:0] node49090;
	wire [4-1:0] node49091;
	wire [4-1:0] node49095;
	wire [4-1:0] node49096;
	wire [4-1:0] node49097;
	wire [4-1:0] node49098;
	wire [4-1:0] node49099;
	wire [4-1:0] node49102;
	wire [4-1:0] node49105;
	wire [4-1:0] node49106;
	wire [4-1:0] node49110;
	wire [4-1:0] node49111;
	wire [4-1:0] node49112;
	wire [4-1:0] node49116;
	wire [4-1:0] node49117;
	wire [4-1:0] node49121;
	wire [4-1:0] node49122;
	wire [4-1:0] node49123;
	wire [4-1:0] node49124;
	wire [4-1:0] node49128;
	wire [4-1:0] node49129;
	wire [4-1:0] node49133;
	wire [4-1:0] node49134;
	wire [4-1:0] node49135;
	wire [4-1:0] node49139;
	wire [4-1:0] node49140;
	wire [4-1:0] node49144;
	wire [4-1:0] node49145;
	wire [4-1:0] node49146;
	wire [4-1:0] node49147;
	wire [4-1:0] node49148;
	wire [4-1:0] node49149;
	wire [4-1:0] node49150;
	wire [4-1:0] node49153;
	wire [4-1:0] node49156;
	wire [4-1:0] node49157;
	wire [4-1:0] node49160;
	wire [4-1:0] node49163;
	wire [4-1:0] node49164;
	wire [4-1:0] node49165;
	wire [4-1:0] node49168;
	wire [4-1:0] node49171;
	wire [4-1:0] node49172;
	wire [4-1:0] node49175;
	wire [4-1:0] node49178;
	wire [4-1:0] node49179;
	wire [4-1:0] node49180;
	wire [4-1:0] node49181;
	wire [4-1:0] node49184;
	wire [4-1:0] node49187;
	wire [4-1:0] node49188;
	wire [4-1:0] node49191;
	wire [4-1:0] node49194;
	wire [4-1:0] node49195;
	wire [4-1:0] node49196;
	wire [4-1:0] node49199;
	wire [4-1:0] node49202;
	wire [4-1:0] node49203;
	wire [4-1:0] node49206;
	wire [4-1:0] node49209;
	wire [4-1:0] node49210;
	wire [4-1:0] node49211;
	wire [4-1:0] node49212;
	wire [4-1:0] node49213;
	wire [4-1:0] node49216;
	wire [4-1:0] node49219;
	wire [4-1:0] node49220;
	wire [4-1:0] node49223;
	wire [4-1:0] node49226;
	wire [4-1:0] node49227;
	wire [4-1:0] node49228;
	wire [4-1:0] node49231;
	wire [4-1:0] node49234;
	wire [4-1:0] node49235;
	wire [4-1:0] node49238;
	wire [4-1:0] node49241;
	wire [4-1:0] node49242;
	wire [4-1:0] node49243;
	wire [4-1:0] node49244;
	wire [4-1:0] node49247;
	wire [4-1:0] node49250;
	wire [4-1:0] node49251;
	wire [4-1:0] node49254;
	wire [4-1:0] node49257;
	wire [4-1:0] node49258;
	wire [4-1:0] node49259;
	wire [4-1:0] node49262;
	wire [4-1:0] node49265;
	wire [4-1:0] node49266;
	wire [4-1:0] node49269;
	wire [4-1:0] node49272;
	wire [4-1:0] node49273;
	wire [4-1:0] node49274;
	wire [4-1:0] node49275;
	wire [4-1:0] node49276;
	wire [4-1:0] node49277;
	wire [4-1:0] node49280;
	wire [4-1:0] node49283;
	wire [4-1:0] node49284;
	wire [4-1:0] node49287;
	wire [4-1:0] node49290;
	wire [4-1:0] node49291;
	wire [4-1:0] node49292;
	wire [4-1:0] node49295;
	wire [4-1:0] node49298;
	wire [4-1:0] node49299;
	wire [4-1:0] node49303;
	wire [4-1:0] node49304;
	wire [4-1:0] node49305;
	wire [4-1:0] node49306;
	wire [4-1:0] node49309;
	wire [4-1:0] node49312;
	wire [4-1:0] node49313;
	wire [4-1:0] node49316;
	wire [4-1:0] node49319;
	wire [4-1:0] node49320;
	wire [4-1:0] node49321;
	wire [4-1:0] node49324;
	wire [4-1:0] node49327;
	wire [4-1:0] node49329;
	wire [4-1:0] node49332;
	wire [4-1:0] node49333;
	wire [4-1:0] node49334;
	wire [4-1:0] node49335;
	wire [4-1:0] node49336;
	wire [4-1:0] node49339;
	wire [4-1:0] node49342;
	wire [4-1:0] node49343;
	wire [4-1:0] node49347;
	wire [4-1:0] node49348;
	wire [4-1:0] node49349;
	wire [4-1:0] node49352;
	wire [4-1:0] node49355;
	wire [4-1:0] node49356;
	wire [4-1:0] node49359;
	wire [4-1:0] node49362;
	wire [4-1:0] node49363;
	wire [4-1:0] node49364;
	wire [4-1:0] node49365;
	wire [4-1:0] node49368;
	wire [4-1:0] node49371;
	wire [4-1:0] node49372;
	wire [4-1:0] node49375;
	wire [4-1:0] node49378;
	wire [4-1:0] node49379;
	wire [4-1:0] node49380;
	wire [4-1:0] node49383;
	wire [4-1:0] node49386;
	wire [4-1:0] node49387;
	wire [4-1:0] node49390;
	wire [4-1:0] node49393;
	wire [4-1:0] node49394;
	wire [4-1:0] node49395;
	wire [4-1:0] node49396;
	wire [4-1:0] node49397;
	wire [4-1:0] node49398;
	wire [4-1:0] node49399;
	wire [4-1:0] node49400;
	wire [4-1:0] node49401;
	wire [4-1:0] node49404;
	wire [4-1:0] node49407;
	wire [4-1:0] node49408;
	wire [4-1:0] node49411;
	wire [4-1:0] node49414;
	wire [4-1:0] node49415;
	wire [4-1:0] node49416;
	wire [4-1:0] node49419;
	wire [4-1:0] node49422;
	wire [4-1:0] node49423;
	wire [4-1:0] node49426;
	wire [4-1:0] node49429;
	wire [4-1:0] node49430;
	wire [4-1:0] node49431;
	wire [4-1:0] node49432;
	wire [4-1:0] node49435;
	wire [4-1:0] node49438;
	wire [4-1:0] node49439;
	wire [4-1:0] node49443;
	wire [4-1:0] node49444;
	wire [4-1:0] node49446;
	wire [4-1:0] node49449;
	wire [4-1:0] node49450;
	wire [4-1:0] node49453;
	wire [4-1:0] node49456;
	wire [4-1:0] node49457;
	wire [4-1:0] node49458;
	wire [4-1:0] node49459;
	wire [4-1:0] node49460;
	wire [4-1:0] node49463;
	wire [4-1:0] node49466;
	wire [4-1:0] node49467;
	wire [4-1:0] node49470;
	wire [4-1:0] node49473;
	wire [4-1:0] node49474;
	wire [4-1:0] node49475;
	wire [4-1:0] node49478;
	wire [4-1:0] node49481;
	wire [4-1:0] node49482;
	wire [4-1:0] node49485;
	wire [4-1:0] node49488;
	wire [4-1:0] node49489;
	wire [4-1:0] node49490;
	wire [4-1:0] node49491;
	wire [4-1:0] node49495;
	wire [4-1:0] node49496;
	wire [4-1:0] node49500;
	wire [4-1:0] node49501;
	wire [4-1:0] node49502;
	wire [4-1:0] node49506;
	wire [4-1:0] node49507;
	wire [4-1:0] node49511;
	wire [4-1:0] node49512;
	wire [4-1:0] node49513;
	wire [4-1:0] node49514;
	wire [4-1:0] node49515;
	wire [4-1:0] node49516;
	wire [4-1:0] node49520;
	wire [4-1:0] node49521;
	wire [4-1:0] node49525;
	wire [4-1:0] node49526;
	wire [4-1:0] node49527;
	wire [4-1:0] node49530;
	wire [4-1:0] node49533;
	wire [4-1:0] node49534;
	wire [4-1:0] node49537;
	wire [4-1:0] node49540;
	wire [4-1:0] node49541;
	wire [4-1:0] node49542;
	wire [4-1:0] node49543;
	wire [4-1:0] node49547;
	wire [4-1:0] node49548;
	wire [4-1:0] node49552;
	wire [4-1:0] node49553;
	wire [4-1:0] node49556;
	wire [4-1:0] node49557;
	wire [4-1:0] node49561;
	wire [4-1:0] node49562;
	wire [4-1:0] node49563;
	wire [4-1:0] node49564;
	wire [4-1:0] node49565;
	wire [4-1:0] node49568;
	wire [4-1:0] node49571;
	wire [4-1:0] node49573;
	wire [4-1:0] node49576;
	wire [4-1:0] node49577;
	wire [4-1:0] node49578;
	wire [4-1:0] node49581;
	wire [4-1:0] node49584;
	wire [4-1:0] node49585;
	wire [4-1:0] node49588;
	wire [4-1:0] node49591;
	wire [4-1:0] node49592;
	wire [4-1:0] node49593;
	wire [4-1:0] node49594;
	wire [4-1:0] node49597;
	wire [4-1:0] node49600;
	wire [4-1:0] node49601;
	wire [4-1:0] node49604;
	wire [4-1:0] node49607;
	wire [4-1:0] node49608;
	wire [4-1:0] node49611;
	wire [4-1:0] node49614;
	wire [4-1:0] node49615;
	wire [4-1:0] node49616;
	wire [4-1:0] node49617;
	wire [4-1:0] node49618;
	wire [4-1:0] node49619;
	wire [4-1:0] node49620;
	wire [4-1:0] node49623;
	wire [4-1:0] node49626;
	wire [4-1:0] node49627;
	wire [4-1:0] node49630;
	wire [4-1:0] node49633;
	wire [4-1:0] node49634;
	wire [4-1:0] node49635;
	wire [4-1:0] node49638;
	wire [4-1:0] node49641;
	wire [4-1:0] node49642;
	wire [4-1:0] node49645;
	wire [4-1:0] node49648;
	wire [4-1:0] node49649;
	wire [4-1:0] node49650;
	wire [4-1:0] node49651;
	wire [4-1:0] node49655;
	wire [4-1:0] node49656;
	wire [4-1:0] node49660;
	wire [4-1:0] node49661;
	wire [4-1:0] node49662;
	wire [4-1:0] node49666;
	wire [4-1:0] node49667;
	wire [4-1:0] node49671;
	wire [4-1:0] node49672;
	wire [4-1:0] node49673;
	wire [4-1:0] node49674;
	wire [4-1:0] node49675;
	wire [4-1:0] node49678;
	wire [4-1:0] node49681;
	wire [4-1:0] node49683;
	wire [4-1:0] node49686;
	wire [4-1:0] node49687;
	wire [4-1:0] node49688;
	wire [4-1:0] node49692;
	wire [4-1:0] node49693;
	wire [4-1:0] node49696;
	wire [4-1:0] node49699;
	wire [4-1:0] node49700;
	wire [4-1:0] node49701;
	wire [4-1:0] node49704;
	wire [4-1:0] node49705;
	wire [4-1:0] node49709;
	wire [4-1:0] node49710;
	wire [4-1:0] node49711;
	wire [4-1:0] node49715;
	wire [4-1:0] node49716;
	wire [4-1:0] node49720;
	wire [4-1:0] node49721;
	wire [4-1:0] node49722;
	wire [4-1:0] node49723;
	wire [4-1:0] node49724;
	wire [4-1:0] node49725;
	wire [4-1:0] node49728;
	wire [4-1:0] node49731;
	wire [4-1:0] node49732;
	wire [4-1:0] node49735;
	wire [4-1:0] node49738;
	wire [4-1:0] node49739;
	wire [4-1:0] node49740;
	wire [4-1:0] node49744;
	wire [4-1:0] node49745;
	wire [4-1:0] node49749;
	wire [4-1:0] node49750;
	wire [4-1:0] node49751;
	wire [4-1:0] node49752;
	wire [4-1:0] node49755;
	wire [4-1:0] node49758;
	wire [4-1:0] node49759;
	wire [4-1:0] node49762;
	wire [4-1:0] node49765;
	wire [4-1:0] node49766;
	wire [4-1:0] node49767;
	wire [4-1:0] node49770;
	wire [4-1:0] node49773;
	wire [4-1:0] node49776;
	wire [4-1:0] node49777;
	wire [4-1:0] node49778;
	wire [4-1:0] node49779;
	wire [4-1:0] node49780;
	wire [4-1:0] node49783;
	wire [4-1:0] node49786;
	wire [4-1:0] node49787;
	wire [4-1:0] node49790;
	wire [4-1:0] node49793;
	wire [4-1:0] node49794;
	wire [4-1:0] node49795;
	wire [4-1:0] node49798;
	wire [4-1:0] node49801;
	wire [4-1:0] node49802;
	wire [4-1:0] node49805;
	wire [4-1:0] node49808;
	wire [4-1:0] node49809;
	wire [4-1:0] node49810;
	wire [4-1:0] node49811;
	wire [4-1:0] node49814;
	wire [4-1:0] node49817;
	wire [4-1:0] node49819;
	wire [4-1:0] node49822;
	wire [4-1:0] node49823;
	wire [4-1:0] node49826;
	wire [4-1:0] node49829;
	wire [4-1:0] node49830;
	wire [4-1:0] node49831;
	wire [4-1:0] node49832;
	wire [4-1:0] node49833;
	wire [4-1:0] node49834;
	wire [4-1:0] node49835;
	wire [4-1:0] node49836;
	wire [4-1:0] node49839;
	wire [4-1:0] node49842;
	wire [4-1:0] node49843;
	wire [4-1:0] node49847;
	wire [4-1:0] node49848;
	wire [4-1:0] node49849;
	wire [4-1:0] node49852;
	wire [4-1:0] node49855;
	wire [4-1:0] node49856;
	wire [4-1:0] node49859;
	wire [4-1:0] node49862;
	wire [4-1:0] node49863;
	wire [4-1:0] node49864;
	wire [4-1:0] node49865;
	wire [4-1:0] node49869;
	wire [4-1:0] node49870;
	wire [4-1:0] node49874;
	wire [4-1:0] node49875;
	wire [4-1:0] node49876;
	wire [4-1:0] node49880;
	wire [4-1:0] node49881;
	wire [4-1:0] node49885;
	wire [4-1:0] node49886;
	wire [4-1:0] node49887;
	wire [4-1:0] node49888;
	wire [4-1:0] node49889;
	wire [4-1:0] node49892;
	wire [4-1:0] node49895;
	wire [4-1:0] node49896;
	wire [4-1:0] node49899;
	wire [4-1:0] node49902;
	wire [4-1:0] node49903;
	wire [4-1:0] node49904;
	wire [4-1:0] node49907;
	wire [4-1:0] node49910;
	wire [4-1:0] node49911;
	wire [4-1:0] node49914;
	wire [4-1:0] node49917;
	wire [4-1:0] node49918;
	wire [4-1:0] node49919;
	wire [4-1:0] node49920;
	wire [4-1:0] node49924;
	wire [4-1:0] node49925;
	wire [4-1:0] node49928;
	wire [4-1:0] node49931;
	wire [4-1:0] node49932;
	wire [4-1:0] node49933;
	wire [4-1:0] node49937;
	wire [4-1:0] node49938;
	wire [4-1:0] node49941;
	wire [4-1:0] node49944;
	wire [4-1:0] node49945;
	wire [4-1:0] node49946;
	wire [4-1:0] node49947;
	wire [4-1:0] node49948;
	wire [4-1:0] node49949;
	wire [4-1:0] node49953;
	wire [4-1:0] node49954;
	wire [4-1:0] node49957;
	wire [4-1:0] node49960;
	wire [4-1:0] node49961;
	wire [4-1:0] node49962;
	wire [4-1:0] node49965;
	wire [4-1:0] node49968;
	wire [4-1:0] node49969;
	wire [4-1:0] node49972;
	wire [4-1:0] node49975;
	wire [4-1:0] node49976;
	wire [4-1:0] node49977;
	wire [4-1:0] node49980;
	wire [4-1:0] node49981;
	wire [4-1:0] node49985;
	wire [4-1:0] node49986;
	wire [4-1:0] node49987;
	wire [4-1:0] node49991;
	wire [4-1:0] node49992;
	wire [4-1:0] node49996;
	wire [4-1:0] node49997;
	wire [4-1:0] node49998;
	wire [4-1:0] node49999;
	wire [4-1:0] node50000;
	wire [4-1:0] node50003;
	wire [4-1:0] node50006;
	wire [4-1:0] node50007;
	wire [4-1:0] node50010;
	wire [4-1:0] node50013;
	wire [4-1:0] node50014;
	wire [4-1:0] node50015;
	wire [4-1:0] node50019;
	wire [4-1:0] node50020;
	wire [4-1:0] node50023;
	wire [4-1:0] node50026;
	wire [4-1:0] node50027;
	wire [4-1:0] node50028;
	wire [4-1:0] node50029;
	wire [4-1:0] node50032;
	wire [4-1:0] node50035;
	wire [4-1:0] node50036;
	wire [4-1:0] node50039;
	wire [4-1:0] node50042;
	wire [4-1:0] node50043;
	wire [4-1:0] node50044;
	wire [4-1:0] node50047;
	wire [4-1:0] node50050;
	wire [4-1:0] node50051;
	wire [4-1:0] node50054;
	wire [4-1:0] node50057;
	wire [4-1:0] node50058;
	wire [4-1:0] node50059;
	wire [4-1:0] node50060;
	wire [4-1:0] node50061;
	wire [4-1:0] node50062;
	wire [4-1:0] node50063;
	wire [4-1:0] node50066;
	wire [4-1:0] node50069;
	wire [4-1:0] node50070;
	wire [4-1:0] node50073;
	wire [4-1:0] node50076;
	wire [4-1:0] node50077;
	wire [4-1:0] node50078;
	wire [4-1:0] node50081;
	wire [4-1:0] node50084;
	wire [4-1:0] node50085;
	wire [4-1:0] node50088;
	wire [4-1:0] node50091;
	wire [4-1:0] node50092;
	wire [4-1:0] node50093;
	wire [4-1:0] node50094;
	wire [4-1:0] node50098;
	wire [4-1:0] node50099;
	wire [4-1:0] node50103;
	wire [4-1:0] node50104;
	wire [4-1:0] node50105;
	wire [4-1:0] node50109;
	wire [4-1:0] node50110;
	wire [4-1:0] node50114;
	wire [4-1:0] node50115;
	wire [4-1:0] node50116;
	wire [4-1:0] node50117;
	wire [4-1:0] node50119;
	wire [4-1:0] node50122;
	wire [4-1:0] node50123;
	wire [4-1:0] node50126;
	wire [4-1:0] node50129;
	wire [4-1:0] node50130;
	wire [4-1:0] node50132;
	wire [4-1:0] node50135;
	wire [4-1:0] node50138;
	wire [4-1:0] node50139;
	wire [4-1:0] node50140;
	wire [4-1:0] node50141;
	wire [4-1:0] node50145;
	wire [4-1:0] node50146;
	wire [4-1:0] node50149;
	wire [4-1:0] node50152;
	wire [4-1:0] node50153;
	wire [4-1:0] node50156;
	wire [4-1:0] node50159;
	wire [4-1:0] node50160;
	wire [4-1:0] node50161;
	wire [4-1:0] node50162;
	wire [4-1:0] node50163;
	wire [4-1:0] node50165;
	wire [4-1:0] node50168;
	wire [4-1:0] node50169;
	wire [4-1:0] node50172;
	wire [4-1:0] node50175;
	wire [4-1:0] node50176;
	wire [4-1:0] node50178;
	wire [4-1:0] node50181;
	wire [4-1:0] node50182;
	wire [4-1:0] node50185;
	wire [4-1:0] node50188;
	wire [4-1:0] node50189;
	wire [4-1:0] node50190;
	wire [4-1:0] node50191;
	wire [4-1:0] node50194;
	wire [4-1:0] node50197;
	wire [4-1:0] node50198;
	wire [4-1:0] node50202;
	wire [4-1:0] node50203;
	wire [4-1:0] node50204;
	wire [4-1:0] node50207;
	wire [4-1:0] node50210;
	wire [4-1:0] node50211;
	wire [4-1:0] node50214;
	wire [4-1:0] node50217;
	wire [4-1:0] node50218;
	wire [4-1:0] node50219;
	wire [4-1:0] node50220;
	wire [4-1:0] node50221;
	wire [4-1:0] node50224;
	wire [4-1:0] node50227;
	wire [4-1:0] node50228;
	wire [4-1:0] node50231;
	wire [4-1:0] node50234;
	wire [4-1:0] node50235;
	wire [4-1:0] node50237;
	wire [4-1:0] node50240;
	wire [4-1:0] node50242;
	wire [4-1:0] node50245;
	wire [4-1:0] node50246;
	wire [4-1:0] node50247;
	wire [4-1:0] node50248;
	wire [4-1:0] node50251;
	wire [4-1:0] node50254;
	wire [4-1:0] node50255;
	wire [4-1:0] node50258;
	wire [4-1:0] node50261;
	wire [4-1:0] node50262;
	wire [4-1:0] node50265;
	wire [4-1:0] node50268;
	wire [4-1:0] node50269;
	wire [4-1:0] node50270;
	wire [4-1:0] node50271;
	wire [4-1:0] node50272;
	wire [4-1:0] node50273;
	wire [4-1:0] node50274;
	wire [4-1:0] node50275;
	wire [4-1:0] node50276;
	wire [4-1:0] node50277;
	wire [4-1:0] node50278;
	wire [4-1:0] node50279;
	wire [4-1:0] node50282;
	wire [4-1:0] node50285;
	wire [4-1:0] node50286;
	wire [4-1:0] node50289;
	wire [4-1:0] node50292;
	wire [4-1:0] node50293;
	wire [4-1:0] node50295;
	wire [4-1:0] node50298;
	wire [4-1:0] node50299;
	wire [4-1:0] node50302;
	wire [4-1:0] node50305;
	wire [4-1:0] node50306;
	wire [4-1:0] node50307;
	wire [4-1:0] node50308;
	wire [4-1:0] node50311;
	wire [4-1:0] node50314;
	wire [4-1:0] node50316;
	wire [4-1:0] node50319;
	wire [4-1:0] node50320;
	wire [4-1:0] node50321;
	wire [4-1:0] node50325;
	wire [4-1:0] node50326;
	wire [4-1:0] node50329;
	wire [4-1:0] node50332;
	wire [4-1:0] node50333;
	wire [4-1:0] node50334;
	wire [4-1:0] node50335;
	wire [4-1:0] node50336;
	wire [4-1:0] node50339;
	wire [4-1:0] node50342;
	wire [4-1:0] node50343;
	wire [4-1:0] node50346;
	wire [4-1:0] node50349;
	wire [4-1:0] node50350;
	wire [4-1:0] node50351;
	wire [4-1:0] node50354;
	wire [4-1:0] node50357;
	wire [4-1:0] node50358;
	wire [4-1:0] node50361;
	wire [4-1:0] node50364;
	wire [4-1:0] node50365;
	wire [4-1:0] node50366;
	wire [4-1:0] node50367;
	wire [4-1:0] node50371;
	wire [4-1:0] node50372;
	wire [4-1:0] node50376;
	wire [4-1:0] node50377;
	wire [4-1:0] node50378;
	wire [4-1:0] node50382;
	wire [4-1:0] node50383;
	wire [4-1:0] node50387;
	wire [4-1:0] node50388;
	wire [4-1:0] node50389;
	wire [4-1:0] node50390;
	wire [4-1:0] node50391;
	wire [4-1:0] node50392;
	wire [4-1:0] node50395;
	wire [4-1:0] node50398;
	wire [4-1:0] node50399;
	wire [4-1:0] node50402;
	wire [4-1:0] node50405;
	wire [4-1:0] node50406;
	wire [4-1:0] node50407;
	wire [4-1:0] node50410;
	wire [4-1:0] node50413;
	wire [4-1:0] node50414;
	wire [4-1:0] node50418;
	wire [4-1:0] node50419;
	wire [4-1:0] node50420;
	wire [4-1:0] node50421;
	wire [4-1:0] node50425;
	wire [4-1:0] node50426;
	wire [4-1:0] node50430;
	wire [4-1:0] node50431;
	wire [4-1:0] node50432;
	wire [4-1:0] node50436;
	wire [4-1:0] node50437;
	wire [4-1:0] node50441;
	wire [4-1:0] node50442;
	wire [4-1:0] node50443;
	wire [4-1:0] node50444;
	wire [4-1:0] node50445;
	wire [4-1:0] node50448;
	wire [4-1:0] node50451;
	wire [4-1:0] node50452;
	wire [4-1:0] node50456;
	wire [4-1:0] node50457;
	wire [4-1:0] node50458;
	wire [4-1:0] node50462;
	wire [4-1:0] node50463;
	wire [4-1:0] node50466;
	wire [4-1:0] node50469;
	wire [4-1:0] node50470;
	wire [4-1:0] node50471;
	wire [4-1:0] node50472;
	wire [4-1:0] node50476;
	wire [4-1:0] node50477;
	wire [4-1:0] node50481;
	wire [4-1:0] node50482;
	wire [4-1:0] node50483;
	wire [4-1:0] node50487;
	wire [4-1:0] node50488;
	wire [4-1:0] node50492;
	wire [4-1:0] node50493;
	wire [4-1:0] node50494;
	wire [4-1:0] node50495;
	wire [4-1:0] node50496;
	wire [4-1:0] node50497;
	wire [4-1:0] node50498;
	wire [4-1:0] node50501;
	wire [4-1:0] node50504;
	wire [4-1:0] node50505;
	wire [4-1:0] node50508;
	wire [4-1:0] node50511;
	wire [4-1:0] node50512;
	wire [4-1:0] node50515;
	wire [4-1:0] node50516;
	wire [4-1:0] node50519;
	wire [4-1:0] node50522;
	wire [4-1:0] node50523;
	wire [4-1:0] node50524;
	wire [4-1:0] node50525;
	wire [4-1:0] node50529;
	wire [4-1:0] node50530;
	wire [4-1:0] node50534;
	wire [4-1:0] node50535;
	wire [4-1:0] node50536;
	wire [4-1:0] node50540;
	wire [4-1:0] node50541;
	wire [4-1:0] node50545;
	wire [4-1:0] node50546;
	wire [4-1:0] node50547;
	wire [4-1:0] node50548;
	wire [4-1:0] node50549;
	wire [4-1:0] node50552;
	wire [4-1:0] node50555;
	wire [4-1:0] node50556;
	wire [4-1:0] node50559;
	wire [4-1:0] node50562;
	wire [4-1:0] node50563;
	wire [4-1:0] node50564;
	wire [4-1:0] node50567;
	wire [4-1:0] node50570;
	wire [4-1:0] node50571;
	wire [4-1:0] node50574;
	wire [4-1:0] node50577;
	wire [4-1:0] node50578;
	wire [4-1:0] node50579;
	wire [4-1:0] node50580;
	wire [4-1:0] node50583;
	wire [4-1:0] node50586;
	wire [4-1:0] node50587;
	wire [4-1:0] node50590;
	wire [4-1:0] node50593;
	wire [4-1:0] node50594;
	wire [4-1:0] node50595;
	wire [4-1:0] node50598;
	wire [4-1:0] node50601;
	wire [4-1:0] node50602;
	wire [4-1:0] node50605;
	wire [4-1:0] node50608;
	wire [4-1:0] node50609;
	wire [4-1:0] node50610;
	wire [4-1:0] node50611;
	wire [4-1:0] node50612;
	wire [4-1:0] node50614;
	wire [4-1:0] node50617;
	wire [4-1:0] node50618;
	wire [4-1:0] node50621;
	wire [4-1:0] node50624;
	wire [4-1:0] node50625;
	wire [4-1:0] node50626;
	wire [4-1:0] node50629;
	wire [4-1:0] node50632;
	wire [4-1:0] node50633;
	wire [4-1:0] node50636;
	wire [4-1:0] node50639;
	wire [4-1:0] node50640;
	wire [4-1:0] node50641;
	wire [4-1:0] node50642;
	wire [4-1:0] node50645;
	wire [4-1:0] node50648;
	wire [4-1:0] node50649;
	wire [4-1:0] node50652;
	wire [4-1:0] node50655;
	wire [4-1:0] node50656;
	wire [4-1:0] node50657;
	wire [4-1:0] node50660;
	wire [4-1:0] node50663;
	wire [4-1:0] node50664;
	wire [4-1:0] node50667;
	wire [4-1:0] node50670;
	wire [4-1:0] node50671;
	wire [4-1:0] node50672;
	wire [4-1:0] node50673;
	wire [4-1:0] node50674;
	wire [4-1:0] node50677;
	wire [4-1:0] node50680;
	wire [4-1:0] node50681;
	wire [4-1:0] node50684;
	wire [4-1:0] node50687;
	wire [4-1:0] node50688;
	wire [4-1:0] node50690;
	wire [4-1:0] node50693;
	wire [4-1:0] node50694;
	wire [4-1:0] node50697;
	wire [4-1:0] node50700;
	wire [4-1:0] node50701;
	wire [4-1:0] node50702;
	wire [4-1:0] node50703;
	wire [4-1:0] node50707;
	wire [4-1:0] node50708;
	wire [4-1:0] node50712;
	wire [4-1:0] node50713;
	wire [4-1:0] node50714;
	wire [4-1:0] node50718;
	wire [4-1:0] node50719;
	wire [4-1:0] node50723;
	wire [4-1:0] node50724;
	wire [4-1:0] node50725;
	wire [4-1:0] node50726;
	wire [4-1:0] node50727;
	wire [4-1:0] node50728;
	wire [4-1:0] node50729;
	wire [4-1:0] node50730;
	wire [4-1:0] node50733;
	wire [4-1:0] node50736;
	wire [4-1:0] node50737;
	wire [4-1:0] node50740;
	wire [4-1:0] node50743;
	wire [4-1:0] node50744;
	wire [4-1:0] node50745;
	wire [4-1:0] node50749;
	wire [4-1:0] node50750;
	wire [4-1:0] node50754;
	wire [4-1:0] node50755;
	wire [4-1:0] node50756;
	wire [4-1:0] node50757;
	wire [4-1:0] node50760;
	wire [4-1:0] node50763;
	wire [4-1:0] node50764;
	wire [4-1:0] node50767;
	wire [4-1:0] node50770;
	wire [4-1:0] node50771;
	wire [4-1:0] node50772;
	wire [4-1:0] node50775;
	wire [4-1:0] node50778;
	wire [4-1:0] node50779;
	wire [4-1:0] node50782;
	wire [4-1:0] node50785;
	wire [4-1:0] node50786;
	wire [4-1:0] node50787;
	wire [4-1:0] node50788;
	wire [4-1:0] node50789;
	wire [4-1:0] node50792;
	wire [4-1:0] node50795;
	wire [4-1:0] node50796;
	wire [4-1:0] node50799;
	wire [4-1:0] node50802;
	wire [4-1:0] node50803;
	wire [4-1:0] node50804;
	wire [4-1:0] node50807;
	wire [4-1:0] node50810;
	wire [4-1:0] node50811;
	wire [4-1:0] node50815;
	wire [4-1:0] node50816;
	wire [4-1:0] node50817;
	wire [4-1:0] node50818;
	wire [4-1:0] node50822;
	wire [4-1:0] node50823;
	wire [4-1:0] node50827;
	wire [4-1:0] node50828;
	wire [4-1:0] node50829;
	wire [4-1:0] node50833;
	wire [4-1:0] node50834;
	wire [4-1:0] node50838;
	wire [4-1:0] node50839;
	wire [4-1:0] node50840;
	wire [4-1:0] node50841;
	wire [4-1:0] node50842;
	wire [4-1:0] node50843;
	wire [4-1:0] node50846;
	wire [4-1:0] node50849;
	wire [4-1:0] node50850;
	wire [4-1:0] node50854;
	wire [4-1:0] node50855;
	wire [4-1:0] node50856;
	wire [4-1:0] node50860;
	wire [4-1:0] node50861;
	wire [4-1:0] node50864;
	wire [4-1:0] node50867;
	wire [4-1:0] node50868;
	wire [4-1:0] node50869;
	wire [4-1:0] node50870;
	wire [4-1:0] node50874;
	wire [4-1:0] node50875;
	wire [4-1:0] node50879;
	wire [4-1:0] node50880;
	wire [4-1:0] node50881;
	wire [4-1:0] node50885;
	wire [4-1:0] node50886;
	wire [4-1:0] node50890;
	wire [4-1:0] node50891;
	wire [4-1:0] node50892;
	wire [4-1:0] node50893;
	wire [4-1:0] node50894;
	wire [4-1:0] node50897;
	wire [4-1:0] node50900;
	wire [4-1:0] node50901;
	wire [4-1:0] node50904;
	wire [4-1:0] node50907;
	wire [4-1:0] node50908;
	wire [4-1:0] node50909;
	wire [4-1:0] node50912;
	wire [4-1:0] node50915;
	wire [4-1:0] node50916;
	wire [4-1:0] node50919;
	wire [4-1:0] node50922;
	wire [4-1:0] node50923;
	wire [4-1:0] node50924;
	wire [4-1:0] node50925;
	wire [4-1:0] node50929;
	wire [4-1:0] node50930;
	wire [4-1:0] node50934;
	wire [4-1:0] node50935;
	wire [4-1:0] node50936;
	wire [4-1:0] node50940;
	wire [4-1:0] node50941;
	wire [4-1:0] node50945;
	wire [4-1:0] node50946;
	wire [4-1:0] node50947;
	wire [4-1:0] node50948;
	wire [4-1:0] node50949;
	wire [4-1:0] node50950;
	wire [4-1:0] node50951;
	wire [4-1:0] node50954;
	wire [4-1:0] node50957;
	wire [4-1:0] node50958;
	wire [4-1:0] node50961;
	wire [4-1:0] node50964;
	wire [4-1:0] node50965;
	wire [4-1:0] node50966;
	wire [4-1:0] node50969;
	wire [4-1:0] node50972;
	wire [4-1:0] node50974;
	wire [4-1:0] node50977;
	wire [4-1:0] node50978;
	wire [4-1:0] node50979;
	wire [4-1:0] node50980;
	wire [4-1:0] node50983;
	wire [4-1:0] node50986;
	wire [4-1:0] node50988;
	wire [4-1:0] node50991;
	wire [4-1:0] node50992;
	wire [4-1:0] node50993;
	wire [4-1:0] node50996;
	wire [4-1:0] node50999;
	wire [4-1:0] node51000;
	wire [4-1:0] node51003;
	wire [4-1:0] node51006;
	wire [4-1:0] node51007;
	wire [4-1:0] node51008;
	wire [4-1:0] node51009;
	wire [4-1:0] node51010;
	wire [4-1:0] node51013;
	wire [4-1:0] node51016;
	wire [4-1:0] node51017;
	wire [4-1:0] node51020;
	wire [4-1:0] node51023;
	wire [4-1:0] node51024;
	wire [4-1:0] node51025;
	wire [4-1:0] node51028;
	wire [4-1:0] node51031;
	wire [4-1:0] node51032;
	wire [4-1:0] node51036;
	wire [4-1:0] node51037;
	wire [4-1:0] node51038;
	wire [4-1:0] node51039;
	wire [4-1:0] node51042;
	wire [4-1:0] node51045;
	wire [4-1:0] node51046;
	wire [4-1:0] node51049;
	wire [4-1:0] node51052;
	wire [4-1:0] node51053;
	wire [4-1:0] node51054;
	wire [4-1:0] node51057;
	wire [4-1:0] node51060;
	wire [4-1:0] node51061;
	wire [4-1:0] node51064;
	wire [4-1:0] node51067;
	wire [4-1:0] node51068;
	wire [4-1:0] node51069;
	wire [4-1:0] node51070;
	wire [4-1:0] node51071;
	wire [4-1:0] node51072;
	wire [4-1:0] node51075;
	wire [4-1:0] node51078;
	wire [4-1:0] node51080;
	wire [4-1:0] node51083;
	wire [4-1:0] node51084;
	wire [4-1:0] node51085;
	wire [4-1:0] node51088;
	wire [4-1:0] node51091;
	wire [4-1:0] node51092;
	wire [4-1:0] node51095;
	wire [4-1:0] node51098;
	wire [4-1:0] node51099;
	wire [4-1:0] node51100;
	wire [4-1:0] node51101;
	wire [4-1:0] node51104;
	wire [4-1:0] node51107;
	wire [4-1:0] node51108;
	wire [4-1:0] node51111;
	wire [4-1:0] node51114;
	wire [4-1:0] node51115;
	wire [4-1:0] node51117;
	wire [4-1:0] node51120;
	wire [4-1:0] node51121;
	wire [4-1:0] node51124;
	wire [4-1:0] node51127;
	wire [4-1:0] node51128;
	wire [4-1:0] node51129;
	wire [4-1:0] node51130;
	wire [4-1:0] node51131;
	wire [4-1:0] node51134;
	wire [4-1:0] node51137;
	wire [4-1:0] node51139;
	wire [4-1:0] node51142;
	wire [4-1:0] node51143;
	wire [4-1:0] node51144;
	wire [4-1:0] node51147;
	wire [4-1:0] node51150;
	wire [4-1:0] node51151;
	wire [4-1:0] node51154;
	wire [4-1:0] node51157;
	wire [4-1:0] node51158;
	wire [4-1:0] node51159;
	wire [4-1:0] node51160;
	wire [4-1:0] node51164;
	wire [4-1:0] node51166;
	wire [4-1:0] node51169;
	wire [4-1:0] node51170;
	wire [4-1:0] node51171;
	wire [4-1:0] node51174;
	wire [4-1:0] node51177;
	wire [4-1:0] node51178;
	wire [4-1:0] node51181;
	wire [4-1:0] node51184;
	wire [4-1:0] node51185;
	wire [4-1:0] node51186;
	wire [4-1:0] node51187;
	wire [4-1:0] node51188;
	wire [4-1:0] node51189;
	wire [4-1:0] node51190;
	wire [4-1:0] node51191;
	wire [4-1:0] node51192;
	wire [4-1:0] node51196;
	wire [4-1:0] node51197;
	wire [4-1:0] node51201;
	wire [4-1:0] node51202;
	wire [4-1:0] node51203;
	wire [4-1:0] node51206;
	wire [4-1:0] node51209;
	wire [4-1:0] node51210;
	wire [4-1:0] node51213;
	wire [4-1:0] node51216;
	wire [4-1:0] node51217;
	wire [4-1:0] node51218;
	wire [4-1:0] node51219;
	wire [4-1:0] node51222;
	wire [4-1:0] node51225;
	wire [4-1:0] node51226;
	wire [4-1:0] node51229;
	wire [4-1:0] node51232;
	wire [4-1:0] node51233;
	wire [4-1:0] node51234;
	wire [4-1:0] node51238;
	wire [4-1:0] node51239;
	wire [4-1:0] node51242;
	wire [4-1:0] node51245;
	wire [4-1:0] node51246;
	wire [4-1:0] node51247;
	wire [4-1:0] node51248;
	wire [4-1:0] node51249;
	wire [4-1:0] node51252;
	wire [4-1:0] node51255;
	wire [4-1:0] node51256;
	wire [4-1:0] node51259;
	wire [4-1:0] node51262;
	wire [4-1:0] node51263;
	wire [4-1:0] node51265;
	wire [4-1:0] node51268;
	wire [4-1:0] node51269;
	wire [4-1:0] node51272;
	wire [4-1:0] node51275;
	wire [4-1:0] node51276;
	wire [4-1:0] node51277;
	wire [4-1:0] node51278;
	wire [4-1:0] node51281;
	wire [4-1:0] node51284;
	wire [4-1:0] node51285;
	wire [4-1:0] node51288;
	wire [4-1:0] node51291;
	wire [4-1:0] node51292;
	wire [4-1:0] node51293;
	wire [4-1:0] node51296;
	wire [4-1:0] node51299;
	wire [4-1:0] node51300;
	wire [4-1:0] node51303;
	wire [4-1:0] node51306;
	wire [4-1:0] node51307;
	wire [4-1:0] node51308;
	wire [4-1:0] node51309;
	wire [4-1:0] node51310;
	wire [4-1:0] node51311;
	wire [4-1:0] node51314;
	wire [4-1:0] node51317;
	wire [4-1:0] node51318;
	wire [4-1:0] node51321;
	wire [4-1:0] node51324;
	wire [4-1:0] node51325;
	wire [4-1:0] node51326;
	wire [4-1:0] node51329;
	wire [4-1:0] node51332;
	wire [4-1:0] node51333;
	wire [4-1:0] node51336;
	wire [4-1:0] node51339;
	wire [4-1:0] node51340;
	wire [4-1:0] node51341;
	wire [4-1:0] node51342;
	wire [4-1:0] node51345;
	wire [4-1:0] node51348;
	wire [4-1:0] node51349;
	wire [4-1:0] node51352;
	wire [4-1:0] node51355;
	wire [4-1:0] node51356;
	wire [4-1:0] node51357;
	wire [4-1:0] node51360;
	wire [4-1:0] node51363;
	wire [4-1:0] node51364;
	wire [4-1:0] node51367;
	wire [4-1:0] node51370;
	wire [4-1:0] node51371;
	wire [4-1:0] node51372;
	wire [4-1:0] node51373;
	wire [4-1:0] node51374;
	wire [4-1:0] node51377;
	wire [4-1:0] node51380;
	wire [4-1:0] node51381;
	wire [4-1:0] node51384;
	wire [4-1:0] node51387;
	wire [4-1:0] node51388;
	wire [4-1:0] node51389;
	wire [4-1:0] node51392;
	wire [4-1:0] node51395;
	wire [4-1:0] node51396;
	wire [4-1:0] node51399;
	wire [4-1:0] node51402;
	wire [4-1:0] node51403;
	wire [4-1:0] node51404;
	wire [4-1:0] node51405;
	wire [4-1:0] node51408;
	wire [4-1:0] node51411;
	wire [4-1:0] node51412;
	wire [4-1:0] node51415;
	wire [4-1:0] node51418;
	wire [4-1:0] node51419;
	wire [4-1:0] node51420;
	wire [4-1:0] node51423;
	wire [4-1:0] node51426;
	wire [4-1:0] node51427;
	wire [4-1:0] node51430;
	wire [4-1:0] node51433;
	wire [4-1:0] node51434;
	wire [4-1:0] node51435;
	wire [4-1:0] node51436;
	wire [4-1:0] node51437;
	wire [4-1:0] node51438;
	wire [4-1:0] node51439;
	wire [4-1:0] node51442;
	wire [4-1:0] node51445;
	wire [4-1:0] node51446;
	wire [4-1:0] node51449;
	wire [4-1:0] node51452;
	wire [4-1:0] node51453;
	wire [4-1:0] node51454;
	wire [4-1:0] node51457;
	wire [4-1:0] node51460;
	wire [4-1:0] node51461;
	wire [4-1:0] node51464;
	wire [4-1:0] node51467;
	wire [4-1:0] node51468;
	wire [4-1:0] node51469;
	wire [4-1:0] node51470;
	wire [4-1:0] node51473;
	wire [4-1:0] node51476;
	wire [4-1:0] node51477;
	wire [4-1:0] node51480;
	wire [4-1:0] node51483;
	wire [4-1:0] node51484;
	wire [4-1:0] node51487;
	wire [4-1:0] node51490;
	wire [4-1:0] node51491;
	wire [4-1:0] node51492;
	wire [4-1:0] node51493;
	wire [4-1:0] node51494;
	wire [4-1:0] node51497;
	wire [4-1:0] node51500;
	wire [4-1:0] node51501;
	wire [4-1:0] node51504;
	wire [4-1:0] node51507;
	wire [4-1:0] node51508;
	wire [4-1:0] node51510;
	wire [4-1:0] node51513;
	wire [4-1:0] node51514;
	wire [4-1:0] node51517;
	wire [4-1:0] node51520;
	wire [4-1:0] node51521;
	wire [4-1:0] node51522;
	wire [4-1:0] node51523;
	wire [4-1:0] node51527;
	wire [4-1:0] node51528;
	wire [4-1:0] node51532;
	wire [4-1:0] node51533;
	wire [4-1:0] node51534;
	wire [4-1:0] node51538;
	wire [4-1:0] node51539;
	wire [4-1:0] node51543;
	wire [4-1:0] node51544;
	wire [4-1:0] node51545;
	wire [4-1:0] node51546;
	wire [4-1:0] node51547;
	wire [4-1:0] node51548;
	wire [4-1:0] node51551;
	wire [4-1:0] node51554;
	wire [4-1:0] node51555;
	wire [4-1:0] node51558;
	wire [4-1:0] node51561;
	wire [4-1:0] node51562;
	wire [4-1:0] node51563;
	wire [4-1:0] node51566;
	wire [4-1:0] node51569;
	wire [4-1:0] node51570;
	wire [4-1:0] node51573;
	wire [4-1:0] node51576;
	wire [4-1:0] node51577;
	wire [4-1:0] node51578;
	wire [4-1:0] node51579;
	wire [4-1:0] node51582;
	wire [4-1:0] node51585;
	wire [4-1:0] node51586;
	wire [4-1:0] node51589;
	wire [4-1:0] node51592;
	wire [4-1:0] node51593;
	wire [4-1:0] node51594;
	wire [4-1:0] node51597;
	wire [4-1:0] node51600;
	wire [4-1:0] node51601;
	wire [4-1:0] node51604;
	wire [4-1:0] node51607;
	wire [4-1:0] node51608;
	wire [4-1:0] node51609;
	wire [4-1:0] node51610;
	wire [4-1:0] node51611;
	wire [4-1:0] node51614;
	wire [4-1:0] node51617;
	wire [4-1:0] node51618;
	wire [4-1:0] node51621;
	wire [4-1:0] node51624;
	wire [4-1:0] node51625;
	wire [4-1:0] node51627;
	wire [4-1:0] node51630;
	wire [4-1:0] node51631;
	wire [4-1:0] node51634;
	wire [4-1:0] node51637;
	wire [4-1:0] node51638;
	wire [4-1:0] node51639;
	wire [4-1:0] node51640;
	wire [4-1:0] node51643;
	wire [4-1:0] node51646;
	wire [4-1:0] node51647;
	wire [4-1:0] node51650;
	wire [4-1:0] node51653;
	wire [4-1:0] node51654;
	wire [4-1:0] node51655;
	wire [4-1:0] node51658;
	wire [4-1:0] node51661;
	wire [4-1:0] node51662;
	wire [4-1:0] node51665;
	wire [4-1:0] node51668;
	wire [4-1:0] node51669;
	wire [4-1:0] node51670;
	wire [4-1:0] node51671;
	wire [4-1:0] node51672;
	wire [4-1:0] node51673;
	wire [4-1:0] node51674;
	wire [4-1:0] node51675;
	wire [4-1:0] node51678;
	wire [4-1:0] node51681;
	wire [4-1:0] node51682;
	wire [4-1:0] node51685;
	wire [4-1:0] node51688;
	wire [4-1:0] node51689;
	wire [4-1:0] node51690;
	wire [4-1:0] node51693;
	wire [4-1:0] node51696;
	wire [4-1:0] node51697;
	wire [4-1:0] node51700;
	wire [4-1:0] node51703;
	wire [4-1:0] node51704;
	wire [4-1:0] node51705;
	wire [4-1:0] node51706;
	wire [4-1:0] node51709;
	wire [4-1:0] node51712;
	wire [4-1:0] node51713;
	wire [4-1:0] node51716;
	wire [4-1:0] node51719;
	wire [4-1:0] node51720;
	wire [4-1:0] node51722;
	wire [4-1:0] node51725;
	wire [4-1:0] node51726;
	wire [4-1:0] node51729;
	wire [4-1:0] node51732;
	wire [4-1:0] node51733;
	wire [4-1:0] node51734;
	wire [4-1:0] node51735;
	wire [4-1:0] node51736;
	wire [4-1:0] node51739;
	wire [4-1:0] node51742;
	wire [4-1:0] node51743;
	wire [4-1:0] node51746;
	wire [4-1:0] node51749;
	wire [4-1:0] node51750;
	wire [4-1:0] node51751;
	wire [4-1:0] node51755;
	wire [4-1:0] node51756;
	wire [4-1:0] node51759;
	wire [4-1:0] node51762;
	wire [4-1:0] node51763;
	wire [4-1:0] node51764;
	wire [4-1:0] node51765;
	wire [4-1:0] node51769;
	wire [4-1:0] node51770;
	wire [4-1:0] node51774;
	wire [4-1:0] node51775;
	wire [4-1:0] node51776;
	wire [4-1:0] node51780;
	wire [4-1:0] node51781;
	wire [4-1:0] node51785;
	wire [4-1:0] node51786;
	wire [4-1:0] node51787;
	wire [4-1:0] node51788;
	wire [4-1:0] node51789;
	wire [4-1:0] node51791;
	wire [4-1:0] node51794;
	wire [4-1:0] node51796;
	wire [4-1:0] node51799;
	wire [4-1:0] node51800;
	wire [4-1:0] node51801;
	wire [4-1:0] node51805;
	wire [4-1:0] node51806;
	wire [4-1:0] node51809;
	wire [4-1:0] node51812;
	wire [4-1:0] node51813;
	wire [4-1:0] node51814;
	wire [4-1:0] node51815;
	wire [4-1:0] node51818;
	wire [4-1:0] node51821;
	wire [4-1:0] node51822;
	wire [4-1:0] node51825;
	wire [4-1:0] node51828;
	wire [4-1:0] node51829;
	wire [4-1:0] node51830;
	wire [4-1:0] node51833;
	wire [4-1:0] node51836;
	wire [4-1:0] node51837;
	wire [4-1:0] node51840;
	wire [4-1:0] node51843;
	wire [4-1:0] node51844;
	wire [4-1:0] node51845;
	wire [4-1:0] node51846;
	wire [4-1:0] node51847;
	wire [4-1:0] node51850;
	wire [4-1:0] node51853;
	wire [4-1:0] node51854;
	wire [4-1:0] node51857;
	wire [4-1:0] node51860;
	wire [4-1:0] node51861;
	wire [4-1:0] node51862;
	wire [4-1:0] node51865;
	wire [4-1:0] node51868;
	wire [4-1:0] node51869;
	wire [4-1:0] node51873;
	wire [4-1:0] node51874;
	wire [4-1:0] node51875;
	wire [4-1:0] node51876;
	wire [4-1:0] node51880;
	wire [4-1:0] node51881;
	wire [4-1:0] node51885;
	wire [4-1:0] node51886;
	wire [4-1:0] node51887;
	wire [4-1:0] node51891;
	wire [4-1:0] node51892;
	wire [4-1:0] node51896;
	wire [4-1:0] node51897;
	wire [4-1:0] node51898;
	wire [4-1:0] node51899;
	wire [4-1:0] node51900;
	wire [4-1:0] node51901;
	wire [4-1:0] node51902;
	wire [4-1:0] node51905;
	wire [4-1:0] node51908;
	wire [4-1:0] node51909;
	wire [4-1:0] node51912;
	wire [4-1:0] node51915;
	wire [4-1:0] node51916;
	wire [4-1:0] node51918;
	wire [4-1:0] node51921;
	wire [4-1:0] node51922;
	wire [4-1:0] node51925;
	wire [4-1:0] node51928;
	wire [4-1:0] node51929;
	wire [4-1:0] node51930;
	wire [4-1:0] node51931;
	wire [4-1:0] node51934;
	wire [4-1:0] node51937;
	wire [4-1:0] node51938;
	wire [4-1:0] node51941;
	wire [4-1:0] node51944;
	wire [4-1:0] node51945;
	wire [4-1:0] node51946;
	wire [4-1:0] node51949;
	wire [4-1:0] node51952;
	wire [4-1:0] node51953;
	wire [4-1:0] node51956;
	wire [4-1:0] node51959;
	wire [4-1:0] node51960;
	wire [4-1:0] node51961;
	wire [4-1:0] node51962;
	wire [4-1:0] node51964;
	wire [4-1:0] node51967;
	wire [4-1:0] node51968;
	wire [4-1:0] node51972;
	wire [4-1:0] node51973;
	wire [4-1:0] node51974;
	wire [4-1:0] node51977;
	wire [4-1:0] node51980;
	wire [4-1:0] node51981;
	wire [4-1:0] node51984;
	wire [4-1:0] node51987;
	wire [4-1:0] node51988;
	wire [4-1:0] node51989;
	wire [4-1:0] node51990;
	wire [4-1:0] node51993;
	wire [4-1:0] node51996;
	wire [4-1:0] node51997;
	wire [4-1:0] node52000;
	wire [4-1:0] node52003;
	wire [4-1:0] node52004;
	wire [4-1:0] node52005;
	wire [4-1:0] node52008;
	wire [4-1:0] node52011;
	wire [4-1:0] node52012;
	wire [4-1:0] node52015;
	wire [4-1:0] node52018;
	wire [4-1:0] node52019;
	wire [4-1:0] node52020;
	wire [4-1:0] node52021;
	wire [4-1:0] node52022;
	wire [4-1:0] node52023;
	wire [4-1:0] node52026;
	wire [4-1:0] node52029;
	wire [4-1:0] node52030;
	wire [4-1:0] node52033;
	wire [4-1:0] node52036;
	wire [4-1:0] node52037;
	wire [4-1:0] node52038;
	wire [4-1:0] node52041;
	wire [4-1:0] node52044;
	wire [4-1:0] node52045;
	wire [4-1:0] node52048;
	wire [4-1:0] node52051;
	wire [4-1:0] node52052;
	wire [4-1:0] node52053;
	wire [4-1:0] node52054;
	wire [4-1:0] node52057;
	wire [4-1:0] node52060;
	wire [4-1:0] node52061;
	wire [4-1:0] node52064;
	wire [4-1:0] node52067;
	wire [4-1:0] node52068;
	wire [4-1:0] node52069;
	wire [4-1:0] node52072;
	wire [4-1:0] node52075;
	wire [4-1:0] node52076;
	wire [4-1:0] node52079;
	wire [4-1:0] node52082;
	wire [4-1:0] node52083;
	wire [4-1:0] node52084;
	wire [4-1:0] node52085;
	wire [4-1:0] node52086;
	wire [4-1:0] node52089;
	wire [4-1:0] node52092;
	wire [4-1:0] node52093;
	wire [4-1:0] node52096;
	wire [4-1:0] node52099;
	wire [4-1:0] node52100;
	wire [4-1:0] node52101;
	wire [4-1:0] node52104;
	wire [4-1:0] node52107;
	wire [4-1:0] node52108;
	wire [4-1:0] node52111;
	wire [4-1:0] node52114;
	wire [4-1:0] node52115;
	wire [4-1:0] node52116;
	wire [4-1:0] node52117;
	wire [4-1:0] node52120;
	wire [4-1:0] node52123;
	wire [4-1:0] node52124;
	wire [4-1:0] node52127;
	wire [4-1:0] node52130;
	wire [4-1:0] node52131;
	wire [4-1:0] node52132;
	wire [4-1:0] node52135;
	wire [4-1:0] node52138;
	wire [4-1:0] node52139;
	wire [4-1:0] node52142;
	wire [4-1:0] node52145;
	wire [4-1:0] node52146;
	wire [4-1:0] node52147;
	wire [4-1:0] node52148;
	wire [4-1:0] node52149;
	wire [4-1:0] node52150;
	wire [4-1:0] node52151;
	wire [4-1:0] node52152;
	wire [4-1:0] node52153;
	wire [4-1:0] node52154;
	wire [4-1:0] node52157;
	wire [4-1:0] node52160;
	wire [4-1:0] node52161;
	wire [4-1:0] node52164;
	wire [4-1:0] node52167;
	wire [4-1:0] node52168;
	wire [4-1:0] node52169;
	wire [4-1:0] node52173;
	wire [4-1:0] node52174;
	wire [4-1:0] node52177;
	wire [4-1:0] node52180;
	wire [4-1:0] node52181;
	wire [4-1:0] node52182;
	wire [4-1:0] node52183;
	wire [4-1:0] node52186;
	wire [4-1:0] node52189;
	wire [4-1:0] node52190;
	wire [4-1:0] node52193;
	wire [4-1:0] node52196;
	wire [4-1:0] node52197;
	wire [4-1:0] node52200;
	wire [4-1:0] node52203;
	wire [4-1:0] node52204;
	wire [4-1:0] node52205;
	wire [4-1:0] node52206;
	wire [4-1:0] node52207;
	wire [4-1:0] node52210;
	wire [4-1:0] node52213;
	wire [4-1:0] node52214;
	wire [4-1:0] node52217;
	wire [4-1:0] node52220;
	wire [4-1:0] node52221;
	wire [4-1:0] node52222;
	wire [4-1:0] node52226;
	wire [4-1:0] node52228;
	wire [4-1:0] node52231;
	wire [4-1:0] node52232;
	wire [4-1:0] node52233;
	wire [4-1:0] node52234;
	wire [4-1:0] node52238;
	wire [4-1:0] node52239;
	wire [4-1:0] node52243;
	wire [4-1:0] node52244;
	wire [4-1:0] node52245;
	wire [4-1:0] node52249;
	wire [4-1:0] node52250;
	wire [4-1:0] node52254;
	wire [4-1:0] node52255;
	wire [4-1:0] node52256;
	wire [4-1:0] node52257;
	wire [4-1:0] node52258;
	wire [4-1:0] node52259;
	wire [4-1:0] node52262;
	wire [4-1:0] node52265;
	wire [4-1:0] node52267;
	wire [4-1:0] node52270;
	wire [4-1:0] node52271;
	wire [4-1:0] node52272;
	wire [4-1:0] node52276;
	wire [4-1:0] node52277;
	wire [4-1:0] node52280;
	wire [4-1:0] node52283;
	wire [4-1:0] node52284;
	wire [4-1:0] node52285;
	wire [4-1:0] node52286;
	wire [4-1:0] node52290;
	wire [4-1:0] node52291;
	wire [4-1:0] node52295;
	wire [4-1:0] node52296;
	wire [4-1:0] node52297;
	wire [4-1:0] node52301;
	wire [4-1:0] node52302;
	wire [4-1:0] node52306;
	wire [4-1:0] node52307;
	wire [4-1:0] node52308;
	wire [4-1:0] node52309;
	wire [4-1:0] node52310;
	wire [4-1:0] node52313;
	wire [4-1:0] node52316;
	wire [4-1:0] node52317;
	wire [4-1:0] node52320;
	wire [4-1:0] node52323;
	wire [4-1:0] node52324;
	wire [4-1:0] node52326;
	wire [4-1:0] node52329;
	wire [4-1:0] node52330;
	wire [4-1:0] node52334;
	wire [4-1:0] node52335;
	wire [4-1:0] node52336;
	wire [4-1:0] node52337;
	wire [4-1:0] node52341;
	wire [4-1:0] node52342;
	wire [4-1:0] node52346;
	wire [4-1:0] node52347;
	wire [4-1:0] node52348;
	wire [4-1:0] node52352;
	wire [4-1:0] node52353;
	wire [4-1:0] node52357;
	wire [4-1:0] node52358;
	wire [4-1:0] node52359;
	wire [4-1:0] node52360;
	wire [4-1:0] node52361;
	wire [4-1:0] node52362;
	wire [4-1:0] node52364;
	wire [4-1:0] node52367;
	wire [4-1:0] node52369;
	wire [4-1:0] node52372;
	wire [4-1:0] node52373;
	wire [4-1:0] node52374;
	wire [4-1:0] node52378;
	wire [4-1:0] node52379;
	wire [4-1:0] node52382;
	wire [4-1:0] node52385;
	wire [4-1:0] node52386;
	wire [4-1:0] node52387;
	wire [4-1:0] node52388;
	wire [4-1:0] node52391;
	wire [4-1:0] node52394;
	wire [4-1:0] node52395;
	wire [4-1:0] node52398;
	wire [4-1:0] node52401;
	wire [4-1:0] node52402;
	wire [4-1:0] node52403;
	wire [4-1:0] node52406;
	wire [4-1:0] node52409;
	wire [4-1:0] node52410;
	wire [4-1:0] node52413;
	wire [4-1:0] node52416;
	wire [4-1:0] node52417;
	wire [4-1:0] node52418;
	wire [4-1:0] node52419;
	wire [4-1:0] node52421;
	wire [4-1:0] node52424;
	wire [4-1:0] node52425;
	wire [4-1:0] node52428;
	wire [4-1:0] node52431;
	wire [4-1:0] node52432;
	wire [4-1:0] node52433;
	wire [4-1:0] node52436;
	wire [4-1:0] node52439;
	wire [4-1:0] node52441;
	wire [4-1:0] node52444;
	wire [4-1:0] node52445;
	wire [4-1:0] node52446;
	wire [4-1:0] node52447;
	wire [4-1:0] node52450;
	wire [4-1:0] node52453;
	wire [4-1:0] node52454;
	wire [4-1:0] node52458;
	wire [4-1:0] node52459;
	wire [4-1:0] node52462;
	wire [4-1:0] node52465;
	wire [4-1:0] node52466;
	wire [4-1:0] node52467;
	wire [4-1:0] node52468;
	wire [4-1:0] node52469;
	wire [4-1:0] node52470;
	wire [4-1:0] node52473;
	wire [4-1:0] node52476;
	wire [4-1:0] node52477;
	wire [4-1:0] node52480;
	wire [4-1:0] node52483;
	wire [4-1:0] node52484;
	wire [4-1:0] node52485;
	wire [4-1:0] node52488;
	wire [4-1:0] node52491;
	wire [4-1:0] node52492;
	wire [4-1:0] node52496;
	wire [4-1:0] node52497;
	wire [4-1:0] node52498;
	wire [4-1:0] node52499;
	wire [4-1:0] node52503;
	wire [4-1:0] node52504;
	wire [4-1:0] node52508;
	wire [4-1:0] node52509;
	wire [4-1:0] node52510;
	wire [4-1:0] node52514;
	wire [4-1:0] node52515;
	wire [4-1:0] node52519;
	wire [4-1:0] node52520;
	wire [4-1:0] node52521;
	wire [4-1:0] node52522;
	wire [4-1:0] node52523;
	wire [4-1:0] node52526;
	wire [4-1:0] node52529;
	wire [4-1:0] node52530;
	wire [4-1:0] node52533;
	wire [4-1:0] node52536;
	wire [4-1:0] node52537;
	wire [4-1:0] node52538;
	wire [4-1:0] node52541;
	wire [4-1:0] node52544;
	wire [4-1:0] node52545;
	wire [4-1:0] node52549;
	wire [4-1:0] node52550;
	wire [4-1:0] node52551;
	wire [4-1:0] node52552;
	wire [4-1:0] node52556;
	wire [4-1:0] node52557;
	wire [4-1:0] node52561;
	wire [4-1:0] node52562;
	wire [4-1:0] node52563;
	wire [4-1:0] node52567;
	wire [4-1:0] node52568;
	wire [4-1:0] node52572;
	wire [4-1:0] node52573;
	wire [4-1:0] node52574;
	wire [4-1:0] node52575;
	wire [4-1:0] node52576;
	wire [4-1:0] node52577;
	wire [4-1:0] node52578;
	wire [4-1:0] node52579;
	wire [4-1:0] node52582;
	wire [4-1:0] node52585;
	wire [4-1:0] node52587;
	wire [4-1:0] node52590;
	wire [4-1:0] node52591;
	wire [4-1:0] node52592;
	wire [4-1:0] node52595;
	wire [4-1:0] node52598;
	wire [4-1:0] node52599;
	wire [4-1:0] node52602;
	wire [4-1:0] node52605;
	wire [4-1:0] node52606;
	wire [4-1:0] node52607;
	wire [4-1:0] node52608;
	wire [4-1:0] node52611;
	wire [4-1:0] node52614;
	wire [4-1:0] node52615;
	wire [4-1:0] node52618;
	wire [4-1:0] node52621;
	wire [4-1:0] node52622;
	wire [4-1:0] node52625;
	wire [4-1:0] node52628;
	wire [4-1:0] node52629;
	wire [4-1:0] node52630;
	wire [4-1:0] node52631;
	wire [4-1:0] node52632;
	wire [4-1:0] node52635;
	wire [4-1:0] node52638;
	wire [4-1:0] node52639;
	wire [4-1:0] node52642;
	wire [4-1:0] node52645;
	wire [4-1:0] node52646;
	wire [4-1:0] node52647;
	wire [4-1:0] node52651;
	wire [4-1:0] node52652;
	wire [4-1:0] node52655;
	wire [4-1:0] node52658;
	wire [4-1:0] node52659;
	wire [4-1:0] node52660;
	wire [4-1:0] node52661;
	wire [4-1:0] node52664;
	wire [4-1:0] node52667;
	wire [4-1:0] node52668;
	wire [4-1:0] node52671;
	wire [4-1:0] node52674;
	wire [4-1:0] node52675;
	wire [4-1:0] node52677;
	wire [4-1:0] node52680;
	wire [4-1:0] node52681;
	wire [4-1:0] node52684;
	wire [4-1:0] node52687;
	wire [4-1:0] node52688;
	wire [4-1:0] node52689;
	wire [4-1:0] node52690;
	wire [4-1:0] node52691;
	wire [4-1:0] node52692;
	wire [4-1:0] node52696;
	wire [4-1:0] node52697;
	wire [4-1:0] node52700;
	wire [4-1:0] node52703;
	wire [4-1:0] node52704;
	wire [4-1:0] node52705;
	wire [4-1:0] node52708;
	wire [4-1:0] node52711;
	wire [4-1:0] node52712;
	wire [4-1:0] node52716;
	wire [4-1:0] node52717;
	wire [4-1:0] node52718;
	wire [4-1:0] node52719;
	wire [4-1:0] node52723;
	wire [4-1:0] node52724;
	wire [4-1:0] node52728;
	wire [4-1:0] node52729;
	wire [4-1:0] node52730;
	wire [4-1:0] node52734;
	wire [4-1:0] node52735;
	wire [4-1:0] node52739;
	wire [4-1:0] node52740;
	wire [4-1:0] node52741;
	wire [4-1:0] node52742;
	wire [4-1:0] node52743;
	wire [4-1:0] node52746;
	wire [4-1:0] node52749;
	wire [4-1:0] node52750;
	wire [4-1:0] node52754;
	wire [4-1:0] node52755;
	wire [4-1:0] node52756;
	wire [4-1:0] node52759;
	wire [4-1:0] node52762;
	wire [4-1:0] node52763;
	wire [4-1:0] node52766;
	wire [4-1:0] node52769;
	wire [4-1:0] node52770;
	wire [4-1:0] node52771;
	wire [4-1:0] node52772;
	wire [4-1:0] node52775;
	wire [4-1:0] node52778;
	wire [4-1:0] node52779;
	wire [4-1:0] node52782;
	wire [4-1:0] node52785;
	wire [4-1:0] node52786;
	wire [4-1:0] node52787;
	wire [4-1:0] node52790;
	wire [4-1:0] node52793;
	wire [4-1:0] node52794;
	wire [4-1:0] node52797;
	wire [4-1:0] node52800;
	wire [4-1:0] node52801;
	wire [4-1:0] node52802;
	wire [4-1:0] node52803;
	wire [4-1:0] node52804;
	wire [4-1:0] node52805;
	wire [4-1:0] node52806;
	wire [4-1:0] node52809;
	wire [4-1:0] node52812;
	wire [4-1:0] node52813;
	wire [4-1:0] node52817;
	wire [4-1:0] node52818;
	wire [4-1:0] node52819;
	wire [4-1:0] node52823;
	wire [4-1:0] node52824;
	wire [4-1:0] node52827;
	wire [4-1:0] node52830;
	wire [4-1:0] node52831;
	wire [4-1:0] node52832;
	wire [4-1:0] node52833;
	wire [4-1:0] node52836;
	wire [4-1:0] node52839;
	wire [4-1:0] node52840;
	wire [4-1:0] node52843;
	wire [4-1:0] node52846;
	wire [4-1:0] node52847;
	wire [4-1:0] node52848;
	wire [4-1:0] node52851;
	wire [4-1:0] node52854;
	wire [4-1:0] node52855;
	wire [4-1:0] node52858;
	wire [4-1:0] node52861;
	wire [4-1:0] node52862;
	wire [4-1:0] node52863;
	wire [4-1:0] node52864;
	wire [4-1:0] node52865;
	wire [4-1:0] node52868;
	wire [4-1:0] node52871;
	wire [4-1:0] node52872;
	wire [4-1:0] node52875;
	wire [4-1:0] node52878;
	wire [4-1:0] node52879;
	wire [4-1:0] node52880;
	wire [4-1:0] node52883;
	wire [4-1:0] node52886;
	wire [4-1:0] node52887;
	wire [4-1:0] node52890;
	wire [4-1:0] node52893;
	wire [4-1:0] node52894;
	wire [4-1:0] node52895;
	wire [4-1:0] node52896;
	wire [4-1:0] node52899;
	wire [4-1:0] node52902;
	wire [4-1:0] node52903;
	wire [4-1:0] node52906;
	wire [4-1:0] node52909;
	wire [4-1:0] node52910;
	wire [4-1:0] node52911;
	wire [4-1:0] node52914;
	wire [4-1:0] node52917;
	wire [4-1:0] node52918;
	wire [4-1:0] node52921;
	wire [4-1:0] node52924;
	wire [4-1:0] node52925;
	wire [4-1:0] node52926;
	wire [4-1:0] node52927;
	wire [4-1:0] node52928;
	wire [4-1:0] node52929;
	wire [4-1:0] node52932;
	wire [4-1:0] node52935;
	wire [4-1:0] node52936;
	wire [4-1:0] node52939;
	wire [4-1:0] node52942;
	wire [4-1:0] node52943;
	wire [4-1:0] node52946;
	wire [4-1:0] node52949;
	wire [4-1:0] node52950;
	wire [4-1:0] node52951;
	wire [4-1:0] node52953;
	wire [4-1:0] node52956;
	wire [4-1:0] node52957;
	wire [4-1:0] node52960;
	wire [4-1:0] node52963;
	wire [4-1:0] node52964;
	wire [4-1:0] node52967;
	wire [4-1:0] node52970;
	wire [4-1:0] node52971;
	wire [4-1:0] node52972;
	wire [4-1:0] node52973;
	wire [4-1:0] node52974;
	wire [4-1:0] node52977;
	wire [4-1:0] node52980;
	wire [4-1:0] node52982;
	wire [4-1:0] node52985;
	wire [4-1:0] node52986;
	wire [4-1:0] node52987;
	wire [4-1:0] node52990;
	wire [4-1:0] node52993;
	wire [4-1:0] node52994;
	wire [4-1:0] node52997;
	wire [4-1:0] node53000;
	wire [4-1:0] node53001;
	wire [4-1:0] node53002;
	wire [4-1:0] node53003;
	wire [4-1:0] node53006;
	wire [4-1:0] node53009;
	wire [4-1:0] node53010;
	wire [4-1:0] node53013;
	wire [4-1:0] node53016;
	wire [4-1:0] node53017;
	wire [4-1:0] node53018;
	wire [4-1:0] node53021;
	wire [4-1:0] node53024;
	wire [4-1:0] node53025;
	wire [4-1:0] node53028;
	wire [4-1:0] node53031;
	wire [4-1:0] node53032;
	wire [4-1:0] node53033;
	wire [4-1:0] node53034;
	wire [4-1:0] node53035;
	wire [4-1:0] node53036;
	wire [4-1:0] node53037;
	wire [4-1:0] node53038;
	wire [4-1:0] node53039;
	wire [4-1:0] node53043;
	wire [4-1:0] node53044;
	wire [4-1:0] node53047;
	wire [4-1:0] node53050;
	wire [4-1:0] node53051;
	wire [4-1:0] node53052;
	wire [4-1:0] node53055;
	wire [4-1:0] node53058;
	wire [4-1:0] node53059;
	wire [4-1:0] node53062;
	wire [4-1:0] node53065;
	wire [4-1:0] node53066;
	wire [4-1:0] node53067;
	wire [4-1:0] node53068;
	wire [4-1:0] node53071;
	wire [4-1:0] node53074;
	wire [4-1:0] node53075;
	wire [4-1:0] node53078;
	wire [4-1:0] node53081;
	wire [4-1:0] node53082;
	wire [4-1:0] node53084;
	wire [4-1:0] node53087;
	wire [4-1:0] node53088;
	wire [4-1:0] node53091;
	wire [4-1:0] node53094;
	wire [4-1:0] node53095;
	wire [4-1:0] node53096;
	wire [4-1:0] node53097;
	wire [4-1:0] node53098;
	wire [4-1:0] node53101;
	wire [4-1:0] node53104;
	wire [4-1:0] node53105;
	wire [4-1:0] node53108;
	wire [4-1:0] node53111;
	wire [4-1:0] node53112;
	wire [4-1:0] node53113;
	wire [4-1:0] node53117;
	wire [4-1:0] node53120;
	wire [4-1:0] node53121;
	wire [4-1:0] node53122;
	wire [4-1:0] node53124;
	wire [4-1:0] node53127;
	wire [4-1:0] node53128;
	wire [4-1:0] node53131;
	wire [4-1:0] node53134;
	wire [4-1:0] node53135;
	wire [4-1:0] node53136;
	wire [4-1:0] node53139;
	wire [4-1:0] node53142;
	wire [4-1:0] node53143;
	wire [4-1:0] node53146;
	wire [4-1:0] node53149;
	wire [4-1:0] node53150;
	wire [4-1:0] node53151;
	wire [4-1:0] node53152;
	wire [4-1:0] node53153;
	wire [4-1:0] node53154;
	wire [4-1:0] node53158;
	wire [4-1:0] node53159;
	wire [4-1:0] node53162;
	wire [4-1:0] node53165;
	wire [4-1:0] node53166;
	wire [4-1:0] node53167;
	wire [4-1:0] node53170;
	wire [4-1:0] node53173;
	wire [4-1:0] node53174;
	wire [4-1:0] node53177;
	wire [4-1:0] node53180;
	wire [4-1:0] node53181;
	wire [4-1:0] node53182;
	wire [4-1:0] node53183;
	wire [4-1:0] node53187;
	wire [4-1:0] node53188;
	wire [4-1:0] node53192;
	wire [4-1:0] node53193;
	wire [4-1:0] node53194;
	wire [4-1:0] node53198;
	wire [4-1:0] node53199;
	wire [4-1:0] node53203;
	wire [4-1:0] node53204;
	wire [4-1:0] node53205;
	wire [4-1:0] node53206;
	wire [4-1:0] node53207;
	wire [4-1:0] node53211;
	wire [4-1:0] node53212;
	wire [4-1:0] node53215;
	wire [4-1:0] node53218;
	wire [4-1:0] node53219;
	wire [4-1:0] node53220;
	wire [4-1:0] node53224;
	wire [4-1:0] node53225;
	wire [4-1:0] node53228;
	wire [4-1:0] node53231;
	wire [4-1:0] node53232;
	wire [4-1:0] node53233;
	wire [4-1:0] node53234;
	wire [4-1:0] node53238;
	wire [4-1:0] node53239;
	wire [4-1:0] node53243;
	wire [4-1:0] node53244;
	wire [4-1:0] node53245;
	wire [4-1:0] node53249;
	wire [4-1:0] node53250;
	wire [4-1:0] node53254;
	wire [4-1:0] node53255;
	wire [4-1:0] node53256;
	wire [4-1:0] node53257;
	wire [4-1:0] node53258;
	wire [4-1:0] node53259;
	wire [4-1:0] node53261;
	wire [4-1:0] node53264;
	wire [4-1:0] node53265;
	wire [4-1:0] node53268;
	wire [4-1:0] node53271;
	wire [4-1:0] node53272;
	wire [4-1:0] node53273;
	wire [4-1:0] node53276;
	wire [4-1:0] node53279;
	wire [4-1:0] node53281;
	wire [4-1:0] node53284;
	wire [4-1:0] node53285;
	wire [4-1:0] node53286;
	wire [4-1:0] node53287;
	wire [4-1:0] node53290;
	wire [4-1:0] node53293;
	wire [4-1:0] node53294;
	wire [4-1:0] node53298;
	wire [4-1:0] node53299;
	wire [4-1:0] node53300;
	wire [4-1:0] node53303;
	wire [4-1:0] node53306;
	wire [4-1:0] node53308;
	wire [4-1:0] node53311;
	wire [4-1:0] node53312;
	wire [4-1:0] node53313;
	wire [4-1:0] node53314;
	wire [4-1:0] node53315;
	wire [4-1:0] node53318;
	wire [4-1:0] node53321;
	wire [4-1:0] node53322;
	wire [4-1:0] node53325;
	wire [4-1:0] node53328;
	wire [4-1:0] node53329;
	wire [4-1:0] node53330;
	wire [4-1:0] node53334;
	wire [4-1:0] node53335;
	wire [4-1:0] node53338;
	wire [4-1:0] node53341;
	wire [4-1:0] node53342;
	wire [4-1:0] node53343;
	wire [4-1:0] node53344;
	wire [4-1:0] node53347;
	wire [4-1:0] node53350;
	wire [4-1:0] node53351;
	wire [4-1:0] node53354;
	wire [4-1:0] node53357;
	wire [4-1:0] node53358;
	wire [4-1:0] node53359;
	wire [4-1:0] node53362;
	wire [4-1:0] node53365;
	wire [4-1:0] node53366;
	wire [4-1:0] node53369;
	wire [4-1:0] node53372;
	wire [4-1:0] node53373;
	wire [4-1:0] node53374;
	wire [4-1:0] node53375;
	wire [4-1:0] node53376;
	wire [4-1:0] node53377;
	wire [4-1:0] node53380;
	wire [4-1:0] node53383;
	wire [4-1:0] node53384;
	wire [4-1:0] node53387;
	wire [4-1:0] node53390;
	wire [4-1:0] node53391;
	wire [4-1:0] node53393;
	wire [4-1:0] node53396;
	wire [4-1:0] node53397;
	wire [4-1:0] node53400;
	wire [4-1:0] node53403;
	wire [4-1:0] node53404;
	wire [4-1:0] node53405;
	wire [4-1:0] node53406;
	wire [4-1:0] node53410;
	wire [4-1:0] node53411;
	wire [4-1:0] node53415;
	wire [4-1:0] node53416;
	wire [4-1:0] node53417;
	wire [4-1:0] node53421;
	wire [4-1:0] node53422;
	wire [4-1:0] node53426;
	wire [4-1:0] node53427;
	wire [4-1:0] node53428;
	wire [4-1:0] node53429;
	wire [4-1:0] node53432;
	wire [4-1:0] node53433;
	wire [4-1:0] node53437;
	wire [4-1:0] node53438;
	wire [4-1:0] node53439;
	wire [4-1:0] node53442;
	wire [4-1:0] node53445;
	wire [4-1:0] node53447;
	wire [4-1:0] node53450;
	wire [4-1:0] node53451;
	wire [4-1:0] node53452;
	wire [4-1:0] node53453;
	wire [4-1:0] node53458;
	wire [4-1:0] node53459;
	wire [4-1:0] node53460;
	wire [4-1:0] node53464;
	wire [4-1:0] node53465;
	wire [4-1:0] node53469;
	wire [4-1:0] node53470;
	wire [4-1:0] node53471;
	wire [4-1:0] node53472;
	wire [4-1:0] node53473;
	wire [4-1:0] node53474;
	wire [4-1:0] node53475;
	wire [4-1:0] node53477;
	wire [4-1:0] node53480;
	wire [4-1:0] node53481;
	wire [4-1:0] node53484;
	wire [4-1:0] node53487;
	wire [4-1:0] node53488;
	wire [4-1:0] node53489;
	wire [4-1:0] node53492;
	wire [4-1:0] node53495;
	wire [4-1:0] node53496;
	wire [4-1:0] node53499;
	wire [4-1:0] node53502;
	wire [4-1:0] node53503;
	wire [4-1:0] node53504;
	wire [4-1:0] node53505;
	wire [4-1:0] node53509;
	wire [4-1:0] node53510;
	wire [4-1:0] node53514;
	wire [4-1:0] node53515;
	wire [4-1:0] node53516;
	wire [4-1:0] node53520;
	wire [4-1:0] node53521;
	wire [4-1:0] node53525;
	wire [4-1:0] node53526;
	wire [4-1:0] node53527;
	wire [4-1:0] node53528;
	wire [4-1:0] node53529;
	wire [4-1:0] node53532;
	wire [4-1:0] node53535;
	wire [4-1:0] node53536;
	wire [4-1:0] node53539;
	wire [4-1:0] node53542;
	wire [4-1:0] node53543;
	wire [4-1:0] node53545;
	wire [4-1:0] node53548;
	wire [4-1:0] node53550;
	wire [4-1:0] node53553;
	wire [4-1:0] node53554;
	wire [4-1:0] node53555;
	wire [4-1:0] node53556;
	wire [4-1:0] node53560;
	wire [4-1:0] node53561;
	wire [4-1:0] node53565;
	wire [4-1:0] node53566;
	wire [4-1:0] node53567;
	wire [4-1:0] node53571;
	wire [4-1:0] node53572;
	wire [4-1:0] node53576;
	wire [4-1:0] node53577;
	wire [4-1:0] node53578;
	wire [4-1:0] node53579;
	wire [4-1:0] node53580;
	wire [4-1:0] node53581;
	wire [4-1:0] node53584;
	wire [4-1:0] node53587;
	wire [4-1:0] node53589;
	wire [4-1:0] node53592;
	wire [4-1:0] node53593;
	wire [4-1:0] node53594;
	wire [4-1:0] node53597;
	wire [4-1:0] node53600;
	wire [4-1:0] node53602;
	wire [4-1:0] node53605;
	wire [4-1:0] node53606;
	wire [4-1:0] node53607;
	wire [4-1:0] node53608;
	wire [4-1:0] node53611;
	wire [4-1:0] node53614;
	wire [4-1:0] node53615;
	wire [4-1:0] node53618;
	wire [4-1:0] node53621;
	wire [4-1:0] node53622;
	wire [4-1:0] node53623;
	wire [4-1:0] node53626;
	wire [4-1:0] node53629;
	wire [4-1:0] node53630;
	wire [4-1:0] node53633;
	wire [4-1:0] node53636;
	wire [4-1:0] node53637;
	wire [4-1:0] node53638;
	wire [4-1:0] node53639;
	wire [4-1:0] node53640;
	wire [4-1:0] node53644;
	wire [4-1:0] node53645;
	wire [4-1:0] node53648;
	wire [4-1:0] node53651;
	wire [4-1:0] node53652;
	wire [4-1:0] node53653;
	wire [4-1:0] node53656;
	wire [4-1:0] node53659;
	wire [4-1:0] node53660;
	wire [4-1:0] node53664;
	wire [4-1:0] node53665;
	wire [4-1:0] node53666;
	wire [4-1:0] node53667;
	wire [4-1:0] node53670;
	wire [4-1:0] node53673;
	wire [4-1:0] node53675;
	wire [4-1:0] node53678;
	wire [4-1:0] node53679;
	wire [4-1:0] node53680;
	wire [4-1:0] node53683;
	wire [4-1:0] node53686;
	wire [4-1:0] node53687;
	wire [4-1:0] node53690;
	wire [4-1:0] node53693;
	wire [4-1:0] node53694;
	wire [4-1:0] node53695;
	wire [4-1:0] node53696;
	wire [4-1:0] node53697;
	wire [4-1:0] node53698;
	wire [4-1:0] node53700;
	wire [4-1:0] node53703;
	wire [4-1:0] node53706;
	wire [4-1:0] node53707;
	wire [4-1:0] node53708;
	wire [4-1:0] node53711;
	wire [4-1:0] node53714;
	wire [4-1:0] node53715;
	wire [4-1:0] node53719;
	wire [4-1:0] node53720;
	wire [4-1:0] node53721;
	wire [4-1:0] node53722;
	wire [4-1:0] node53725;
	wire [4-1:0] node53728;
	wire [4-1:0] node53729;
	wire [4-1:0] node53732;
	wire [4-1:0] node53735;
	wire [4-1:0] node53736;
	wire [4-1:0] node53737;
	wire [4-1:0] node53740;
	wire [4-1:0] node53743;
	wire [4-1:0] node53744;
	wire [4-1:0] node53747;
	wire [4-1:0] node53750;
	wire [4-1:0] node53751;
	wire [4-1:0] node53752;
	wire [4-1:0] node53753;
	wire [4-1:0] node53754;
	wire [4-1:0] node53757;
	wire [4-1:0] node53760;
	wire [4-1:0] node53761;
	wire [4-1:0] node53764;
	wire [4-1:0] node53767;
	wire [4-1:0] node53768;
	wire [4-1:0] node53769;
	wire [4-1:0] node53772;
	wire [4-1:0] node53775;
	wire [4-1:0] node53776;
	wire [4-1:0] node53779;
	wire [4-1:0] node53782;
	wire [4-1:0] node53783;
	wire [4-1:0] node53784;
	wire [4-1:0] node53785;
	wire [4-1:0] node53788;
	wire [4-1:0] node53791;
	wire [4-1:0] node53792;
	wire [4-1:0] node53795;
	wire [4-1:0] node53798;
	wire [4-1:0] node53799;
	wire [4-1:0] node53800;
	wire [4-1:0] node53803;
	wire [4-1:0] node53806;
	wire [4-1:0] node53807;
	wire [4-1:0] node53810;
	wire [4-1:0] node53813;
	wire [4-1:0] node53814;
	wire [4-1:0] node53815;
	wire [4-1:0] node53816;
	wire [4-1:0] node53817;
	wire [4-1:0] node53818;
	wire [4-1:0] node53821;
	wire [4-1:0] node53824;
	wire [4-1:0] node53825;
	wire [4-1:0] node53828;
	wire [4-1:0] node53831;
	wire [4-1:0] node53832;
	wire [4-1:0] node53834;
	wire [4-1:0] node53837;
	wire [4-1:0] node53838;
	wire [4-1:0] node53841;
	wire [4-1:0] node53844;
	wire [4-1:0] node53845;
	wire [4-1:0] node53846;
	wire [4-1:0] node53847;
	wire [4-1:0] node53850;
	wire [4-1:0] node53853;
	wire [4-1:0] node53854;
	wire [4-1:0] node53857;
	wire [4-1:0] node53860;
	wire [4-1:0] node53861;
	wire [4-1:0] node53862;
	wire [4-1:0] node53865;
	wire [4-1:0] node53868;
	wire [4-1:0] node53869;
	wire [4-1:0] node53872;
	wire [4-1:0] node53875;
	wire [4-1:0] node53876;
	wire [4-1:0] node53877;
	wire [4-1:0] node53878;
	wire [4-1:0] node53879;
	wire [4-1:0] node53882;
	wire [4-1:0] node53885;
	wire [4-1:0] node53886;
	wire [4-1:0] node53889;
	wire [4-1:0] node53892;
	wire [4-1:0] node53893;
	wire [4-1:0] node53894;
	wire [4-1:0] node53897;
	wire [4-1:0] node53900;
	wire [4-1:0] node53901;
	wire [4-1:0] node53904;
	wire [4-1:0] node53907;
	wire [4-1:0] node53908;
	wire [4-1:0] node53909;
	wire [4-1:0] node53911;
	wire [4-1:0] node53914;
	wire [4-1:0] node53915;
	wire [4-1:0] node53918;
	wire [4-1:0] node53921;
	wire [4-1:0] node53922;
	wire [4-1:0] node53924;
	wire [4-1:0] node53927;
	wire [4-1:0] node53928;
	wire [4-1:0] node53931;
	wire [4-1:0] node53934;
	wire [4-1:0] node53935;
	wire [4-1:0] node53936;
	wire [4-1:0] node53937;
	wire [4-1:0] node53938;
	wire [4-1:0] node53939;
	wire [4-1:0] node53940;
	wire [4-1:0] node53941;
	wire [4-1:0] node53942;
	wire [4-1:0] node53943;
	wire [4-1:0] node53944;
	wire [4-1:0] node53947;
	wire [4-1:0] node53950;
	wire [4-1:0] node53951;
	wire [4-1:0] node53954;
	wire [4-1:0] node53957;
	wire [4-1:0] node53958;
	wire [4-1:0] node53959;
	wire [4-1:0] node53962;
	wire [4-1:0] node53965;
	wire [4-1:0] node53966;
	wire [4-1:0] node53969;
	wire [4-1:0] node53972;
	wire [4-1:0] node53973;
	wire [4-1:0] node53974;
	wire [4-1:0] node53975;
	wire [4-1:0] node53978;
	wire [4-1:0] node53981;
	wire [4-1:0] node53982;
	wire [4-1:0] node53985;
	wire [4-1:0] node53988;
	wire [4-1:0] node53989;
	wire [4-1:0] node53990;
	wire [4-1:0] node53993;
	wire [4-1:0] node53996;
	wire [4-1:0] node53997;
	wire [4-1:0] node54000;
	wire [4-1:0] node54003;
	wire [4-1:0] node54004;
	wire [4-1:0] node54005;
	wire [4-1:0] node54006;
	wire [4-1:0] node54007;
	wire [4-1:0] node54011;
	wire [4-1:0] node54012;
	wire [4-1:0] node54015;
	wire [4-1:0] node54018;
	wire [4-1:0] node54019;
	wire [4-1:0] node54021;
	wire [4-1:0] node54024;
	wire [4-1:0] node54025;
	wire [4-1:0] node54028;
	wire [4-1:0] node54031;
	wire [4-1:0] node54032;
	wire [4-1:0] node54033;
	wire [4-1:0] node54034;
	wire [4-1:0] node54037;
	wire [4-1:0] node54040;
	wire [4-1:0] node54042;
	wire [4-1:0] node54045;
	wire [4-1:0] node54046;
	wire [4-1:0] node54047;
	wire [4-1:0] node54050;
	wire [4-1:0] node54053;
	wire [4-1:0] node54054;
	wire [4-1:0] node54057;
	wire [4-1:0] node54060;
	wire [4-1:0] node54061;
	wire [4-1:0] node54062;
	wire [4-1:0] node54063;
	wire [4-1:0] node54064;
	wire [4-1:0] node54065;
	wire [4-1:0] node54068;
	wire [4-1:0] node54072;
	wire [4-1:0] node54073;
	wire [4-1:0] node54074;
	wire [4-1:0] node54077;
	wire [4-1:0] node54080;
	wire [4-1:0] node54082;
	wire [4-1:0] node54085;
	wire [4-1:0] node54086;
	wire [4-1:0] node54087;
	wire [4-1:0] node54088;
	wire [4-1:0] node54091;
	wire [4-1:0] node54094;
	wire [4-1:0] node54095;
	wire [4-1:0] node54098;
	wire [4-1:0] node54101;
	wire [4-1:0] node54102;
	wire [4-1:0] node54105;
	wire [4-1:0] node54108;
	wire [4-1:0] node54109;
	wire [4-1:0] node54110;
	wire [4-1:0] node54111;
	wire [4-1:0] node54112;
	wire [4-1:0] node54115;
	wire [4-1:0] node54118;
	wire [4-1:0] node54119;
	wire [4-1:0] node54122;
	wire [4-1:0] node54125;
	wire [4-1:0] node54126;
	wire [4-1:0] node54128;
	wire [4-1:0] node54131;
	wire [4-1:0] node54132;
	wire [4-1:0] node54136;
	wire [4-1:0] node54137;
	wire [4-1:0] node54138;
	wire [4-1:0] node54139;
	wire [4-1:0] node54142;
	wire [4-1:0] node54145;
	wire [4-1:0] node54146;
	wire [4-1:0] node54149;
	wire [4-1:0] node54152;
	wire [4-1:0] node54153;
	wire [4-1:0] node54156;
	wire [4-1:0] node54159;
	wire [4-1:0] node54160;
	wire [4-1:0] node54161;
	wire [4-1:0] node54162;
	wire [4-1:0] node54163;
	wire [4-1:0] node54164;
	wire [4-1:0] node54166;
	wire [4-1:0] node54169;
	wire [4-1:0] node54170;
	wire [4-1:0] node54173;
	wire [4-1:0] node54176;
	wire [4-1:0] node54177;
	wire [4-1:0] node54178;
	wire [4-1:0] node54181;
	wire [4-1:0] node54184;
	wire [4-1:0] node54186;
	wire [4-1:0] node54189;
	wire [4-1:0] node54190;
	wire [4-1:0] node54191;
	wire [4-1:0] node54192;
	wire [4-1:0] node54196;
	wire [4-1:0] node54197;
	wire [4-1:0] node54200;
	wire [4-1:0] node54203;
	wire [4-1:0] node54204;
	wire [4-1:0] node54207;
	wire [4-1:0] node54210;
	wire [4-1:0] node54211;
	wire [4-1:0] node54212;
	wire [4-1:0] node54213;
	wire [4-1:0] node54214;
	wire [4-1:0] node54217;
	wire [4-1:0] node54220;
	wire [4-1:0] node54221;
	wire [4-1:0] node54224;
	wire [4-1:0] node54227;
	wire [4-1:0] node54228;
	wire [4-1:0] node54229;
	wire [4-1:0] node54232;
	wire [4-1:0] node54235;
	wire [4-1:0] node54236;
	wire [4-1:0] node54239;
	wire [4-1:0] node54242;
	wire [4-1:0] node54243;
	wire [4-1:0] node54244;
	wire [4-1:0] node54245;
	wire [4-1:0] node54249;
	wire [4-1:0] node54250;
	wire [4-1:0] node54254;
	wire [4-1:0] node54255;
	wire [4-1:0] node54256;
	wire [4-1:0] node54260;
	wire [4-1:0] node54261;
	wire [4-1:0] node54265;
	wire [4-1:0] node54266;
	wire [4-1:0] node54267;
	wire [4-1:0] node54268;
	wire [4-1:0] node54269;
	wire [4-1:0] node54270;
	wire [4-1:0] node54273;
	wire [4-1:0] node54276;
	wire [4-1:0] node54277;
	wire [4-1:0] node54280;
	wire [4-1:0] node54283;
	wire [4-1:0] node54284;
	wire [4-1:0] node54286;
	wire [4-1:0] node54289;
	wire [4-1:0] node54290;
	wire [4-1:0] node54293;
	wire [4-1:0] node54296;
	wire [4-1:0] node54297;
	wire [4-1:0] node54298;
	wire [4-1:0] node54299;
	wire [4-1:0] node54302;
	wire [4-1:0] node54305;
	wire [4-1:0] node54306;
	wire [4-1:0] node54309;
	wire [4-1:0] node54312;
	wire [4-1:0] node54313;
	wire [4-1:0] node54314;
	wire [4-1:0] node54317;
	wire [4-1:0] node54320;
	wire [4-1:0] node54321;
	wire [4-1:0] node54324;
	wire [4-1:0] node54327;
	wire [4-1:0] node54328;
	wire [4-1:0] node54329;
	wire [4-1:0] node54330;
	wire [4-1:0] node54331;
	wire [4-1:0] node54334;
	wire [4-1:0] node54337;
	wire [4-1:0] node54338;
	wire [4-1:0] node54341;
	wire [4-1:0] node54344;
	wire [4-1:0] node54345;
	wire [4-1:0] node54346;
	wire [4-1:0] node54350;
	wire [4-1:0] node54352;
	wire [4-1:0] node54355;
	wire [4-1:0] node54356;
	wire [4-1:0] node54357;
	wire [4-1:0] node54358;
	wire [4-1:0] node54361;
	wire [4-1:0] node54364;
	wire [4-1:0] node54365;
	wire [4-1:0] node54368;
	wire [4-1:0] node54371;
	wire [4-1:0] node54372;
	wire [4-1:0] node54373;
	wire [4-1:0] node54376;
	wire [4-1:0] node54379;
	wire [4-1:0] node54380;
	wire [4-1:0] node54383;
	wire [4-1:0] node54386;
	wire [4-1:0] node54387;
	wire [4-1:0] node54388;
	wire [4-1:0] node54389;
	wire [4-1:0] node54390;
	wire [4-1:0] node54391;
	wire [4-1:0] node54392;
	wire [4-1:0] node54393;
	wire [4-1:0] node54396;
	wire [4-1:0] node54399;
	wire [4-1:0] node54400;
	wire [4-1:0] node54403;
	wire [4-1:0] node54406;
	wire [4-1:0] node54407;
	wire [4-1:0] node54408;
	wire [4-1:0] node54411;
	wire [4-1:0] node54414;
	wire [4-1:0] node54415;
	wire [4-1:0] node54418;
	wire [4-1:0] node54421;
	wire [4-1:0] node54422;
	wire [4-1:0] node54423;
	wire [4-1:0] node54424;
	wire [4-1:0] node54427;
	wire [4-1:0] node54430;
	wire [4-1:0] node54431;
	wire [4-1:0] node54434;
	wire [4-1:0] node54437;
	wire [4-1:0] node54438;
	wire [4-1:0] node54439;
	wire [4-1:0] node54442;
	wire [4-1:0] node54445;
	wire [4-1:0] node54446;
	wire [4-1:0] node54449;
	wire [4-1:0] node54452;
	wire [4-1:0] node54453;
	wire [4-1:0] node54454;
	wire [4-1:0] node54455;
	wire [4-1:0] node54456;
	wire [4-1:0] node54459;
	wire [4-1:0] node54462;
	wire [4-1:0] node54463;
	wire [4-1:0] node54466;
	wire [4-1:0] node54469;
	wire [4-1:0] node54470;
	wire [4-1:0] node54471;
	wire [4-1:0] node54474;
	wire [4-1:0] node54477;
	wire [4-1:0] node54480;
	wire [4-1:0] node54481;
	wire [4-1:0] node54482;
	wire [4-1:0] node54483;
	wire [4-1:0] node54486;
	wire [4-1:0] node54489;
	wire [4-1:0] node54490;
	wire [4-1:0] node54493;
	wire [4-1:0] node54496;
	wire [4-1:0] node54497;
	wire [4-1:0] node54498;
	wire [4-1:0] node54501;
	wire [4-1:0] node54504;
	wire [4-1:0] node54505;
	wire [4-1:0] node54508;
	wire [4-1:0] node54511;
	wire [4-1:0] node54512;
	wire [4-1:0] node54513;
	wire [4-1:0] node54514;
	wire [4-1:0] node54515;
	wire [4-1:0] node54516;
	wire [4-1:0] node54519;
	wire [4-1:0] node54522;
	wire [4-1:0] node54523;
	wire [4-1:0] node54526;
	wire [4-1:0] node54529;
	wire [4-1:0] node54530;
	wire [4-1:0] node54531;
	wire [4-1:0] node54534;
	wire [4-1:0] node54537;
	wire [4-1:0] node54538;
	wire [4-1:0] node54541;
	wire [4-1:0] node54544;
	wire [4-1:0] node54545;
	wire [4-1:0] node54546;
	wire [4-1:0] node54547;
	wire [4-1:0] node54550;
	wire [4-1:0] node54553;
	wire [4-1:0] node54554;
	wire [4-1:0] node54557;
	wire [4-1:0] node54560;
	wire [4-1:0] node54561;
	wire [4-1:0] node54564;
	wire [4-1:0] node54567;
	wire [4-1:0] node54568;
	wire [4-1:0] node54569;
	wire [4-1:0] node54570;
	wire [4-1:0] node54571;
	wire [4-1:0] node54575;
	wire [4-1:0] node54576;
	wire [4-1:0] node54579;
	wire [4-1:0] node54582;
	wire [4-1:0] node54583;
	wire [4-1:0] node54585;
	wire [4-1:0] node54588;
	wire [4-1:0] node54589;
	wire [4-1:0] node54592;
	wire [4-1:0] node54595;
	wire [4-1:0] node54596;
	wire [4-1:0] node54597;
	wire [4-1:0] node54598;
	wire [4-1:0] node54601;
	wire [4-1:0] node54604;
	wire [4-1:0] node54605;
	wire [4-1:0] node54608;
	wire [4-1:0] node54611;
	wire [4-1:0] node54612;
	wire [4-1:0] node54614;
	wire [4-1:0] node54617;
	wire [4-1:0] node54618;
	wire [4-1:0] node54621;
	wire [4-1:0] node54624;
	wire [4-1:0] node54625;
	wire [4-1:0] node54626;
	wire [4-1:0] node54627;
	wire [4-1:0] node54628;
	wire [4-1:0] node54629;
	wire [4-1:0] node54630;
	wire [4-1:0] node54634;
	wire [4-1:0] node54635;
	wire [4-1:0] node54638;
	wire [4-1:0] node54641;
	wire [4-1:0] node54642;
	wire [4-1:0] node54644;
	wire [4-1:0] node54647;
	wire [4-1:0] node54649;
	wire [4-1:0] node54652;
	wire [4-1:0] node54653;
	wire [4-1:0] node54654;
	wire [4-1:0] node54655;
	wire [4-1:0] node54660;
	wire [4-1:0] node54661;
	wire [4-1:0] node54662;
	wire [4-1:0] node54666;
	wire [4-1:0] node54667;
	wire [4-1:0] node54671;
	wire [4-1:0] node54672;
	wire [4-1:0] node54673;
	wire [4-1:0] node54674;
	wire [4-1:0] node54675;
	wire [4-1:0] node54679;
	wire [4-1:0] node54680;
	wire [4-1:0] node54684;
	wire [4-1:0] node54685;
	wire [4-1:0] node54686;
	wire [4-1:0] node54690;
	wire [4-1:0] node54691;
	wire [4-1:0] node54695;
	wire [4-1:0] node54696;
	wire [4-1:0] node54697;
	wire [4-1:0] node54698;
	wire [4-1:0] node54702;
	wire [4-1:0] node54703;
	wire [4-1:0] node54707;
	wire [4-1:0] node54708;
	wire [4-1:0] node54709;
	wire [4-1:0] node54713;
	wire [4-1:0] node54714;
	wire [4-1:0] node54718;
	wire [4-1:0] node54719;
	wire [4-1:0] node54720;
	wire [4-1:0] node54721;
	wire [4-1:0] node54722;
	wire [4-1:0] node54723;
	wire [4-1:0] node54726;
	wire [4-1:0] node54729;
	wire [4-1:0] node54730;
	wire [4-1:0] node54734;
	wire [4-1:0] node54735;
	wire [4-1:0] node54737;
	wire [4-1:0] node54740;
	wire [4-1:0] node54741;
	wire [4-1:0] node54744;
	wire [4-1:0] node54747;
	wire [4-1:0] node54748;
	wire [4-1:0] node54749;
	wire [4-1:0] node54750;
	wire [4-1:0] node54754;
	wire [4-1:0] node54755;
	wire [4-1:0] node54759;
	wire [4-1:0] node54760;
	wire [4-1:0] node54761;
	wire [4-1:0] node54765;
	wire [4-1:0] node54766;
	wire [4-1:0] node54770;
	wire [4-1:0] node54771;
	wire [4-1:0] node54772;
	wire [4-1:0] node54773;
	wire [4-1:0] node54774;
	wire [4-1:0] node54777;
	wire [4-1:0] node54780;
	wire [4-1:0] node54781;
	wire [4-1:0] node54784;
	wire [4-1:0] node54787;
	wire [4-1:0] node54788;
	wire [4-1:0] node54789;
	wire [4-1:0] node54792;
	wire [4-1:0] node54795;
	wire [4-1:0] node54797;
	wire [4-1:0] node54800;
	wire [4-1:0] node54801;
	wire [4-1:0] node54802;
	wire [4-1:0] node54803;
	wire [4-1:0] node54806;
	wire [4-1:0] node54809;
	wire [4-1:0] node54810;
	wire [4-1:0] node54813;
	wire [4-1:0] node54816;
	wire [4-1:0] node54817;
	wire [4-1:0] node54818;
	wire [4-1:0] node54821;
	wire [4-1:0] node54824;
	wire [4-1:0] node54825;
	wire [4-1:0] node54829;
	wire [4-1:0] node54830;
	wire [4-1:0] node54831;
	wire [4-1:0] node54832;
	wire [4-1:0] node54833;
	wire [4-1:0] node54834;
	wire [4-1:0] node54835;
	wire [4-1:0] node54836;
	wire [4-1:0] node54837;
	wire [4-1:0] node54840;
	wire [4-1:0] node54843;
	wire [4-1:0] node54844;
	wire [4-1:0] node54847;
	wire [4-1:0] node54850;
	wire [4-1:0] node54851;
	wire [4-1:0] node54852;
	wire [4-1:0] node54855;
	wire [4-1:0] node54858;
	wire [4-1:0] node54859;
	wire [4-1:0] node54862;
	wire [4-1:0] node54865;
	wire [4-1:0] node54866;
	wire [4-1:0] node54867;
	wire [4-1:0] node54868;
	wire [4-1:0] node54871;
	wire [4-1:0] node54874;
	wire [4-1:0] node54875;
	wire [4-1:0] node54878;
	wire [4-1:0] node54881;
	wire [4-1:0] node54882;
	wire [4-1:0] node54883;
	wire [4-1:0] node54886;
	wire [4-1:0] node54889;
	wire [4-1:0] node54890;
	wire [4-1:0] node54893;
	wire [4-1:0] node54896;
	wire [4-1:0] node54897;
	wire [4-1:0] node54898;
	wire [4-1:0] node54899;
	wire [4-1:0] node54900;
	wire [4-1:0] node54903;
	wire [4-1:0] node54906;
	wire [4-1:0] node54908;
	wire [4-1:0] node54911;
	wire [4-1:0] node54912;
	wire [4-1:0] node54913;
	wire [4-1:0] node54916;
	wire [4-1:0] node54919;
	wire [4-1:0] node54921;
	wire [4-1:0] node54924;
	wire [4-1:0] node54925;
	wire [4-1:0] node54926;
	wire [4-1:0] node54927;
	wire [4-1:0] node54930;
	wire [4-1:0] node54933;
	wire [4-1:0] node54934;
	wire [4-1:0] node54937;
	wire [4-1:0] node54940;
	wire [4-1:0] node54941;
	wire [4-1:0] node54942;
	wire [4-1:0] node54945;
	wire [4-1:0] node54948;
	wire [4-1:0] node54950;
	wire [4-1:0] node54953;
	wire [4-1:0] node54954;
	wire [4-1:0] node54955;
	wire [4-1:0] node54956;
	wire [4-1:0] node54957;
	wire [4-1:0] node54958;
	wire [4-1:0] node54962;
	wire [4-1:0] node54963;
	wire [4-1:0] node54967;
	wire [4-1:0] node54968;
	wire [4-1:0] node54969;
	wire [4-1:0] node54973;
	wire [4-1:0] node54974;
	wire [4-1:0] node54978;
	wire [4-1:0] node54979;
	wire [4-1:0] node54980;
	wire [4-1:0] node54981;
	wire [4-1:0] node54985;
	wire [4-1:0] node54986;
	wire [4-1:0] node54990;
	wire [4-1:0] node54991;
	wire [4-1:0] node54992;
	wire [4-1:0] node54996;
	wire [4-1:0] node54997;
	wire [4-1:0] node55001;
	wire [4-1:0] node55002;
	wire [4-1:0] node55003;
	wire [4-1:0] node55004;
	wire [4-1:0] node55005;
	wire [4-1:0] node55009;
	wire [4-1:0] node55010;
	wire [4-1:0] node55014;
	wire [4-1:0] node55015;
	wire [4-1:0] node55016;
	wire [4-1:0] node55020;
	wire [4-1:0] node55021;
	wire [4-1:0] node55025;
	wire [4-1:0] node55026;
	wire [4-1:0] node55027;
	wire [4-1:0] node55028;
	wire [4-1:0] node55032;
	wire [4-1:0] node55033;
	wire [4-1:0] node55037;
	wire [4-1:0] node55038;
	wire [4-1:0] node55039;
	wire [4-1:0] node55043;
	wire [4-1:0] node55044;
	wire [4-1:0] node55048;
	wire [4-1:0] node55049;
	wire [4-1:0] node55050;
	wire [4-1:0] node55051;
	wire [4-1:0] node55052;
	wire [4-1:0] node55053;
	wire [4-1:0] node55054;
	wire [4-1:0] node55057;
	wire [4-1:0] node55060;
	wire [4-1:0] node55061;
	wire [4-1:0] node55064;
	wire [4-1:0] node55067;
	wire [4-1:0] node55068;
	wire [4-1:0] node55069;
	wire [4-1:0] node55072;
	wire [4-1:0] node55075;
	wire [4-1:0] node55076;
	wire [4-1:0] node55079;
	wire [4-1:0] node55082;
	wire [4-1:0] node55083;
	wire [4-1:0] node55084;
	wire [4-1:0] node55085;
	wire [4-1:0] node55088;
	wire [4-1:0] node55091;
	wire [4-1:0] node55092;
	wire [4-1:0] node55095;
	wire [4-1:0] node55098;
	wire [4-1:0] node55099;
	wire [4-1:0] node55100;
	wire [4-1:0] node55103;
	wire [4-1:0] node55106;
	wire [4-1:0] node55107;
	wire [4-1:0] node55110;
	wire [4-1:0] node55113;
	wire [4-1:0] node55114;
	wire [4-1:0] node55115;
	wire [4-1:0] node55116;
	wire [4-1:0] node55117;
	wire [4-1:0] node55120;
	wire [4-1:0] node55123;
	wire [4-1:0] node55125;
	wire [4-1:0] node55128;
	wire [4-1:0] node55129;
	wire [4-1:0] node55131;
	wire [4-1:0] node55134;
	wire [4-1:0] node55135;
	wire [4-1:0] node55138;
	wire [4-1:0] node55141;
	wire [4-1:0] node55142;
	wire [4-1:0] node55143;
	wire [4-1:0] node55144;
	wire [4-1:0] node55148;
	wire [4-1:0] node55150;
	wire [4-1:0] node55153;
	wire [4-1:0] node55154;
	wire [4-1:0] node55155;
	wire [4-1:0] node55159;
	wire [4-1:0] node55161;
	wire [4-1:0] node55164;
	wire [4-1:0] node55165;
	wire [4-1:0] node55166;
	wire [4-1:0] node55167;
	wire [4-1:0] node55168;
	wire [4-1:0] node55170;
	wire [4-1:0] node55173;
	wire [4-1:0] node55174;
	wire [4-1:0] node55177;
	wire [4-1:0] node55180;
	wire [4-1:0] node55181;
	wire [4-1:0] node55184;
	wire [4-1:0] node55187;
	wire [4-1:0] node55188;
	wire [4-1:0] node55189;
	wire [4-1:0] node55190;
	wire [4-1:0] node55193;
	wire [4-1:0] node55196;
	wire [4-1:0] node55197;
	wire [4-1:0] node55200;
	wire [4-1:0] node55203;
	wire [4-1:0] node55204;
	wire [4-1:0] node55207;
	wire [4-1:0] node55210;
	wire [4-1:0] node55211;
	wire [4-1:0] node55212;
	wire [4-1:0] node55213;
	wire [4-1:0] node55214;
	wire [4-1:0] node55217;
	wire [4-1:0] node55220;
	wire [4-1:0] node55221;
	wire [4-1:0] node55224;
	wire [4-1:0] node55227;
	wire [4-1:0] node55228;
	wire [4-1:0] node55229;
	wire [4-1:0] node55232;
	wire [4-1:0] node55235;
	wire [4-1:0] node55236;
	wire [4-1:0] node55239;
	wire [4-1:0] node55242;
	wire [4-1:0] node55243;
	wire [4-1:0] node55244;
	wire [4-1:0] node55245;
	wire [4-1:0] node55248;
	wire [4-1:0] node55251;
	wire [4-1:0] node55252;
	wire [4-1:0] node55255;
	wire [4-1:0] node55258;
	wire [4-1:0] node55259;
	wire [4-1:0] node55260;
	wire [4-1:0] node55263;
	wire [4-1:0] node55266;
	wire [4-1:0] node55267;
	wire [4-1:0] node55270;
	wire [4-1:0] node55273;
	wire [4-1:0] node55274;
	wire [4-1:0] node55275;
	wire [4-1:0] node55276;
	wire [4-1:0] node55277;
	wire [4-1:0] node55278;
	wire [4-1:0] node55279;
	wire [4-1:0] node55280;
	wire [4-1:0] node55283;
	wire [4-1:0] node55286;
	wire [4-1:0] node55287;
	wire [4-1:0] node55290;
	wire [4-1:0] node55293;
	wire [4-1:0] node55294;
	wire [4-1:0] node55295;
	wire [4-1:0] node55298;
	wire [4-1:0] node55301;
	wire [4-1:0] node55302;
	wire [4-1:0] node55305;
	wire [4-1:0] node55308;
	wire [4-1:0] node55309;
	wire [4-1:0] node55310;
	wire [4-1:0] node55312;
	wire [4-1:0] node55315;
	wire [4-1:0] node55316;
	wire [4-1:0] node55319;
	wire [4-1:0] node55322;
	wire [4-1:0] node55323;
	wire [4-1:0] node55324;
	wire [4-1:0] node55327;
	wire [4-1:0] node55330;
	wire [4-1:0] node55331;
	wire [4-1:0] node55334;
	wire [4-1:0] node55337;
	wire [4-1:0] node55338;
	wire [4-1:0] node55339;
	wire [4-1:0] node55340;
	wire [4-1:0] node55341;
	wire [4-1:0] node55344;
	wire [4-1:0] node55347;
	wire [4-1:0] node55348;
	wire [4-1:0] node55351;
	wire [4-1:0] node55354;
	wire [4-1:0] node55355;
	wire [4-1:0] node55356;
	wire [4-1:0] node55359;
	wire [4-1:0] node55362;
	wire [4-1:0] node55363;
	wire [4-1:0] node55367;
	wire [4-1:0] node55368;
	wire [4-1:0] node55369;
	wire [4-1:0] node55370;
	wire [4-1:0] node55373;
	wire [4-1:0] node55376;
	wire [4-1:0] node55377;
	wire [4-1:0] node55380;
	wire [4-1:0] node55383;
	wire [4-1:0] node55384;
	wire [4-1:0] node55385;
	wire [4-1:0] node55388;
	wire [4-1:0] node55391;
	wire [4-1:0] node55392;
	wire [4-1:0] node55395;
	wire [4-1:0] node55398;
	wire [4-1:0] node55399;
	wire [4-1:0] node55400;
	wire [4-1:0] node55401;
	wire [4-1:0] node55402;
	wire [4-1:0] node55403;
	wire [4-1:0] node55406;
	wire [4-1:0] node55409;
	wire [4-1:0] node55410;
	wire [4-1:0] node55413;
	wire [4-1:0] node55416;
	wire [4-1:0] node55417;
	wire [4-1:0] node55418;
	wire [4-1:0] node55421;
	wire [4-1:0] node55424;
	wire [4-1:0] node55425;
	wire [4-1:0] node55429;
	wire [4-1:0] node55430;
	wire [4-1:0] node55431;
	wire [4-1:0] node55432;
	wire [4-1:0] node55435;
	wire [4-1:0] node55438;
	wire [4-1:0] node55439;
	wire [4-1:0] node55442;
	wire [4-1:0] node55445;
	wire [4-1:0] node55446;
	wire [4-1:0] node55447;
	wire [4-1:0] node55450;
	wire [4-1:0] node55453;
	wire [4-1:0] node55454;
	wire [4-1:0] node55457;
	wire [4-1:0] node55460;
	wire [4-1:0] node55461;
	wire [4-1:0] node55462;
	wire [4-1:0] node55463;
	wire [4-1:0] node55464;
	wire [4-1:0] node55467;
	wire [4-1:0] node55470;
	wire [4-1:0] node55471;
	wire [4-1:0] node55474;
	wire [4-1:0] node55477;
	wire [4-1:0] node55478;
	wire [4-1:0] node55479;
	wire [4-1:0] node55482;
	wire [4-1:0] node55485;
	wire [4-1:0] node55486;
	wire [4-1:0] node55489;
	wire [4-1:0] node55492;
	wire [4-1:0] node55493;
	wire [4-1:0] node55494;
	wire [4-1:0] node55495;
	wire [4-1:0] node55498;
	wire [4-1:0] node55501;
	wire [4-1:0] node55502;
	wire [4-1:0] node55505;
	wire [4-1:0] node55508;
	wire [4-1:0] node55509;
	wire [4-1:0] node55510;
	wire [4-1:0] node55513;
	wire [4-1:0] node55516;
	wire [4-1:0] node55517;
	wire [4-1:0] node55520;
	wire [4-1:0] node55523;
	wire [4-1:0] node55524;
	wire [4-1:0] node55525;
	wire [4-1:0] node55526;
	wire [4-1:0] node55527;
	wire [4-1:0] node55528;
	wire [4-1:0] node55529;
	wire [4-1:0] node55532;
	wire [4-1:0] node55535;
	wire [4-1:0] node55536;
	wire [4-1:0] node55539;
	wire [4-1:0] node55542;
	wire [4-1:0] node55543;
	wire [4-1:0] node55544;
	wire [4-1:0] node55547;
	wire [4-1:0] node55550;
	wire [4-1:0] node55551;
	wire [4-1:0] node55554;
	wire [4-1:0] node55557;
	wire [4-1:0] node55558;
	wire [4-1:0] node55559;
	wire [4-1:0] node55560;
	wire [4-1:0] node55563;
	wire [4-1:0] node55566;
	wire [4-1:0] node55567;
	wire [4-1:0] node55570;
	wire [4-1:0] node55573;
	wire [4-1:0] node55574;
	wire [4-1:0] node55575;
	wire [4-1:0] node55579;
	wire [4-1:0] node55580;
	wire [4-1:0] node55583;
	wire [4-1:0] node55586;
	wire [4-1:0] node55587;
	wire [4-1:0] node55588;
	wire [4-1:0] node55589;
	wire [4-1:0] node55590;
	wire [4-1:0] node55593;
	wire [4-1:0] node55596;
	wire [4-1:0] node55597;
	wire [4-1:0] node55600;
	wire [4-1:0] node55603;
	wire [4-1:0] node55604;
	wire [4-1:0] node55605;
	wire [4-1:0] node55608;
	wire [4-1:0] node55611;
	wire [4-1:0] node55612;
	wire [4-1:0] node55615;
	wire [4-1:0] node55618;
	wire [4-1:0] node55619;
	wire [4-1:0] node55620;
	wire [4-1:0] node55621;
	wire [4-1:0] node55624;
	wire [4-1:0] node55627;
	wire [4-1:0] node55628;
	wire [4-1:0] node55631;
	wire [4-1:0] node55634;
	wire [4-1:0] node55635;
	wire [4-1:0] node55636;
	wire [4-1:0] node55640;
	wire [4-1:0] node55641;
	wire [4-1:0] node55644;
	wire [4-1:0] node55647;
	wire [4-1:0] node55648;
	wire [4-1:0] node55649;
	wire [4-1:0] node55650;
	wire [4-1:0] node55651;
	wire [4-1:0] node55652;
	wire [4-1:0] node55655;
	wire [4-1:0] node55658;
	wire [4-1:0] node55659;
	wire [4-1:0] node55662;
	wire [4-1:0] node55665;
	wire [4-1:0] node55666;
	wire [4-1:0] node55667;
	wire [4-1:0] node55670;
	wire [4-1:0] node55673;
	wire [4-1:0] node55674;
	wire [4-1:0] node55677;
	wire [4-1:0] node55680;
	wire [4-1:0] node55681;
	wire [4-1:0] node55682;
	wire [4-1:0] node55683;
	wire [4-1:0] node55686;
	wire [4-1:0] node55689;
	wire [4-1:0] node55690;
	wire [4-1:0] node55694;
	wire [4-1:0] node55695;
	wire [4-1:0] node55696;
	wire [4-1:0] node55699;
	wire [4-1:0] node55702;
	wire [4-1:0] node55703;
	wire [4-1:0] node55706;
	wire [4-1:0] node55709;
	wire [4-1:0] node55710;
	wire [4-1:0] node55711;
	wire [4-1:0] node55712;
	wire [4-1:0] node55713;
	wire [4-1:0] node55716;
	wire [4-1:0] node55719;
	wire [4-1:0] node55720;
	wire [4-1:0] node55723;
	wire [4-1:0] node55726;
	wire [4-1:0] node55727;
	wire [4-1:0] node55730;
	wire [4-1:0] node55733;
	wire [4-1:0] node55734;
	wire [4-1:0] node55735;
	wire [4-1:0] node55736;
	wire [4-1:0] node55739;
	wire [4-1:0] node55742;
	wire [4-1:0] node55743;
	wire [4-1:0] node55746;
	wire [4-1:0] node55749;
	wire [4-1:0] node55750;
	wire [4-1:0] node55753;
	wire [4-1:0] node55756;
	wire [4-1:0] node55757;
	wire [4-1:0] node55758;
	wire [4-1:0] node55759;
	wire [4-1:0] node55760;
	wire [4-1:0] node55761;
	wire [4-1:0] node55762;
	wire [4-1:0] node55763;
	wire [4-1:0] node55764;
	wire [4-1:0] node55765;
	wire [4-1:0] node55768;
	wire [4-1:0] node55771;
	wire [4-1:0] node55772;
	wire [4-1:0] node55775;
	wire [4-1:0] node55778;
	wire [4-1:0] node55779;
	wire [4-1:0] node55780;
	wire [4-1:0] node55783;
	wire [4-1:0] node55786;
	wire [4-1:0] node55787;
	wire [4-1:0] node55791;
	wire [4-1:0] node55792;
	wire [4-1:0] node55793;
	wire [4-1:0] node55794;
	wire [4-1:0] node55797;
	wire [4-1:0] node55800;
	wire [4-1:0] node55801;
	wire [4-1:0] node55804;
	wire [4-1:0] node55807;
	wire [4-1:0] node55808;
	wire [4-1:0] node55809;
	wire [4-1:0] node55812;
	wire [4-1:0] node55815;
	wire [4-1:0] node55816;
	wire [4-1:0] node55819;
	wire [4-1:0] node55822;
	wire [4-1:0] node55823;
	wire [4-1:0] node55824;
	wire [4-1:0] node55825;
	wire [4-1:0] node55826;
	wire [4-1:0] node55829;
	wire [4-1:0] node55832;
	wire [4-1:0] node55833;
	wire [4-1:0] node55836;
	wire [4-1:0] node55839;
	wire [4-1:0] node55840;
	wire [4-1:0] node55841;
	wire [4-1:0] node55844;
	wire [4-1:0] node55847;
	wire [4-1:0] node55848;
	wire [4-1:0] node55851;
	wire [4-1:0] node55854;
	wire [4-1:0] node55855;
	wire [4-1:0] node55856;
	wire [4-1:0] node55857;
	wire [4-1:0] node55860;
	wire [4-1:0] node55863;
	wire [4-1:0] node55864;
	wire [4-1:0] node55867;
	wire [4-1:0] node55870;
	wire [4-1:0] node55871;
	wire [4-1:0] node55872;
	wire [4-1:0] node55875;
	wire [4-1:0] node55878;
	wire [4-1:0] node55879;
	wire [4-1:0] node55882;
	wire [4-1:0] node55885;
	wire [4-1:0] node55886;
	wire [4-1:0] node55887;
	wire [4-1:0] node55888;
	wire [4-1:0] node55889;
	wire [4-1:0] node55890;
	wire [4-1:0] node55893;
	wire [4-1:0] node55896;
	wire [4-1:0] node55897;
	wire [4-1:0] node55900;
	wire [4-1:0] node55903;
	wire [4-1:0] node55904;
	wire [4-1:0] node55906;
	wire [4-1:0] node55909;
	wire [4-1:0] node55910;
	wire [4-1:0] node55913;
	wire [4-1:0] node55916;
	wire [4-1:0] node55917;
	wire [4-1:0] node55918;
	wire [4-1:0] node55919;
	wire [4-1:0] node55922;
	wire [4-1:0] node55925;
	wire [4-1:0] node55926;
	wire [4-1:0] node55930;
	wire [4-1:0] node55931;
	wire [4-1:0] node55932;
	wire [4-1:0] node55935;
	wire [4-1:0] node55938;
	wire [4-1:0] node55939;
	wire [4-1:0] node55942;
	wire [4-1:0] node55945;
	wire [4-1:0] node55946;
	wire [4-1:0] node55947;
	wire [4-1:0] node55948;
	wire [4-1:0] node55949;
	wire [4-1:0] node55952;
	wire [4-1:0] node55955;
	wire [4-1:0] node55956;
	wire [4-1:0] node55959;
	wire [4-1:0] node55962;
	wire [4-1:0] node55963;
	wire [4-1:0] node55964;
	wire [4-1:0] node55967;
	wire [4-1:0] node55970;
	wire [4-1:0] node55971;
	wire [4-1:0] node55974;
	wire [4-1:0] node55977;
	wire [4-1:0] node55978;
	wire [4-1:0] node55979;
	wire [4-1:0] node55980;
	wire [4-1:0] node55983;
	wire [4-1:0] node55986;
	wire [4-1:0] node55988;
	wire [4-1:0] node55991;
	wire [4-1:0] node55992;
	wire [4-1:0] node55994;
	wire [4-1:0] node55997;
	wire [4-1:0] node55998;
	wire [4-1:0] node56001;
	wire [4-1:0] node56004;
	wire [4-1:0] node56005;
	wire [4-1:0] node56006;
	wire [4-1:0] node56007;
	wire [4-1:0] node56008;
	wire [4-1:0] node56009;
	wire [4-1:0] node56010;
	wire [4-1:0] node56013;
	wire [4-1:0] node56016;
	wire [4-1:0] node56017;
	wire [4-1:0] node56020;
	wire [4-1:0] node56023;
	wire [4-1:0] node56024;
	wire [4-1:0] node56025;
	wire [4-1:0] node56028;
	wire [4-1:0] node56031;
	wire [4-1:0] node56032;
	wire [4-1:0] node56035;
	wire [4-1:0] node56038;
	wire [4-1:0] node56039;
	wire [4-1:0] node56040;
	wire [4-1:0] node56041;
	wire [4-1:0] node56044;
	wire [4-1:0] node56047;
	wire [4-1:0] node56048;
	wire [4-1:0] node56051;
	wire [4-1:0] node56054;
	wire [4-1:0] node56055;
	wire [4-1:0] node56058;
	wire [4-1:0] node56061;
	wire [4-1:0] node56062;
	wire [4-1:0] node56063;
	wire [4-1:0] node56064;
	wire [4-1:0] node56065;
	wire [4-1:0] node56068;
	wire [4-1:0] node56071;
	wire [4-1:0] node56072;
	wire [4-1:0] node56075;
	wire [4-1:0] node56078;
	wire [4-1:0] node56079;
	wire [4-1:0] node56080;
	wire [4-1:0] node56083;
	wire [4-1:0] node56086;
	wire [4-1:0] node56087;
	wire [4-1:0] node56090;
	wire [4-1:0] node56093;
	wire [4-1:0] node56094;
	wire [4-1:0] node56095;
	wire [4-1:0] node56096;
	wire [4-1:0] node56099;
	wire [4-1:0] node56102;
	wire [4-1:0] node56103;
	wire [4-1:0] node56106;
	wire [4-1:0] node56109;
	wire [4-1:0] node56110;
	wire [4-1:0] node56111;
	wire [4-1:0] node56114;
	wire [4-1:0] node56117;
	wire [4-1:0] node56118;
	wire [4-1:0] node56121;
	wire [4-1:0] node56124;
	wire [4-1:0] node56125;
	wire [4-1:0] node56126;
	wire [4-1:0] node56127;
	wire [4-1:0] node56128;
	wire [4-1:0] node56129;
	wire [4-1:0] node56132;
	wire [4-1:0] node56135;
	wire [4-1:0] node56136;
	wire [4-1:0] node56139;
	wire [4-1:0] node56142;
	wire [4-1:0] node56143;
	wire [4-1:0] node56144;
	wire [4-1:0] node56147;
	wire [4-1:0] node56150;
	wire [4-1:0] node56152;
	wire [4-1:0] node56155;
	wire [4-1:0] node56156;
	wire [4-1:0] node56157;
	wire [4-1:0] node56158;
	wire [4-1:0] node56161;
	wire [4-1:0] node56164;
	wire [4-1:0] node56165;
	wire [4-1:0] node56168;
	wire [4-1:0] node56171;
	wire [4-1:0] node56172;
	wire [4-1:0] node56173;
	wire [4-1:0] node56176;
	wire [4-1:0] node56179;
	wire [4-1:0] node56180;
	wire [4-1:0] node56184;
	wire [4-1:0] node56185;
	wire [4-1:0] node56186;
	wire [4-1:0] node56187;
	wire [4-1:0] node56188;
	wire [4-1:0] node56191;
	wire [4-1:0] node56194;
	wire [4-1:0] node56195;
	wire [4-1:0] node56198;
	wire [4-1:0] node56201;
	wire [4-1:0] node56202;
	wire [4-1:0] node56205;
	wire [4-1:0] node56208;
	wire [4-1:0] node56209;
	wire [4-1:0] node56210;
	wire [4-1:0] node56211;
	wire [4-1:0] node56214;
	wire [4-1:0] node56217;
	wire [4-1:0] node56218;
	wire [4-1:0] node56221;
	wire [4-1:0] node56224;
	wire [4-1:0] node56225;
	wire [4-1:0] node56228;
	wire [4-1:0] node56231;
	wire [4-1:0] node56232;
	wire [4-1:0] node56233;
	wire [4-1:0] node56234;
	wire [4-1:0] node56235;
	wire [4-1:0] node56236;
	wire [4-1:0] node56237;
	wire [4-1:0] node56238;
	wire [4-1:0] node56242;
	wire [4-1:0] node56244;
	wire [4-1:0] node56247;
	wire [4-1:0] node56248;
	wire [4-1:0] node56249;
	wire [4-1:0] node56252;
	wire [4-1:0] node56255;
	wire [4-1:0] node56256;
	wire [4-1:0] node56259;
	wire [4-1:0] node56262;
	wire [4-1:0] node56263;
	wire [4-1:0] node56264;
	wire [4-1:0] node56265;
	wire [4-1:0] node56268;
	wire [4-1:0] node56271;
	wire [4-1:0] node56272;
	wire [4-1:0] node56275;
	wire [4-1:0] node56278;
	wire [4-1:0] node56279;
	wire [4-1:0] node56280;
	wire [4-1:0] node56283;
	wire [4-1:0] node56286;
	wire [4-1:0] node56287;
	wire [4-1:0] node56290;
	wire [4-1:0] node56293;
	wire [4-1:0] node56294;
	wire [4-1:0] node56295;
	wire [4-1:0] node56296;
	wire [4-1:0] node56297;
	wire [4-1:0] node56300;
	wire [4-1:0] node56303;
	wire [4-1:0] node56304;
	wire [4-1:0] node56307;
	wire [4-1:0] node56310;
	wire [4-1:0] node56311;
	wire [4-1:0] node56312;
	wire [4-1:0] node56316;
	wire [4-1:0] node56317;
	wire [4-1:0] node56320;
	wire [4-1:0] node56323;
	wire [4-1:0] node56324;
	wire [4-1:0] node56325;
	wire [4-1:0] node56326;
	wire [4-1:0] node56330;
	wire [4-1:0] node56331;
	wire [4-1:0] node56334;
	wire [4-1:0] node56337;
	wire [4-1:0] node56338;
	wire [4-1:0] node56339;
	wire [4-1:0] node56342;
	wire [4-1:0] node56345;
	wire [4-1:0] node56346;
	wire [4-1:0] node56349;
	wire [4-1:0] node56352;
	wire [4-1:0] node56353;
	wire [4-1:0] node56354;
	wire [4-1:0] node56355;
	wire [4-1:0] node56356;
	wire [4-1:0] node56357;
	wire [4-1:0] node56361;
	wire [4-1:0] node56362;
	wire [4-1:0] node56366;
	wire [4-1:0] node56367;
	wire [4-1:0] node56368;
	wire [4-1:0] node56372;
	wire [4-1:0] node56373;
	wire [4-1:0] node56377;
	wire [4-1:0] node56378;
	wire [4-1:0] node56379;
	wire [4-1:0] node56380;
	wire [4-1:0] node56384;
	wire [4-1:0] node56385;
	wire [4-1:0] node56389;
	wire [4-1:0] node56390;
	wire [4-1:0] node56391;
	wire [4-1:0] node56395;
	wire [4-1:0] node56396;
	wire [4-1:0] node56400;
	wire [4-1:0] node56401;
	wire [4-1:0] node56402;
	wire [4-1:0] node56403;
	wire [4-1:0] node56404;
	wire [4-1:0] node56407;
	wire [4-1:0] node56410;
	wire [4-1:0] node56411;
	wire [4-1:0] node56414;
	wire [4-1:0] node56417;
	wire [4-1:0] node56418;
	wire [4-1:0] node56419;
	wire [4-1:0] node56422;
	wire [4-1:0] node56425;
	wire [4-1:0] node56426;
	wire [4-1:0] node56430;
	wire [4-1:0] node56431;
	wire [4-1:0] node56432;
	wire [4-1:0] node56434;
	wire [4-1:0] node56437;
	wire [4-1:0] node56438;
	wire [4-1:0] node56441;
	wire [4-1:0] node56444;
	wire [4-1:0] node56445;
	wire [4-1:0] node56448;
	wire [4-1:0] node56451;
	wire [4-1:0] node56452;
	wire [4-1:0] node56453;
	wire [4-1:0] node56454;
	wire [4-1:0] node56455;
	wire [4-1:0] node56456;
	wire [4-1:0] node56459;
	wire [4-1:0] node56462;
	wire [4-1:0] node56463;
	wire [4-1:0] node56464;
	wire [4-1:0] node56467;
	wire [4-1:0] node56470;
	wire [4-1:0] node56471;
	wire [4-1:0] node56474;
	wire [4-1:0] node56477;
	wire [4-1:0] node56478;
	wire [4-1:0] node56481;
	wire [4-1:0] node56484;
	wire [4-1:0] node56485;
	wire [4-1:0] node56486;
	wire [4-1:0] node56487;
	wire [4-1:0] node56491;
	wire [4-1:0] node56492;
	wire [4-1:0] node56496;
	wire [4-1:0] node56497;
	wire [4-1:0] node56498;
	wire [4-1:0] node56502;
	wire [4-1:0] node56503;
	wire [4-1:0] node56507;
	wire [4-1:0] node56508;
	wire [4-1:0] node56509;
	wire [4-1:0] node56510;
	wire [4-1:0] node56511;
	wire [4-1:0] node56515;
	wire [4-1:0] node56516;
	wire [4-1:0] node56520;
	wire [4-1:0] node56521;
	wire [4-1:0] node56522;
	wire [4-1:0] node56526;
	wire [4-1:0] node56527;
	wire [4-1:0] node56531;
	wire [4-1:0] node56532;
	wire [4-1:0] node56533;
	wire [4-1:0] node56534;
	wire [4-1:0] node56538;
	wire [4-1:0] node56539;
	wire [4-1:0] node56543;
	wire [4-1:0] node56544;
	wire [4-1:0] node56545;
	wire [4-1:0] node56549;
	wire [4-1:0] node56550;
	wire [4-1:0] node56554;
	wire [4-1:0] node56555;
	wire [4-1:0] node56556;
	wire [4-1:0] node56557;
	wire [4-1:0] node56558;
	wire [4-1:0] node56559;
	wire [4-1:0] node56560;
	wire [4-1:0] node56561;
	wire [4-1:0] node56562;
	wire [4-1:0] node56565;
	wire [4-1:0] node56568;
	wire [4-1:0] node56569;
	wire [4-1:0] node56572;
	wire [4-1:0] node56575;
	wire [4-1:0] node56576;
	wire [4-1:0] node56577;
	wire [4-1:0] node56580;
	wire [4-1:0] node56583;
	wire [4-1:0] node56584;
	wire [4-1:0] node56587;
	wire [4-1:0] node56590;
	wire [4-1:0] node56591;
	wire [4-1:0] node56592;
	wire [4-1:0] node56593;
	wire [4-1:0] node56596;
	wire [4-1:0] node56599;
	wire [4-1:0] node56600;
	wire [4-1:0] node56603;
	wire [4-1:0] node56606;
	wire [4-1:0] node56607;
	wire [4-1:0] node56608;
	wire [4-1:0] node56611;
	wire [4-1:0] node56614;
	wire [4-1:0] node56615;
	wire [4-1:0] node56618;
	wire [4-1:0] node56621;
	wire [4-1:0] node56622;
	wire [4-1:0] node56623;
	wire [4-1:0] node56624;
	wire [4-1:0] node56625;
	wire [4-1:0] node56628;
	wire [4-1:0] node56631;
	wire [4-1:0] node56632;
	wire [4-1:0] node56635;
	wire [4-1:0] node56638;
	wire [4-1:0] node56639;
	wire [4-1:0] node56640;
	wire [4-1:0] node56643;
	wire [4-1:0] node56646;
	wire [4-1:0] node56647;
	wire [4-1:0] node56650;
	wire [4-1:0] node56653;
	wire [4-1:0] node56654;
	wire [4-1:0] node56655;
	wire [4-1:0] node56656;
	wire [4-1:0] node56659;
	wire [4-1:0] node56662;
	wire [4-1:0] node56663;
	wire [4-1:0] node56666;
	wire [4-1:0] node56669;
	wire [4-1:0] node56670;
	wire [4-1:0] node56671;
	wire [4-1:0] node56674;
	wire [4-1:0] node56677;
	wire [4-1:0] node56678;
	wire [4-1:0] node56681;
	wire [4-1:0] node56684;
	wire [4-1:0] node56685;
	wire [4-1:0] node56686;
	wire [4-1:0] node56687;
	wire [4-1:0] node56688;
	wire [4-1:0] node56689;
	wire [4-1:0] node56692;
	wire [4-1:0] node56695;
	wire [4-1:0] node56696;
	wire [4-1:0] node56699;
	wire [4-1:0] node56702;
	wire [4-1:0] node56703;
	wire [4-1:0] node56706;
	wire [4-1:0] node56709;
	wire [4-1:0] node56710;
	wire [4-1:0] node56711;
	wire [4-1:0] node56712;
	wire [4-1:0] node56716;
	wire [4-1:0] node56717;
	wire [4-1:0] node56721;
	wire [4-1:0] node56722;
	wire [4-1:0] node56723;
	wire [4-1:0] node56727;
	wire [4-1:0] node56728;
	wire [4-1:0] node56732;
	wire [4-1:0] node56733;
	wire [4-1:0] node56734;
	wire [4-1:0] node56735;
	wire [4-1:0] node56736;
	wire [4-1:0] node56740;
	wire [4-1:0] node56741;
	wire [4-1:0] node56745;
	wire [4-1:0] node56746;
	wire [4-1:0] node56747;
	wire [4-1:0] node56751;
	wire [4-1:0] node56752;
	wire [4-1:0] node56756;
	wire [4-1:0] node56757;
	wire [4-1:0] node56758;
	wire [4-1:0] node56759;
	wire [4-1:0] node56763;
	wire [4-1:0] node56766;
	wire [4-1:0] node56767;
	wire [4-1:0] node56768;
	wire [4-1:0] node56772;
	wire [4-1:0] node56773;
	wire [4-1:0] node56777;
	wire [4-1:0] node56778;
	wire [4-1:0] node56779;
	wire [4-1:0] node56780;
	wire [4-1:0] node56781;
	wire [4-1:0] node56782;
	wire [4-1:0] node56785;
	wire [4-1:0] node56788;
	wire [4-1:0] node56789;
	wire [4-1:0] node56792;
	wire [4-1:0] node56795;
	wire [4-1:0] node56796;
	wire [4-1:0] node56797;
	wire [4-1:0] node56798;
	wire [4-1:0] node56801;
	wire [4-1:0] node56804;
	wire [4-1:0] node56805;
	wire [4-1:0] node56808;
	wire [4-1:0] node56811;
	wire [4-1:0] node56812;
	wire [4-1:0] node56815;
	wire [4-1:0] node56818;
	wire [4-1:0] node56819;
	wire [4-1:0] node56820;
	wire [4-1:0] node56821;
	wire [4-1:0] node56822;
	wire [4-1:0] node56825;
	wire [4-1:0] node56828;
	wire [4-1:0] node56829;
	wire [4-1:0] node56832;
	wire [4-1:0] node56835;
	wire [4-1:0] node56836;
	wire [4-1:0] node56839;
	wire [4-1:0] node56842;
	wire [4-1:0] node56843;
	wire [4-1:0] node56846;
	wire [4-1:0] node56849;
	wire [4-1:0] node56850;
	wire [4-1:0] node56851;
	wire [4-1:0] node56852;
	wire [4-1:0] node56853;
	wire [4-1:0] node56856;
	wire [4-1:0] node56859;
	wire [4-1:0] node56860;
	wire [4-1:0] node56863;
	wire [4-1:0] node56866;
	wire [4-1:0] node56867;
	wire [4-1:0] node56868;
	wire [4-1:0] node56869;
	wire [4-1:0] node56872;
	wire [4-1:0] node56875;
	wire [4-1:0] node56877;
	wire [4-1:0] node56880;
	wire [4-1:0] node56881;
	wire [4-1:0] node56882;
	wire [4-1:0] node56885;
	wire [4-1:0] node56888;
	wire [4-1:0] node56889;
	wire [4-1:0] node56892;
	wire [4-1:0] node56895;
	wire [4-1:0] node56896;
	wire [4-1:0] node56897;
	wire [4-1:0] node56898;
	wire [4-1:0] node56899;
	wire [4-1:0] node56902;
	wire [4-1:0] node56905;
	wire [4-1:0] node56906;
	wire [4-1:0] node56909;
	wire [4-1:0] node56912;
	wire [4-1:0] node56913;
	wire [4-1:0] node56916;
	wire [4-1:0] node56919;
	wire [4-1:0] node56920;
	wire [4-1:0] node56921;
	wire [4-1:0] node56924;
	wire [4-1:0] node56927;
	wire [4-1:0] node56928;
	wire [4-1:0] node56931;
	wire [4-1:0] node56934;
	wire [4-1:0] node56935;
	wire [4-1:0] node56936;
	wire [4-1:0] node56937;
	wire [4-1:0] node56938;
	wire [4-1:0] node56939;
	wire [4-1:0] node56940;
	wire [4-1:0] node56941;
	wire [4-1:0] node56944;
	wire [4-1:0] node56947;
	wire [4-1:0] node56949;
	wire [4-1:0] node56952;
	wire [4-1:0] node56953;
	wire [4-1:0] node56956;
	wire [4-1:0] node56959;
	wire [4-1:0] node56960;
	wire [4-1:0] node56961;
	wire [4-1:0] node56962;
	wire [4-1:0] node56965;
	wire [4-1:0] node56968;
	wire [4-1:0] node56969;
	wire [4-1:0] node56972;
	wire [4-1:0] node56975;
	wire [4-1:0] node56976;
	wire [4-1:0] node56979;
	wire [4-1:0] node56982;
	wire [4-1:0] node56983;
	wire [4-1:0] node56984;
	wire [4-1:0] node56985;
	wire [4-1:0] node56986;
	wire [4-1:0] node56989;
	wire [4-1:0] node56992;
	wire [4-1:0] node56993;
	wire [4-1:0] node56996;
	wire [4-1:0] node56999;
	wire [4-1:0] node57000;
	wire [4-1:0] node57003;
	wire [4-1:0] node57006;
	wire [4-1:0] node57007;
	wire [4-1:0] node57008;
	wire [4-1:0] node57009;
	wire [4-1:0] node57012;
	wire [4-1:0] node57015;
	wire [4-1:0] node57016;
	wire [4-1:0] node57019;
	wire [4-1:0] node57022;
	wire [4-1:0] node57023;
	wire [4-1:0] node57024;
	wire [4-1:0] node57027;
	wire [4-1:0] node57030;
	wire [4-1:0] node57031;
	wire [4-1:0] node57034;
	wire [4-1:0] node57037;
	wire [4-1:0] node57038;
	wire [4-1:0] node57039;
	wire [4-1:0] node57040;
	wire [4-1:0] node57041;
	wire [4-1:0] node57042;
	wire [4-1:0] node57045;
	wire [4-1:0] node57048;
	wire [4-1:0] node57049;
	wire [4-1:0] node57053;
	wire [4-1:0] node57054;
	wire [4-1:0] node57055;
	wire [4-1:0] node57058;
	wire [4-1:0] node57061;
	wire [4-1:0] node57062;
	wire [4-1:0] node57065;
	wire [4-1:0] node57068;
	wire [4-1:0] node57069;
	wire [4-1:0] node57070;
	wire [4-1:0] node57071;
	wire [4-1:0] node57074;
	wire [4-1:0] node57077;
	wire [4-1:0] node57078;
	wire [4-1:0] node57081;
	wire [4-1:0] node57084;
	wire [4-1:0] node57085;
	wire [4-1:0] node57086;
	wire [4-1:0] node57090;
	wire [4-1:0] node57091;
	wire [4-1:0] node57094;
	wire [4-1:0] node57097;
	wire [4-1:0] node57098;
	wire [4-1:0] node57099;
	wire [4-1:0] node57100;
	wire [4-1:0] node57101;
	wire [4-1:0] node57105;
	wire [4-1:0] node57106;
	wire [4-1:0] node57109;
	wire [4-1:0] node57112;
	wire [4-1:0] node57113;
	wire [4-1:0] node57116;
	wire [4-1:0] node57119;
	wire [4-1:0] node57120;
	wire [4-1:0] node57121;
	wire [4-1:0] node57124;
	wire [4-1:0] node57127;
	wire [4-1:0] node57128;
	wire [4-1:0] node57131;
	wire [4-1:0] node57134;
	wire [4-1:0] node57135;
	wire [4-1:0] node57136;
	wire [4-1:0] node57137;
	wire [4-1:0] node57138;
	wire [4-1:0] node57139;
	wire [4-1:0] node57140;
	wire [4-1:0] node57143;
	wire [4-1:0] node57146;
	wire [4-1:0] node57147;
	wire [4-1:0] node57150;
	wire [4-1:0] node57153;
	wire [4-1:0] node57154;
	wire [4-1:0] node57155;
	wire [4-1:0] node57158;
	wire [4-1:0] node57161;
	wire [4-1:0] node57162;
	wire [4-1:0] node57165;
	wire [4-1:0] node57168;
	wire [4-1:0] node57169;
	wire [4-1:0] node57170;
	wire [4-1:0] node57171;
	wire [4-1:0] node57174;
	wire [4-1:0] node57177;
	wire [4-1:0] node57178;
	wire [4-1:0] node57181;
	wire [4-1:0] node57184;
	wire [4-1:0] node57185;
	wire [4-1:0] node57188;
	wire [4-1:0] node57191;
	wire [4-1:0] node57192;
	wire [4-1:0] node57193;
	wire [4-1:0] node57194;
	wire [4-1:0] node57195;
	wire [4-1:0] node57198;
	wire [4-1:0] node57201;
	wire [4-1:0] node57202;
	wire [4-1:0] node57205;
	wire [4-1:0] node57208;
	wire [4-1:0] node57209;
	wire [4-1:0] node57210;
	wire [4-1:0] node57213;
	wire [4-1:0] node57216;
	wire [4-1:0] node57217;
	wire [4-1:0] node57220;
	wire [4-1:0] node57223;
	wire [4-1:0] node57224;
	wire [4-1:0] node57227;
	wire [4-1:0] node57230;
	wire [4-1:0] node57231;
	wire [4-1:0] node57232;
	wire [4-1:0] node57233;
	wire [4-1:0] node57234;
	wire [4-1:0] node57235;
	wire [4-1:0] node57238;
	wire [4-1:0] node57241;
	wire [4-1:0] node57243;
	wire [4-1:0] node57246;
	wire [4-1:0] node57247;
	wire [4-1:0] node57250;
	wire [4-1:0] node57253;
	wire [4-1:0] node57254;
	wire [4-1:0] node57255;
	wire [4-1:0] node57256;
	wire [4-1:0] node57259;
	wire [4-1:0] node57262;
	wire [4-1:0] node57263;
	wire [4-1:0] node57266;
	wire [4-1:0] node57269;
	wire [4-1:0] node57270;
	wire [4-1:0] node57271;
	wire [4-1:0] node57274;
	wire [4-1:0] node57277;
	wire [4-1:0] node57278;
	wire [4-1:0] node57281;
	wire [4-1:0] node57284;
	wire [4-1:0] node57285;
	wire [4-1:0] node57286;
	wire [4-1:0] node57287;
	wire [4-1:0] node57290;
	wire [4-1:0] node57293;
	wire [4-1:0] node57294;
	wire [4-1:0] node57295;
	wire [4-1:0] node57298;
	wire [4-1:0] node57301;
	wire [4-1:0] node57303;
	wire [4-1:0] node57306;
	wire [4-1:0] node57307;
	wire [4-1:0] node57310;

	assign outp = (inp[9]) ? node28536 : node1;
		assign node1 = (inp[4]) ? node14259 : node2;
			assign node2 = (inp[10]) ? node7166 : node3;
				assign node3 = (inp[12]) ? node3511 : node4;
					assign node4 = (inp[15]) ? node1710 : node5;
						assign node5 = (inp[0]) ? node833 : node6;
							assign node6 = (inp[3]) ? node404 : node7;
								assign node7 = (inp[7]) ? node179 : node8;
									assign node8 = (inp[8]) ? node80 : node9;
										assign node9 = (inp[2]) ? node57 : node10;
											assign node10 = (inp[14]) ? node34 : node11;
												assign node11 = (inp[6]) ? node23 : node12;
													assign node12 = (inp[11]) ? node18 : node13;
														assign node13 = (inp[13]) ? node15 : 4'b1111;
															assign node15 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node18 = (inp[1]) ? node20 : 4'b0111;
															assign node20 = (inp[13]) ? 4'b1111 : 4'b0111;
													assign node23 = (inp[11]) ? node29 : node24;
														assign node24 = (inp[13]) ? node26 : 4'b0111;
															assign node26 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node29 = (inp[13]) ? node31 : 4'b1111;
															assign node31 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node34 = (inp[13]) ? node42 : node35;
													assign node35 = (inp[6]) ? node39 : node36;
														assign node36 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node39 = (inp[11]) ? 4'b1110 : 4'b0110;
													assign node42 = (inp[1]) ? node50 : node43;
														assign node43 = (inp[11]) ? node47 : node44;
															assign node44 = (inp[6]) ? 4'b0110 : 4'b1110;
															assign node47 = (inp[6]) ? 4'b1110 : 4'b0110;
														assign node50 = (inp[6]) ? node54 : node51;
															assign node51 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node54 = (inp[11]) ? 4'b0110 : 4'b1110;
											assign node57 = (inp[11]) ? node69 : node58;
												assign node58 = (inp[6]) ? node64 : node59;
													assign node59 = (inp[1]) ? node61 : 4'b1110;
														assign node61 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node64 = (inp[1]) ? node66 : 4'b0110;
														assign node66 = (inp[13]) ? 4'b1110 : 4'b0110;
												assign node69 = (inp[6]) ? node75 : node70;
													assign node70 = (inp[13]) ? node72 : 4'b0110;
														assign node72 = (inp[1]) ? 4'b1110 : 4'b0110;
													assign node75 = (inp[13]) ? node77 : 4'b1110;
														assign node77 = (inp[1]) ? 4'b0110 : 4'b1110;
										assign node80 = (inp[14]) ? node128 : node81;
											assign node81 = (inp[2]) ? node101 : node82;
												assign node82 = (inp[6]) ? node94 : node83;
													assign node83 = (inp[11]) ? node89 : node84;
														assign node84 = (inp[13]) ? node86 : 4'b1110;
															assign node86 = (inp[1]) ? 4'b0110 : 4'b1110;
														assign node89 = (inp[13]) ? node91 : 4'b0110;
															assign node91 = (inp[1]) ? 4'b1110 : 4'b0110;
													assign node94 = (inp[11]) ? 4'b1110 : node95;
														assign node95 = (inp[1]) ? node97 : 4'b0110;
															assign node97 = (inp[13]) ? 4'b1110 : 4'b0110;
												assign node101 = (inp[5]) ? node115 : node102;
													assign node102 = (inp[6]) ? node110 : node103;
														assign node103 = (inp[11]) ? node107 : node104;
															assign node104 = (inp[1]) ? 4'b0111 : 4'b1111;
															assign node107 = (inp[13]) ? 4'b1111 : 4'b0111;
														assign node110 = (inp[11]) ? 4'b0111 : node111;
															assign node111 = (inp[1]) ? 4'b1111 : 4'b0111;
													assign node115 = (inp[1]) ? node123 : node116;
														assign node116 = (inp[11]) ? node120 : node117;
															assign node117 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node120 = (inp[6]) ? 4'b0111 : 4'b0111;
														assign node123 = (inp[13]) ? 4'b1111 : node124;
															assign node124 = (inp[6]) ? 4'b0111 : 4'b0111;
											assign node128 = (inp[5]) ? node156 : node129;
												assign node129 = (inp[2]) ? node143 : node130;
													assign node130 = (inp[6]) ? node138 : node131;
														assign node131 = (inp[11]) ? node135 : node132;
															assign node132 = (inp[1]) ? 4'b0111 : 4'b1111;
															assign node135 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node138 = (inp[11]) ? 4'b0111 : node139;
															assign node139 = (inp[13]) ? 4'b1111 : 4'b0111;
													assign node143 = (inp[1]) ? node151 : node144;
														assign node144 = (inp[13]) ? node148 : node145;
															assign node145 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node148 = (inp[11]) ? 4'b0111 : 4'b0111;
														assign node151 = (inp[6]) ? 4'b1111 : node152;
															assign node152 = (inp[11]) ? 4'b1111 : 4'b0111;
												assign node156 = (inp[6]) ? node168 : node157;
													assign node157 = (inp[11]) ? node163 : node158;
														assign node158 = (inp[13]) ? 4'b0111 : node159;
															assign node159 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node163 = (inp[1]) ? 4'b1111 : node164;
															assign node164 = (inp[13]) ? 4'b1111 : 4'b0111;
													assign node168 = (inp[11]) ? node174 : node169;
														assign node169 = (inp[13]) ? 4'b1111 : node170;
															assign node170 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node174 = (inp[13]) ? 4'b0111 : node175;
															assign node175 = (inp[1]) ? 4'b0111 : 4'b1111;
									assign node179 = (inp[8]) ? node287 : node180;
										assign node180 = (inp[2]) ? node234 : node181;
											assign node181 = (inp[14]) ? node205 : node182;
												assign node182 = (inp[11]) ? node194 : node183;
													assign node183 = (inp[6]) ? node189 : node184;
														assign node184 = (inp[13]) ? node186 : 4'b1110;
															assign node186 = (inp[1]) ? 4'b0110 : 4'b1110;
														assign node189 = (inp[13]) ? node191 : 4'b0110;
															assign node191 = (inp[1]) ? 4'b1110 : 4'b0110;
													assign node194 = (inp[6]) ? node200 : node195;
														assign node195 = (inp[13]) ? node197 : 4'b0110;
															assign node197 = (inp[1]) ? 4'b1110 : 4'b0110;
														assign node200 = (inp[13]) ? node202 : 4'b1110;
															assign node202 = (inp[1]) ? 4'b0110 : 4'b1110;
												assign node205 = (inp[13]) ? node221 : node206;
													assign node206 = (inp[11]) ? node214 : node207;
														assign node207 = (inp[5]) ? node211 : node208;
															assign node208 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node211 = (inp[1]) ? 4'b0111 : 4'b0111;
														assign node214 = (inp[5]) ? node218 : node215;
															assign node215 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node218 = (inp[6]) ? 4'b0111 : 4'b0111;
													assign node221 = (inp[1]) ? node229 : node222;
														assign node222 = (inp[5]) ? node226 : node223;
															assign node223 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node226 = (inp[11]) ? 4'b0111 : 4'b0111;
														assign node229 = (inp[6]) ? 4'b0111 : node230;
															assign node230 = (inp[11]) ? 4'b1111 : 4'b0111;
											assign node234 = (inp[13]) ? node264 : node235;
												assign node235 = (inp[14]) ? node251 : node236;
													assign node236 = (inp[11]) ? node244 : node237;
														assign node237 = (inp[6]) ? node241 : node238;
															assign node238 = (inp[1]) ? 4'b0111 : 4'b1111;
															assign node241 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node244 = (inp[6]) ? node248 : node245;
															assign node245 = (inp[1]) ? 4'b1111 : 4'b0111;
															assign node248 = (inp[1]) ? 4'b0111 : 4'b1111;
													assign node251 = (inp[5]) ? node259 : node252;
														assign node252 = (inp[11]) ? node256 : node253;
															assign node253 = (inp[1]) ? 4'b0111 : 4'b0111;
															assign node256 = (inp[6]) ? 4'b0111 : 4'b0111;
														assign node259 = (inp[6]) ? node261 : 4'b0111;
															assign node261 = (inp[11]) ? 4'b0111 : 4'b0111;
												assign node264 = (inp[5]) ? node272 : node265;
													assign node265 = (inp[6]) ? node269 : node266;
														assign node266 = (inp[11]) ? 4'b1111 : 4'b0111;
														assign node269 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node272 = (inp[1]) ? node280 : node273;
														assign node273 = (inp[11]) ? node277 : node274;
															assign node274 = (inp[6]) ? 4'b1111 : 4'b0111;
															assign node277 = (inp[6]) ? 4'b0111 : 4'b1111;
														assign node280 = (inp[6]) ? node284 : node281;
															assign node281 = (inp[11]) ? 4'b1111 : 4'b0111;
															assign node284 = (inp[11]) ? 4'b0111 : 4'b1111;
										assign node287 = (inp[14]) ? node343 : node288;
											assign node288 = (inp[2]) ? node320 : node289;
												assign node289 = (inp[13]) ? node305 : node290;
													assign node290 = (inp[1]) ? node298 : node291;
														assign node291 = (inp[5]) ? node295 : node292;
															assign node292 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node295 = (inp[11]) ? 4'b0111 : 4'b0111;
														assign node298 = (inp[5]) ? node302 : node299;
															assign node299 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node302 = (inp[6]) ? 4'b0111 : 4'b0111;
													assign node305 = (inp[1]) ? node313 : node306;
														assign node306 = (inp[5]) ? node310 : node307;
															assign node307 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node310 = (inp[6]) ? 4'b0111 : 4'b0111;
														assign node313 = (inp[6]) ? node317 : node314;
															assign node314 = (inp[11]) ? 4'b1111 : 4'b0111;
															assign node317 = (inp[11]) ? 4'b0111 : 4'b1111;
												assign node320 = (inp[1]) ? node336 : node321;
													assign node321 = (inp[13]) ? node329 : node322;
														assign node322 = (inp[6]) ? node326 : node323;
															assign node323 = (inp[11]) ? 4'b0110 : 4'b1110;
															assign node326 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node329 = (inp[11]) ? node333 : node330;
															assign node330 = (inp[6]) ? 4'b1110 : 4'b0110;
															assign node333 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node336 = (inp[6]) ? node340 : node337;
														assign node337 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node340 = (inp[11]) ? 4'b0110 : 4'b1110;
											assign node343 = (inp[1]) ? node375 : node344;
												assign node344 = (inp[5]) ? node360 : node345;
													assign node345 = (inp[11]) ? node353 : node346;
														assign node346 = (inp[13]) ? node350 : node347;
															assign node347 = (inp[6]) ? 4'b0110 : 4'b1110;
															assign node350 = (inp[6]) ? 4'b1110 : 4'b0110;
														assign node353 = (inp[2]) ? node357 : node354;
															assign node354 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node357 = (inp[13]) ? 4'b0110 : 4'b0110;
													assign node360 = (inp[11]) ? node368 : node361;
														assign node361 = (inp[13]) ? node365 : node362;
															assign node362 = (inp[6]) ? 4'b0110 : 4'b1110;
															assign node365 = (inp[6]) ? 4'b1110 : 4'b0110;
														assign node368 = (inp[6]) ? node372 : node369;
															assign node369 = (inp[13]) ? 4'b1110 : 4'b0110;
															assign node372 = (inp[13]) ? 4'b0110 : 4'b1110;
												assign node375 = (inp[5]) ? node389 : node376;
													assign node376 = (inp[2]) ? node384 : node377;
														assign node377 = (inp[13]) ? node381 : node378;
															assign node378 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node381 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node384 = (inp[13]) ? node386 : 4'b0110;
															assign node386 = (inp[11]) ? 4'b0110 : 4'b0110;
													assign node389 = (inp[13]) ? node397 : node390;
														assign node390 = (inp[6]) ? node394 : node391;
															assign node391 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node394 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node397 = (inp[11]) ? node401 : node398;
															assign node398 = (inp[6]) ? 4'b1110 : 4'b0110;
															assign node401 = (inp[6]) ? 4'b0110 : 4'b1110;
								assign node404 = (inp[5]) ? node622 : node405;
									assign node405 = (inp[11]) ? node523 : node406;
										assign node406 = (inp[6]) ? node466 : node407;
											assign node407 = (inp[13]) ? node439 : node408;
												assign node408 = (inp[1]) ? node424 : node409;
													assign node409 = (inp[2]) ? node417 : node410;
														assign node410 = (inp[8]) ? node414 : node411;
															assign node411 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node414 = (inp[14]) ? 4'b1110 : 4'b1110;
														assign node417 = (inp[7]) ? node421 : node418;
															assign node418 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node421 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node424 = (inp[7]) ? node432 : node425;
														assign node425 = (inp[8]) ? node429 : node426;
															assign node426 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node429 = (inp[14]) ? 4'b0111 : 4'b1110;
														assign node432 = (inp[8]) ? node436 : node433;
															assign node433 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node436 = (inp[14]) ? 4'b0110 : 4'b0110;
												assign node439 = (inp[1]) ? node453 : node440;
													assign node440 = (inp[7]) ? node448 : node441;
														assign node441 = (inp[8]) ? node445 : node442;
															assign node442 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node445 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node448 = (inp[8]) ? 4'b0110 : node449;
															assign node449 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node453 = (inp[7]) ? node459 : node454;
														assign node454 = (inp[14]) ? 4'b0111 : node455;
															assign node455 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node459 = (inp[8]) ? node463 : node460;
															assign node460 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node463 = (inp[14]) ? 4'b0110 : 4'b0110;
											assign node466 = (inp[13]) ? node494 : node467;
												assign node467 = (inp[1]) ? node483 : node468;
													assign node468 = (inp[8]) ? node476 : node469;
														assign node469 = (inp[7]) ? node473 : node470;
															assign node470 = (inp[2]) ? 4'b0110 : 4'b0110;
															assign node473 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node476 = (inp[7]) ? node480 : node477;
															assign node477 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node480 = (inp[2]) ? 4'b0110 : 4'b0110;
													assign node483 = (inp[8]) ? node491 : node484;
														assign node484 = (inp[7]) ? node488 : node485;
															assign node485 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node488 = (inp[2]) ? 4'b1111 : 4'b0110;
														assign node491 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node494 = (inp[1]) ? node510 : node495;
													assign node495 = (inp[7]) ? node503 : node496;
														assign node496 = (inp[8]) ? node500 : node497;
															assign node497 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node500 = (inp[2]) ? 4'b1111 : 4'b0110;
														assign node503 = (inp[8]) ? node507 : node504;
															assign node504 = (inp[14]) ? 4'b1111 : 4'b0110;
															assign node507 = (inp[14]) ? 4'b1110 : 4'b1110;
													assign node510 = (inp[7]) ? node516 : node511;
														assign node511 = (inp[8]) ? node513 : 4'b1110;
															assign node513 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node516 = (inp[8]) ? node520 : node517;
															assign node517 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node520 = (inp[14]) ? 4'b1110 : 4'b1110;
										assign node523 = (inp[7]) ? node575 : node524;
											assign node524 = (inp[8]) ? node552 : node525;
												assign node525 = (inp[14]) ? node541 : node526;
													assign node526 = (inp[2]) ? node534 : node527;
														assign node527 = (inp[6]) ? node531 : node528;
															assign node528 = (inp[1]) ? 4'b0111 : 4'b0111;
															assign node531 = (inp[13]) ? 4'b0111 : 4'b1111;
														assign node534 = (inp[6]) ? node538 : node535;
															assign node535 = (inp[1]) ? 4'b0110 : 4'b0110;
															assign node538 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node541 = (inp[6]) ? node547 : node542;
														assign node542 = (inp[13]) ? node544 : 4'b0110;
															assign node544 = (inp[1]) ? 4'b1110 : 4'b0110;
														assign node547 = (inp[13]) ? node549 : 4'b1110;
															assign node549 = (inp[1]) ? 4'b0110 : 4'b1110;
												assign node552 = (inp[14]) ? node564 : node553;
													assign node553 = (inp[2]) ? node559 : node554;
														assign node554 = (inp[6]) ? node556 : 4'b0110;
															assign node556 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node559 = (inp[6]) ? node561 : 4'b1111;
															assign node561 = (inp[13]) ? 4'b0111 : 4'b0111;
													assign node564 = (inp[6]) ? node570 : node565;
														assign node565 = (inp[1]) ? 4'b1111 : node566;
															assign node566 = (inp[13]) ? 4'b1111 : 4'b0111;
														assign node570 = (inp[13]) ? 4'b0111 : node571;
															assign node571 = (inp[1]) ? 4'b0111 : 4'b1111;
											assign node575 = (inp[8]) ? node603 : node576;
												assign node576 = (inp[14]) ? node592 : node577;
													assign node577 = (inp[2]) ? node585 : node578;
														assign node578 = (inp[6]) ? node582 : node579;
															assign node579 = (inp[13]) ? 4'b0110 : 4'b0110;
															assign node582 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node585 = (inp[6]) ? node589 : node586;
															assign node586 = (inp[13]) ? 4'b1111 : 4'b0111;
															assign node589 = (inp[1]) ? 4'b0111 : 4'b1111;
													assign node592 = (inp[6]) ? node598 : node593;
														assign node593 = (inp[13]) ? 4'b1111 : node594;
															assign node594 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node598 = (inp[13]) ? 4'b0111 : node599;
															assign node599 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node603 = (inp[6]) ? node615 : node604;
													assign node604 = (inp[1]) ? node610 : node605;
														assign node605 = (inp[13]) ? 4'b1110 : node606;
															assign node606 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node610 = (inp[2]) ? 4'b1110 : node611;
															assign node611 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node615 = (inp[1]) ? 4'b0110 : node616;
														assign node616 = (inp[13]) ? 4'b0110 : node617;
															assign node617 = (inp[2]) ? 4'b1110 : 4'b1110;
									assign node622 = (inp[8]) ? node726 : node623;
										assign node623 = (inp[7]) ? node679 : node624;
											assign node624 = (inp[2]) ? node656 : node625;
												assign node625 = (inp[14]) ? node641 : node626;
													assign node626 = (inp[13]) ? node634 : node627;
														assign node627 = (inp[6]) ? node631 : node628;
															assign node628 = (inp[11]) ? 4'b0101 : 4'b1101;
															assign node631 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node634 = (inp[1]) ? node638 : node635;
															assign node635 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node638 = (inp[11]) ? 4'b0101 : 4'b0101;
													assign node641 = (inp[13]) ? node649 : node642;
														assign node642 = (inp[1]) ? node646 : node643;
															assign node643 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node646 = (inp[6]) ? 4'b0100 : 4'b0100;
														assign node649 = (inp[1]) ? node653 : node650;
															assign node650 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node653 = (inp[11]) ? 4'b0100 : 4'b0100;
												assign node656 = (inp[6]) ? node668 : node657;
													assign node657 = (inp[11]) ? node663 : node658;
														assign node658 = (inp[1]) ? node660 : 4'b1100;
															assign node660 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node663 = (inp[1]) ? node665 : 4'b0100;
															assign node665 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node668 = (inp[11]) ? node674 : node669;
														assign node669 = (inp[13]) ? node671 : 4'b0100;
															assign node671 = (inp[1]) ? 4'b1100 : 4'b0100;
														assign node674 = (inp[1]) ? node676 : 4'b1100;
															assign node676 = (inp[13]) ? 4'b0100 : 4'b1100;
											assign node679 = (inp[2]) ? node705 : node680;
												assign node680 = (inp[14]) ? node694 : node681;
													assign node681 = (inp[11]) ? node687 : node682;
														assign node682 = (inp[6]) ? node684 : 4'b1100;
															assign node684 = (inp[1]) ? 4'b1100 : 4'b0100;
														assign node687 = (inp[6]) ? node691 : node688;
															assign node688 = (inp[13]) ? 4'b0100 : 4'b0100;
															assign node691 = (inp[1]) ? 4'b0100 : 4'b1100;
													assign node694 = (inp[11]) ? node700 : node695;
														assign node695 = (inp[1]) ? 4'b0101 : node696;
															assign node696 = (inp[13]) ? 4'b0101 : 4'b0101;
														assign node700 = (inp[6]) ? 4'b0101 : node701;
															assign node701 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node705 = (inp[1]) ? node719 : node706;
													assign node706 = (inp[14]) ? node714 : node707;
														assign node707 = (inp[11]) ? node711 : node708;
															assign node708 = (inp[13]) ? 4'b0101 : 4'b0101;
															assign node711 = (inp[6]) ? 4'b0101 : 4'b0101;
														assign node714 = (inp[11]) ? node716 : 4'b1101;
															assign node716 = (inp[6]) ? 4'b0101 : 4'b0101;
													assign node719 = (inp[11]) ? node723 : node720;
														assign node720 = (inp[6]) ? 4'b1101 : 4'b0101;
														assign node723 = (inp[6]) ? 4'b0101 : 4'b1101;
										assign node726 = (inp[7]) ? node774 : node727;
											assign node727 = (inp[2]) ? node757 : node728;
												assign node728 = (inp[14]) ? node744 : node729;
													assign node729 = (inp[13]) ? node737 : node730;
														assign node730 = (inp[1]) ? node734 : node731;
															assign node731 = (inp[11]) ? 4'b0100 : 4'b0100;
															assign node734 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node737 = (inp[11]) ? node741 : node738;
															assign node738 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node741 = (inp[6]) ? 4'b0100 : 4'b0100;
													assign node744 = (inp[13]) ? node750 : node745;
														assign node745 = (inp[6]) ? 4'b1101 : node746;
															assign node746 = (inp[1]) ? 4'b0101 : 4'b0101;
														assign node750 = (inp[6]) ? node754 : node751;
															assign node751 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node754 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node757 = (inp[11]) ? node765 : node758;
													assign node758 = (inp[6]) ? 4'b1101 : node759;
														assign node759 = (inp[13]) ? 4'b0101 : node760;
															assign node760 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node765 = (inp[6]) ? node769 : node766;
														assign node766 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node769 = (inp[13]) ? 4'b0101 : node770;
															assign node770 = (inp[1]) ? 4'b0101 : 4'b1101;
											assign node774 = (inp[14]) ? node802 : node775;
												assign node775 = (inp[2]) ? node789 : node776;
													assign node776 = (inp[11]) ? node784 : node777;
														assign node777 = (inp[6]) ? node781 : node778;
															assign node778 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node781 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node784 = (inp[6]) ? 4'b0101 : node785;
															assign node785 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node789 = (inp[13]) ? node795 : node790;
														assign node790 = (inp[1]) ? node792 : 4'b0100;
															assign node792 = (inp[6]) ? 4'b0100 : 4'b0100;
														assign node795 = (inp[6]) ? node799 : node796;
															assign node796 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node799 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node802 = (inp[2]) ? node818 : node803;
													assign node803 = (inp[1]) ? node811 : node804;
														assign node804 = (inp[13]) ? node808 : node805;
															assign node805 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node808 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node811 = (inp[11]) ? node815 : node812;
															assign node812 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node815 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node818 = (inp[6]) ? node826 : node819;
														assign node819 = (inp[11]) ? node823 : node820;
															assign node820 = (inp[13]) ? 4'b0100 : 4'b0100;
															assign node823 = (inp[1]) ? 4'b1100 : 4'b0100;
														assign node826 = (inp[11]) ? node830 : node827;
															assign node827 = (inp[13]) ? 4'b1100 : 4'b0100;
															assign node830 = (inp[13]) ? 4'b0100 : 4'b0100;
							assign node833 = (inp[3]) ? node1259 : node834;
								assign node834 = (inp[13]) ? node1048 : node835;
									assign node835 = (inp[6]) ? node945 : node836;
										assign node836 = (inp[11]) ? node892 : node837;
											assign node837 = (inp[1]) ? node869 : node838;
												assign node838 = (inp[14]) ? node854 : node839;
													assign node839 = (inp[2]) ? node847 : node840;
														assign node840 = (inp[5]) ? node844 : node841;
															assign node841 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node844 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node847 = (inp[7]) ? node851 : node848;
															assign node848 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node851 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node854 = (inp[2]) ? node862 : node855;
														assign node855 = (inp[8]) ? node859 : node856;
															assign node856 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node859 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node862 = (inp[5]) ? node866 : node863;
															assign node863 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node866 = (inp[8]) ? 4'b1100 : 4'b1100;
												assign node869 = (inp[7]) ? node881 : node870;
													assign node870 = (inp[8]) ? node876 : node871;
														assign node871 = (inp[14]) ? 4'b1100 : node872;
															assign node872 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node876 = (inp[14]) ? 4'b0101 : node877;
															assign node877 = (inp[2]) ? 4'b0101 : 4'b1100;
													assign node881 = (inp[8]) ? node887 : node882;
														assign node882 = (inp[2]) ? 4'b0101 : node883;
															assign node883 = (inp[14]) ? 4'b0101 : 4'b1100;
														assign node887 = (inp[14]) ? 4'b0100 : node888;
															assign node888 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node892 = (inp[1]) ? node922 : node893;
												assign node893 = (inp[5]) ? node909 : node894;
													assign node894 = (inp[7]) ? node902 : node895;
														assign node895 = (inp[8]) ? node899 : node896;
															assign node896 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node899 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node902 = (inp[8]) ? node906 : node903;
															assign node903 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node906 = (inp[2]) ? 4'b0100 : 4'b0100;
													assign node909 = (inp[8]) ? node917 : node910;
														assign node910 = (inp[7]) ? node914 : node911;
															assign node911 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node914 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node917 = (inp[7]) ? node919 : 4'b0101;
															assign node919 = (inp[2]) ? 4'b0100 : 4'b0100;
												assign node922 = (inp[14]) ? node938 : node923;
													assign node923 = (inp[2]) ? node931 : node924;
														assign node924 = (inp[7]) ? node928 : node925;
															assign node925 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node928 = (inp[8]) ? 4'b1101 : 4'b0100;
														assign node931 = (inp[7]) ? node935 : node932;
															assign node932 = (inp[8]) ? 4'b1101 : 4'b0100;
															assign node935 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node938 = (inp[8]) ? node942 : node939;
														assign node939 = (inp[7]) ? 4'b1101 : 4'b0100;
														assign node942 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node945 = (inp[11]) ? node1001 : node946;
											assign node946 = (inp[1]) ? node978 : node947;
												assign node947 = (inp[14]) ? node963 : node948;
													assign node948 = (inp[7]) ? node956 : node949;
														assign node949 = (inp[8]) ? node953 : node950;
															assign node950 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node953 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node956 = (inp[8]) ? node960 : node957;
															assign node957 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node960 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node963 = (inp[5]) ? node971 : node964;
														assign node964 = (inp[7]) ? node968 : node965;
															assign node965 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node968 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node971 = (inp[8]) ? node975 : node972;
															assign node972 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node975 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node978 = (inp[8]) ? node990 : node979;
													assign node979 = (inp[7]) ? node985 : node980;
														assign node980 = (inp[2]) ? 4'b0100 : node981;
															assign node981 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node985 = (inp[2]) ? 4'b1101 : node986;
															assign node986 = (inp[14]) ? 4'b1101 : 4'b0100;
													assign node990 = (inp[7]) ? node996 : node991;
														assign node991 = (inp[2]) ? 4'b1101 : node992;
															assign node992 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node996 = (inp[14]) ? 4'b1100 : node997;
															assign node997 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node1001 = (inp[1]) ? node1025 : node1002;
												assign node1002 = (inp[7]) ? node1014 : node1003;
													assign node1003 = (inp[8]) ? node1009 : node1004;
														assign node1004 = (inp[14]) ? 4'b1100 : node1005;
															assign node1005 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node1009 = (inp[2]) ? 4'b1101 : node1010;
															assign node1010 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node1014 = (inp[8]) ? node1020 : node1015;
														assign node1015 = (inp[2]) ? 4'b1101 : node1016;
															assign node1016 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node1020 = (inp[14]) ? 4'b1100 : node1021;
															assign node1021 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node1025 = (inp[8]) ? node1037 : node1026;
													assign node1026 = (inp[7]) ? node1032 : node1027;
														assign node1027 = (inp[2]) ? 4'b1100 : node1028;
															assign node1028 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node1032 = (inp[14]) ? 4'b0101 : node1033;
															assign node1033 = (inp[2]) ? 4'b0101 : 4'b1100;
													assign node1037 = (inp[7]) ? node1043 : node1038;
														assign node1038 = (inp[14]) ? 4'b0101 : node1039;
															assign node1039 = (inp[2]) ? 4'b0101 : 4'b1100;
														assign node1043 = (inp[2]) ? 4'b0100 : node1044;
															assign node1044 = (inp[14]) ? 4'b0100 : 4'b0101;
									assign node1048 = (inp[6]) ? node1150 : node1049;
										assign node1049 = (inp[11]) ? node1097 : node1050;
											assign node1050 = (inp[1]) ? node1074 : node1051;
												assign node1051 = (inp[8]) ? node1063 : node1052;
													assign node1052 = (inp[7]) ? node1058 : node1053;
														assign node1053 = (inp[2]) ? 4'b1100 : node1054;
															assign node1054 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node1058 = (inp[14]) ? 4'b0101 : node1059;
															assign node1059 = (inp[2]) ? 4'b0101 : 4'b1100;
													assign node1063 = (inp[7]) ? node1069 : node1064;
														assign node1064 = (inp[2]) ? 4'b0101 : node1065;
															assign node1065 = (inp[14]) ? 4'b0101 : 4'b1100;
														assign node1069 = (inp[14]) ? 4'b0100 : node1070;
															assign node1070 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node1074 = (inp[7]) ? node1086 : node1075;
													assign node1075 = (inp[8]) ? node1081 : node1076;
														assign node1076 = (inp[14]) ? 4'b0100 : node1077;
															assign node1077 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node1081 = (inp[14]) ? 4'b0101 : node1082;
															assign node1082 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node1086 = (inp[8]) ? node1092 : node1087;
														assign node1087 = (inp[2]) ? 4'b0101 : node1088;
															assign node1088 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node1092 = (inp[2]) ? 4'b0100 : node1093;
															assign node1093 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node1097 = (inp[1]) ? node1121 : node1098;
												assign node1098 = (inp[7]) ? node1110 : node1099;
													assign node1099 = (inp[8]) ? node1105 : node1100;
														assign node1100 = (inp[2]) ? 4'b0100 : node1101;
															assign node1101 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node1105 = (inp[2]) ? 4'b1101 : node1106;
															assign node1106 = (inp[14]) ? 4'b1101 : 4'b0100;
													assign node1110 = (inp[8]) ? node1116 : node1111;
														assign node1111 = (inp[14]) ? 4'b1101 : node1112;
															assign node1112 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node1116 = (inp[14]) ? 4'b1100 : node1117;
															assign node1117 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node1121 = (inp[2]) ? node1137 : node1122;
													assign node1122 = (inp[8]) ? node1130 : node1123;
														assign node1123 = (inp[5]) ? node1127 : node1124;
															assign node1124 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node1127 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node1130 = (inp[14]) ? node1134 : node1131;
															assign node1131 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node1134 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node1137 = (inp[5]) ? node1143 : node1138;
														assign node1138 = (inp[14]) ? 4'b1101 : node1139;
															assign node1139 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node1143 = (inp[7]) ? node1147 : node1144;
															assign node1144 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node1147 = (inp[8]) ? 4'b1100 : 4'b1101;
										assign node1150 = (inp[11]) ? node1204 : node1151;
											assign node1151 = (inp[1]) ? node1175 : node1152;
												assign node1152 = (inp[8]) ? node1164 : node1153;
													assign node1153 = (inp[7]) ? node1159 : node1154;
														assign node1154 = (inp[2]) ? 4'b0100 : node1155;
															assign node1155 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node1159 = (inp[14]) ? 4'b1101 : node1160;
															assign node1160 = (inp[2]) ? 4'b1101 : 4'b0100;
													assign node1164 = (inp[7]) ? node1170 : node1165;
														assign node1165 = (inp[14]) ? 4'b1101 : node1166;
															assign node1166 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node1170 = (inp[14]) ? 4'b1100 : node1171;
															assign node1171 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node1175 = (inp[5]) ? node1191 : node1176;
													assign node1176 = (inp[2]) ? node1184 : node1177;
														assign node1177 = (inp[7]) ? node1181 : node1178;
															assign node1178 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node1181 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node1184 = (inp[14]) ? node1188 : node1185;
															assign node1185 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node1188 = (inp[7]) ? 4'b1100 : 4'b1100;
													assign node1191 = (inp[14]) ? node1197 : node1192;
														assign node1192 = (inp[8]) ? 4'b1100 : node1193;
															assign node1193 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node1197 = (inp[8]) ? node1201 : node1198;
															assign node1198 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node1201 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node1204 = (inp[1]) ? node1228 : node1205;
												assign node1205 = (inp[8]) ? node1217 : node1206;
													assign node1206 = (inp[7]) ? node1212 : node1207;
														assign node1207 = (inp[14]) ? 4'b1100 : node1208;
															assign node1208 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node1212 = (inp[14]) ? 4'b0101 : node1213;
															assign node1213 = (inp[2]) ? 4'b0101 : 4'b1100;
													assign node1217 = (inp[7]) ? node1223 : node1218;
														assign node1218 = (inp[2]) ? 4'b0101 : node1219;
															assign node1219 = (inp[14]) ? 4'b0101 : 4'b1100;
														assign node1223 = (inp[2]) ? 4'b0100 : node1224;
															assign node1224 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node1228 = (inp[2]) ? node1244 : node1229;
													assign node1229 = (inp[7]) ? node1237 : node1230;
														assign node1230 = (inp[14]) ? node1234 : node1231;
															assign node1231 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node1234 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node1237 = (inp[14]) ? node1241 : node1238;
															assign node1238 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node1241 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node1244 = (inp[14]) ? node1252 : node1245;
														assign node1245 = (inp[8]) ? node1249 : node1246;
															assign node1246 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node1249 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node1252 = (inp[7]) ? node1256 : node1253;
															assign node1253 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node1256 = (inp[8]) ? 4'b0100 : 4'b0101;
								assign node1259 = (inp[5]) ? node1497 : node1260;
									assign node1260 = (inp[6]) ? node1378 : node1261;
										assign node1261 = (inp[11]) ? node1321 : node1262;
											assign node1262 = (inp[1]) ? node1290 : node1263;
												assign node1263 = (inp[13]) ? node1277 : node1264;
													assign node1264 = (inp[14]) ? node1270 : node1265;
														assign node1265 = (inp[2]) ? node1267 : 4'b1100;
															assign node1267 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node1270 = (inp[2]) ? node1274 : node1271;
															assign node1271 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node1274 = (inp[7]) ? 4'b1100 : 4'b1100;
													assign node1277 = (inp[8]) ? node1285 : node1278;
														assign node1278 = (inp[7]) ? node1282 : node1279;
															assign node1279 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node1282 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node1285 = (inp[7]) ? node1287 : 4'b0101;
															assign node1287 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node1290 = (inp[13]) ? node1306 : node1291;
													assign node1291 = (inp[7]) ? node1299 : node1292;
														assign node1292 = (inp[8]) ? node1296 : node1293;
															assign node1293 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node1296 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node1299 = (inp[8]) ? node1303 : node1300;
															assign node1300 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node1303 = (inp[2]) ? 4'b0100 : 4'b0100;
													assign node1306 = (inp[14]) ? node1314 : node1307;
														assign node1307 = (inp[8]) ? node1311 : node1308;
															assign node1308 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node1311 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node1314 = (inp[7]) ? node1318 : node1315;
															assign node1315 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node1318 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node1321 = (inp[13]) ? node1347 : node1322;
												assign node1322 = (inp[1]) ? node1334 : node1323;
													assign node1323 = (inp[8]) ? node1329 : node1324;
														assign node1324 = (inp[7]) ? 4'b0101 : node1325;
															assign node1325 = (inp[2]) ? 4'b0100 : 4'b0100;
														assign node1329 = (inp[14]) ? 4'b0100 : node1330;
															assign node1330 = (inp[2]) ? 4'b0100 : 4'b0100;
													assign node1334 = (inp[7]) ? node1342 : node1335;
														assign node1335 = (inp[8]) ? node1339 : node1336;
															assign node1336 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node1339 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node1342 = (inp[14]) ? node1344 : 4'b0100;
															assign node1344 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node1347 = (inp[1]) ? node1363 : node1348;
													assign node1348 = (inp[7]) ? node1356 : node1349;
														assign node1349 = (inp[8]) ? node1353 : node1350;
															assign node1350 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node1353 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node1356 = (inp[8]) ? node1360 : node1357;
															assign node1357 = (inp[2]) ? 4'b1101 : 4'b0100;
															assign node1360 = (inp[14]) ? 4'b1100 : 4'b1100;
													assign node1363 = (inp[2]) ? node1371 : node1364;
														assign node1364 = (inp[7]) ? node1368 : node1365;
															assign node1365 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node1368 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node1371 = (inp[8]) ? node1375 : node1372;
															assign node1372 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node1375 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node1378 = (inp[11]) ? node1438 : node1379;
											assign node1379 = (inp[1]) ? node1407 : node1380;
												assign node1380 = (inp[13]) ? node1394 : node1381;
													assign node1381 = (inp[8]) ? node1389 : node1382;
														assign node1382 = (inp[7]) ? node1386 : node1383;
															assign node1383 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node1386 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node1389 = (inp[7]) ? node1391 : 4'b0101;
															assign node1391 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node1394 = (inp[7]) ? node1402 : node1395;
														assign node1395 = (inp[8]) ? node1399 : node1396;
															assign node1396 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node1399 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node1402 = (inp[8]) ? node1404 : 4'b1101;
															assign node1404 = (inp[14]) ? 4'b1100 : 4'b1100;
												assign node1407 = (inp[13]) ? node1423 : node1408;
													assign node1408 = (inp[8]) ? node1416 : node1409;
														assign node1409 = (inp[7]) ? node1413 : node1410;
															assign node1410 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node1413 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node1416 = (inp[7]) ? node1420 : node1417;
															assign node1417 = (inp[2]) ? 4'b1101 : 4'b0100;
															assign node1420 = (inp[14]) ? 4'b1100 : 4'b1100;
													assign node1423 = (inp[2]) ? node1431 : node1424;
														assign node1424 = (inp[14]) ? node1428 : node1425;
															assign node1425 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node1428 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node1431 = (inp[14]) ? node1435 : node1432;
															assign node1432 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node1435 = (inp[7]) ? 4'b1100 : 4'b1100;
											assign node1438 = (inp[1]) ? node1470 : node1439;
												assign node1439 = (inp[13]) ? node1455 : node1440;
													assign node1440 = (inp[8]) ? node1448 : node1441;
														assign node1441 = (inp[7]) ? node1445 : node1442;
															assign node1442 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node1445 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node1448 = (inp[7]) ? node1452 : node1449;
															assign node1449 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node1452 = (inp[2]) ? 4'b1100 : 4'b1100;
													assign node1455 = (inp[7]) ? node1463 : node1456;
														assign node1456 = (inp[8]) ? node1460 : node1457;
															assign node1457 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node1460 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node1463 = (inp[8]) ? node1467 : node1464;
															assign node1464 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node1467 = (inp[2]) ? 4'b0100 : 4'b0100;
												assign node1470 = (inp[13]) ? node1484 : node1471;
													assign node1471 = (inp[8]) ? node1477 : node1472;
														assign node1472 = (inp[7]) ? node1474 : 4'b1100;
															assign node1474 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node1477 = (inp[7]) ? node1481 : node1478;
															assign node1478 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node1481 = (inp[2]) ? 4'b0100 : 4'b0100;
													assign node1484 = (inp[14]) ? node1490 : node1485;
														assign node1485 = (inp[2]) ? node1487 : 4'b0101;
															assign node1487 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node1490 = (inp[2]) ? node1494 : node1491;
															assign node1491 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node1494 = (inp[7]) ? 4'b0100 : 4'b0100;
									assign node1497 = (inp[7]) ? node1601 : node1498;
										assign node1498 = (inp[8]) ? node1552 : node1499;
											assign node1499 = (inp[2]) ? node1529 : node1500;
												assign node1500 = (inp[14]) ? node1514 : node1501;
													assign node1501 = (inp[6]) ? node1509 : node1502;
														assign node1502 = (inp[11]) ? node1506 : node1503;
															assign node1503 = (inp[13]) ? 4'b0111 : 4'b1111;
															assign node1506 = (inp[1]) ? 4'b0111 : 4'b0111;
														assign node1509 = (inp[11]) ? node1511 : 4'b0111;
															assign node1511 = (inp[1]) ? 4'b0111 : 4'b1111;
													assign node1514 = (inp[13]) ? node1522 : node1515;
														assign node1515 = (inp[11]) ? node1519 : node1516;
															assign node1516 = (inp[6]) ? 4'b0110 : 4'b1110;
															assign node1519 = (inp[6]) ? 4'b1110 : 4'b0110;
														assign node1522 = (inp[1]) ? node1526 : node1523;
															assign node1523 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node1526 = (inp[11]) ? 4'b0110 : 4'b0110;
												assign node1529 = (inp[13]) ? node1537 : node1530;
													assign node1530 = (inp[11]) ? node1534 : node1531;
														assign node1531 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node1534 = (inp[6]) ? 4'b1110 : 4'b0110;
													assign node1537 = (inp[6]) ? node1545 : node1538;
														assign node1538 = (inp[14]) ? node1542 : node1539;
															assign node1539 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node1542 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node1545 = (inp[1]) ? node1549 : node1546;
															assign node1546 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node1549 = (inp[11]) ? 4'b0110 : 4'b1110;
											assign node1552 = (inp[2]) ? node1578 : node1553;
												assign node1553 = (inp[14]) ? node1565 : node1554;
													assign node1554 = (inp[6]) ? node1558 : node1555;
														assign node1555 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node1558 = (inp[11]) ? node1562 : node1559;
															assign node1559 = (inp[13]) ? 4'b0110 : 4'b0110;
															assign node1562 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node1565 = (inp[1]) ? node1571 : node1566;
														assign node1566 = (inp[13]) ? node1568 : 4'b0111;
															assign node1568 = (inp[6]) ? 4'b0111 : 4'b0111;
														assign node1571 = (inp[11]) ? node1575 : node1572;
															assign node1572 = (inp[6]) ? 4'b1111 : 4'b0111;
															assign node1575 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node1578 = (inp[6]) ? node1590 : node1579;
													assign node1579 = (inp[11]) ? node1585 : node1580;
														assign node1580 = (inp[13]) ? 4'b0111 : node1581;
															assign node1581 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node1585 = (inp[1]) ? 4'b1111 : node1586;
															assign node1586 = (inp[13]) ? 4'b1111 : 4'b0111;
													assign node1590 = (inp[11]) ? node1596 : node1591;
														assign node1591 = (inp[1]) ? 4'b1111 : node1592;
															assign node1592 = (inp[13]) ? 4'b1111 : 4'b0111;
														assign node1596 = (inp[1]) ? 4'b0111 : node1597;
															assign node1597 = (inp[13]) ? 4'b0111 : 4'b1111;
										assign node1601 = (inp[8]) ? node1655 : node1602;
											assign node1602 = (inp[14]) ? node1632 : node1603;
												assign node1603 = (inp[2]) ? node1617 : node1604;
													assign node1604 = (inp[11]) ? node1610 : node1605;
														assign node1605 = (inp[6]) ? node1607 : 4'b1110;
															assign node1607 = (inp[1]) ? 4'b1110 : 4'b0110;
														assign node1610 = (inp[6]) ? node1614 : node1611;
															assign node1611 = (inp[13]) ? 4'b1110 : 4'b0110;
															assign node1614 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node1617 = (inp[1]) ? node1625 : node1618;
														assign node1618 = (inp[11]) ? node1622 : node1619;
															assign node1619 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node1622 = (inp[13]) ? 4'b0111 : 4'b0111;
														assign node1625 = (inp[13]) ? node1629 : node1626;
															assign node1626 = (inp[11]) ? 4'b1111 : 4'b0111;
															assign node1629 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node1632 = (inp[11]) ? node1644 : node1633;
													assign node1633 = (inp[6]) ? node1639 : node1634;
														assign node1634 = (inp[13]) ? 4'b0111 : node1635;
															assign node1635 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node1639 = (inp[1]) ? 4'b1111 : node1640;
															assign node1640 = (inp[13]) ? 4'b1111 : 4'b0111;
													assign node1644 = (inp[6]) ? node1650 : node1645;
														assign node1645 = (inp[13]) ? 4'b1111 : node1646;
															assign node1646 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node1650 = (inp[1]) ? 4'b0111 : node1651;
															assign node1651 = (inp[13]) ? 4'b0111 : 4'b1111;
											assign node1655 = (inp[2]) ? node1687 : node1656;
												assign node1656 = (inp[14]) ? node1672 : node1657;
													assign node1657 = (inp[11]) ? node1665 : node1658;
														assign node1658 = (inp[6]) ? node1662 : node1659;
															assign node1659 = (inp[1]) ? 4'b0111 : 4'b1111;
															assign node1662 = (inp[13]) ? 4'b1111 : 4'b0111;
														assign node1665 = (inp[6]) ? node1669 : node1666;
															assign node1666 = (inp[13]) ? 4'b1111 : 4'b0111;
															assign node1669 = (inp[1]) ? 4'b0111 : 4'b0111;
													assign node1672 = (inp[1]) ? node1680 : node1673;
														assign node1673 = (inp[13]) ? node1677 : node1674;
															assign node1674 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node1677 = (inp[6]) ? 4'b0110 : 4'b0110;
														assign node1680 = (inp[13]) ? node1684 : node1681;
															assign node1681 = (inp[6]) ? 4'b0110 : 4'b1110;
															assign node1684 = (inp[11]) ? 4'b0110 : 4'b0110;
												assign node1687 = (inp[11]) ? node1699 : node1688;
													assign node1688 = (inp[6]) ? node1694 : node1689;
														assign node1689 = (inp[13]) ? 4'b0110 : node1690;
															assign node1690 = (inp[1]) ? 4'b0110 : 4'b1110;
														assign node1694 = (inp[1]) ? 4'b1110 : node1695;
															assign node1695 = (inp[13]) ? 4'b1110 : 4'b0110;
													assign node1699 = (inp[6]) ? node1705 : node1700;
														assign node1700 = (inp[1]) ? 4'b1110 : node1701;
															assign node1701 = (inp[13]) ? 4'b1110 : 4'b0110;
														assign node1705 = (inp[1]) ? 4'b0110 : node1706;
															assign node1706 = (inp[13]) ? 4'b0110 : 4'b1110;
						assign node1710 = (inp[0]) ? node2618 : node1711;
							assign node1711 = (inp[3]) ? node2137 : node1712;
								assign node1712 = (inp[13]) ? node1962 : node1713;
									assign node1713 = (inp[5]) ? node1837 : node1714;
										assign node1714 = (inp[2]) ? node1774 : node1715;
											assign node1715 = (inp[8]) ? node1745 : node1716;
												assign node1716 = (inp[7]) ? node1730 : node1717;
													assign node1717 = (inp[14]) ? node1725 : node1718;
														assign node1718 = (inp[11]) ? node1722 : node1719;
															assign node1719 = (inp[6]) ? 4'b0101 : 4'b1101;
															assign node1722 = (inp[6]) ? 4'b1101 : 4'b0101;
														assign node1725 = (inp[1]) ? 4'b1100 : node1726;
															assign node1726 = (inp[6]) ? 4'b0100 : 4'b0100;
													assign node1730 = (inp[14]) ? node1738 : node1731;
														assign node1731 = (inp[1]) ? node1735 : node1732;
															assign node1732 = (inp[11]) ? 4'b0100 : 4'b0100;
															assign node1735 = (inp[6]) ? 4'b0100 : 4'b0100;
														assign node1738 = (inp[6]) ? node1742 : node1739;
															assign node1739 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node1742 = (inp[11]) ? 4'b1101 : 4'b0101;
												assign node1745 = (inp[14]) ? node1761 : node1746;
													assign node1746 = (inp[7]) ? node1754 : node1747;
														assign node1747 = (inp[1]) ? node1751 : node1748;
															assign node1748 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node1751 = (inp[6]) ? 4'b0100 : 4'b0100;
														assign node1754 = (inp[6]) ? node1758 : node1755;
															assign node1755 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node1758 = (inp[11]) ? 4'b0101 : 4'b0101;
													assign node1761 = (inp[7]) ? node1769 : node1762;
														assign node1762 = (inp[1]) ? node1766 : node1763;
															assign node1763 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node1766 = (inp[11]) ? 4'b0101 : 4'b0101;
														assign node1769 = (inp[11]) ? 4'b1100 : node1770;
															assign node1770 = (inp[6]) ? 4'b0100 : 4'b0100;
											assign node1774 = (inp[6]) ? node1806 : node1775;
												assign node1775 = (inp[11]) ? node1791 : node1776;
													assign node1776 = (inp[1]) ? node1784 : node1777;
														assign node1777 = (inp[8]) ? node1781 : node1778;
															assign node1778 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node1781 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node1784 = (inp[8]) ? node1788 : node1785;
															assign node1785 = (inp[7]) ? 4'b0101 : 4'b1100;
															assign node1788 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node1791 = (inp[1]) ? node1799 : node1792;
														assign node1792 = (inp[8]) ? node1796 : node1793;
															assign node1793 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node1796 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node1799 = (inp[7]) ? node1803 : node1800;
															assign node1800 = (inp[8]) ? 4'b1101 : 4'b0100;
															assign node1803 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node1806 = (inp[11]) ? node1822 : node1807;
													assign node1807 = (inp[1]) ? node1815 : node1808;
														assign node1808 = (inp[8]) ? node1812 : node1809;
															assign node1809 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node1812 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node1815 = (inp[8]) ? node1819 : node1816;
															assign node1816 = (inp[7]) ? 4'b1101 : 4'b0100;
															assign node1819 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node1822 = (inp[1]) ? node1830 : node1823;
														assign node1823 = (inp[14]) ? node1827 : node1824;
															assign node1824 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node1827 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node1830 = (inp[7]) ? node1834 : node1831;
															assign node1831 = (inp[8]) ? 4'b0101 : 4'b1100;
															assign node1834 = (inp[8]) ? 4'b0100 : 4'b0101;
										assign node1837 = (inp[8]) ? node1899 : node1838;
											assign node1838 = (inp[7]) ? node1868 : node1839;
												assign node1839 = (inp[2]) ? node1855 : node1840;
													assign node1840 = (inp[14]) ? node1848 : node1841;
														assign node1841 = (inp[6]) ? node1845 : node1842;
															assign node1842 = (inp[11]) ? 4'b0101 : 4'b1101;
															assign node1845 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node1848 = (inp[11]) ? node1852 : node1849;
															assign node1849 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node1852 = (inp[6]) ? 4'b1100 : 4'b0100;
													assign node1855 = (inp[1]) ? node1863 : node1856;
														assign node1856 = (inp[11]) ? node1860 : node1857;
															assign node1857 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node1860 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node1863 = (inp[6]) ? node1865 : 4'b0100;
															assign node1865 = (inp[11]) ? 4'b1100 : 4'b0100;
												assign node1868 = (inp[2]) ? node1884 : node1869;
													assign node1869 = (inp[14]) ? node1877 : node1870;
														assign node1870 = (inp[1]) ? node1874 : node1871;
															assign node1871 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node1874 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node1877 = (inp[1]) ? node1881 : node1878;
															assign node1878 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node1881 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node1884 = (inp[6]) ? node1892 : node1885;
														assign node1885 = (inp[1]) ? node1889 : node1886;
															assign node1886 = (inp[11]) ? 4'b0101 : 4'b1101;
															assign node1889 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node1892 = (inp[14]) ? node1896 : node1893;
															assign node1893 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node1896 = (inp[11]) ? 4'b0101 : 4'b0101;
											assign node1899 = (inp[7]) ? node1931 : node1900;
												assign node1900 = (inp[2]) ? node1916 : node1901;
													assign node1901 = (inp[14]) ? node1909 : node1902;
														assign node1902 = (inp[11]) ? node1906 : node1903;
															assign node1903 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node1906 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node1909 = (inp[1]) ? node1913 : node1910;
															assign node1910 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node1913 = (inp[11]) ? 4'b0101 : 4'b0101;
													assign node1916 = (inp[1]) ? node1924 : node1917;
														assign node1917 = (inp[6]) ? node1921 : node1918;
															assign node1918 = (inp[11]) ? 4'b0101 : 4'b1101;
															assign node1921 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node1924 = (inp[14]) ? node1928 : node1925;
															assign node1925 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node1928 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node1931 = (inp[2]) ? node1947 : node1932;
													assign node1932 = (inp[14]) ? node1940 : node1933;
														assign node1933 = (inp[1]) ? node1937 : node1934;
															assign node1934 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node1937 = (inp[6]) ? 4'b0101 : 4'b0101;
														assign node1940 = (inp[1]) ? node1944 : node1941;
															assign node1941 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node1944 = (inp[6]) ? 4'b0100 : 4'b0100;
													assign node1947 = (inp[11]) ? node1955 : node1948;
														assign node1948 = (inp[14]) ? node1952 : node1949;
															assign node1949 = (inp[1]) ? 4'b0100 : 4'b0100;
															assign node1952 = (inp[6]) ? 4'b0100 : 4'b0100;
														assign node1955 = (inp[14]) ? node1959 : node1956;
															assign node1956 = (inp[1]) ? 4'b0100 : 4'b1100;
															assign node1959 = (inp[6]) ? 4'b1100 : 4'b0100;
									assign node1962 = (inp[7]) ? node2082 : node1963;
										assign node1963 = (inp[8]) ? node2027 : node1964;
											assign node1964 = (inp[14]) ? node1996 : node1965;
												assign node1965 = (inp[2]) ? node1981 : node1966;
													assign node1966 = (inp[5]) ? node1974 : node1967;
														assign node1967 = (inp[6]) ? node1971 : node1968;
															assign node1968 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node1971 = (inp[1]) ? 4'b0101 : 4'b0101;
														assign node1974 = (inp[6]) ? node1978 : node1975;
															assign node1975 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node1978 = (inp[1]) ? 4'b0101 : 4'b0101;
													assign node1981 = (inp[11]) ? node1989 : node1982;
														assign node1982 = (inp[5]) ? node1986 : node1983;
															assign node1983 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node1986 = (inp[1]) ? 4'b0100 : 4'b0100;
														assign node1989 = (inp[1]) ? node1993 : node1990;
															assign node1990 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node1993 = (inp[6]) ? 4'b0100 : 4'b1100;
												assign node1996 = (inp[2]) ? node2012 : node1997;
													assign node1997 = (inp[5]) ? node2005 : node1998;
														assign node1998 = (inp[1]) ? node2002 : node1999;
															assign node1999 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node2002 = (inp[6]) ? 4'b0100 : 4'b0100;
														assign node2005 = (inp[1]) ? node2009 : node2006;
															assign node2006 = (inp[11]) ? 4'b0100 : 4'b0100;
															assign node2009 = (inp[6]) ? 4'b0100 : 4'b0100;
													assign node2012 = (inp[11]) ? node2020 : node2013;
														assign node2013 = (inp[6]) ? node2017 : node2014;
															assign node2014 = (inp[1]) ? 4'b0100 : 4'b1100;
															assign node2017 = (inp[1]) ? 4'b1100 : 4'b0100;
														assign node2020 = (inp[1]) ? node2024 : node2021;
															assign node2021 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node2024 = (inp[6]) ? 4'b0100 : 4'b1100;
											assign node2027 = (inp[2]) ? node2059 : node2028;
												assign node2028 = (inp[14]) ? node2044 : node2029;
													assign node2029 = (inp[11]) ? node2037 : node2030;
														assign node2030 = (inp[1]) ? node2034 : node2031;
															assign node2031 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node2034 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node2037 = (inp[5]) ? node2041 : node2038;
															assign node2038 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node2041 = (inp[1]) ? 4'b0100 : 4'b0100;
													assign node2044 = (inp[5]) ? node2052 : node2045;
														assign node2045 = (inp[6]) ? node2049 : node2046;
															assign node2046 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node2049 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node2052 = (inp[1]) ? node2056 : node2053;
															assign node2053 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node2056 = (inp[11]) ? 4'b0101 : 4'b0101;
												assign node2059 = (inp[5]) ? node2067 : node2060;
													assign node2060 = (inp[11]) ? node2064 : node2061;
														assign node2061 = (inp[6]) ? 4'b1101 : 4'b0101;
														assign node2064 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node2067 = (inp[1]) ? node2075 : node2068;
														assign node2068 = (inp[14]) ? node2072 : node2069;
															assign node2069 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node2072 = (inp[6]) ? 4'b0101 : 4'b0101;
														assign node2075 = (inp[14]) ? node2079 : node2076;
															assign node2076 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node2079 = (inp[6]) ? 4'b0101 : 4'b0101;
										assign node2082 = (inp[8]) ? node2114 : node2083;
											assign node2083 = (inp[14]) ? node2107 : node2084;
												assign node2084 = (inp[2]) ? node2100 : node2085;
													assign node2085 = (inp[1]) ? node2093 : node2086;
														assign node2086 = (inp[5]) ? node2090 : node2087;
															assign node2087 = (inp[11]) ? 4'b0100 : 4'b0100;
															assign node2090 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node2093 = (inp[6]) ? node2097 : node2094;
															assign node2094 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node2097 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node2100 = (inp[6]) ? node2104 : node2101;
														assign node2101 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node2104 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node2107 = (inp[6]) ? node2111 : node2108;
													assign node2108 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node2111 = (inp[11]) ? 4'b0101 : 4'b1101;
											assign node2114 = (inp[2]) ? node2130 : node2115;
												assign node2115 = (inp[14]) ? node2123 : node2116;
													assign node2116 = (inp[6]) ? node2120 : node2117;
														assign node2117 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node2120 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node2123 = (inp[11]) ? node2127 : node2124;
														assign node2124 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node2127 = (inp[6]) ? 4'b0100 : 4'b1100;
												assign node2130 = (inp[6]) ? node2134 : node2131;
													assign node2131 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node2134 = (inp[11]) ? 4'b0100 : 4'b1100;
								assign node2137 = (inp[5]) ? node2375 : node2138;
									assign node2138 = (inp[11]) ? node2260 : node2139;
										assign node2139 = (inp[6]) ? node2201 : node2140;
											assign node2140 = (inp[1]) ? node2172 : node2141;
												assign node2141 = (inp[13]) ? node2157 : node2142;
													assign node2142 = (inp[8]) ? node2150 : node2143;
														assign node2143 = (inp[7]) ? node2147 : node2144;
															assign node2144 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node2147 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node2150 = (inp[7]) ? node2154 : node2151;
															assign node2151 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node2154 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node2157 = (inp[7]) ? node2165 : node2158;
														assign node2158 = (inp[8]) ? node2162 : node2159;
															assign node2159 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node2162 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node2165 = (inp[8]) ? node2169 : node2166;
															assign node2166 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node2169 = (inp[2]) ? 4'b0100 : 4'b0100;
												assign node2172 = (inp[13]) ? node2188 : node2173;
													assign node2173 = (inp[8]) ? node2181 : node2174;
														assign node2174 = (inp[7]) ? node2178 : node2175;
															assign node2175 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node2178 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node2181 = (inp[7]) ? node2185 : node2182;
															assign node2182 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node2185 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node2188 = (inp[7]) ? node2196 : node2189;
														assign node2189 = (inp[8]) ? node2193 : node2190;
															assign node2190 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node2193 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node2196 = (inp[14]) ? 4'b0100 : node2197;
															assign node2197 = (inp[8]) ? 4'b0100 : 4'b0100;
											assign node2201 = (inp[13]) ? node2233 : node2202;
												assign node2202 = (inp[1]) ? node2218 : node2203;
													assign node2203 = (inp[2]) ? node2211 : node2204;
														assign node2204 = (inp[7]) ? node2208 : node2205;
															assign node2205 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node2208 = (inp[14]) ? 4'b0100 : 4'b0100;
														assign node2211 = (inp[8]) ? node2215 : node2212;
															assign node2212 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node2215 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node2218 = (inp[8]) ? node2226 : node2219;
														assign node2219 = (inp[7]) ? node2223 : node2220;
															assign node2220 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node2223 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node2226 = (inp[7]) ? node2230 : node2227;
															assign node2227 = (inp[14]) ? 4'b1101 : 4'b0100;
															assign node2230 = (inp[14]) ? 4'b1100 : 4'b1100;
												assign node2233 = (inp[1]) ? node2247 : node2234;
													assign node2234 = (inp[7]) ? node2242 : node2235;
														assign node2235 = (inp[8]) ? node2239 : node2236;
															assign node2236 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node2239 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node2242 = (inp[8]) ? node2244 : 4'b1101;
															assign node2244 = (inp[14]) ? 4'b1100 : 4'b1100;
													assign node2247 = (inp[7]) ? node2255 : node2248;
														assign node2248 = (inp[8]) ? node2252 : node2249;
															assign node2249 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node2252 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node2255 = (inp[8]) ? 4'b1100 : node2256;
															assign node2256 = (inp[14]) ? 4'b1101 : 4'b1100;
										assign node2260 = (inp[6]) ? node2320 : node2261;
											assign node2261 = (inp[1]) ? node2291 : node2262;
												assign node2262 = (inp[13]) ? node2278 : node2263;
													assign node2263 = (inp[14]) ? node2271 : node2264;
														assign node2264 = (inp[7]) ? node2268 : node2265;
															assign node2265 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node2268 = (inp[2]) ? 4'b0100 : 4'b0100;
														assign node2271 = (inp[7]) ? node2275 : node2272;
															assign node2272 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node2275 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node2278 = (inp[8]) ? node2286 : node2279;
														assign node2279 = (inp[7]) ? node2283 : node2280;
															assign node2280 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node2283 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node2286 = (inp[14]) ? 4'b1101 : node2287;
															assign node2287 = (inp[2]) ? 4'b1100 : 4'b0100;
												assign node2291 = (inp[13]) ? node2307 : node2292;
													assign node2292 = (inp[8]) ? node2300 : node2293;
														assign node2293 = (inp[7]) ? node2297 : node2294;
															assign node2294 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node2297 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node2300 = (inp[7]) ? node2304 : node2301;
															assign node2301 = (inp[2]) ? 4'b1101 : 4'b0100;
															assign node2304 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node2307 = (inp[2]) ? node2313 : node2308;
														assign node2308 = (inp[7]) ? node2310 : 4'b1101;
															assign node2310 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node2313 = (inp[8]) ? node2317 : node2314;
															assign node2314 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node2317 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node2320 = (inp[1]) ? node2348 : node2321;
												assign node2321 = (inp[13]) ? node2333 : node2322;
													assign node2322 = (inp[8]) ? node2328 : node2323;
														assign node2323 = (inp[7]) ? node2325 : 4'b1100;
															assign node2325 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node2328 = (inp[7]) ? node2330 : 4'b1101;
															assign node2330 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node2333 = (inp[8]) ? node2341 : node2334;
														assign node2334 = (inp[7]) ? node2338 : node2335;
															assign node2335 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node2338 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node2341 = (inp[7]) ? node2345 : node2342;
															assign node2342 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node2345 = (inp[2]) ? 4'b0100 : 4'b0100;
												assign node2348 = (inp[13]) ? node2362 : node2349;
													assign node2349 = (inp[7]) ? node2357 : node2350;
														assign node2350 = (inp[8]) ? node2354 : node2351;
															assign node2351 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node2354 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node2357 = (inp[8]) ? node2359 : 4'b0101;
															assign node2359 = (inp[2]) ? 4'b0100 : 4'b0100;
													assign node2362 = (inp[2]) ? node2370 : node2363;
														assign node2363 = (inp[7]) ? node2367 : node2364;
															assign node2364 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node2367 = (inp[14]) ? 4'b0100 : 4'b0100;
														assign node2370 = (inp[14]) ? node2372 : 4'b0101;
															assign node2372 = (inp[7]) ? 4'b0100 : 4'b0100;
									assign node2375 = (inp[2]) ? node2497 : node2376;
										assign node2376 = (inp[7]) ? node2438 : node2377;
											assign node2377 = (inp[8]) ? node2407 : node2378;
												assign node2378 = (inp[14]) ? node2392 : node2379;
													assign node2379 = (inp[1]) ? node2385 : node2380;
														assign node2380 = (inp[6]) ? 4'b1111 : node2381;
															assign node2381 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node2385 = (inp[13]) ? node2389 : node2386;
															assign node2386 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node2389 = (inp[11]) ? 4'b0111 : 4'b0111;
													assign node2392 = (inp[1]) ? node2400 : node2393;
														assign node2393 = (inp[11]) ? node2397 : node2394;
															assign node2394 = (inp[6]) ? 4'b0110 : 4'b1110;
															assign node2397 = (inp[6]) ? 4'b1110 : 4'b0110;
														assign node2400 = (inp[11]) ? node2404 : node2401;
															assign node2401 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node2404 = (inp[6]) ? 4'b1110 : 4'b0110;
												assign node2407 = (inp[14]) ? node2423 : node2408;
													assign node2408 = (inp[11]) ? node2416 : node2409;
														assign node2409 = (inp[6]) ? node2413 : node2410;
															assign node2410 = (inp[13]) ? 4'b0110 : 4'b1110;
															assign node2413 = (inp[13]) ? 4'b0110 : 4'b0110;
														assign node2416 = (inp[6]) ? node2420 : node2417;
															assign node2417 = (inp[1]) ? 4'b1110 : 4'b0110;
															assign node2420 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node2423 = (inp[11]) ? node2431 : node2424;
														assign node2424 = (inp[6]) ? node2428 : node2425;
															assign node2425 = (inp[1]) ? 4'b0111 : 4'b0111;
															assign node2428 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node2431 = (inp[6]) ? node2435 : node2432;
															assign node2432 = (inp[1]) ? 4'b1111 : 4'b0111;
															assign node2435 = (inp[1]) ? 4'b0111 : 4'b0111;
											assign node2438 = (inp[11]) ? node2468 : node2439;
												assign node2439 = (inp[1]) ? node2455 : node2440;
													assign node2440 = (inp[6]) ? node2448 : node2441;
														assign node2441 = (inp[13]) ? node2445 : node2442;
															assign node2442 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node2445 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node2448 = (inp[13]) ? node2452 : node2449;
															assign node2449 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node2452 = (inp[14]) ? 4'b1110 : 4'b0110;
													assign node2455 = (inp[6]) ? node2463 : node2456;
														assign node2456 = (inp[8]) ? node2460 : node2457;
															assign node2457 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node2460 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node2463 = (inp[14]) ? node2465 : 4'b0110;
															assign node2465 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node2468 = (inp[6]) ? node2484 : node2469;
													assign node2469 = (inp[13]) ? node2477 : node2470;
														assign node2470 = (inp[1]) ? node2474 : node2471;
															assign node2471 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node2474 = (inp[14]) ? 4'b1111 : 4'b0110;
														assign node2477 = (inp[14]) ? node2481 : node2478;
															assign node2478 = (inp[8]) ? 4'b1111 : 4'b0110;
															assign node2481 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node2484 = (inp[13]) ? node2492 : node2485;
														assign node2485 = (inp[1]) ? node2489 : node2486;
															assign node2486 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node2489 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node2492 = (inp[8]) ? node2494 : 4'b0111;
															assign node2494 = (inp[14]) ? 4'b0110 : 4'b0111;
										assign node2497 = (inp[14]) ? node2559 : node2498;
											assign node2498 = (inp[6]) ? node2530 : node2499;
												assign node2499 = (inp[11]) ? node2515 : node2500;
													assign node2500 = (inp[1]) ? node2508 : node2501;
														assign node2501 = (inp[13]) ? node2505 : node2502;
															assign node2502 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node2505 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node2508 = (inp[7]) ? node2512 : node2509;
															assign node2509 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node2512 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node2515 = (inp[1]) ? node2523 : node2516;
														assign node2516 = (inp[13]) ? node2520 : node2517;
															assign node2517 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node2520 = (inp[7]) ? 4'b1111 : 4'b0110;
														assign node2523 = (inp[8]) ? node2527 : node2524;
															assign node2524 = (inp[7]) ? 4'b1111 : 4'b0110;
															assign node2527 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node2530 = (inp[11]) ? node2546 : node2531;
													assign node2531 = (inp[1]) ? node2539 : node2532;
														assign node2532 = (inp[13]) ? node2536 : node2533;
															assign node2533 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node2536 = (inp[7]) ? 4'b1110 : 4'b0110;
														assign node2539 = (inp[7]) ? node2543 : node2540;
															assign node2540 = (inp[8]) ? 4'b1111 : 4'b0110;
															assign node2543 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node2546 = (inp[1]) ? node2552 : node2547;
														assign node2547 = (inp[13]) ? node2549 : 4'b1111;
															assign node2549 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node2552 = (inp[13]) ? node2556 : node2553;
															assign node2553 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node2556 = (inp[8]) ? 4'b0110 : 4'b0110;
											assign node2559 = (inp[7]) ? node2589 : node2560;
												assign node2560 = (inp[8]) ? node2574 : node2561;
													assign node2561 = (inp[11]) ? node2567 : node2562;
														assign node2562 = (inp[6]) ? node2564 : 4'b1110;
															assign node2564 = (inp[1]) ? 4'b1110 : 4'b0110;
														assign node2567 = (inp[6]) ? node2571 : node2568;
															assign node2568 = (inp[1]) ? 4'b0110 : 4'b0110;
															assign node2571 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node2574 = (inp[11]) ? node2582 : node2575;
														assign node2575 = (inp[6]) ? node2579 : node2576;
															assign node2576 = (inp[1]) ? 4'b0111 : 4'b0111;
															assign node2579 = (inp[13]) ? 4'b1111 : 4'b0111;
														assign node2582 = (inp[6]) ? node2586 : node2583;
															assign node2583 = (inp[1]) ? 4'b1111 : 4'b0111;
															assign node2586 = (inp[1]) ? 4'b0111 : 4'b0111;
												assign node2589 = (inp[8]) ? node2605 : node2590;
													assign node2590 = (inp[13]) ? node2598 : node2591;
														assign node2591 = (inp[1]) ? node2595 : node2592;
															assign node2592 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node2595 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node2598 = (inp[1]) ? node2602 : node2599;
															assign node2599 = (inp[6]) ? 4'b1111 : 4'b0111;
															assign node2602 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node2605 = (inp[11]) ? node2611 : node2606;
														assign node2606 = (inp[6]) ? 4'b1110 : node2607;
															assign node2607 = (inp[1]) ? 4'b0110 : 4'b1110;
														assign node2611 = (inp[6]) ? node2615 : node2612;
															assign node2612 = (inp[1]) ? 4'b1110 : 4'b0110;
															assign node2615 = (inp[1]) ? 4'b0110 : 4'b0110;
							assign node2618 = (inp[3]) ? node3030 : node2619;
								assign node2619 = (inp[11]) ? node2825 : node2620;
									assign node2620 = (inp[6]) ? node2732 : node2621;
										assign node2621 = (inp[1]) ? node2677 : node2622;
											assign node2622 = (inp[13]) ? node2654 : node2623;
												assign node2623 = (inp[5]) ? node2639 : node2624;
													assign node2624 = (inp[8]) ? node2632 : node2625;
														assign node2625 = (inp[7]) ? node2629 : node2626;
															assign node2626 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node2629 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node2632 = (inp[7]) ? node2636 : node2633;
															assign node2633 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node2636 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node2639 = (inp[8]) ? node2647 : node2640;
														assign node2640 = (inp[7]) ? node2644 : node2641;
															assign node2641 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node2644 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node2647 = (inp[7]) ? node2651 : node2648;
															assign node2648 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node2651 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node2654 = (inp[7]) ? node2666 : node2655;
													assign node2655 = (inp[8]) ? node2661 : node2656;
														assign node2656 = (inp[14]) ? 4'b1110 : node2657;
															assign node2657 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node2661 = (inp[14]) ? 4'b0111 : node2662;
															assign node2662 = (inp[2]) ? 4'b0111 : 4'b1110;
													assign node2666 = (inp[8]) ? node2672 : node2667;
														assign node2667 = (inp[2]) ? 4'b0111 : node2668;
															assign node2668 = (inp[14]) ? 4'b0111 : 4'b1110;
														assign node2672 = (inp[2]) ? 4'b0110 : node2673;
															assign node2673 = (inp[14]) ? 4'b0110 : 4'b0111;
											assign node2677 = (inp[13]) ? node2701 : node2678;
												assign node2678 = (inp[8]) ? node2690 : node2679;
													assign node2679 = (inp[7]) ? node2685 : node2680;
														assign node2680 = (inp[14]) ? 4'b1110 : node2681;
															assign node2681 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node2685 = (inp[2]) ? 4'b0111 : node2686;
															assign node2686 = (inp[14]) ? 4'b0111 : 4'b1110;
													assign node2690 = (inp[7]) ? node2696 : node2691;
														assign node2691 = (inp[14]) ? 4'b0111 : node2692;
															assign node2692 = (inp[2]) ? 4'b0111 : 4'b1110;
														assign node2696 = (inp[14]) ? 4'b0110 : node2697;
															assign node2697 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node2701 = (inp[14]) ? node2717 : node2702;
													assign node2702 = (inp[5]) ? node2710 : node2703;
														assign node2703 = (inp[7]) ? node2707 : node2704;
															assign node2704 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node2707 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node2710 = (inp[2]) ? node2714 : node2711;
															assign node2711 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node2714 = (inp[8]) ? 4'b0110 : 4'b0110;
													assign node2717 = (inp[5]) ? node2725 : node2718;
														assign node2718 = (inp[7]) ? node2722 : node2719;
															assign node2719 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node2722 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node2725 = (inp[7]) ? node2729 : node2726;
															assign node2726 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node2729 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node2732 = (inp[13]) ? node2778 : node2733;
											assign node2733 = (inp[1]) ? node2755 : node2734;
												assign node2734 = (inp[8]) ? node2744 : node2735;
													assign node2735 = (inp[2]) ? 4'b0110 : node2736;
														assign node2736 = (inp[7]) ? node2740 : node2737;
															assign node2737 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node2740 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node2744 = (inp[7]) ? node2750 : node2745;
														assign node2745 = (inp[14]) ? 4'b0111 : node2746;
															assign node2746 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node2750 = (inp[2]) ? 4'b0110 : node2751;
															assign node2751 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node2755 = (inp[7]) ? node2767 : node2756;
													assign node2756 = (inp[8]) ? node2762 : node2757;
														assign node2757 = (inp[2]) ? 4'b0110 : node2758;
															assign node2758 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node2762 = (inp[14]) ? 4'b1111 : node2763;
															assign node2763 = (inp[2]) ? 4'b1111 : 4'b0110;
													assign node2767 = (inp[8]) ? node2773 : node2768;
														assign node2768 = (inp[14]) ? 4'b1111 : node2769;
															assign node2769 = (inp[2]) ? 4'b1111 : 4'b0110;
														assign node2773 = (inp[14]) ? 4'b1110 : node2774;
															assign node2774 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node2778 = (inp[1]) ? node2802 : node2779;
												assign node2779 = (inp[7]) ? node2791 : node2780;
													assign node2780 = (inp[8]) ? node2786 : node2781;
														assign node2781 = (inp[14]) ? 4'b0110 : node2782;
															assign node2782 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node2786 = (inp[14]) ? 4'b1111 : node2787;
															assign node2787 = (inp[2]) ? 4'b1111 : 4'b0110;
													assign node2791 = (inp[8]) ? node2797 : node2792;
														assign node2792 = (inp[2]) ? 4'b1111 : node2793;
															assign node2793 = (inp[14]) ? 4'b1111 : 4'b0110;
														assign node2797 = (inp[14]) ? 4'b1110 : node2798;
															assign node2798 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node2802 = (inp[8]) ? node2814 : node2803;
													assign node2803 = (inp[7]) ? node2809 : node2804;
														assign node2804 = (inp[14]) ? 4'b1110 : node2805;
															assign node2805 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node2809 = (inp[2]) ? 4'b1111 : node2810;
															assign node2810 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node2814 = (inp[7]) ? node2820 : node2815;
														assign node2815 = (inp[5]) ? 4'b1111 : node2816;
															assign node2816 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node2820 = (inp[2]) ? 4'b1110 : node2821;
															assign node2821 = (inp[14]) ? 4'b1110 : 4'b1111;
									assign node2825 = (inp[6]) ? node2931 : node2826;
										assign node2826 = (inp[13]) ? node2882 : node2827;
											assign node2827 = (inp[1]) ? node2859 : node2828;
												assign node2828 = (inp[14]) ? node2844 : node2829;
													assign node2829 = (inp[8]) ? node2837 : node2830;
														assign node2830 = (inp[2]) ? node2834 : node2831;
															assign node2831 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node2834 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node2837 = (inp[7]) ? node2841 : node2838;
															assign node2838 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node2841 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node2844 = (inp[5]) ? node2852 : node2845;
														assign node2845 = (inp[8]) ? node2849 : node2846;
															assign node2846 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node2849 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node2852 = (inp[7]) ? node2856 : node2853;
															assign node2853 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node2856 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node2859 = (inp[8]) ? node2871 : node2860;
													assign node2860 = (inp[7]) ? node2866 : node2861;
														assign node2861 = (inp[14]) ? 4'b0110 : node2862;
															assign node2862 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node2866 = (inp[2]) ? 4'b1111 : node2867;
															assign node2867 = (inp[14]) ? 4'b1111 : 4'b0110;
													assign node2871 = (inp[7]) ? node2877 : node2872;
														assign node2872 = (inp[2]) ? 4'b1111 : node2873;
															assign node2873 = (inp[14]) ? 4'b1111 : 4'b0110;
														assign node2877 = (inp[2]) ? 4'b1110 : node2878;
															assign node2878 = (inp[14]) ? 4'b1110 : 4'b1111;
											assign node2882 = (inp[1]) ? node2906 : node2883;
												assign node2883 = (inp[8]) ? node2895 : node2884;
													assign node2884 = (inp[7]) ? node2890 : node2885;
														assign node2885 = (inp[2]) ? 4'b0110 : node2886;
															assign node2886 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node2890 = (inp[2]) ? 4'b1111 : node2891;
															assign node2891 = (inp[14]) ? 4'b1111 : 4'b0110;
													assign node2895 = (inp[7]) ? node2901 : node2896;
														assign node2896 = (inp[2]) ? 4'b1111 : node2897;
															assign node2897 = (inp[14]) ? 4'b1111 : 4'b0110;
														assign node2901 = (inp[2]) ? 4'b1110 : node2902;
															assign node2902 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node2906 = (inp[2]) ? node2920 : node2907;
													assign node2907 = (inp[8]) ? node2915 : node2908;
														assign node2908 = (inp[5]) ? node2912 : node2909;
															assign node2909 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node2912 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node2915 = (inp[5]) ? 4'b1110 : node2916;
															assign node2916 = (inp[7]) ? 4'b1110 : 4'b1110;
													assign node2920 = (inp[14]) ? node2926 : node2921;
														assign node2921 = (inp[8]) ? 4'b1111 : node2922;
															assign node2922 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node2926 = (inp[7]) ? node2928 : 4'b1111;
															assign node2928 = (inp[8]) ? 4'b1110 : 4'b1111;
										assign node2931 = (inp[13]) ? node2975 : node2932;
											assign node2932 = (inp[1]) ? node2952 : node2933;
												assign node2933 = (inp[7]) ? node2941 : node2934;
													assign node2934 = (inp[8]) ? 4'b1111 : node2935;
														assign node2935 = (inp[2]) ? 4'b1110 : node2936;
															assign node2936 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node2941 = (inp[8]) ? node2947 : node2942;
														assign node2942 = (inp[2]) ? 4'b1111 : node2943;
															assign node2943 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node2947 = (inp[14]) ? 4'b1110 : node2948;
															assign node2948 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node2952 = (inp[7]) ? node2964 : node2953;
													assign node2953 = (inp[8]) ? node2959 : node2954;
														assign node2954 = (inp[14]) ? 4'b1110 : node2955;
															assign node2955 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node2959 = (inp[2]) ? 4'b0111 : node2960;
															assign node2960 = (inp[14]) ? 4'b0111 : 4'b1110;
													assign node2964 = (inp[8]) ? node2970 : node2965;
														assign node2965 = (inp[14]) ? 4'b0111 : node2966;
															assign node2966 = (inp[2]) ? 4'b0111 : 4'b1110;
														assign node2970 = (inp[2]) ? 4'b0110 : node2971;
															assign node2971 = (inp[14]) ? 4'b0110 : 4'b0111;
											assign node2975 = (inp[1]) ? node2999 : node2976;
												assign node2976 = (inp[7]) ? node2988 : node2977;
													assign node2977 = (inp[8]) ? node2983 : node2978;
														assign node2978 = (inp[14]) ? 4'b1110 : node2979;
															assign node2979 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node2983 = (inp[14]) ? 4'b0111 : node2984;
															assign node2984 = (inp[2]) ? 4'b0111 : 4'b1110;
													assign node2988 = (inp[8]) ? node2994 : node2989;
														assign node2989 = (inp[2]) ? 4'b0111 : node2990;
															assign node2990 = (inp[14]) ? 4'b0111 : 4'b1110;
														assign node2994 = (inp[2]) ? 4'b0110 : node2995;
															assign node2995 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node2999 = (inp[5]) ? node3015 : node3000;
													assign node3000 = (inp[14]) ? node3008 : node3001;
														assign node3001 = (inp[7]) ? node3005 : node3002;
															assign node3002 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node3005 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node3008 = (inp[7]) ? node3012 : node3009;
															assign node3009 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node3012 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node3015 = (inp[8]) ? node3023 : node3016;
														assign node3016 = (inp[7]) ? node3020 : node3017;
															assign node3017 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node3020 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node3023 = (inp[7]) ? node3027 : node3024;
															assign node3024 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node3027 = (inp[2]) ? 4'b0110 : 4'b0110;
								assign node3030 = (inp[5]) ? node3270 : node3031;
									assign node3031 = (inp[13]) ? node3157 : node3032;
										assign node3032 = (inp[14]) ? node3096 : node3033;
											assign node3033 = (inp[8]) ? node3065 : node3034;
												assign node3034 = (inp[6]) ? node3050 : node3035;
													assign node3035 = (inp[11]) ? node3043 : node3036;
														assign node3036 = (inp[1]) ? node3040 : node3037;
															assign node3037 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node3040 = (inp[2]) ? 4'b0110 : 4'b1110;
														assign node3043 = (inp[2]) ? node3047 : node3044;
															assign node3044 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node3047 = (inp[7]) ? 4'b1111 : 4'b0110;
													assign node3050 = (inp[11]) ? node3058 : node3051;
														assign node3051 = (inp[2]) ? node3055 : node3052;
															assign node3052 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node3055 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node3058 = (inp[1]) ? node3062 : node3059;
															assign node3059 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node3062 = (inp[2]) ? 4'b0111 : 4'b1110;
												assign node3065 = (inp[11]) ? node3081 : node3066;
													assign node3066 = (inp[6]) ? node3074 : node3067;
														assign node3067 = (inp[1]) ? node3071 : node3068;
															assign node3068 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node3071 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node3074 = (inp[1]) ? node3078 : node3075;
															assign node3075 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node3078 = (inp[2]) ? 4'b1110 : 4'b0110;
													assign node3081 = (inp[6]) ? node3089 : node3082;
														assign node3082 = (inp[1]) ? node3086 : node3083;
															assign node3083 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node3086 = (inp[7]) ? 4'b1110 : 4'b0110;
														assign node3089 = (inp[1]) ? node3093 : node3090;
															assign node3090 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node3093 = (inp[2]) ? 4'b0110 : 4'b0110;
											assign node3096 = (inp[2]) ? node3126 : node3097;
												assign node3097 = (inp[11]) ? node3111 : node3098;
													assign node3098 = (inp[6]) ? node3106 : node3099;
														assign node3099 = (inp[1]) ? node3103 : node3100;
															assign node3100 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node3103 = (inp[7]) ? 4'b0110 : 4'b1110;
														assign node3106 = (inp[1]) ? node3108 : 4'b0110;
															assign node3108 = (inp[7]) ? 4'b1110 : 4'b0110;
													assign node3111 = (inp[6]) ? node3119 : node3112;
														assign node3112 = (inp[1]) ? node3116 : node3113;
															assign node3113 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node3116 = (inp[8]) ? 4'b1110 : 4'b0110;
														assign node3119 = (inp[1]) ? node3123 : node3120;
															assign node3120 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node3123 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node3126 = (inp[8]) ? node3142 : node3127;
													assign node3127 = (inp[7]) ? node3135 : node3128;
														assign node3128 = (inp[1]) ? node3132 : node3129;
															assign node3129 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node3132 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node3135 = (inp[11]) ? node3139 : node3136;
															assign node3136 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node3139 = (inp[6]) ? 4'b0111 : 4'b0111;
													assign node3142 = (inp[7]) ? node3150 : node3143;
														assign node3143 = (inp[11]) ? node3147 : node3144;
															assign node3144 = (inp[1]) ? 4'b1111 : 4'b0111;
															assign node3147 = (inp[1]) ? 4'b0111 : 4'b0111;
														assign node3150 = (inp[1]) ? node3154 : node3151;
															assign node3151 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node3154 = (inp[11]) ? 4'b0110 : 4'b0110;
										assign node3157 = (inp[11]) ? node3211 : node3158;
											assign node3158 = (inp[6]) ? node3184 : node3159;
												assign node3159 = (inp[1]) ? node3171 : node3160;
													assign node3160 = (inp[8]) ? node3166 : node3161;
														assign node3161 = (inp[2]) ? 4'b1110 : node3162;
															assign node3162 = (inp[14]) ? 4'b0110 : 4'b1110;
														assign node3166 = (inp[14]) ? 4'b0111 : node3167;
															assign node3167 = (inp[2]) ? 4'b0110 : 4'b0110;
													assign node3171 = (inp[14]) ? node3177 : node3172;
														assign node3172 = (inp[8]) ? node3174 : 4'b0111;
															assign node3174 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node3177 = (inp[2]) ? node3181 : node3178;
															assign node3178 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node3181 = (inp[8]) ? 4'b0110 : 4'b0110;
												assign node3184 = (inp[1]) ? node3198 : node3185;
													assign node3185 = (inp[7]) ? node3193 : node3186;
														assign node3186 = (inp[8]) ? node3190 : node3187;
															assign node3187 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node3190 = (inp[2]) ? 4'b1111 : 4'b0110;
														assign node3193 = (inp[8]) ? node3195 : 4'b1111;
															assign node3195 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node3198 = (inp[14]) ? node3206 : node3199;
														assign node3199 = (inp[8]) ? node3203 : node3200;
															assign node3200 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node3203 = (inp[2]) ? 4'b1110 : 4'b1110;
														assign node3206 = (inp[7]) ? 4'b1111 : node3207;
															assign node3207 = (inp[8]) ? 4'b1111 : 4'b1110;
											assign node3211 = (inp[6]) ? node3243 : node3212;
												assign node3212 = (inp[1]) ? node3228 : node3213;
													assign node3213 = (inp[7]) ? node3221 : node3214;
														assign node3214 = (inp[8]) ? node3218 : node3215;
															assign node3215 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node3218 = (inp[2]) ? 4'b1111 : 4'b0110;
														assign node3221 = (inp[8]) ? node3225 : node3222;
															assign node3222 = (inp[14]) ? 4'b1111 : 4'b0110;
															assign node3225 = (inp[2]) ? 4'b1110 : 4'b1110;
													assign node3228 = (inp[8]) ? node3236 : node3229;
														assign node3229 = (inp[7]) ? node3233 : node3230;
															assign node3230 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node3233 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node3236 = (inp[7]) ? node3240 : node3237;
															assign node3237 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node3240 = (inp[14]) ? 4'b1110 : 4'b1110;
												assign node3243 = (inp[1]) ? node3257 : node3244;
													assign node3244 = (inp[7]) ? node3250 : node3245;
														assign node3245 = (inp[8]) ? node3247 : 4'b1110;
															assign node3247 = (inp[2]) ? 4'b0111 : 4'b1110;
														assign node3250 = (inp[8]) ? node3254 : node3251;
															assign node3251 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node3254 = (inp[2]) ? 4'b0110 : 4'b0110;
													assign node3257 = (inp[14]) ? node3263 : node3258;
														assign node3258 = (inp[7]) ? 4'b0110 : node3259;
															assign node3259 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node3263 = (inp[8]) ? node3267 : node3264;
															assign node3264 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node3267 = (inp[7]) ? 4'b0110 : 4'b0111;
									assign node3270 = (inp[6]) ? node3388 : node3271;
										assign node3271 = (inp[11]) ? node3331 : node3272;
											assign node3272 = (inp[13]) ? node3302 : node3273;
												assign node3273 = (inp[1]) ? node3287 : node3274;
													assign node3274 = (inp[8]) ? node3282 : node3275;
														assign node3275 = (inp[7]) ? node3279 : node3276;
															assign node3276 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node3279 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node3282 = (inp[7]) ? node3284 : 4'b1101;
															assign node3284 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node3287 = (inp[8]) ? node3295 : node3288;
														assign node3288 = (inp[7]) ? node3292 : node3289;
															assign node3289 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node3292 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node3295 = (inp[7]) ? node3299 : node3296;
															assign node3296 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node3299 = (inp[14]) ? 4'b0100 : 4'b0100;
												assign node3302 = (inp[1]) ? node3318 : node3303;
													assign node3303 = (inp[7]) ? node3311 : node3304;
														assign node3304 = (inp[8]) ? node3308 : node3305;
															assign node3305 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node3308 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node3311 = (inp[8]) ? node3315 : node3312;
															assign node3312 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node3315 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node3318 = (inp[2]) ? node3324 : node3319;
														assign node3319 = (inp[14]) ? node3321 : 4'b0100;
															assign node3321 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node3324 = (inp[14]) ? node3328 : node3325;
															assign node3325 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node3328 = (inp[8]) ? 4'b0100 : 4'b0100;
											assign node3331 = (inp[13]) ? node3357 : node3332;
												assign node3332 = (inp[1]) ? node3344 : node3333;
													assign node3333 = (inp[7]) ? node3341 : node3334;
														assign node3334 = (inp[8]) ? node3338 : node3335;
															assign node3335 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node3338 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node3341 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node3344 = (inp[8]) ? node3352 : node3345;
														assign node3345 = (inp[7]) ? node3349 : node3346;
															assign node3346 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node3349 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node3352 = (inp[14]) ? 4'b1101 : node3353;
															assign node3353 = (inp[2]) ? 4'b1100 : 4'b0100;
												assign node3357 = (inp[1]) ? node3373 : node3358;
													assign node3358 = (inp[8]) ? node3366 : node3359;
														assign node3359 = (inp[7]) ? node3363 : node3360;
															assign node3360 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node3363 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node3366 = (inp[7]) ? node3370 : node3367;
															assign node3367 = (inp[2]) ? 4'b1101 : 4'b0100;
															assign node3370 = (inp[14]) ? 4'b1100 : 4'b1100;
													assign node3373 = (inp[14]) ? node3381 : node3374;
														assign node3374 = (inp[8]) ? node3378 : node3375;
															assign node3375 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node3378 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node3381 = (inp[8]) ? node3385 : node3382;
															assign node3382 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node3385 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node3388 = (inp[11]) ? node3450 : node3389;
											assign node3389 = (inp[13]) ? node3421 : node3390;
												assign node3390 = (inp[1]) ? node3406 : node3391;
													assign node3391 = (inp[7]) ? node3399 : node3392;
														assign node3392 = (inp[8]) ? node3396 : node3393;
															assign node3393 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node3396 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node3399 = (inp[8]) ? node3403 : node3400;
															assign node3400 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node3403 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node3406 = (inp[8]) ? node3414 : node3407;
														assign node3407 = (inp[7]) ? node3411 : node3408;
															assign node3408 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node3411 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node3414 = (inp[7]) ? node3418 : node3415;
															assign node3415 = (inp[2]) ? 4'b1101 : 4'b0100;
															assign node3418 = (inp[14]) ? 4'b1100 : 4'b1100;
												assign node3421 = (inp[1]) ? node3435 : node3422;
													assign node3422 = (inp[7]) ? node3428 : node3423;
														assign node3423 = (inp[8]) ? node3425 : 4'b0100;
															assign node3425 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node3428 = (inp[8]) ? node3432 : node3429;
															assign node3429 = (inp[14]) ? 4'b1101 : 4'b0100;
															assign node3432 = (inp[2]) ? 4'b1100 : 4'b1100;
													assign node3435 = (inp[2]) ? node3443 : node3436;
														assign node3436 = (inp[7]) ? node3440 : node3437;
															assign node3437 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node3440 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node3443 = (inp[14]) ? node3447 : node3444;
															assign node3444 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node3447 = (inp[8]) ? 4'b1100 : 4'b1100;
											assign node3450 = (inp[1]) ? node3482 : node3451;
												assign node3451 = (inp[13]) ? node3467 : node3452;
													assign node3452 = (inp[7]) ? node3460 : node3453;
														assign node3453 = (inp[8]) ? node3457 : node3454;
															assign node3454 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node3457 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node3460 = (inp[8]) ? node3464 : node3461;
															assign node3461 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node3464 = (inp[14]) ? 4'b1100 : 4'b1100;
													assign node3467 = (inp[8]) ? node3475 : node3468;
														assign node3468 = (inp[7]) ? node3472 : node3469;
															assign node3469 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node3472 = (inp[2]) ? 4'b0101 : 4'b1100;
														assign node3475 = (inp[7]) ? node3479 : node3476;
															assign node3476 = (inp[14]) ? 4'b0101 : 4'b1100;
															assign node3479 = (inp[2]) ? 4'b0100 : 4'b0100;
												assign node3482 = (inp[13]) ? node3498 : node3483;
													assign node3483 = (inp[7]) ? node3491 : node3484;
														assign node3484 = (inp[8]) ? node3488 : node3485;
															assign node3485 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node3488 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node3491 = (inp[8]) ? node3495 : node3492;
															assign node3492 = (inp[14]) ? 4'b0101 : 4'b1100;
															assign node3495 = (inp[2]) ? 4'b0100 : 4'b0100;
													assign node3498 = (inp[7]) ? node3506 : node3499;
														assign node3499 = (inp[8]) ? node3503 : node3500;
															assign node3500 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node3503 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node3506 = (inp[8]) ? 4'b0100 : node3507;
															assign node3507 = (inp[2]) ? 4'b0101 : 4'b0100;
					assign node3511 = (inp[11]) ? node5327 : node3512;
						assign node3512 = (inp[6]) ? node4440 : node3513;
							assign node3513 = (inp[1]) ? node3981 : node3514;
								assign node3514 = (inp[13]) ? node3746 : node3515;
									assign node3515 = (inp[5]) ? node3623 : node3516;
										assign node3516 = (inp[7]) ? node3572 : node3517;
											assign node3517 = (inp[8]) ? node3541 : node3518;
												assign node3518 = (inp[2]) ? node3534 : node3519;
													assign node3519 = (inp[14]) ? node3527 : node3520;
														assign node3520 = (inp[3]) ? node3524 : node3521;
															assign node3521 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node3524 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node3527 = (inp[3]) ? node3531 : node3528;
															assign node3528 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node3531 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node3534 = (inp[15]) ? node3538 : node3535;
														assign node3535 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node3538 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node3541 = (inp[14]) ? node3557 : node3542;
													assign node3542 = (inp[2]) ? node3550 : node3543;
														assign node3543 = (inp[3]) ? node3547 : node3544;
															assign node3544 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node3547 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node3550 = (inp[15]) ? node3554 : node3551;
															assign node3551 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node3554 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node3557 = (inp[2]) ? node3565 : node3558;
														assign node3558 = (inp[15]) ? node3562 : node3559;
															assign node3559 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node3562 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node3565 = (inp[0]) ? node3569 : node3566;
															assign node3566 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node3569 = (inp[15]) ? 4'b1111 : 4'b1101;
											assign node3572 = (inp[8]) ? node3592 : node3573;
												assign node3573 = (inp[2]) ? node3585 : node3574;
													assign node3574 = (inp[14]) ? node3580 : node3575;
														assign node3575 = (inp[3]) ? 4'b1100 : node3576;
															assign node3576 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node3580 = (inp[0]) ? node3582 : 4'b1111;
															assign node3582 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node3585 = (inp[0]) ? node3589 : node3586;
														assign node3586 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node3589 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node3592 = (inp[14]) ? node3608 : node3593;
													assign node3593 = (inp[2]) ? node3601 : node3594;
														assign node3594 = (inp[3]) ? node3598 : node3595;
															assign node3595 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node3598 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node3601 = (inp[3]) ? node3605 : node3602;
															assign node3602 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node3605 = (inp[0]) ? 4'b1100 : 4'b1100;
													assign node3608 = (inp[2]) ? node3616 : node3609;
														assign node3609 = (inp[15]) ? node3613 : node3610;
															assign node3610 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node3613 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node3616 = (inp[15]) ? node3620 : node3617;
															assign node3617 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node3620 = (inp[0]) ? 4'b1110 : 4'b1100;
										assign node3623 = (inp[14]) ? node3685 : node3624;
											assign node3624 = (inp[8]) ? node3654 : node3625;
												assign node3625 = (inp[7]) ? node3641 : node3626;
													assign node3626 = (inp[2]) ? node3634 : node3627;
														assign node3627 = (inp[3]) ? node3631 : node3628;
															assign node3628 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node3631 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node3634 = (inp[0]) ? node3638 : node3635;
															assign node3635 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node3638 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node3641 = (inp[2]) ? node3649 : node3642;
														assign node3642 = (inp[0]) ? node3646 : node3643;
															assign node3643 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node3646 = (inp[3]) ? 4'b1100 : 4'b1100;
														assign node3649 = (inp[0]) ? node3651 : 4'b1101;
															assign node3651 = (inp[15]) ? 4'b1101 : 4'b1101;
												assign node3654 = (inp[0]) ? node3670 : node3655;
													assign node3655 = (inp[15]) ? node3663 : node3656;
														assign node3656 = (inp[3]) ? node3660 : node3657;
															assign node3657 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node3660 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node3663 = (inp[3]) ? node3667 : node3664;
															assign node3664 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node3667 = (inp[7]) ? 4'b1110 : 4'b1110;
													assign node3670 = (inp[15]) ? node3678 : node3671;
														assign node3671 = (inp[3]) ? node3675 : node3672;
															assign node3672 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node3675 = (inp[2]) ? 4'b1110 : 4'b1110;
														assign node3678 = (inp[3]) ? node3682 : node3679;
															assign node3679 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node3682 = (inp[2]) ? 4'b1100 : 4'b1100;
											assign node3685 = (inp[8]) ? node3717 : node3686;
												assign node3686 = (inp[7]) ? node3702 : node3687;
													assign node3687 = (inp[3]) ? node3695 : node3688;
														assign node3688 = (inp[15]) ? node3692 : node3689;
															assign node3689 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node3692 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node3695 = (inp[2]) ? node3699 : node3696;
															assign node3696 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node3699 = (inp[0]) ? 4'b1100 : 4'b1100;
													assign node3702 = (inp[15]) ? node3710 : node3703;
														assign node3703 = (inp[2]) ? node3707 : node3704;
															assign node3704 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node3707 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node3710 = (inp[0]) ? node3714 : node3711;
															assign node3711 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node3714 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node3717 = (inp[7]) ? node3731 : node3718;
													assign node3718 = (inp[0]) ? node3724 : node3719;
														assign node3719 = (inp[15]) ? node3721 : 4'b1101;
															assign node3721 = (inp[2]) ? 4'b1101 : 4'b1111;
														assign node3724 = (inp[15]) ? node3728 : node3725;
															assign node3725 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node3728 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node3731 = (inp[0]) ? node3739 : node3732;
														assign node3732 = (inp[3]) ? node3736 : node3733;
															assign node3733 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node3736 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node3739 = (inp[3]) ? node3743 : node3740;
															assign node3740 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node3743 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node3746 = (inp[8]) ? node3872 : node3747;
										assign node3747 = (inp[7]) ? node3809 : node3748;
											assign node3748 = (inp[2]) ? node3778 : node3749;
												assign node3749 = (inp[14]) ? node3765 : node3750;
													assign node3750 = (inp[5]) ? node3758 : node3751;
														assign node3751 = (inp[15]) ? node3755 : node3752;
															assign node3752 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node3755 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node3758 = (inp[3]) ? node3762 : node3759;
															assign node3759 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node3762 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node3765 = (inp[15]) ? node3771 : node3766;
														assign node3766 = (inp[5]) ? node3768 : 4'b1100;
															assign node3768 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node3771 = (inp[0]) ? node3775 : node3772;
															assign node3772 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node3775 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node3778 = (inp[3]) ? node3794 : node3779;
													assign node3779 = (inp[5]) ? node3787 : node3780;
														assign node3780 = (inp[14]) ? node3784 : node3781;
															assign node3781 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node3784 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node3787 = (inp[14]) ? node3791 : node3788;
															assign node3788 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node3791 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node3794 = (inp[14]) ? node3802 : node3795;
														assign node3795 = (inp[0]) ? node3799 : node3796;
															assign node3796 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node3799 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node3802 = (inp[5]) ? node3806 : node3803;
															assign node3803 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node3806 = (inp[0]) ? 4'b1100 : 4'b1100;
											assign node3809 = (inp[14]) ? node3841 : node3810;
												assign node3810 = (inp[2]) ? node3826 : node3811;
													assign node3811 = (inp[3]) ? node3819 : node3812;
														assign node3812 = (inp[0]) ? node3816 : node3813;
															assign node3813 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node3816 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node3819 = (inp[0]) ? node3823 : node3820;
															assign node3820 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node3823 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node3826 = (inp[15]) ? node3834 : node3827;
														assign node3827 = (inp[0]) ? node3831 : node3828;
															assign node3828 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node3831 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node3834 = (inp[0]) ? node3838 : node3835;
															assign node3835 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node3838 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node3841 = (inp[5]) ? node3857 : node3842;
													assign node3842 = (inp[2]) ? node3850 : node3843;
														assign node3843 = (inp[0]) ? node3847 : node3844;
															assign node3844 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node3847 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node3850 = (inp[0]) ? node3854 : node3851;
															assign node3851 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node3854 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node3857 = (inp[0]) ? node3865 : node3858;
														assign node3858 = (inp[15]) ? node3862 : node3859;
															assign node3859 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node3862 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node3865 = (inp[2]) ? node3869 : node3866;
															assign node3866 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node3869 = (inp[3]) ? 4'b0101 : 4'b0101;
										assign node3872 = (inp[7]) ? node3928 : node3873;
											assign node3873 = (inp[14]) ? node3905 : node3874;
												assign node3874 = (inp[2]) ? node3890 : node3875;
													assign node3875 = (inp[3]) ? node3883 : node3876;
														assign node3876 = (inp[0]) ? node3880 : node3877;
															assign node3877 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node3880 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node3883 = (inp[0]) ? node3887 : node3884;
															assign node3884 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node3887 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node3890 = (inp[3]) ? node3898 : node3891;
														assign node3891 = (inp[0]) ? node3895 : node3892;
															assign node3892 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node3895 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node3898 = (inp[5]) ? node3902 : node3899;
															assign node3899 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node3902 = (inp[0]) ? 4'b0101 : 4'b0101;
												assign node3905 = (inp[5]) ? node3913 : node3906;
													assign node3906 = (inp[15]) ? node3910 : node3907;
														assign node3907 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node3910 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node3913 = (inp[0]) ? node3921 : node3914;
														assign node3914 = (inp[2]) ? node3918 : node3915;
															assign node3915 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node3918 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node3921 = (inp[15]) ? node3925 : node3922;
															assign node3922 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node3925 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node3928 = (inp[2]) ? node3960 : node3929;
												assign node3929 = (inp[14]) ? node3945 : node3930;
													assign node3930 = (inp[3]) ? node3938 : node3931;
														assign node3931 = (inp[0]) ? node3935 : node3932;
															assign node3932 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node3935 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node3938 = (inp[0]) ? node3942 : node3939;
															assign node3939 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node3942 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node3945 = (inp[3]) ? node3953 : node3946;
														assign node3946 = (inp[15]) ? node3950 : node3947;
															assign node3947 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node3950 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node3953 = (inp[0]) ? node3957 : node3954;
															assign node3954 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node3957 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node3960 = (inp[0]) ? node3972 : node3961;
													assign node3961 = (inp[15]) ? node3967 : node3962;
														assign node3962 = (inp[3]) ? node3964 : 4'b0110;
															assign node3964 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node3967 = (inp[5]) ? node3969 : 4'b0100;
															assign node3969 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node3972 = (inp[15]) ? node3978 : node3973;
														assign node3973 = (inp[5]) ? node3975 : 4'b0100;
															assign node3975 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node3978 = (inp[3]) ? 4'b0100 : 4'b0110;
								assign node3981 = (inp[13]) ? node4211 : node3982;
									assign node3982 = (inp[8]) ? node4100 : node3983;
										assign node3983 = (inp[7]) ? node4047 : node3984;
											assign node3984 = (inp[2]) ? node4016 : node3985;
												assign node3985 = (inp[14]) ? node4001 : node3986;
													assign node3986 = (inp[15]) ? node3994 : node3987;
														assign node3987 = (inp[0]) ? node3991 : node3988;
															assign node3988 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node3991 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node3994 = (inp[0]) ? node3998 : node3995;
															assign node3995 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node3998 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node4001 = (inp[5]) ? node4009 : node4002;
														assign node4002 = (inp[3]) ? node4006 : node4003;
															assign node4003 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node4006 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node4009 = (inp[15]) ? node4013 : node4010;
															assign node4010 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node4013 = (inp[3]) ? 4'b1100 : 4'b1100;
												assign node4016 = (inp[14]) ? node4032 : node4017;
													assign node4017 = (inp[3]) ? node4025 : node4018;
														assign node4018 = (inp[5]) ? node4022 : node4019;
															assign node4019 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node4022 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node4025 = (inp[5]) ? node4029 : node4026;
															assign node4026 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node4029 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node4032 = (inp[3]) ? node4040 : node4033;
														assign node4033 = (inp[5]) ? node4037 : node4034;
															assign node4034 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node4037 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node4040 = (inp[15]) ? node4044 : node4041;
															assign node4041 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node4044 = (inp[0]) ? 4'b1100 : 4'b1100;
											assign node4047 = (inp[14]) ? node4077 : node4048;
												assign node4048 = (inp[2]) ? node4064 : node4049;
													assign node4049 = (inp[3]) ? node4057 : node4050;
														assign node4050 = (inp[5]) ? node4054 : node4051;
															assign node4051 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node4054 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node4057 = (inp[0]) ? node4061 : node4058;
															assign node4058 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node4061 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node4064 = (inp[0]) ? node4070 : node4065;
														assign node4065 = (inp[15]) ? 4'b0101 : node4066;
															assign node4066 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node4070 = (inp[15]) ? node4074 : node4071;
															assign node4071 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node4074 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node4077 = (inp[3]) ? node4085 : node4078;
													assign node4078 = (inp[0]) ? node4082 : node4079;
														assign node4079 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node4082 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node4085 = (inp[0]) ? node4093 : node4086;
														assign node4086 = (inp[15]) ? node4090 : node4087;
															assign node4087 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node4090 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node4093 = (inp[5]) ? node4097 : node4094;
															assign node4094 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node4097 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node4100 = (inp[7]) ? node4152 : node4101;
											assign node4101 = (inp[2]) ? node4129 : node4102;
												assign node4102 = (inp[14]) ? node4116 : node4103;
													assign node4103 = (inp[15]) ? node4111 : node4104;
														assign node4104 = (inp[0]) ? node4108 : node4105;
															assign node4105 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node4108 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node4111 = (inp[0]) ? 4'b1110 : node4112;
															assign node4112 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node4116 = (inp[5]) ? node4124 : node4117;
														assign node4117 = (inp[15]) ? node4121 : node4118;
															assign node4118 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node4121 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node4124 = (inp[3]) ? 4'b0101 : node4125;
															assign node4125 = (inp[0]) ? 4'b0101 : 4'b0101;
												assign node4129 = (inp[15]) ? node4141 : node4130;
													assign node4130 = (inp[0]) ? node4136 : node4131;
														assign node4131 = (inp[3]) ? node4133 : 4'b0111;
															assign node4133 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node4136 = (inp[5]) ? node4138 : 4'b0101;
															assign node4138 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node4141 = (inp[0]) ? node4147 : node4142;
														assign node4142 = (inp[3]) ? node4144 : 4'b0101;
															assign node4144 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node4147 = (inp[5]) ? node4149 : 4'b0111;
															assign node4149 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node4152 = (inp[2]) ? node4182 : node4153;
												assign node4153 = (inp[14]) ? node4167 : node4154;
													assign node4154 = (inp[15]) ? node4162 : node4155;
														assign node4155 = (inp[0]) ? node4159 : node4156;
															assign node4156 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node4159 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node4162 = (inp[0]) ? 4'b0111 : node4163;
															assign node4163 = (inp[3]) ? 4'b0101 : 4'b0101;
													assign node4167 = (inp[0]) ? node4175 : node4168;
														assign node4168 = (inp[15]) ? node4172 : node4169;
															assign node4169 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node4172 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node4175 = (inp[15]) ? node4179 : node4176;
															assign node4176 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node4179 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node4182 = (inp[14]) ? node4198 : node4183;
													assign node4183 = (inp[15]) ? node4191 : node4184;
														assign node4184 = (inp[0]) ? node4188 : node4185;
															assign node4185 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node4188 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node4191 = (inp[0]) ? node4195 : node4192;
															assign node4192 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node4195 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node4198 = (inp[3]) ? node4206 : node4199;
														assign node4199 = (inp[0]) ? node4203 : node4200;
															assign node4200 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node4203 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node4206 = (inp[0]) ? node4208 : 4'b0100;
															assign node4208 = (inp[15]) ? 4'b0100 : 4'b0100;
									assign node4211 = (inp[5]) ? node4319 : node4212;
										assign node4212 = (inp[14]) ? node4276 : node4213;
											assign node4213 = (inp[8]) ? node4245 : node4214;
												assign node4214 = (inp[7]) ? node4230 : node4215;
													assign node4215 = (inp[2]) ? node4223 : node4216;
														assign node4216 = (inp[0]) ? node4220 : node4217;
															assign node4217 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node4220 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node4223 = (inp[3]) ? node4227 : node4224;
															assign node4224 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node4227 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node4230 = (inp[2]) ? node4238 : node4231;
														assign node4231 = (inp[15]) ? node4235 : node4232;
															assign node4232 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node4235 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node4238 = (inp[15]) ? node4242 : node4239;
															assign node4239 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node4242 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node4245 = (inp[7]) ? node4261 : node4246;
													assign node4246 = (inp[2]) ? node4254 : node4247;
														assign node4247 = (inp[0]) ? node4251 : node4248;
															assign node4248 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node4251 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node4254 = (inp[3]) ? node4258 : node4255;
															assign node4255 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node4258 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node4261 = (inp[2]) ? node4269 : node4262;
														assign node4262 = (inp[3]) ? node4266 : node4263;
															assign node4263 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node4266 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node4269 = (inp[15]) ? node4273 : node4270;
															assign node4270 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node4273 = (inp[0]) ? 4'b0110 : 4'b0100;
											assign node4276 = (inp[0]) ? node4304 : node4277;
												assign node4277 = (inp[15]) ? node4291 : node4278;
													assign node4278 = (inp[2]) ? node4284 : node4279;
														assign node4279 = (inp[3]) ? 4'b0110 : node4280;
															assign node4280 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node4284 = (inp[8]) ? node4288 : node4285;
															assign node4285 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node4288 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node4291 = (inp[2]) ? node4299 : node4292;
														assign node4292 = (inp[3]) ? node4296 : node4293;
															assign node4293 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node4296 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node4299 = (inp[3]) ? 4'b0100 : node4300;
															assign node4300 = (inp[7]) ? 4'b0100 : 4'b0100;
												assign node4304 = (inp[15]) ? node4312 : node4305;
													assign node4305 = (inp[8]) ? node4309 : node4306;
														assign node4306 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node4309 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node4312 = (inp[8]) ? node4316 : node4313;
														assign node4313 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node4316 = (inp[7]) ? 4'b0110 : 4'b0111;
										assign node4319 = (inp[7]) ? node4377 : node4320;
											assign node4320 = (inp[8]) ? node4348 : node4321;
												assign node4321 = (inp[14]) ? node4335 : node4322;
													assign node4322 = (inp[2]) ? node4330 : node4323;
														assign node4323 = (inp[3]) ? node4327 : node4324;
															assign node4324 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node4327 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node4330 = (inp[15]) ? 4'b0100 : node4331;
															assign node4331 = (inp[3]) ? 4'b0100 : 4'b0100;
													assign node4335 = (inp[2]) ? node4341 : node4336;
														assign node4336 = (inp[0]) ? 4'b0110 : node4337;
															assign node4337 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node4341 = (inp[3]) ? node4345 : node4342;
															assign node4342 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node4345 = (inp[15]) ? 4'b0100 : 4'b0100;
												assign node4348 = (inp[2]) ? node4362 : node4349;
													assign node4349 = (inp[14]) ? node4355 : node4350;
														assign node4350 = (inp[3]) ? 4'b0110 : node4351;
															assign node4351 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node4355 = (inp[3]) ? node4359 : node4356;
															assign node4356 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node4359 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node4362 = (inp[15]) ? node4370 : node4363;
														assign node4363 = (inp[0]) ? node4367 : node4364;
															assign node4364 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node4367 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node4370 = (inp[14]) ? node4374 : node4371;
															assign node4371 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node4374 = (inp[3]) ? 4'b0101 : 4'b0101;
											assign node4377 = (inp[8]) ? node4409 : node4378;
												assign node4378 = (inp[2]) ? node4394 : node4379;
													assign node4379 = (inp[14]) ? node4387 : node4380;
														assign node4380 = (inp[15]) ? node4384 : node4381;
															assign node4381 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node4384 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node4387 = (inp[15]) ? node4391 : node4388;
															assign node4388 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node4391 = (inp[0]) ? 4'b0101 : 4'b0101;
													assign node4394 = (inp[14]) ? node4402 : node4395;
														assign node4395 = (inp[3]) ? node4399 : node4396;
															assign node4396 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node4399 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node4402 = (inp[15]) ? node4406 : node4403;
															assign node4403 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node4406 = (inp[0]) ? 4'b0101 : 4'b0101;
												assign node4409 = (inp[2]) ? node4425 : node4410;
													assign node4410 = (inp[14]) ? node4418 : node4411;
														assign node4411 = (inp[15]) ? node4415 : node4412;
															assign node4412 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node4415 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node4418 = (inp[3]) ? node4422 : node4419;
															assign node4419 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node4422 = (inp[0]) ? 4'b0100 : 4'b0100;
													assign node4425 = (inp[14]) ? node4433 : node4426;
														assign node4426 = (inp[3]) ? node4430 : node4427;
															assign node4427 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node4430 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node4433 = (inp[0]) ? node4437 : node4434;
															assign node4434 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node4437 = (inp[3]) ? 4'b0100 : 4'b0100;
							assign node4440 = (inp[13]) ? node4880 : node4441;
								assign node4441 = (inp[1]) ? node4663 : node4442;
									assign node4442 = (inp[8]) ? node4562 : node4443;
										assign node4443 = (inp[7]) ? node4499 : node4444;
											assign node4444 = (inp[2]) ? node4476 : node4445;
												assign node4445 = (inp[14]) ? node4461 : node4446;
													assign node4446 = (inp[3]) ? node4454 : node4447;
														assign node4447 = (inp[15]) ? node4451 : node4448;
															assign node4448 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node4451 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node4454 = (inp[0]) ? node4458 : node4455;
															assign node4455 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node4458 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node4461 = (inp[5]) ? node4469 : node4462;
														assign node4462 = (inp[0]) ? node4466 : node4463;
															assign node4463 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node4466 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node4469 = (inp[3]) ? node4473 : node4470;
															assign node4470 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node4473 = (inp[0]) ? 4'b0100 : 4'b0100;
												assign node4476 = (inp[15]) ? node4488 : node4477;
													assign node4477 = (inp[0]) ? node4483 : node4478;
														assign node4478 = (inp[5]) ? node4480 : 4'b0110;
															assign node4480 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node4483 = (inp[3]) ? node4485 : 4'b0100;
															assign node4485 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node4488 = (inp[0]) ? node4494 : node4489;
														assign node4489 = (inp[3]) ? node4491 : 4'b0100;
															assign node4491 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node4494 = (inp[5]) ? node4496 : 4'b0110;
															assign node4496 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node4499 = (inp[2]) ? node4531 : node4500;
												assign node4500 = (inp[14]) ? node4516 : node4501;
													assign node4501 = (inp[0]) ? node4509 : node4502;
														assign node4502 = (inp[15]) ? node4506 : node4503;
															assign node4503 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node4506 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node4509 = (inp[15]) ? node4513 : node4510;
															assign node4510 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node4513 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node4516 = (inp[15]) ? node4524 : node4517;
														assign node4517 = (inp[0]) ? node4521 : node4518;
															assign node4518 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node4521 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node4524 = (inp[0]) ? node4528 : node4525;
															assign node4525 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node4528 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node4531 = (inp[3]) ? node4547 : node4532;
													assign node4532 = (inp[5]) ? node4540 : node4533;
														assign node4533 = (inp[0]) ? node4537 : node4534;
															assign node4534 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node4537 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node4540 = (inp[14]) ? node4544 : node4541;
															assign node4541 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node4544 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node4547 = (inp[15]) ? node4555 : node4548;
														assign node4548 = (inp[0]) ? node4552 : node4549;
															assign node4549 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node4552 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node4555 = (inp[5]) ? node4559 : node4556;
															assign node4556 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node4559 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node4562 = (inp[7]) ? node4612 : node4563;
											assign node4563 = (inp[2]) ? node4589 : node4564;
												assign node4564 = (inp[14]) ? node4580 : node4565;
													assign node4565 = (inp[3]) ? node4573 : node4566;
														assign node4566 = (inp[5]) ? node4570 : node4567;
															assign node4567 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node4570 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node4573 = (inp[0]) ? node4577 : node4574;
															assign node4574 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node4577 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node4580 = (inp[0]) ? node4584 : node4581;
														assign node4581 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node4584 = (inp[15]) ? 4'b0111 : node4585;
															assign node4585 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node4589 = (inp[3]) ? node4597 : node4590;
													assign node4590 = (inp[15]) ? node4594 : node4591;
														assign node4591 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node4594 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node4597 = (inp[5]) ? node4605 : node4598;
														assign node4598 = (inp[0]) ? node4602 : node4599;
															assign node4599 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node4602 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node4605 = (inp[14]) ? node4609 : node4606;
															assign node4606 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node4609 = (inp[15]) ? 4'b0101 : 4'b0101;
											assign node4612 = (inp[14]) ? node4640 : node4613;
												assign node4613 = (inp[2]) ? node4629 : node4614;
													assign node4614 = (inp[5]) ? node4622 : node4615;
														assign node4615 = (inp[0]) ? node4619 : node4616;
															assign node4616 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node4619 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node4622 = (inp[0]) ? node4626 : node4623;
															assign node4623 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node4626 = (inp[3]) ? 4'b0101 : 4'b0101;
													assign node4629 = (inp[0]) ? node4637 : node4630;
														assign node4630 = (inp[15]) ? node4634 : node4631;
															assign node4631 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node4634 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node4637 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node4640 = (inp[0]) ? node4652 : node4641;
													assign node4641 = (inp[15]) ? node4647 : node4642;
														assign node4642 = (inp[5]) ? node4644 : 4'b0110;
															assign node4644 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node4647 = (inp[3]) ? node4649 : 4'b0100;
															assign node4649 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node4652 = (inp[15]) ? node4658 : node4653;
														assign node4653 = (inp[5]) ? node4655 : 4'b0100;
															assign node4655 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node4658 = (inp[5]) ? node4660 : 4'b0110;
															assign node4660 = (inp[3]) ? 4'b0100 : 4'b0110;
									assign node4663 = (inp[7]) ? node4773 : node4664;
										assign node4664 = (inp[8]) ? node4720 : node4665;
											assign node4665 = (inp[14]) ? node4697 : node4666;
												assign node4666 = (inp[2]) ? node4682 : node4667;
													assign node4667 = (inp[5]) ? node4675 : node4668;
														assign node4668 = (inp[3]) ? node4672 : node4669;
															assign node4669 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node4672 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node4675 = (inp[3]) ? node4679 : node4676;
															assign node4676 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node4679 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node4682 = (inp[5]) ? node4690 : node4683;
														assign node4683 = (inp[3]) ? node4687 : node4684;
															assign node4684 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node4687 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node4690 = (inp[0]) ? node4694 : node4691;
															assign node4691 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node4694 = (inp[15]) ? 4'b0100 : 4'b0100;
												assign node4697 = (inp[15]) ? node4709 : node4698;
													assign node4698 = (inp[0]) ? node4704 : node4699;
														assign node4699 = (inp[5]) ? node4701 : 4'b0110;
															assign node4701 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node4704 = (inp[3]) ? node4706 : 4'b0100;
															assign node4706 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node4709 = (inp[0]) ? node4715 : node4710;
														assign node4710 = (inp[5]) ? node4712 : 4'b0100;
															assign node4712 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node4715 = (inp[3]) ? node4717 : 4'b0110;
															assign node4717 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node4720 = (inp[14]) ? node4750 : node4721;
												assign node4721 = (inp[2]) ? node4737 : node4722;
													assign node4722 = (inp[15]) ? node4730 : node4723;
														assign node4723 = (inp[0]) ? node4727 : node4724;
															assign node4724 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node4727 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node4730 = (inp[0]) ? node4734 : node4731;
															assign node4731 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node4734 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node4737 = (inp[0]) ? node4745 : node4738;
														assign node4738 = (inp[15]) ? node4742 : node4739;
															assign node4739 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node4742 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node4745 = (inp[15]) ? 4'b1011 : node4746;
															assign node4746 = (inp[3]) ? 4'b1001 : 4'b1001;
												assign node4750 = (inp[0]) ? node4762 : node4751;
													assign node4751 = (inp[15]) ? node4757 : node4752;
														assign node4752 = (inp[5]) ? node4754 : 4'b1011;
															assign node4754 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node4757 = (inp[3]) ? node4759 : 4'b1001;
															assign node4759 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node4762 = (inp[15]) ? node4768 : node4763;
														assign node4763 = (inp[3]) ? node4765 : 4'b1001;
															assign node4765 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node4768 = (inp[5]) ? node4770 : 4'b1011;
															assign node4770 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node4773 = (inp[8]) ? node4827 : node4774;
											assign node4774 = (inp[14]) ? node4804 : node4775;
												assign node4775 = (inp[2]) ? node4791 : node4776;
													assign node4776 = (inp[5]) ? node4784 : node4777;
														assign node4777 = (inp[0]) ? node4781 : node4778;
															assign node4778 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node4781 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node4784 = (inp[0]) ? node4788 : node4785;
															assign node4785 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node4788 = (inp[3]) ? 4'b0100 : 4'b0100;
													assign node4791 = (inp[3]) ? node4797 : node4792;
														assign node4792 = (inp[15]) ? 4'b1001 : node4793;
															assign node4793 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node4797 = (inp[15]) ? node4801 : node4798;
															assign node4798 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node4801 = (inp[5]) ? 4'b1001 : 4'b1001;
												assign node4804 = (inp[0]) ? node4816 : node4805;
													assign node4805 = (inp[15]) ? node4811 : node4806;
														assign node4806 = (inp[3]) ? node4808 : 4'b1011;
															assign node4808 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node4811 = (inp[5]) ? node4813 : 4'b1001;
															assign node4813 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node4816 = (inp[15]) ? node4822 : node4817;
														assign node4817 = (inp[3]) ? node4819 : 4'b1001;
															assign node4819 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node4822 = (inp[5]) ? node4824 : 4'b1011;
															assign node4824 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node4827 = (inp[2]) ? node4857 : node4828;
												assign node4828 = (inp[14]) ? node4842 : node4829;
													assign node4829 = (inp[5]) ? node4837 : node4830;
														assign node4830 = (inp[0]) ? node4834 : node4831;
															assign node4831 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node4834 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node4837 = (inp[15]) ? 4'b1011 : node4838;
															assign node4838 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node4842 = (inp[5]) ? node4850 : node4843;
														assign node4843 = (inp[15]) ? node4847 : node4844;
															assign node4844 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node4847 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node4850 = (inp[15]) ? node4854 : node4851;
															assign node4851 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node4854 = (inp[3]) ? 4'b1000 : 4'b1000;
												assign node4857 = (inp[3]) ? node4865 : node4858;
													assign node4858 = (inp[15]) ? node4862 : node4859;
														assign node4859 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node4862 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node4865 = (inp[5]) ? node4873 : node4866;
														assign node4866 = (inp[15]) ? node4870 : node4867;
															assign node4867 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node4870 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node4873 = (inp[0]) ? node4877 : node4874;
															assign node4874 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node4877 = (inp[15]) ? 4'b1000 : 4'b1010;
								assign node4880 = (inp[1]) ? node5100 : node4881;
									assign node4881 = (inp[7]) ? node4995 : node4882;
										assign node4882 = (inp[8]) ? node4942 : node4883;
											assign node4883 = (inp[2]) ? node4911 : node4884;
												assign node4884 = (inp[14]) ? node4898 : node4885;
													assign node4885 = (inp[5]) ? node4893 : node4886;
														assign node4886 = (inp[0]) ? node4890 : node4887;
															assign node4887 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node4890 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node4893 = (inp[3]) ? node4895 : 4'b0101;
															assign node4895 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node4898 = (inp[0]) ? node4904 : node4899;
														assign node4899 = (inp[15]) ? 4'b0100 : node4900;
															assign node4900 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node4904 = (inp[15]) ? node4908 : node4905;
															assign node4905 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node4908 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node4911 = (inp[3]) ? node4927 : node4912;
													assign node4912 = (inp[5]) ? node4920 : node4913;
														assign node4913 = (inp[14]) ? node4917 : node4914;
															assign node4914 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node4917 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node4920 = (inp[15]) ? node4924 : node4921;
															assign node4921 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node4924 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node4927 = (inp[5]) ? node4935 : node4928;
														assign node4928 = (inp[0]) ? node4932 : node4929;
															assign node4929 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node4932 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node4935 = (inp[14]) ? node4939 : node4936;
															assign node4936 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node4939 = (inp[15]) ? 4'b0100 : 4'b0100;
											assign node4942 = (inp[14]) ? node4972 : node4943;
												assign node4943 = (inp[2]) ? node4957 : node4944;
													assign node4944 = (inp[0]) ? node4952 : node4945;
														assign node4945 = (inp[15]) ? node4949 : node4946;
															assign node4946 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node4949 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node4952 = (inp[15]) ? 4'b0110 : node4953;
															assign node4953 = (inp[3]) ? 4'b0100 : 4'b0100;
													assign node4957 = (inp[5]) ? node4965 : node4958;
														assign node4958 = (inp[3]) ? node4962 : node4959;
															assign node4959 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node4962 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node4965 = (inp[0]) ? node4969 : node4966;
															assign node4966 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node4969 = (inp[3]) ? 4'b1001 : 4'b1001;
												assign node4972 = (inp[0]) ? node4984 : node4973;
													assign node4973 = (inp[15]) ? node4979 : node4974;
														assign node4974 = (inp[5]) ? node4976 : 4'b1011;
															assign node4976 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node4979 = (inp[3]) ? node4981 : 4'b1001;
															assign node4981 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node4984 = (inp[15]) ? node4990 : node4985;
														assign node4985 = (inp[5]) ? node4987 : 4'b1001;
															assign node4987 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node4990 = (inp[3]) ? node4992 : 4'b1011;
															assign node4992 = (inp[5]) ? 4'b1001 : 4'b1011;
										assign node4995 = (inp[8]) ? node5049 : node4996;
											assign node4996 = (inp[14]) ? node5026 : node4997;
												assign node4997 = (inp[2]) ? node5013 : node4998;
													assign node4998 = (inp[5]) ? node5006 : node4999;
														assign node4999 = (inp[0]) ? node5003 : node5000;
															assign node5000 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node5003 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node5006 = (inp[0]) ? node5010 : node5007;
															assign node5007 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node5010 = (inp[3]) ? 4'b0100 : 4'b0100;
													assign node5013 = (inp[0]) ? node5019 : node5014;
														assign node5014 = (inp[15]) ? node5016 : 4'b1011;
															assign node5016 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node5019 = (inp[15]) ? node5023 : node5020;
															assign node5020 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node5023 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node5026 = (inp[0]) ? node5038 : node5027;
													assign node5027 = (inp[15]) ? node5033 : node5028;
														assign node5028 = (inp[3]) ? node5030 : 4'b1011;
															assign node5030 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node5033 = (inp[5]) ? node5035 : 4'b1001;
															assign node5035 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node5038 = (inp[15]) ? node5044 : node5039;
														assign node5039 = (inp[3]) ? node5041 : 4'b1001;
															assign node5041 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node5044 = (inp[5]) ? node5046 : 4'b1011;
															assign node5046 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node5049 = (inp[2]) ? node5079 : node5050;
												assign node5050 = (inp[14]) ? node5066 : node5051;
													assign node5051 = (inp[15]) ? node5059 : node5052;
														assign node5052 = (inp[0]) ? node5056 : node5053;
															assign node5053 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node5056 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node5059 = (inp[0]) ? node5063 : node5060;
															assign node5060 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node5063 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node5066 = (inp[5]) ? node5072 : node5067;
														assign node5067 = (inp[3]) ? node5069 : 4'b1000;
															assign node5069 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node5072 = (inp[3]) ? node5076 : node5073;
															assign node5073 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node5076 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node5079 = (inp[3]) ? node5087 : node5080;
													assign node5080 = (inp[15]) ? node5084 : node5081;
														assign node5081 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node5084 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node5087 = (inp[5]) ? node5093 : node5088;
														assign node5088 = (inp[14]) ? 4'b1010 : node5089;
															assign node5089 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node5093 = (inp[14]) ? node5097 : node5094;
															assign node5094 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node5097 = (inp[0]) ? 4'b1000 : 4'b1000;
									assign node5100 = (inp[5]) ? node5208 : node5101;
										assign node5101 = (inp[7]) ? node5155 : node5102;
											assign node5102 = (inp[8]) ? node5132 : node5103;
												assign node5103 = (inp[2]) ? node5119 : node5104;
													assign node5104 = (inp[14]) ? node5112 : node5105;
														assign node5105 = (inp[0]) ? node5109 : node5106;
															assign node5106 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node5109 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node5112 = (inp[15]) ? node5116 : node5113;
															assign node5113 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node5116 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node5119 = (inp[3]) ? node5127 : node5120;
														assign node5120 = (inp[0]) ? node5124 : node5121;
															assign node5121 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node5124 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node5127 = (inp[14]) ? 4'b1000 : node5128;
															assign node5128 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node5132 = (inp[14]) ? node5148 : node5133;
													assign node5133 = (inp[2]) ? node5141 : node5134;
														assign node5134 = (inp[3]) ? node5138 : node5135;
															assign node5135 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node5138 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node5141 = (inp[3]) ? node5145 : node5142;
															assign node5142 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node5145 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node5148 = (inp[0]) ? node5152 : node5149;
														assign node5149 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node5152 = (inp[15]) ? 4'b1011 : 4'b1001;
											assign node5155 = (inp[8]) ? node5179 : node5156;
												assign node5156 = (inp[2]) ? node5172 : node5157;
													assign node5157 = (inp[14]) ? node5165 : node5158;
														assign node5158 = (inp[0]) ? node5162 : node5159;
															assign node5159 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node5162 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node5165 = (inp[0]) ? node5169 : node5166;
															assign node5166 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node5169 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node5172 = (inp[15]) ? node5176 : node5173;
														assign node5173 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node5176 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node5179 = (inp[2]) ? node5193 : node5180;
													assign node5180 = (inp[14]) ? node5188 : node5181;
														assign node5181 = (inp[0]) ? node5185 : node5182;
															assign node5182 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node5185 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node5188 = (inp[3]) ? 4'b1010 : node5189;
															assign node5189 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node5193 = (inp[14]) ? node5201 : node5194;
														assign node5194 = (inp[3]) ? node5198 : node5195;
															assign node5195 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node5198 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node5201 = (inp[3]) ? node5205 : node5202;
															assign node5202 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node5205 = (inp[15]) ? 4'b1000 : 4'b1000;
										assign node5208 = (inp[7]) ? node5268 : node5209;
											assign node5209 = (inp[8]) ? node5239 : node5210;
												assign node5210 = (inp[2]) ? node5226 : node5211;
													assign node5211 = (inp[14]) ? node5219 : node5212;
														assign node5212 = (inp[15]) ? node5216 : node5213;
															assign node5213 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node5216 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node5219 = (inp[15]) ? node5223 : node5220;
															assign node5220 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node5223 = (inp[3]) ? 4'b1000 : 4'b1000;
													assign node5226 = (inp[14]) ? node5234 : node5227;
														assign node5227 = (inp[15]) ? node5231 : node5228;
															assign node5228 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node5231 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node5234 = (inp[15]) ? 4'b1000 : node5235;
															assign node5235 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node5239 = (inp[14]) ? node5253 : node5240;
													assign node5240 = (inp[2]) ? node5246 : node5241;
														assign node5241 = (inp[15]) ? node5243 : 4'b1000;
															assign node5243 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node5246 = (inp[3]) ? node5250 : node5247;
															assign node5247 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node5250 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node5253 = (inp[3]) ? node5261 : node5254;
														assign node5254 = (inp[0]) ? node5258 : node5255;
															assign node5255 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node5258 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node5261 = (inp[2]) ? node5265 : node5262;
															assign node5262 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node5265 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node5268 = (inp[8]) ? node5296 : node5269;
												assign node5269 = (inp[2]) ? node5283 : node5270;
													assign node5270 = (inp[14]) ? node5278 : node5271;
														assign node5271 = (inp[3]) ? node5275 : node5272;
															assign node5272 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node5275 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node5278 = (inp[15]) ? node5280 : 4'b1011;
															assign node5280 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node5283 = (inp[3]) ? node5291 : node5284;
														assign node5284 = (inp[15]) ? node5288 : node5285;
															assign node5285 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node5288 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node5291 = (inp[14]) ? node5293 : 4'b1011;
															assign node5293 = (inp[0]) ? 4'b1001 : 4'b1001;
												assign node5296 = (inp[14]) ? node5312 : node5297;
													assign node5297 = (inp[2]) ? node5305 : node5298;
														assign node5298 = (inp[0]) ? node5302 : node5299;
															assign node5299 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node5302 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node5305 = (inp[0]) ? node5309 : node5306;
															assign node5306 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node5309 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node5312 = (inp[3]) ? node5320 : node5313;
														assign node5313 = (inp[2]) ? node5317 : node5314;
															assign node5314 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node5317 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node5320 = (inp[2]) ? node5324 : node5321;
															assign node5321 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node5324 = (inp[15]) ? 4'b1000 : 4'b1000;
						assign node5327 = (inp[6]) ? node6233 : node5328;
							assign node5328 = (inp[13]) ? node5770 : node5329;
								assign node5329 = (inp[1]) ? node5549 : node5330;
									assign node5330 = (inp[15]) ? node5442 : node5331;
										assign node5331 = (inp[0]) ? node5387 : node5332;
											assign node5332 = (inp[3]) ? node5358 : node5333;
												assign node5333 = (inp[14]) ? node5343 : node5334;
													assign node5334 = (inp[8]) ? node5336 : 4'b0110;
														assign node5336 = (inp[7]) ? node5340 : node5337;
															assign node5337 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node5340 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node5343 = (inp[5]) ? node5351 : node5344;
														assign node5344 = (inp[8]) ? node5348 : node5345;
															assign node5345 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node5348 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node5351 = (inp[8]) ? node5355 : node5352;
															assign node5352 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node5355 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node5358 = (inp[5]) ? node5372 : node5359;
													assign node5359 = (inp[14]) ? node5365 : node5360;
														assign node5360 = (inp[8]) ? 4'b0111 : node5361;
															assign node5361 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node5365 = (inp[8]) ? node5369 : node5366;
															assign node5366 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node5369 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node5372 = (inp[14]) ? node5380 : node5373;
														assign node5373 = (inp[8]) ? node5377 : node5374;
															assign node5374 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node5377 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node5380 = (inp[7]) ? node5384 : node5381;
															assign node5381 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node5384 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node5387 = (inp[3]) ? node5411 : node5388;
												assign node5388 = (inp[7]) ? node5400 : node5389;
													assign node5389 = (inp[8]) ? node5395 : node5390;
														assign node5390 = (inp[14]) ? 4'b0100 : node5391;
															assign node5391 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node5395 = (inp[14]) ? 4'b0101 : node5396;
															assign node5396 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node5400 = (inp[8]) ? node5406 : node5401;
														assign node5401 = (inp[2]) ? 4'b0101 : node5402;
															assign node5402 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node5406 = (inp[2]) ? 4'b0100 : node5407;
															assign node5407 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node5411 = (inp[5]) ? node5427 : node5412;
													assign node5412 = (inp[8]) ? node5420 : node5413;
														assign node5413 = (inp[7]) ? node5417 : node5414;
															assign node5414 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node5417 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node5420 = (inp[14]) ? node5424 : node5421;
															assign node5421 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node5424 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node5427 = (inp[7]) ? node5435 : node5428;
														assign node5428 = (inp[8]) ? node5432 : node5429;
															assign node5429 = (inp[2]) ? 4'b0110 : 4'b0110;
															assign node5432 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node5435 = (inp[8]) ? node5439 : node5436;
															assign node5436 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node5439 = (inp[14]) ? 4'b0110 : 4'b0110;
										assign node5442 = (inp[0]) ? node5496 : node5443;
											assign node5443 = (inp[3]) ? node5467 : node5444;
												assign node5444 = (inp[7]) ? node5456 : node5445;
													assign node5445 = (inp[8]) ? node5451 : node5446;
														assign node5446 = (inp[2]) ? 4'b0100 : node5447;
															assign node5447 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node5451 = (inp[2]) ? 4'b0101 : node5452;
															assign node5452 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node5456 = (inp[8]) ? node5462 : node5457;
														assign node5457 = (inp[14]) ? 4'b0101 : node5458;
															assign node5458 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node5462 = (inp[14]) ? 4'b0100 : node5463;
															assign node5463 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node5467 = (inp[5]) ? node5481 : node5468;
													assign node5468 = (inp[14]) ? node5476 : node5469;
														assign node5469 = (inp[2]) ? node5473 : node5470;
															assign node5470 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node5473 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node5476 = (inp[2]) ? node5478 : 4'b0101;
															assign node5478 = (inp[8]) ? 4'b0100 : 4'b0100;
													assign node5481 = (inp[2]) ? node5489 : node5482;
														assign node5482 = (inp[8]) ? node5486 : node5483;
															assign node5483 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node5486 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node5489 = (inp[14]) ? node5493 : node5490;
															assign node5490 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node5493 = (inp[8]) ? 4'b0110 : 4'b0110;
											assign node5496 = (inp[3]) ? node5520 : node5497;
												assign node5497 = (inp[2]) ? node5513 : node5498;
													assign node5498 = (inp[5]) ? node5506 : node5499;
														assign node5499 = (inp[8]) ? node5503 : node5500;
															assign node5500 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node5503 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node5506 = (inp[7]) ? node5510 : node5507;
															assign node5507 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node5510 = (inp[14]) ? 4'b0110 : 4'b0110;
													assign node5513 = (inp[8]) ? node5517 : node5514;
														assign node5514 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node5517 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node5520 = (inp[5]) ? node5536 : node5521;
													assign node5521 = (inp[7]) ? node5529 : node5522;
														assign node5522 = (inp[8]) ? node5526 : node5523;
															assign node5523 = (inp[2]) ? 4'b0110 : 4'b0110;
															assign node5526 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node5529 = (inp[8]) ? node5533 : node5530;
															assign node5530 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node5533 = (inp[14]) ? 4'b0110 : 4'b0110;
													assign node5536 = (inp[14]) ? node5542 : node5537;
														assign node5537 = (inp[7]) ? 4'b0101 : node5538;
															assign node5538 = (inp[2]) ? 4'b0100 : 4'b0100;
														assign node5542 = (inp[2]) ? node5546 : node5543;
															assign node5543 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node5546 = (inp[7]) ? 4'b0100 : 4'b0100;
									assign node5549 = (inp[7]) ? node5655 : node5550;
										assign node5550 = (inp[8]) ? node5602 : node5551;
											assign node5551 = (inp[14]) ? node5579 : node5552;
												assign node5552 = (inp[2]) ? node5564 : node5553;
													assign node5553 = (inp[0]) ? node5559 : node5554;
														assign node5554 = (inp[15]) ? node5556 : 4'b0111;
															assign node5556 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node5559 = (inp[15]) ? node5561 : 4'b0101;
															assign node5561 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node5564 = (inp[5]) ? node5572 : node5565;
														assign node5565 = (inp[0]) ? node5569 : node5566;
															assign node5566 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node5569 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node5572 = (inp[15]) ? node5576 : node5573;
															assign node5573 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node5576 = (inp[3]) ? 4'b0100 : 4'b0100;
												assign node5579 = (inp[0]) ? node5591 : node5580;
													assign node5580 = (inp[15]) ? node5586 : node5581;
														assign node5581 = (inp[3]) ? node5583 : 4'b0110;
															assign node5583 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node5586 = (inp[5]) ? node5588 : 4'b0100;
															assign node5588 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node5591 = (inp[15]) ? node5597 : node5592;
														assign node5592 = (inp[5]) ? node5594 : 4'b0100;
															assign node5594 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node5597 = (inp[3]) ? node5599 : 4'b0110;
															assign node5599 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node5602 = (inp[14]) ? node5632 : node5603;
												assign node5603 = (inp[2]) ? node5619 : node5604;
													assign node5604 = (inp[5]) ? node5612 : node5605;
														assign node5605 = (inp[3]) ? node5609 : node5606;
															assign node5606 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node5609 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node5612 = (inp[3]) ? node5616 : node5613;
															assign node5613 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node5616 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node5619 = (inp[3]) ? node5627 : node5620;
														assign node5620 = (inp[15]) ? node5624 : node5621;
															assign node5621 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node5624 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node5627 = (inp[15]) ? node5629 : 4'b1001;
															assign node5629 = (inp[0]) ? 4'b1001 : 4'b1001;
												assign node5632 = (inp[5]) ? node5640 : node5633;
													assign node5633 = (inp[15]) ? node5637 : node5634;
														assign node5634 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node5637 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node5640 = (inp[2]) ? node5648 : node5641;
														assign node5641 = (inp[15]) ? node5645 : node5642;
															assign node5642 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node5645 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node5648 = (inp[15]) ? node5652 : node5649;
															assign node5649 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node5652 = (inp[3]) ? 4'b1001 : 4'b1001;
										assign node5655 = (inp[8]) ? node5709 : node5656;
											assign node5656 = (inp[14]) ? node5686 : node5657;
												assign node5657 = (inp[2]) ? node5673 : node5658;
													assign node5658 = (inp[5]) ? node5666 : node5659;
														assign node5659 = (inp[0]) ? node5663 : node5660;
															assign node5660 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node5663 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node5666 = (inp[0]) ? node5670 : node5667;
															assign node5667 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node5670 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node5673 = (inp[5]) ? node5681 : node5674;
														assign node5674 = (inp[0]) ? node5678 : node5675;
															assign node5675 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node5678 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node5681 = (inp[0]) ? node5683 : 4'b1001;
															assign node5683 = (inp[3]) ? 4'b1001 : 4'b1001;
												assign node5686 = (inp[15]) ? node5698 : node5687;
													assign node5687 = (inp[0]) ? node5693 : node5688;
														assign node5688 = (inp[5]) ? node5690 : 4'b1011;
															assign node5690 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node5693 = (inp[5]) ? node5695 : 4'b1001;
															assign node5695 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node5698 = (inp[0]) ? node5704 : node5699;
														assign node5699 = (inp[3]) ? node5701 : 4'b1001;
															assign node5701 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node5704 = (inp[5]) ? node5706 : 4'b1011;
															assign node5706 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node5709 = (inp[2]) ? node5739 : node5710;
												assign node5710 = (inp[14]) ? node5724 : node5711;
													assign node5711 = (inp[0]) ? node5717 : node5712;
														assign node5712 = (inp[15]) ? node5714 : 4'b1011;
															assign node5714 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node5717 = (inp[15]) ? node5721 : node5718;
															assign node5718 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node5721 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node5724 = (inp[5]) ? node5732 : node5725;
														assign node5725 = (inp[0]) ? node5729 : node5726;
															assign node5726 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node5729 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node5732 = (inp[3]) ? node5736 : node5733;
															assign node5733 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node5736 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node5739 = (inp[14]) ? node5755 : node5740;
													assign node5740 = (inp[3]) ? node5748 : node5741;
														assign node5741 = (inp[0]) ? node5745 : node5742;
															assign node5742 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node5745 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node5748 = (inp[5]) ? node5752 : node5749;
															assign node5749 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node5752 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node5755 = (inp[15]) ? node5763 : node5756;
														assign node5756 = (inp[0]) ? node5760 : node5757;
															assign node5757 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node5760 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node5763 = (inp[0]) ? node5767 : node5764;
															assign node5764 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node5767 = (inp[5]) ? 4'b1000 : 4'b1010;
								assign node5770 = (inp[1]) ? node6008 : node5771;
									assign node5771 = (inp[7]) ? node5887 : node5772;
										assign node5772 = (inp[8]) ? node5828 : node5773;
											assign node5773 = (inp[2]) ? node5805 : node5774;
												assign node5774 = (inp[14]) ? node5790 : node5775;
													assign node5775 = (inp[15]) ? node5783 : node5776;
														assign node5776 = (inp[0]) ? node5780 : node5777;
															assign node5777 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node5780 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node5783 = (inp[0]) ? node5787 : node5784;
															assign node5784 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node5787 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node5790 = (inp[3]) ? node5798 : node5791;
														assign node5791 = (inp[0]) ? node5795 : node5792;
															assign node5792 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node5795 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node5798 = (inp[15]) ? node5802 : node5799;
															assign node5799 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node5802 = (inp[0]) ? 4'b0100 : 4'b0100;
												assign node5805 = (inp[0]) ? node5817 : node5806;
													assign node5806 = (inp[15]) ? node5812 : node5807;
														assign node5807 = (inp[3]) ? node5809 : 4'b0110;
															assign node5809 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node5812 = (inp[5]) ? node5814 : 4'b0100;
															assign node5814 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node5817 = (inp[15]) ? node5823 : node5818;
														assign node5818 = (inp[3]) ? node5820 : 4'b0100;
															assign node5820 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node5823 = (inp[3]) ? node5825 : 4'b0110;
															assign node5825 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node5828 = (inp[14]) ? node5856 : node5829;
												assign node5829 = (inp[2]) ? node5845 : node5830;
													assign node5830 = (inp[5]) ? node5838 : node5831;
														assign node5831 = (inp[3]) ? node5835 : node5832;
															assign node5832 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node5835 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node5838 = (inp[0]) ? node5842 : node5839;
															assign node5839 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node5842 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node5845 = (inp[5]) ? node5851 : node5846;
														assign node5846 = (inp[0]) ? node5848 : 4'b1011;
															assign node5848 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node5851 = (inp[15]) ? 4'b1001 : node5852;
															assign node5852 = (inp[0]) ? 4'b1001 : 4'b1001;
												assign node5856 = (inp[5]) ? node5872 : node5857;
													assign node5857 = (inp[3]) ? node5865 : node5858;
														assign node5858 = (inp[0]) ? node5862 : node5859;
															assign node5859 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node5862 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node5865 = (inp[0]) ? node5869 : node5866;
															assign node5866 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node5869 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node5872 = (inp[15]) ? node5880 : node5873;
														assign node5873 = (inp[3]) ? node5877 : node5874;
															assign node5874 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node5877 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node5880 = (inp[3]) ? node5884 : node5881;
															assign node5881 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node5884 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node5887 = (inp[8]) ? node5949 : node5888;
											assign node5888 = (inp[2]) ? node5918 : node5889;
												assign node5889 = (inp[14]) ? node5903 : node5890;
													assign node5890 = (inp[0]) ? node5896 : node5891;
														assign node5891 = (inp[15]) ? node5893 : 4'b0110;
															assign node5893 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node5896 = (inp[15]) ? node5900 : node5897;
															assign node5897 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node5900 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node5903 = (inp[3]) ? node5911 : node5904;
														assign node5904 = (inp[0]) ? node5908 : node5905;
															assign node5905 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node5908 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node5911 = (inp[5]) ? node5915 : node5912;
															assign node5912 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node5915 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node5918 = (inp[5]) ? node5934 : node5919;
													assign node5919 = (inp[3]) ? node5927 : node5920;
														assign node5920 = (inp[0]) ? node5924 : node5921;
															assign node5921 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node5924 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node5927 = (inp[14]) ? node5931 : node5928;
															assign node5928 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node5931 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node5934 = (inp[15]) ? node5942 : node5935;
														assign node5935 = (inp[3]) ? node5939 : node5936;
															assign node5936 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node5939 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node5942 = (inp[14]) ? node5946 : node5943;
															assign node5943 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node5946 = (inp[0]) ? 4'b1001 : 4'b1001;
											assign node5949 = (inp[2]) ? node5979 : node5950;
												assign node5950 = (inp[14]) ? node5966 : node5951;
													assign node5951 = (inp[15]) ? node5959 : node5952;
														assign node5952 = (inp[0]) ? node5956 : node5953;
															assign node5953 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node5956 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node5959 = (inp[0]) ? node5963 : node5960;
															assign node5960 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node5963 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node5966 = (inp[0]) ? node5974 : node5967;
														assign node5967 = (inp[15]) ? node5971 : node5968;
															assign node5968 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node5971 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node5974 = (inp[15]) ? node5976 : 4'b1000;
															assign node5976 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node5979 = (inp[14]) ? node5995 : node5980;
													assign node5980 = (inp[15]) ? node5988 : node5981;
														assign node5981 = (inp[0]) ? node5985 : node5982;
															assign node5982 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node5985 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node5988 = (inp[0]) ? node5992 : node5989;
															assign node5989 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node5992 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node5995 = (inp[3]) ? node6001 : node5996;
														assign node5996 = (inp[0]) ? 4'b1010 : node5997;
															assign node5997 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node6001 = (inp[5]) ? node6005 : node6002;
															assign node6002 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node6005 = (inp[0]) ? 4'b1000 : 4'b1000;
									assign node6008 = (inp[7]) ? node6118 : node6009;
										assign node6009 = (inp[8]) ? node6059 : node6010;
											assign node6010 = (inp[14]) ? node6036 : node6011;
												assign node6011 = (inp[2]) ? node6025 : node6012;
													assign node6012 = (inp[5]) ? node6018 : node6013;
														assign node6013 = (inp[3]) ? node6015 : 4'b1011;
															assign node6015 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node6018 = (inp[0]) ? node6022 : node6019;
															assign node6019 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node6022 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node6025 = (inp[15]) ? node6029 : node6026;
														assign node6026 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node6029 = (inp[0]) ? node6033 : node6030;
															assign node6030 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node6033 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node6036 = (inp[15]) ? node6046 : node6037;
													assign node6037 = (inp[0]) ? node6041 : node6038;
														assign node6038 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node6041 = (inp[5]) ? node6043 : 4'b1000;
															assign node6043 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node6046 = (inp[2]) ? node6054 : node6047;
														assign node6047 = (inp[0]) ? node6051 : node6048;
															assign node6048 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node6051 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node6054 = (inp[3]) ? node6056 : 4'b1010;
															assign node6056 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node6059 = (inp[2]) ? node6087 : node6060;
												assign node6060 = (inp[14]) ? node6074 : node6061;
													assign node6061 = (inp[3]) ? node6067 : node6062;
														assign node6062 = (inp[15]) ? node6064 : 4'b1010;
															assign node6064 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node6067 = (inp[0]) ? node6071 : node6068;
															assign node6068 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node6071 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node6074 = (inp[0]) ? node6080 : node6075;
														assign node6075 = (inp[15]) ? node6077 : 4'b1011;
															assign node6077 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node6080 = (inp[15]) ? node6084 : node6081;
															assign node6081 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node6084 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node6087 = (inp[14]) ? node6103 : node6088;
													assign node6088 = (inp[0]) ? node6096 : node6089;
														assign node6089 = (inp[15]) ? node6093 : node6090;
															assign node6090 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node6093 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node6096 = (inp[15]) ? node6100 : node6097;
															assign node6097 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node6100 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node6103 = (inp[15]) ? node6111 : node6104;
														assign node6104 = (inp[0]) ? node6108 : node6105;
															assign node6105 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node6108 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node6111 = (inp[0]) ? node6115 : node6112;
															assign node6112 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node6115 = (inp[5]) ? 4'b1001 : 4'b1011;
										assign node6118 = (inp[8]) ? node6172 : node6119;
											assign node6119 = (inp[2]) ? node6149 : node6120;
												assign node6120 = (inp[14]) ? node6136 : node6121;
													assign node6121 = (inp[5]) ? node6129 : node6122;
														assign node6122 = (inp[0]) ? node6126 : node6123;
															assign node6123 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node6126 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node6129 = (inp[3]) ? node6133 : node6130;
															assign node6130 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node6133 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node6136 = (inp[0]) ? node6142 : node6137;
														assign node6137 = (inp[15]) ? 4'b1001 : node6138;
															assign node6138 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node6142 = (inp[15]) ? node6146 : node6143;
															assign node6143 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node6146 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node6149 = (inp[15]) ? node6161 : node6150;
													assign node6150 = (inp[0]) ? node6156 : node6151;
														assign node6151 = (inp[5]) ? node6153 : 4'b1011;
															assign node6153 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node6156 = (inp[5]) ? node6158 : 4'b1001;
															assign node6158 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node6161 = (inp[0]) ? node6167 : node6162;
														assign node6162 = (inp[3]) ? node6164 : 4'b1001;
															assign node6164 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node6167 = (inp[3]) ? node6169 : 4'b1011;
															assign node6169 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node6172 = (inp[14]) ? node6204 : node6173;
												assign node6173 = (inp[2]) ? node6189 : node6174;
													assign node6174 = (inp[3]) ? node6182 : node6175;
														assign node6175 = (inp[0]) ? node6179 : node6176;
															assign node6176 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node6179 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node6182 = (inp[15]) ? node6186 : node6183;
															assign node6183 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node6186 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node6189 = (inp[15]) ? node6197 : node6190;
														assign node6190 = (inp[0]) ? node6194 : node6191;
															assign node6191 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node6194 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node6197 = (inp[0]) ? node6201 : node6198;
															assign node6198 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node6201 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node6204 = (inp[2]) ? node6220 : node6205;
													assign node6205 = (inp[3]) ? node6213 : node6206;
														assign node6206 = (inp[0]) ? node6210 : node6207;
															assign node6207 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node6210 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node6213 = (inp[15]) ? node6217 : node6214;
															assign node6214 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node6217 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node6220 = (inp[3]) ? node6228 : node6221;
														assign node6221 = (inp[5]) ? node6225 : node6222;
															assign node6222 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node6225 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node6228 = (inp[0]) ? 4'b1010 : node6229;
															assign node6229 = (inp[15]) ? 4'b1000 : 4'b1000;
							assign node6233 = (inp[1]) ? node6693 : node6234;
								assign node6234 = (inp[13]) ? node6454 : node6235;
									assign node6235 = (inp[5]) ? node6331 : node6236;
										assign node6236 = (inp[2]) ? node6300 : node6237;
											assign node6237 = (inp[7]) ? node6269 : node6238;
												assign node6238 = (inp[14]) ? node6254 : node6239;
													assign node6239 = (inp[8]) ? node6247 : node6240;
														assign node6240 = (inp[15]) ? node6244 : node6241;
															assign node6241 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node6244 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node6247 = (inp[0]) ? node6251 : node6248;
															assign node6248 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node6251 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node6254 = (inp[8]) ? node6262 : node6255;
														assign node6255 = (inp[15]) ? node6259 : node6256;
															assign node6256 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node6259 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node6262 = (inp[3]) ? node6266 : node6263;
															assign node6263 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node6266 = (inp[15]) ? 4'b1001 : 4'b1001;
												assign node6269 = (inp[3]) ? node6285 : node6270;
													assign node6270 = (inp[14]) ? node6278 : node6271;
														assign node6271 = (inp[8]) ? node6275 : node6272;
															assign node6272 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node6275 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node6278 = (inp[8]) ? node6282 : node6279;
															assign node6279 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node6282 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node6285 = (inp[0]) ? node6293 : node6286;
														assign node6286 = (inp[15]) ? node6290 : node6287;
															assign node6287 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node6290 = (inp[14]) ? 4'b1000 : 4'b1000;
														assign node6293 = (inp[15]) ? node6297 : node6294;
															assign node6294 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node6297 = (inp[14]) ? 4'b1010 : 4'b1010;
											assign node6300 = (inp[15]) ? node6316 : node6301;
												assign node6301 = (inp[0]) ? node6309 : node6302;
													assign node6302 = (inp[8]) ? node6306 : node6303;
														assign node6303 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node6306 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node6309 = (inp[7]) ? node6313 : node6310;
														assign node6310 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node6313 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node6316 = (inp[0]) ? node6324 : node6317;
													assign node6317 = (inp[7]) ? node6321 : node6318;
														assign node6318 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node6321 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node6324 = (inp[8]) ? node6328 : node6325;
														assign node6325 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node6328 = (inp[7]) ? 4'b1010 : 4'b1011;
										assign node6331 = (inp[3]) ? node6393 : node6332;
											assign node6332 = (inp[8]) ? node6364 : node6333;
												assign node6333 = (inp[7]) ? node6349 : node6334;
													assign node6334 = (inp[2]) ? node6342 : node6335;
														assign node6335 = (inp[14]) ? node6339 : node6336;
															assign node6336 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node6339 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node6342 = (inp[15]) ? node6346 : node6343;
															assign node6343 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node6346 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node6349 = (inp[14]) ? node6357 : node6350;
														assign node6350 = (inp[2]) ? node6354 : node6351;
															assign node6351 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node6354 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node6357 = (inp[0]) ? node6361 : node6358;
															assign node6358 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node6361 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node6364 = (inp[7]) ? node6380 : node6365;
													assign node6365 = (inp[14]) ? node6373 : node6366;
														assign node6366 = (inp[2]) ? node6370 : node6367;
															assign node6367 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node6370 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node6373 = (inp[0]) ? node6377 : node6374;
															assign node6374 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node6377 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node6380 = (inp[2]) ? node6388 : node6381;
														assign node6381 = (inp[14]) ? node6385 : node6382;
															assign node6382 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node6385 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node6388 = (inp[14]) ? 4'b1000 : node6389;
															assign node6389 = (inp[15]) ? 4'b1000 : 4'b1000;
											assign node6393 = (inp[7]) ? node6423 : node6394;
												assign node6394 = (inp[8]) ? node6410 : node6395;
													assign node6395 = (inp[14]) ? node6403 : node6396;
														assign node6396 = (inp[2]) ? node6400 : node6397;
															assign node6397 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node6400 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node6403 = (inp[15]) ? node6407 : node6404;
															assign node6404 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node6407 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node6410 = (inp[2]) ? node6418 : node6411;
														assign node6411 = (inp[14]) ? node6415 : node6412;
															assign node6412 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node6415 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node6418 = (inp[14]) ? 4'b1001 : node6419;
															assign node6419 = (inp[0]) ? 4'b1001 : 4'b1001;
												assign node6423 = (inp[8]) ? node6439 : node6424;
													assign node6424 = (inp[2]) ? node6432 : node6425;
														assign node6425 = (inp[14]) ? node6429 : node6426;
															assign node6426 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node6429 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node6432 = (inp[15]) ? node6436 : node6433;
															assign node6433 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node6436 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node6439 = (inp[2]) ? node6447 : node6440;
														assign node6440 = (inp[14]) ? node6444 : node6441;
															assign node6441 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node6444 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node6447 = (inp[15]) ? node6451 : node6448;
															assign node6448 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node6451 = (inp[0]) ? 4'b1000 : 4'b1010;
									assign node6454 = (inp[8]) ? node6572 : node6455;
										assign node6455 = (inp[7]) ? node6515 : node6456;
											assign node6456 = (inp[14]) ? node6486 : node6457;
												assign node6457 = (inp[2]) ? node6471 : node6458;
													assign node6458 = (inp[15]) ? node6464 : node6459;
														assign node6459 = (inp[0]) ? node6461 : 4'b1011;
															assign node6461 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node6464 = (inp[0]) ? node6468 : node6465;
															assign node6465 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node6468 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node6471 = (inp[0]) ? node6479 : node6472;
														assign node6472 = (inp[15]) ? node6476 : node6473;
															assign node6473 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node6476 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node6479 = (inp[15]) ? node6483 : node6480;
															assign node6480 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node6483 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node6486 = (inp[5]) ? node6500 : node6487;
													assign node6487 = (inp[3]) ? node6495 : node6488;
														assign node6488 = (inp[15]) ? node6492 : node6489;
															assign node6489 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node6492 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node6495 = (inp[2]) ? 4'b1010 : node6496;
															assign node6496 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node6500 = (inp[0]) ? node6508 : node6501;
														assign node6501 = (inp[2]) ? node6505 : node6502;
															assign node6502 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node6505 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node6508 = (inp[3]) ? node6512 : node6509;
															assign node6509 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node6512 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node6515 = (inp[14]) ? node6543 : node6516;
												assign node6516 = (inp[2]) ? node6532 : node6517;
													assign node6517 = (inp[0]) ? node6525 : node6518;
														assign node6518 = (inp[15]) ? node6522 : node6519;
															assign node6519 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node6522 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node6525 = (inp[15]) ? node6529 : node6526;
															assign node6526 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node6529 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node6532 = (inp[15]) ? node6538 : node6533;
														assign node6533 = (inp[5]) ? node6535 : 4'b0011;
															assign node6535 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node6538 = (inp[0]) ? node6540 : 4'b0001;
															assign node6540 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node6543 = (inp[2]) ? node6557 : node6544;
													assign node6544 = (inp[0]) ? node6552 : node6545;
														assign node6545 = (inp[15]) ? node6549 : node6546;
															assign node6546 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node6549 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node6552 = (inp[15]) ? 4'b0011 : node6553;
															assign node6553 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node6557 = (inp[5]) ? node6565 : node6558;
														assign node6558 = (inp[0]) ? node6562 : node6559;
															assign node6559 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node6562 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node6565 = (inp[15]) ? node6569 : node6566;
															assign node6566 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node6569 = (inp[0]) ? 4'b0001 : 4'b0001;
										assign node6572 = (inp[7]) ? node6634 : node6573;
											assign node6573 = (inp[14]) ? node6603 : node6574;
												assign node6574 = (inp[2]) ? node6590 : node6575;
													assign node6575 = (inp[5]) ? node6583 : node6576;
														assign node6576 = (inp[0]) ? node6580 : node6577;
															assign node6577 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node6580 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node6583 = (inp[3]) ? node6587 : node6584;
															assign node6584 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node6587 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node6590 = (inp[5]) ? node6598 : node6591;
														assign node6591 = (inp[15]) ? node6595 : node6592;
															assign node6592 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node6595 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node6598 = (inp[0]) ? node6600 : 4'b0001;
															assign node6600 = (inp[15]) ? 4'b0001 : 4'b0001;
												assign node6603 = (inp[2]) ? node6619 : node6604;
													assign node6604 = (inp[3]) ? node6612 : node6605;
														assign node6605 = (inp[5]) ? node6609 : node6606;
															assign node6606 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node6609 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node6612 = (inp[5]) ? node6616 : node6613;
															assign node6613 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node6616 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node6619 = (inp[3]) ? node6627 : node6620;
														assign node6620 = (inp[15]) ? node6624 : node6621;
															assign node6621 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node6624 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node6627 = (inp[15]) ? node6631 : node6628;
															assign node6628 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node6631 = (inp[0]) ? 4'b0001 : 4'b0001;
											assign node6634 = (inp[2]) ? node6664 : node6635;
												assign node6635 = (inp[14]) ? node6649 : node6636;
													assign node6636 = (inp[15]) ? node6644 : node6637;
														assign node6637 = (inp[0]) ? node6641 : node6638;
															assign node6638 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node6641 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node6644 = (inp[0]) ? 4'b0011 : node6645;
															assign node6645 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node6649 = (inp[15]) ? node6657 : node6650;
														assign node6650 = (inp[0]) ? node6654 : node6651;
															assign node6651 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node6654 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node6657 = (inp[0]) ? node6661 : node6658;
															assign node6658 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node6661 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node6664 = (inp[14]) ? node6680 : node6665;
													assign node6665 = (inp[15]) ? node6673 : node6666;
														assign node6666 = (inp[0]) ? node6670 : node6667;
															assign node6667 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node6670 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node6673 = (inp[0]) ? node6677 : node6674;
															assign node6674 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node6677 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node6680 = (inp[15]) ? node6688 : node6681;
														assign node6681 = (inp[0]) ? node6685 : node6682;
															assign node6682 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node6685 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node6688 = (inp[0]) ? node6690 : 4'b0000;
															assign node6690 = (inp[5]) ? 4'b0000 : 4'b0010;
								assign node6693 = (inp[13]) ? node6923 : node6694;
									assign node6694 = (inp[7]) ? node6804 : node6695;
										assign node6695 = (inp[8]) ? node6749 : node6696;
											assign node6696 = (inp[2]) ? node6728 : node6697;
												assign node6697 = (inp[14]) ? node6713 : node6698;
													assign node6698 = (inp[0]) ? node6706 : node6699;
														assign node6699 = (inp[15]) ? node6703 : node6700;
															assign node6700 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node6703 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node6706 = (inp[15]) ? node6710 : node6707;
															assign node6707 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node6710 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node6713 = (inp[5]) ? node6721 : node6714;
														assign node6714 = (inp[3]) ? node6718 : node6715;
															assign node6715 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node6718 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node6721 = (inp[3]) ? node6725 : node6722;
															assign node6722 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node6725 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node6728 = (inp[5]) ? node6736 : node6729;
													assign node6729 = (inp[0]) ? node6733 : node6730;
														assign node6730 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node6733 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node6736 = (inp[14]) ? node6742 : node6737;
														assign node6737 = (inp[3]) ? node6739 : 4'b1000;
															assign node6739 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node6742 = (inp[0]) ? node6746 : node6743;
															assign node6743 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node6746 = (inp[3]) ? 4'b1000 : 4'b1000;
											assign node6749 = (inp[14]) ? node6775 : node6750;
												assign node6750 = (inp[2]) ? node6762 : node6751;
													assign node6751 = (inp[15]) ? node6757 : node6752;
														assign node6752 = (inp[0]) ? 4'b1000 : node6753;
															assign node6753 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node6757 = (inp[0]) ? 4'b1010 : node6758;
															assign node6758 = (inp[3]) ? 4'b1000 : 4'b1000;
													assign node6762 = (inp[0]) ? node6768 : node6763;
														assign node6763 = (inp[15]) ? 4'b0001 : node6764;
															assign node6764 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node6768 = (inp[3]) ? node6772 : node6769;
															assign node6769 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node6772 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node6775 = (inp[5]) ? node6791 : node6776;
													assign node6776 = (inp[3]) ? node6784 : node6777;
														assign node6777 = (inp[2]) ? node6781 : node6778;
															assign node6778 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node6781 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node6784 = (inp[15]) ? node6788 : node6785;
															assign node6785 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node6788 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node6791 = (inp[3]) ? node6797 : node6792;
														assign node6792 = (inp[2]) ? node6794 : 4'b0011;
															assign node6794 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node6797 = (inp[2]) ? node6801 : node6798;
															assign node6798 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node6801 = (inp[15]) ? 4'b0001 : 4'b0001;
										assign node6804 = (inp[8]) ? node6860 : node6805;
											assign node6805 = (inp[2]) ? node6837 : node6806;
												assign node6806 = (inp[14]) ? node6822 : node6807;
													assign node6807 = (inp[15]) ? node6815 : node6808;
														assign node6808 = (inp[0]) ? node6812 : node6809;
															assign node6809 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node6812 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node6815 = (inp[0]) ? node6819 : node6816;
															assign node6816 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node6819 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node6822 = (inp[3]) ? node6830 : node6823;
														assign node6823 = (inp[0]) ? node6827 : node6824;
															assign node6824 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node6827 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node6830 = (inp[15]) ? node6834 : node6831;
															assign node6831 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node6834 = (inp[0]) ? 4'b0001 : 4'b0001;
												assign node6837 = (inp[0]) ? node6849 : node6838;
													assign node6838 = (inp[15]) ? node6844 : node6839;
														assign node6839 = (inp[5]) ? node6841 : 4'b0011;
															assign node6841 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node6844 = (inp[5]) ? node6846 : 4'b0001;
															assign node6846 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node6849 = (inp[15]) ? node6855 : node6850;
														assign node6850 = (inp[5]) ? node6852 : 4'b0001;
															assign node6852 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node6855 = (inp[5]) ? node6857 : 4'b0011;
															assign node6857 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node6860 = (inp[2]) ? node6892 : node6861;
												assign node6861 = (inp[14]) ? node6877 : node6862;
													assign node6862 = (inp[5]) ? node6870 : node6863;
														assign node6863 = (inp[3]) ? node6867 : node6864;
															assign node6864 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node6867 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node6870 = (inp[15]) ? node6874 : node6871;
															assign node6871 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node6874 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node6877 = (inp[3]) ? node6885 : node6878;
														assign node6878 = (inp[0]) ? node6882 : node6879;
															assign node6879 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node6882 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node6885 = (inp[0]) ? node6889 : node6886;
															assign node6886 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node6889 = (inp[5]) ? 4'b0000 : 4'b0000;
												assign node6892 = (inp[14]) ? node6908 : node6893;
													assign node6893 = (inp[15]) ? node6901 : node6894;
														assign node6894 = (inp[0]) ? node6898 : node6895;
															assign node6895 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node6898 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node6901 = (inp[0]) ? node6905 : node6902;
															assign node6902 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node6905 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node6908 = (inp[3]) ? node6916 : node6909;
														assign node6909 = (inp[0]) ? node6913 : node6910;
															assign node6910 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node6913 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node6916 = (inp[0]) ? node6920 : node6917;
															assign node6917 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node6920 = (inp[5]) ? 4'b0000 : 4'b0000;
									assign node6923 = (inp[2]) ? node7045 : node6924;
										assign node6924 = (inp[5]) ? node6986 : node6925;
											assign node6925 = (inp[3]) ? node6955 : node6926;
												assign node6926 = (inp[8]) ? node6940 : node6927;
													assign node6927 = (inp[7]) ? node6933 : node6928;
														assign node6928 = (inp[14]) ? 4'b0000 : node6929;
															assign node6929 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node6933 = (inp[14]) ? node6937 : node6934;
															assign node6934 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node6937 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node6940 = (inp[0]) ? node6948 : node6941;
														assign node6941 = (inp[15]) ? node6945 : node6942;
															assign node6942 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node6945 = (inp[7]) ? 4'b0000 : 4'b0000;
														assign node6948 = (inp[15]) ? node6952 : node6949;
															assign node6949 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node6952 = (inp[7]) ? 4'b0010 : 4'b0010;
												assign node6955 = (inp[8]) ? node6971 : node6956;
													assign node6956 = (inp[14]) ? node6964 : node6957;
														assign node6957 = (inp[7]) ? node6961 : node6958;
															assign node6958 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node6961 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node6964 = (inp[7]) ? node6968 : node6965;
															assign node6965 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node6968 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node6971 = (inp[0]) ? node6979 : node6972;
														assign node6972 = (inp[15]) ? node6976 : node6973;
															assign node6973 = (inp[14]) ? 4'b0010 : 4'b0010;
															assign node6976 = (inp[14]) ? 4'b0000 : 4'b0000;
														assign node6979 = (inp[15]) ? node6983 : node6980;
															assign node6980 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node6983 = (inp[14]) ? 4'b0011 : 4'b0010;
											assign node6986 = (inp[14]) ? node7016 : node6987;
												assign node6987 = (inp[0]) ? node7003 : node6988;
													assign node6988 = (inp[3]) ? node6996 : node6989;
														assign node6989 = (inp[15]) ? node6993 : node6990;
															assign node6990 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node6993 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node6996 = (inp[15]) ? node7000 : node6997;
															assign node6997 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node7000 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node7003 = (inp[8]) ? node7011 : node7004;
														assign node7004 = (inp[7]) ? node7008 : node7005;
															assign node7005 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node7008 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node7011 = (inp[7]) ? node7013 : 4'b0010;
															assign node7013 = (inp[3]) ? 4'b0001 : 4'b0001;
												assign node7016 = (inp[3]) ? node7032 : node7017;
													assign node7017 = (inp[8]) ? node7025 : node7018;
														assign node7018 = (inp[7]) ? node7022 : node7019;
															assign node7019 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node7022 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node7025 = (inp[7]) ? node7029 : node7026;
															assign node7026 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node7029 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node7032 = (inp[7]) ? node7038 : node7033;
														assign node7033 = (inp[8]) ? node7035 : 4'b0000;
															assign node7035 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node7038 = (inp[8]) ? node7042 : node7039;
															assign node7039 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node7042 = (inp[0]) ? 4'b0000 : 4'b0000;
										assign node7045 = (inp[14]) ? node7107 : node7046;
											assign node7046 = (inp[0]) ? node7076 : node7047;
												assign node7047 = (inp[15]) ? node7063 : node7048;
													assign node7048 = (inp[3]) ? node7056 : node7049;
														assign node7049 = (inp[5]) ? node7053 : node7050;
															assign node7050 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node7053 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node7056 = (inp[5]) ? node7060 : node7057;
															assign node7057 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node7060 = (inp[7]) ? 4'b0000 : 4'b0000;
													assign node7063 = (inp[5]) ? node7069 : node7064;
														assign node7064 = (inp[8]) ? node7066 : 4'b0001;
															assign node7066 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node7069 = (inp[3]) ? node7073 : node7070;
															assign node7070 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node7073 = (inp[7]) ? 4'b0010 : 4'b0010;
												assign node7076 = (inp[15]) ? node7092 : node7077;
													assign node7077 = (inp[5]) ? node7085 : node7078;
														assign node7078 = (inp[3]) ? node7082 : node7079;
															assign node7079 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node7082 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node7085 = (inp[3]) ? node7089 : node7086;
															assign node7086 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node7089 = (inp[7]) ? 4'b0010 : 4'b0010;
													assign node7092 = (inp[3]) ? node7100 : node7093;
														assign node7093 = (inp[8]) ? node7097 : node7094;
															assign node7094 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node7097 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node7100 = (inp[5]) ? node7104 : node7101;
															assign node7101 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node7104 = (inp[8]) ? 4'b0000 : 4'b0000;
											assign node7107 = (inp[8]) ? node7139 : node7108;
												assign node7108 = (inp[7]) ? node7124 : node7109;
													assign node7109 = (inp[15]) ? node7117 : node7110;
														assign node7110 = (inp[0]) ? node7114 : node7111;
															assign node7111 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node7114 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node7117 = (inp[0]) ? node7121 : node7118;
															assign node7118 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node7121 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node7124 = (inp[0]) ? node7132 : node7125;
														assign node7125 = (inp[15]) ? node7129 : node7126;
															assign node7126 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node7129 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node7132 = (inp[15]) ? node7136 : node7133;
															assign node7133 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node7136 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node7139 = (inp[7]) ? node7153 : node7140;
													assign node7140 = (inp[0]) ? node7146 : node7141;
														assign node7141 = (inp[15]) ? node7143 : 4'b0011;
															assign node7143 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node7146 = (inp[15]) ? node7150 : node7147;
															assign node7147 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node7150 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node7153 = (inp[0]) ? node7161 : node7154;
														assign node7154 = (inp[15]) ? node7158 : node7155;
															assign node7155 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node7158 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node7161 = (inp[15]) ? 4'b0010 : node7162;
															assign node7162 = (inp[5]) ? 4'b0010 : 4'b0000;
				assign node7166 = (inp[12]) ? node10778 : node7167;
					assign node7167 = (inp[6]) ? node8967 : node7168;
						assign node7168 = (inp[11]) ? node8076 : node7169;
							assign node7169 = (inp[13]) ? node7611 : node7170;
								assign node7170 = (inp[1]) ? node7400 : node7171;
									assign node7171 = (inp[3]) ? node7277 : node7172;
										assign node7172 = (inp[14]) ? node7232 : node7173;
											assign node7173 = (inp[0]) ? node7203 : node7174;
												assign node7174 = (inp[15]) ? node7188 : node7175;
													assign node7175 = (inp[7]) ? node7183 : node7176;
														assign node7176 = (inp[2]) ? node7180 : node7177;
															assign node7177 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node7180 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node7183 = (inp[5]) ? node7185 : 4'b1110;
															assign node7185 = (inp[8]) ? 4'b1110 : 4'b1110;
													assign node7188 = (inp[5]) ? node7196 : node7189;
														assign node7189 = (inp[7]) ? node7193 : node7190;
															assign node7190 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node7193 = (inp[2]) ? 4'b1100 : 4'b1100;
														assign node7196 = (inp[7]) ? node7200 : node7197;
															assign node7197 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node7200 = (inp[8]) ? 4'b1100 : 4'b1100;
												assign node7203 = (inp[15]) ? node7219 : node7204;
													assign node7204 = (inp[8]) ? node7212 : node7205;
														assign node7205 = (inp[2]) ? node7209 : node7206;
															assign node7206 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node7209 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node7212 = (inp[2]) ? node7216 : node7213;
															assign node7213 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node7216 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node7219 = (inp[8]) ? node7227 : node7220;
														assign node7220 = (inp[7]) ? node7224 : node7221;
															assign node7221 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node7224 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node7227 = (inp[2]) ? node7229 : 4'b1111;
															assign node7229 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node7232 = (inp[0]) ? node7256 : node7233;
												assign node7233 = (inp[15]) ? node7243 : node7234;
													assign node7234 = (inp[5]) ? node7236 : 4'b1111;
														assign node7236 = (inp[7]) ? node7240 : node7237;
															assign node7237 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node7240 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node7243 = (inp[5]) ? node7251 : node7244;
														assign node7244 = (inp[2]) ? node7248 : node7245;
															assign node7245 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node7248 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node7251 = (inp[2]) ? node7253 : 4'b1101;
															assign node7253 = (inp[7]) ? 4'b1100 : 4'b1100;
												assign node7256 = (inp[15]) ? node7264 : node7257;
													assign node7257 = (inp[8]) ? node7261 : node7258;
														assign node7258 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node7261 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node7264 = (inp[2]) ? node7272 : node7265;
														assign node7265 = (inp[7]) ? node7269 : node7266;
															assign node7266 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node7269 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node7272 = (inp[7]) ? node7274 : 4'b1111;
															assign node7274 = (inp[8]) ? 4'b1110 : 4'b1111;
										assign node7277 = (inp[7]) ? node7339 : node7278;
											assign node7278 = (inp[8]) ? node7310 : node7279;
												assign node7279 = (inp[2]) ? node7295 : node7280;
													assign node7280 = (inp[14]) ? node7288 : node7281;
														assign node7281 = (inp[5]) ? node7285 : node7282;
															assign node7282 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node7285 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node7288 = (inp[15]) ? node7292 : node7289;
															assign node7289 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node7292 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node7295 = (inp[15]) ? node7303 : node7296;
														assign node7296 = (inp[14]) ? node7300 : node7297;
															assign node7297 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node7300 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node7303 = (inp[0]) ? node7307 : node7304;
															assign node7304 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node7307 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node7310 = (inp[2]) ? node7324 : node7311;
													assign node7311 = (inp[14]) ? node7319 : node7312;
														assign node7312 = (inp[15]) ? node7316 : node7313;
															assign node7313 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node7316 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node7319 = (inp[15]) ? node7321 : 4'b1111;
															assign node7321 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node7324 = (inp[15]) ? node7332 : node7325;
														assign node7325 = (inp[14]) ? node7329 : node7326;
															assign node7326 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node7329 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node7332 = (inp[5]) ? node7336 : node7333;
															assign node7333 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node7336 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node7339 = (inp[8]) ? node7371 : node7340;
												assign node7340 = (inp[2]) ? node7356 : node7341;
													assign node7341 = (inp[14]) ? node7349 : node7342;
														assign node7342 = (inp[15]) ? node7346 : node7343;
															assign node7343 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node7346 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node7349 = (inp[15]) ? node7353 : node7350;
															assign node7350 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node7353 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node7356 = (inp[15]) ? node7364 : node7357;
														assign node7357 = (inp[5]) ? node7361 : node7358;
															assign node7358 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node7361 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node7364 = (inp[5]) ? node7368 : node7365;
															assign node7365 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node7368 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node7371 = (inp[14]) ? node7385 : node7372;
													assign node7372 = (inp[2]) ? node7378 : node7373;
														assign node7373 = (inp[15]) ? 4'b1101 : node7374;
															assign node7374 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node7378 = (inp[5]) ? node7382 : node7379;
															assign node7379 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node7382 = (inp[0]) ? 4'b1100 : 4'b1100;
													assign node7385 = (inp[2]) ? node7393 : node7386;
														assign node7386 = (inp[0]) ? node7390 : node7387;
															assign node7387 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node7390 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node7393 = (inp[5]) ? node7397 : node7394;
															assign node7394 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node7397 = (inp[0]) ? 4'b1100 : 4'b1100;
									assign node7400 = (inp[7]) ? node7506 : node7401;
										assign node7401 = (inp[8]) ? node7453 : node7402;
											assign node7402 = (inp[14]) ? node7430 : node7403;
												assign node7403 = (inp[2]) ? node7417 : node7404;
													assign node7404 = (inp[15]) ? node7410 : node7405;
														assign node7405 = (inp[0]) ? 4'b1101 : node7406;
															assign node7406 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node7410 = (inp[0]) ? node7414 : node7411;
															assign node7411 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node7414 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node7417 = (inp[15]) ? node7425 : node7418;
														assign node7418 = (inp[0]) ? node7422 : node7419;
															assign node7419 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node7422 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node7425 = (inp[0]) ? node7427 : 4'b1100;
															assign node7427 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node7430 = (inp[15]) ? node7442 : node7431;
													assign node7431 = (inp[0]) ? node7437 : node7432;
														assign node7432 = (inp[3]) ? node7434 : 4'b1110;
															assign node7434 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node7437 = (inp[5]) ? node7439 : 4'b1100;
															assign node7439 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node7442 = (inp[0]) ? node7448 : node7443;
														assign node7443 = (inp[3]) ? node7445 : 4'b1100;
															assign node7445 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node7448 = (inp[5]) ? node7450 : 4'b1110;
															assign node7450 = (inp[3]) ? 4'b1100 : 4'b1110;
											assign node7453 = (inp[14]) ? node7483 : node7454;
												assign node7454 = (inp[2]) ? node7470 : node7455;
													assign node7455 = (inp[15]) ? node7463 : node7456;
														assign node7456 = (inp[0]) ? node7460 : node7457;
															assign node7457 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node7460 = (inp[3]) ? 4'b1100 : 4'b1100;
														assign node7463 = (inp[0]) ? node7467 : node7464;
															assign node7464 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node7467 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node7470 = (inp[0]) ? node7478 : node7471;
														assign node7471 = (inp[15]) ? node7475 : node7472;
															assign node7472 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node7475 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node7478 = (inp[15]) ? node7480 : 4'b0101;
															assign node7480 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node7483 = (inp[3]) ? node7491 : node7484;
													assign node7484 = (inp[15]) ? node7488 : node7485;
														assign node7485 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node7488 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node7491 = (inp[5]) ? node7499 : node7492;
														assign node7492 = (inp[0]) ? node7496 : node7493;
															assign node7493 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node7496 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node7499 = (inp[2]) ? node7503 : node7500;
															assign node7500 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node7503 = (inp[0]) ? 4'b0101 : 4'b0101;
										assign node7506 = (inp[8]) ? node7560 : node7507;
											assign node7507 = (inp[2]) ? node7537 : node7508;
												assign node7508 = (inp[14]) ? node7524 : node7509;
													assign node7509 = (inp[15]) ? node7517 : node7510;
														assign node7510 = (inp[0]) ? node7514 : node7511;
															assign node7511 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node7514 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node7517 = (inp[0]) ? node7521 : node7518;
															assign node7518 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node7521 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node7524 = (inp[0]) ? node7530 : node7525;
														assign node7525 = (inp[15]) ? 4'b0101 : node7526;
															assign node7526 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node7530 = (inp[15]) ? node7534 : node7531;
															assign node7531 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node7534 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node7537 = (inp[15]) ? node7549 : node7538;
													assign node7538 = (inp[0]) ? node7544 : node7539;
														assign node7539 = (inp[3]) ? node7541 : 4'b0111;
															assign node7541 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node7544 = (inp[3]) ? node7546 : 4'b0101;
															assign node7546 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node7549 = (inp[0]) ? node7555 : node7550;
														assign node7550 = (inp[3]) ? node7552 : 4'b0101;
															assign node7552 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node7555 = (inp[3]) ? node7557 : 4'b0111;
															assign node7557 = (inp[5]) ? 4'b0101 : 4'b0111;
											assign node7560 = (inp[14]) ? node7588 : node7561;
												assign node7561 = (inp[2]) ? node7577 : node7562;
													assign node7562 = (inp[3]) ? node7570 : node7563;
														assign node7563 = (inp[15]) ? node7567 : node7564;
															assign node7564 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node7567 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node7570 = (inp[0]) ? node7574 : node7571;
															assign node7571 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node7574 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node7577 = (inp[0]) ? node7583 : node7578;
														assign node7578 = (inp[15]) ? node7580 : 4'b0110;
															assign node7580 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node7583 = (inp[15]) ? node7585 : 4'b0100;
															assign node7585 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node7588 = (inp[0]) ? node7600 : node7589;
													assign node7589 = (inp[15]) ? node7595 : node7590;
														assign node7590 = (inp[5]) ? node7592 : 4'b0110;
															assign node7592 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node7595 = (inp[3]) ? node7597 : 4'b0100;
															assign node7597 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node7600 = (inp[15]) ? node7606 : node7601;
														assign node7601 = (inp[5]) ? node7603 : 4'b0100;
															assign node7603 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node7606 = (inp[3]) ? node7608 : 4'b0110;
															assign node7608 = (inp[5]) ? 4'b0100 : 4'b0110;
								assign node7611 = (inp[1]) ? node7847 : node7612;
									assign node7612 = (inp[7]) ? node7734 : node7613;
										assign node7613 = (inp[8]) ? node7673 : node7614;
											assign node7614 = (inp[2]) ? node7644 : node7615;
												assign node7615 = (inp[14]) ? node7631 : node7616;
													assign node7616 = (inp[3]) ? node7624 : node7617;
														assign node7617 = (inp[15]) ? node7621 : node7618;
															assign node7618 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node7621 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node7624 = (inp[15]) ? node7628 : node7625;
															assign node7625 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node7628 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node7631 = (inp[5]) ? node7637 : node7632;
														assign node7632 = (inp[3]) ? node7634 : 4'b1110;
															assign node7634 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node7637 = (inp[3]) ? node7641 : node7638;
															assign node7638 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node7641 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node7644 = (inp[14]) ? node7658 : node7645;
													assign node7645 = (inp[5]) ? node7653 : node7646;
														assign node7646 = (inp[0]) ? node7650 : node7647;
															assign node7647 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node7650 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node7653 = (inp[15]) ? node7655 : 4'b1110;
															assign node7655 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node7658 = (inp[3]) ? node7666 : node7659;
														assign node7659 = (inp[5]) ? node7663 : node7660;
															assign node7660 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node7663 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node7666 = (inp[5]) ? node7670 : node7667;
															assign node7667 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node7670 = (inp[0]) ? 4'b1100 : 4'b1100;
											assign node7673 = (inp[14]) ? node7705 : node7674;
												assign node7674 = (inp[2]) ? node7690 : node7675;
													assign node7675 = (inp[3]) ? node7683 : node7676;
														assign node7676 = (inp[15]) ? node7680 : node7677;
															assign node7677 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node7680 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node7683 = (inp[0]) ? node7687 : node7684;
															assign node7684 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node7687 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node7690 = (inp[5]) ? node7698 : node7691;
														assign node7691 = (inp[0]) ? node7695 : node7692;
															assign node7692 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node7695 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node7698 = (inp[3]) ? node7702 : node7699;
															assign node7699 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node7702 = (inp[0]) ? 4'b0101 : 4'b0101;
												assign node7705 = (inp[5]) ? node7721 : node7706;
													assign node7706 = (inp[3]) ? node7714 : node7707;
														assign node7707 = (inp[2]) ? node7711 : node7708;
															assign node7708 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node7711 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node7714 = (inp[15]) ? node7718 : node7715;
															assign node7715 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node7718 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node7721 = (inp[2]) ? node7729 : node7722;
														assign node7722 = (inp[0]) ? node7726 : node7723;
															assign node7723 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node7726 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node7729 = (inp[0]) ? 4'b0101 : node7730;
															assign node7730 = (inp[15]) ? 4'b0101 : 4'b0101;
										assign node7734 = (inp[8]) ? node7786 : node7735;
											assign node7735 = (inp[14]) ? node7763 : node7736;
												assign node7736 = (inp[2]) ? node7750 : node7737;
													assign node7737 = (inp[3]) ? node7745 : node7738;
														assign node7738 = (inp[15]) ? node7742 : node7739;
															assign node7739 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node7742 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node7745 = (inp[5]) ? 4'b1110 : node7746;
															assign node7746 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node7750 = (inp[0]) ? node7756 : node7751;
														assign node7751 = (inp[3]) ? node7753 : 4'b0111;
															assign node7753 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node7756 = (inp[15]) ? node7760 : node7757;
															assign node7757 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node7760 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node7763 = (inp[3]) ? node7771 : node7764;
													assign node7764 = (inp[15]) ? node7768 : node7765;
														assign node7765 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node7768 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node7771 = (inp[0]) ? node7779 : node7772;
														assign node7772 = (inp[15]) ? node7776 : node7773;
															assign node7773 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node7776 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node7779 = (inp[15]) ? node7783 : node7780;
															assign node7780 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node7783 = (inp[5]) ? 4'b0101 : 4'b0111;
											assign node7786 = (inp[2]) ? node7816 : node7787;
												assign node7787 = (inp[14]) ? node7803 : node7788;
													assign node7788 = (inp[3]) ? node7796 : node7789;
														assign node7789 = (inp[5]) ? node7793 : node7790;
															assign node7790 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node7793 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node7796 = (inp[0]) ? node7800 : node7797;
															assign node7797 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node7800 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node7803 = (inp[3]) ? node7809 : node7804;
														assign node7804 = (inp[5]) ? 4'b0110 : node7805;
															assign node7805 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node7809 = (inp[0]) ? node7813 : node7810;
															assign node7810 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node7813 = (inp[15]) ? 4'b0100 : 4'b0100;
												assign node7816 = (inp[3]) ? node7832 : node7817;
													assign node7817 = (inp[14]) ? node7825 : node7818;
														assign node7818 = (inp[0]) ? node7822 : node7819;
															assign node7819 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node7822 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node7825 = (inp[15]) ? node7829 : node7826;
															assign node7826 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node7829 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node7832 = (inp[5]) ? node7840 : node7833;
														assign node7833 = (inp[15]) ? node7837 : node7834;
															assign node7834 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node7837 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node7840 = (inp[0]) ? node7844 : node7841;
															assign node7841 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node7844 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node7847 = (inp[0]) ? node7963 : node7848;
										assign node7848 = (inp[15]) ? node7910 : node7849;
											assign node7849 = (inp[3]) ? node7879 : node7850;
												assign node7850 = (inp[14]) ? node7864 : node7851;
													assign node7851 = (inp[5]) ? node7857 : node7852;
														assign node7852 = (inp[8]) ? node7854 : 4'b0110;
															assign node7854 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node7857 = (inp[7]) ? node7861 : node7858;
															assign node7858 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node7861 = (inp[2]) ? 4'b0110 : 4'b0110;
													assign node7864 = (inp[5]) ? node7872 : node7865;
														assign node7865 = (inp[7]) ? node7869 : node7866;
															assign node7866 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node7869 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node7872 = (inp[2]) ? node7876 : node7873;
															assign node7873 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node7876 = (inp[8]) ? 4'b0110 : 4'b0110;
												assign node7879 = (inp[5]) ? node7895 : node7880;
													assign node7880 = (inp[2]) ? node7888 : node7881;
														assign node7881 = (inp[8]) ? node7885 : node7882;
															assign node7882 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node7885 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node7888 = (inp[8]) ? node7892 : node7889;
															assign node7889 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node7892 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node7895 = (inp[14]) ? node7903 : node7896;
														assign node7896 = (inp[2]) ? node7900 : node7897;
															assign node7897 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node7900 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node7903 = (inp[7]) ? node7907 : node7904;
															assign node7904 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node7907 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node7910 = (inp[5]) ? node7934 : node7911;
												assign node7911 = (inp[14]) ? node7927 : node7912;
													assign node7912 = (inp[3]) ? node7920 : node7913;
														assign node7913 = (inp[2]) ? node7917 : node7914;
															assign node7914 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node7917 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node7920 = (inp[7]) ? node7924 : node7921;
															assign node7921 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node7924 = (inp[2]) ? 4'b0100 : 4'b0100;
													assign node7927 = (inp[7]) ? node7931 : node7928;
														assign node7928 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node7931 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node7934 = (inp[3]) ? node7950 : node7935;
													assign node7935 = (inp[14]) ? node7943 : node7936;
														assign node7936 = (inp[7]) ? node7940 : node7937;
															assign node7937 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node7940 = (inp[2]) ? 4'b0100 : 4'b0100;
														assign node7943 = (inp[2]) ? node7947 : node7944;
															assign node7944 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node7947 = (inp[8]) ? 4'b0100 : 4'b0100;
													assign node7950 = (inp[8]) ? node7956 : node7951;
														assign node7951 = (inp[7]) ? node7953 : 4'b0110;
															assign node7953 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node7956 = (inp[7]) ? node7960 : node7957;
															assign node7957 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node7960 = (inp[14]) ? 4'b0110 : 4'b0111;
										assign node7963 = (inp[15]) ? node8017 : node7964;
											assign node7964 = (inp[3]) ? node7988 : node7965;
												assign node7965 = (inp[2]) ? node7981 : node7966;
													assign node7966 = (inp[14]) ? node7974 : node7967;
														assign node7967 = (inp[7]) ? node7971 : node7968;
															assign node7968 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node7971 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node7974 = (inp[7]) ? node7978 : node7975;
															assign node7975 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node7978 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node7981 = (inp[8]) ? node7985 : node7982;
														assign node7982 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node7985 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node7988 = (inp[5]) ? node8002 : node7989;
													assign node7989 = (inp[14]) ? node7997 : node7990;
														assign node7990 = (inp[7]) ? node7994 : node7991;
															assign node7991 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node7994 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node7997 = (inp[7]) ? node7999 : 4'b0101;
															assign node7999 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node8002 = (inp[14]) ? node8010 : node8003;
														assign node8003 = (inp[2]) ? node8007 : node8004;
															assign node8004 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node8007 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node8010 = (inp[8]) ? node8014 : node8011;
															assign node8011 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node8014 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node8017 = (inp[5]) ? node8049 : node8018;
												assign node8018 = (inp[14]) ? node8034 : node8019;
													assign node8019 = (inp[8]) ? node8027 : node8020;
														assign node8020 = (inp[3]) ? node8024 : node8021;
															assign node8021 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node8024 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node8027 = (inp[2]) ? node8031 : node8028;
															assign node8028 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node8031 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node8034 = (inp[3]) ? node8042 : node8035;
														assign node8035 = (inp[2]) ? node8039 : node8036;
															assign node8036 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node8039 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node8042 = (inp[7]) ? node8046 : node8043;
															assign node8043 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node8046 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node8049 = (inp[3]) ? node8063 : node8050;
													assign node8050 = (inp[7]) ? node8058 : node8051;
														assign node8051 = (inp[8]) ? node8055 : node8052;
															assign node8052 = (inp[2]) ? 4'b0110 : 4'b0110;
															assign node8055 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node8058 = (inp[8]) ? 4'b0110 : node8059;
															assign node8059 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node8063 = (inp[14]) ? node8069 : node8064;
														assign node8064 = (inp[2]) ? 4'b0101 : node8065;
															assign node8065 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node8069 = (inp[8]) ? node8073 : node8070;
															assign node8070 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node8073 = (inp[7]) ? 4'b0100 : 4'b0101;
							assign node8076 = (inp[13]) ? node8518 : node8077;
								assign node8077 = (inp[1]) ? node8297 : node8078;
									assign node8078 = (inp[15]) ? node8192 : node8079;
										assign node8079 = (inp[0]) ? node8141 : node8080;
											assign node8080 = (inp[5]) ? node8112 : node8081;
												assign node8081 = (inp[3]) ? node8097 : node8082;
													assign node8082 = (inp[14]) ? node8090 : node8083;
														assign node8083 = (inp[8]) ? node8087 : node8084;
															assign node8084 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node8087 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node8090 = (inp[7]) ? node8094 : node8091;
															assign node8091 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node8094 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node8097 = (inp[2]) ? node8105 : node8098;
														assign node8098 = (inp[7]) ? node8102 : node8099;
															assign node8099 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node8102 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node8105 = (inp[7]) ? node8109 : node8106;
															assign node8106 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node8109 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node8112 = (inp[3]) ? node8126 : node8113;
													assign node8113 = (inp[8]) ? node8121 : node8114;
														assign node8114 = (inp[7]) ? node8118 : node8115;
															assign node8115 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node8118 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node8121 = (inp[7]) ? node8123 : 4'b0111;
															assign node8123 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node8126 = (inp[8]) ? node8134 : node8127;
														assign node8127 = (inp[7]) ? node8131 : node8128;
															assign node8128 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node8131 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node8134 = (inp[7]) ? node8138 : node8135;
															assign node8135 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node8138 = (inp[2]) ? 4'b0100 : 4'b0100;
											assign node8141 = (inp[5]) ? node8165 : node8142;
												assign node8142 = (inp[14]) ? node8158 : node8143;
													assign node8143 = (inp[2]) ? node8151 : node8144;
														assign node8144 = (inp[8]) ? node8148 : node8145;
															assign node8145 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node8148 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node8151 = (inp[3]) ? node8155 : node8152;
															assign node8152 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node8155 = (inp[8]) ? 4'b0100 : 4'b0100;
													assign node8158 = (inp[8]) ? node8162 : node8159;
														assign node8159 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node8162 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node8165 = (inp[3]) ? node8179 : node8166;
													assign node8166 = (inp[7]) ? node8172 : node8167;
														assign node8167 = (inp[8]) ? node8169 : 4'b0100;
															assign node8169 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node8172 = (inp[8]) ? node8176 : node8173;
															assign node8173 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node8176 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node8179 = (inp[8]) ? node8185 : node8180;
														assign node8180 = (inp[2]) ? 4'b0111 : node8181;
															assign node8181 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node8185 = (inp[7]) ? node8189 : node8186;
															assign node8186 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node8189 = (inp[2]) ? 4'b0110 : 4'b0110;
										assign node8192 = (inp[0]) ? node8246 : node8193;
											assign node8193 = (inp[3]) ? node8217 : node8194;
												assign node8194 = (inp[7]) ? node8206 : node8195;
													assign node8195 = (inp[8]) ? node8201 : node8196;
														assign node8196 = (inp[14]) ? 4'b0100 : node8197;
															assign node8197 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node8201 = (inp[14]) ? 4'b0101 : node8202;
															assign node8202 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node8206 = (inp[8]) ? node8212 : node8207;
														assign node8207 = (inp[14]) ? 4'b0101 : node8208;
															assign node8208 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node8212 = (inp[2]) ? 4'b0100 : node8213;
															assign node8213 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node8217 = (inp[5]) ? node8231 : node8218;
													assign node8218 = (inp[8]) ? node8224 : node8219;
														assign node8219 = (inp[7]) ? 4'b0101 : node8220;
															assign node8220 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node8224 = (inp[7]) ? node8228 : node8225;
															assign node8225 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node8228 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node8231 = (inp[2]) ? node8239 : node8232;
														assign node8232 = (inp[7]) ? node8236 : node8233;
															assign node8233 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node8236 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node8239 = (inp[8]) ? node8243 : node8240;
															assign node8240 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node8243 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node8246 = (inp[5]) ? node8270 : node8247;
												assign node8247 = (inp[8]) ? node8259 : node8248;
													assign node8248 = (inp[7]) ? node8254 : node8249;
														assign node8249 = (inp[2]) ? 4'b0110 : node8250;
															assign node8250 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node8254 = (inp[14]) ? 4'b0111 : node8255;
															assign node8255 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node8259 = (inp[7]) ? node8265 : node8260;
														assign node8260 = (inp[14]) ? 4'b0111 : node8261;
															assign node8261 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node8265 = (inp[14]) ? 4'b0110 : node8266;
															assign node8266 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node8270 = (inp[3]) ? node8284 : node8271;
													assign node8271 = (inp[8]) ? node8279 : node8272;
														assign node8272 = (inp[7]) ? node8276 : node8273;
															assign node8273 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node8276 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node8279 = (inp[7]) ? 4'b0110 : node8280;
															assign node8280 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node8284 = (inp[7]) ? node8292 : node8285;
														assign node8285 = (inp[8]) ? node8289 : node8286;
															assign node8286 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node8289 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node8292 = (inp[8]) ? 4'b0100 : node8293;
															assign node8293 = (inp[14]) ? 4'b0101 : 4'b0100;
									assign node8297 = (inp[7]) ? node8407 : node8298;
										assign node8298 = (inp[8]) ? node8356 : node8299;
											assign node8299 = (inp[14]) ? node8327 : node8300;
												assign node8300 = (inp[2]) ? node8314 : node8301;
													assign node8301 = (inp[15]) ? node8309 : node8302;
														assign node8302 = (inp[0]) ? node8306 : node8303;
															assign node8303 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node8306 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node8309 = (inp[0]) ? node8311 : 4'b0101;
															assign node8311 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node8314 = (inp[3]) ? node8320 : node8315;
														assign node8315 = (inp[0]) ? node8317 : 4'b0110;
															assign node8317 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node8320 = (inp[0]) ? node8324 : node8321;
															assign node8321 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node8324 = (inp[5]) ? 4'b0100 : 4'b0100;
												assign node8327 = (inp[2]) ? node8343 : node8328;
													assign node8328 = (inp[15]) ? node8336 : node8329;
														assign node8329 = (inp[0]) ? node8333 : node8330;
															assign node8330 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node8333 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node8336 = (inp[0]) ? node8340 : node8337;
															assign node8337 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node8340 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node8343 = (inp[3]) ? node8349 : node8344;
														assign node8344 = (inp[0]) ? 4'b0100 : node8345;
															assign node8345 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node8349 = (inp[5]) ? node8353 : node8350;
															assign node8350 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node8353 = (inp[15]) ? 4'b0100 : 4'b0100;
											assign node8356 = (inp[2]) ? node8384 : node8357;
												assign node8357 = (inp[14]) ? node8373 : node8358;
													assign node8358 = (inp[15]) ? node8366 : node8359;
														assign node8359 = (inp[0]) ? node8363 : node8360;
															assign node8360 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node8363 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node8366 = (inp[0]) ? node8370 : node8367;
															assign node8367 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node8370 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node8373 = (inp[3]) ? node8379 : node8374;
														assign node8374 = (inp[5]) ? node8376 : 4'b1011;
															assign node8376 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node8379 = (inp[15]) ? node8381 : 4'b1001;
															assign node8381 = (inp[5]) ? 4'b1001 : 4'b1001;
												assign node8384 = (inp[15]) ? node8396 : node8385;
													assign node8385 = (inp[0]) ? node8391 : node8386;
														assign node8386 = (inp[3]) ? node8388 : 4'b1011;
															assign node8388 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node8391 = (inp[5]) ? node8393 : 4'b1001;
															assign node8393 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node8396 = (inp[0]) ? node8402 : node8397;
														assign node8397 = (inp[5]) ? node8399 : 4'b1001;
															assign node8399 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node8402 = (inp[5]) ? node8404 : 4'b1011;
															assign node8404 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node8407 = (inp[8]) ? node8467 : node8408;
											assign node8408 = (inp[14]) ? node8436 : node8409;
												assign node8409 = (inp[2]) ? node8423 : node8410;
													assign node8410 = (inp[0]) ? node8416 : node8411;
														assign node8411 = (inp[15]) ? node8413 : 4'b0110;
															assign node8413 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node8416 = (inp[15]) ? node8420 : node8417;
															assign node8417 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node8420 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node8423 = (inp[0]) ? node8429 : node8424;
														assign node8424 = (inp[15]) ? node8426 : 4'b1011;
															assign node8426 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node8429 = (inp[15]) ? node8433 : node8430;
															assign node8430 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node8433 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node8436 = (inp[2]) ? node8452 : node8437;
													assign node8437 = (inp[5]) ? node8445 : node8438;
														assign node8438 = (inp[3]) ? node8442 : node8439;
															assign node8439 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node8442 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node8445 = (inp[0]) ? node8449 : node8446;
															assign node8446 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node8449 = (inp[3]) ? 4'b1001 : 4'b1001;
													assign node8452 = (inp[0]) ? node8460 : node8453;
														assign node8453 = (inp[15]) ? node8457 : node8454;
															assign node8454 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node8457 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node8460 = (inp[15]) ? node8464 : node8461;
															assign node8461 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node8464 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node8467 = (inp[14]) ? node8495 : node8468;
												assign node8468 = (inp[2]) ? node8482 : node8469;
													assign node8469 = (inp[3]) ? node8477 : node8470;
														assign node8470 = (inp[0]) ? node8474 : node8471;
															assign node8471 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node8474 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node8477 = (inp[5]) ? 4'b1001 : node8478;
															assign node8478 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node8482 = (inp[3]) ? node8490 : node8483;
														assign node8483 = (inp[5]) ? node8487 : node8484;
															assign node8484 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node8487 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node8490 = (inp[0]) ? 4'b1000 : node8491;
															assign node8491 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node8495 = (inp[15]) ? node8507 : node8496;
													assign node8496 = (inp[0]) ? node8502 : node8497;
														assign node8497 = (inp[3]) ? node8499 : 4'b1010;
															assign node8499 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node8502 = (inp[3]) ? node8504 : 4'b1000;
															assign node8504 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node8507 = (inp[0]) ? node8513 : node8508;
														assign node8508 = (inp[3]) ? node8510 : 4'b1000;
															assign node8510 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node8513 = (inp[3]) ? node8515 : 4'b1010;
															assign node8515 = (inp[5]) ? 4'b1000 : 4'b1010;
								assign node8518 = (inp[1]) ? node8740 : node8519;
									assign node8519 = (inp[8]) ? node8631 : node8520;
										assign node8520 = (inp[7]) ? node8580 : node8521;
											assign node8521 = (inp[2]) ? node8551 : node8522;
												assign node8522 = (inp[14]) ? node8538 : node8523;
													assign node8523 = (inp[3]) ? node8531 : node8524;
														assign node8524 = (inp[5]) ? node8528 : node8525;
															assign node8525 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node8528 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node8531 = (inp[0]) ? node8535 : node8532;
															assign node8532 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node8535 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node8538 = (inp[3]) ? node8544 : node8539;
														assign node8539 = (inp[5]) ? node8541 : 4'b0100;
															assign node8541 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node8544 = (inp[0]) ? node8548 : node8545;
															assign node8545 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node8548 = (inp[5]) ? 4'b0100 : 4'b0100;
												assign node8551 = (inp[14]) ? node8567 : node8552;
													assign node8552 = (inp[5]) ? node8560 : node8553;
														assign node8553 = (inp[0]) ? node8557 : node8554;
															assign node8554 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node8557 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node8560 = (inp[3]) ? node8564 : node8561;
															assign node8561 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node8564 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node8567 = (inp[0]) ? node8575 : node8568;
														assign node8568 = (inp[15]) ? node8572 : node8569;
															assign node8569 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node8572 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node8575 = (inp[15]) ? 4'b0110 : node8576;
															assign node8576 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node8580 = (inp[2]) ? node8608 : node8581;
												assign node8581 = (inp[14]) ? node8595 : node8582;
													assign node8582 = (inp[0]) ? node8590 : node8583;
														assign node8583 = (inp[15]) ? node8587 : node8584;
															assign node8584 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node8587 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node8590 = (inp[5]) ? node8592 : 4'b0110;
															assign node8592 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node8595 = (inp[15]) ? node8603 : node8596;
														assign node8596 = (inp[0]) ? node8600 : node8597;
															assign node8597 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node8600 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node8603 = (inp[3]) ? node8605 : 4'b1001;
															assign node8605 = (inp[5]) ? 4'b1001 : 4'b1001;
												assign node8608 = (inp[0]) ? node8620 : node8609;
													assign node8609 = (inp[15]) ? node8615 : node8610;
														assign node8610 = (inp[3]) ? node8612 : 4'b1011;
															assign node8612 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node8615 = (inp[5]) ? node8617 : 4'b1001;
															assign node8617 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node8620 = (inp[15]) ? node8626 : node8621;
														assign node8621 = (inp[3]) ? node8623 : 4'b1001;
															assign node8623 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node8626 = (inp[3]) ? node8628 : 4'b1011;
															assign node8628 = (inp[5]) ? 4'b1001 : 4'b1011;
										assign node8631 = (inp[7]) ? node8685 : node8632;
											assign node8632 = (inp[2]) ? node8662 : node8633;
												assign node8633 = (inp[14]) ? node8647 : node8634;
													assign node8634 = (inp[3]) ? node8642 : node8635;
														assign node8635 = (inp[15]) ? node8639 : node8636;
															assign node8636 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node8639 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node8642 = (inp[0]) ? 4'b0100 : node8643;
															assign node8643 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node8647 = (inp[0]) ? node8655 : node8648;
														assign node8648 = (inp[15]) ? node8652 : node8649;
															assign node8649 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node8652 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node8655 = (inp[15]) ? node8659 : node8656;
															assign node8656 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node8659 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node8662 = (inp[15]) ? node8674 : node8663;
													assign node8663 = (inp[0]) ? node8669 : node8664;
														assign node8664 = (inp[5]) ? node8666 : 4'b1011;
															assign node8666 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node8669 = (inp[3]) ? node8671 : 4'b1001;
															assign node8671 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node8674 = (inp[0]) ? node8680 : node8675;
														assign node8675 = (inp[3]) ? node8677 : 4'b1001;
															assign node8677 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node8680 = (inp[3]) ? node8682 : 4'b1011;
															assign node8682 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node8685 = (inp[2]) ? node8717 : node8686;
												assign node8686 = (inp[14]) ? node8702 : node8687;
													assign node8687 = (inp[5]) ? node8695 : node8688;
														assign node8688 = (inp[3]) ? node8692 : node8689;
															assign node8689 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node8692 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node8695 = (inp[0]) ? node8699 : node8696;
															assign node8696 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node8699 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node8702 = (inp[0]) ? node8710 : node8703;
														assign node8703 = (inp[15]) ? node8707 : node8704;
															assign node8704 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node8707 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node8710 = (inp[15]) ? node8714 : node8711;
															assign node8711 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node8714 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node8717 = (inp[0]) ? node8729 : node8718;
													assign node8718 = (inp[15]) ? node8724 : node8719;
														assign node8719 = (inp[3]) ? node8721 : 4'b1010;
															assign node8721 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node8724 = (inp[5]) ? node8726 : 4'b1000;
															assign node8726 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node8729 = (inp[15]) ? node8735 : node8730;
														assign node8730 = (inp[5]) ? node8732 : 4'b1000;
															assign node8732 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node8735 = (inp[5]) ? node8737 : 4'b1010;
															assign node8737 = (inp[3]) ? 4'b1000 : 4'b1010;
									assign node8740 = (inp[8]) ? node8860 : node8741;
										assign node8741 = (inp[7]) ? node8801 : node8742;
											assign node8742 = (inp[2]) ? node8772 : node8743;
												assign node8743 = (inp[14]) ? node8757 : node8744;
													assign node8744 = (inp[15]) ? node8752 : node8745;
														assign node8745 = (inp[0]) ? node8749 : node8746;
															assign node8746 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node8749 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node8752 = (inp[3]) ? node8754 : 4'b1011;
															assign node8754 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node8757 = (inp[15]) ? node8765 : node8758;
														assign node8758 = (inp[0]) ? node8762 : node8759;
															assign node8759 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node8762 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node8765 = (inp[0]) ? node8769 : node8766;
															assign node8766 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node8769 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node8772 = (inp[14]) ? node8788 : node8773;
													assign node8773 = (inp[5]) ? node8781 : node8774;
														assign node8774 = (inp[3]) ? node8778 : node8775;
															assign node8775 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node8778 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node8781 = (inp[15]) ? node8785 : node8782;
															assign node8782 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node8785 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node8788 = (inp[5]) ? node8796 : node8789;
														assign node8789 = (inp[15]) ? node8793 : node8790;
															assign node8790 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node8793 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node8796 = (inp[0]) ? node8798 : 4'b1000;
															assign node8798 = (inp[15]) ? 4'b1000 : 4'b1000;
											assign node8801 = (inp[2]) ? node8831 : node8802;
												assign node8802 = (inp[14]) ? node8818 : node8803;
													assign node8803 = (inp[15]) ? node8811 : node8804;
														assign node8804 = (inp[0]) ? node8808 : node8805;
															assign node8805 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node8808 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node8811 = (inp[0]) ? node8815 : node8812;
															assign node8812 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node8815 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node8818 = (inp[5]) ? node8826 : node8819;
														assign node8819 = (inp[0]) ? node8823 : node8820;
															assign node8820 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node8823 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node8826 = (inp[3]) ? 4'b1001 : node8827;
															assign node8827 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node8831 = (inp[3]) ? node8847 : node8832;
													assign node8832 = (inp[5]) ? node8840 : node8833;
														assign node8833 = (inp[15]) ? node8837 : node8834;
															assign node8834 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node8837 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node8840 = (inp[14]) ? node8844 : node8841;
															assign node8841 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node8844 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node8847 = (inp[5]) ? node8855 : node8848;
														assign node8848 = (inp[0]) ? node8852 : node8849;
															assign node8849 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node8852 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node8855 = (inp[15]) ? node8857 : 4'b1011;
															assign node8857 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node8860 = (inp[7]) ? node8908 : node8861;
											assign node8861 = (inp[2]) ? node8887 : node8862;
												assign node8862 = (inp[14]) ? node8874 : node8863;
													assign node8863 = (inp[15]) ? node8869 : node8864;
														assign node8864 = (inp[0]) ? 4'b1000 : node8865;
															assign node8865 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node8869 = (inp[0]) ? 4'b1010 : node8870;
															assign node8870 = (inp[5]) ? 4'b1000 : 4'b1000;
													assign node8874 = (inp[0]) ? node8880 : node8875;
														assign node8875 = (inp[15]) ? 4'b1001 : node8876;
															assign node8876 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node8880 = (inp[15]) ? node8884 : node8881;
															assign node8881 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node8884 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node8887 = (inp[5]) ? node8895 : node8888;
													assign node8888 = (inp[0]) ? node8892 : node8889;
														assign node8889 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node8892 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node8895 = (inp[3]) ? node8903 : node8896;
														assign node8896 = (inp[14]) ? node8900 : node8897;
															assign node8897 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node8900 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node8903 = (inp[14]) ? 4'b1001 : node8904;
															assign node8904 = (inp[15]) ? 4'b1001 : 4'b1001;
											assign node8908 = (inp[14]) ? node8938 : node8909;
												assign node8909 = (inp[2]) ? node8925 : node8910;
													assign node8910 = (inp[5]) ? node8918 : node8911;
														assign node8911 = (inp[3]) ? node8915 : node8912;
															assign node8912 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node8915 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node8918 = (inp[0]) ? node8922 : node8919;
															assign node8919 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node8922 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node8925 = (inp[0]) ? node8931 : node8926;
														assign node8926 = (inp[3]) ? node8928 : 4'b1000;
															assign node8928 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node8931 = (inp[15]) ? node8935 : node8932;
															assign node8932 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node8935 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node8938 = (inp[2]) ? node8952 : node8939;
													assign node8939 = (inp[15]) ? node8945 : node8940;
														assign node8940 = (inp[0]) ? node8942 : 4'b1010;
															assign node8942 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node8945 = (inp[0]) ? node8949 : node8946;
															assign node8946 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node8949 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node8952 = (inp[3]) ? node8960 : node8953;
														assign node8953 = (inp[15]) ? node8957 : node8954;
															assign node8954 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node8957 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node8960 = (inp[15]) ? node8964 : node8961;
															assign node8961 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node8964 = (inp[5]) ? 4'b1000 : 4'b1000;
						assign node8967 = (inp[11]) ? node9891 : node8968;
							assign node8968 = (inp[13]) ? node9440 : node8969;
								assign node8969 = (inp[1]) ? node9203 : node8970;
									assign node8970 = (inp[3]) ? node9078 : node8971;
										assign node8971 = (inp[14]) ? node9031 : node8972;
											assign node8972 = (inp[2]) ? node9002 : node8973;
												assign node8973 = (inp[0]) ? node8989 : node8974;
													assign node8974 = (inp[15]) ? node8982 : node8975;
														assign node8975 = (inp[7]) ? node8979 : node8976;
															assign node8976 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node8979 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node8982 = (inp[7]) ? node8986 : node8983;
															assign node8983 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node8986 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node8989 = (inp[15]) ? node8995 : node8990;
														assign node8990 = (inp[5]) ? 4'b0100 : node8991;
															assign node8991 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node8995 = (inp[7]) ? node8999 : node8996;
															assign node8996 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node8999 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node9002 = (inp[7]) ? node9016 : node9003;
													assign node9003 = (inp[8]) ? node9011 : node9004;
														assign node9004 = (inp[5]) ? node9008 : node9005;
															assign node9005 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node9008 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node9011 = (inp[15]) ? node9013 : 4'b0101;
															assign node9013 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node9016 = (inp[8]) ? node9024 : node9017;
														assign node9017 = (inp[5]) ? node9021 : node9018;
															assign node9018 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node9021 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node9024 = (inp[15]) ? node9028 : node9025;
															assign node9025 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node9028 = (inp[0]) ? 4'b0110 : 4'b0100;
											assign node9031 = (inp[0]) ? node9055 : node9032;
												assign node9032 = (inp[15]) ? node9040 : node9033;
													assign node9033 = (inp[7]) ? node9037 : node9034;
														assign node9034 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node9037 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node9040 = (inp[5]) ? node9048 : node9041;
														assign node9041 = (inp[8]) ? node9045 : node9042;
															assign node9042 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node9045 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node9048 = (inp[7]) ? node9052 : node9049;
															assign node9049 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node9052 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node9055 = (inp[15]) ? node9071 : node9056;
													assign node9056 = (inp[5]) ? node9064 : node9057;
														assign node9057 = (inp[2]) ? node9061 : node9058;
															assign node9058 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node9061 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node9064 = (inp[7]) ? node9068 : node9065;
															assign node9065 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node9068 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node9071 = (inp[8]) ? node9075 : node9072;
														assign node9072 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node9075 = (inp[7]) ? 4'b0110 : 4'b0111;
										assign node9078 = (inp[15]) ? node9140 : node9079;
											assign node9079 = (inp[14]) ? node9111 : node9080;
												assign node9080 = (inp[2]) ? node9096 : node9081;
													assign node9081 = (inp[8]) ? node9089 : node9082;
														assign node9082 = (inp[7]) ? node9086 : node9083;
															assign node9083 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node9086 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node9089 = (inp[7]) ? node9093 : node9090;
															assign node9090 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node9093 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node9096 = (inp[7]) ? node9104 : node9097;
														assign node9097 = (inp[8]) ? node9101 : node9098;
															assign node9098 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node9101 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node9104 = (inp[8]) ? node9108 : node9105;
															assign node9105 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node9108 = (inp[0]) ? 4'b0100 : 4'b0100;
												assign node9111 = (inp[5]) ? node9125 : node9112;
													assign node9112 = (inp[0]) ? node9118 : node9113;
														assign node9113 = (inp[8]) ? node9115 : 4'b0110;
															assign node9115 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node9118 = (inp[7]) ? node9122 : node9119;
															assign node9119 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node9122 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node9125 = (inp[0]) ? node9133 : node9126;
														assign node9126 = (inp[2]) ? node9130 : node9127;
															assign node9127 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node9130 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node9133 = (inp[7]) ? node9137 : node9134;
															assign node9134 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node9137 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node9140 = (inp[7]) ? node9172 : node9141;
												assign node9141 = (inp[8]) ? node9157 : node9142;
													assign node9142 = (inp[14]) ? node9150 : node9143;
														assign node9143 = (inp[2]) ? node9147 : node9144;
															assign node9144 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node9147 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node9150 = (inp[0]) ? node9154 : node9151;
															assign node9151 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node9154 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node9157 = (inp[14]) ? node9165 : node9158;
														assign node9158 = (inp[2]) ? node9162 : node9159;
															assign node9159 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node9162 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node9165 = (inp[2]) ? node9169 : node9166;
															assign node9166 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node9169 = (inp[5]) ? 4'b0101 : 4'b0101;
												assign node9172 = (inp[8]) ? node9188 : node9173;
													assign node9173 = (inp[14]) ? node9181 : node9174;
														assign node9174 = (inp[2]) ? node9178 : node9175;
															assign node9175 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node9178 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node9181 = (inp[5]) ? node9185 : node9182;
															assign node9182 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node9185 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node9188 = (inp[14]) ? node9196 : node9189;
														assign node9189 = (inp[2]) ? node9193 : node9190;
															assign node9190 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node9193 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node9196 = (inp[5]) ? node9200 : node9197;
															assign node9197 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node9200 = (inp[0]) ? 4'b0100 : 4'b0110;
									assign node9203 = (inp[8]) ? node9321 : node9204;
										assign node9204 = (inp[7]) ? node9268 : node9205;
											assign node9205 = (inp[2]) ? node9237 : node9206;
												assign node9206 = (inp[14]) ? node9222 : node9207;
													assign node9207 = (inp[3]) ? node9215 : node9208;
														assign node9208 = (inp[15]) ? node9212 : node9209;
															assign node9209 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node9212 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node9215 = (inp[5]) ? node9219 : node9216;
															assign node9216 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node9219 = (inp[0]) ? 4'b0101 : 4'b0101;
													assign node9222 = (inp[5]) ? node9230 : node9223;
														assign node9223 = (inp[3]) ? node9227 : node9224;
															assign node9224 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node9227 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node9230 = (inp[3]) ? node9234 : node9231;
															assign node9231 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node9234 = (inp[0]) ? 4'b0100 : 4'b0100;
												assign node9237 = (inp[5]) ? node9253 : node9238;
													assign node9238 = (inp[14]) ? node9246 : node9239;
														assign node9239 = (inp[3]) ? node9243 : node9240;
															assign node9240 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node9243 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node9246 = (inp[0]) ? node9250 : node9247;
															assign node9247 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node9250 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node9253 = (inp[0]) ? node9261 : node9254;
														assign node9254 = (inp[15]) ? node9258 : node9255;
															assign node9255 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node9258 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node9261 = (inp[15]) ? node9265 : node9262;
															assign node9262 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node9265 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node9268 = (inp[14]) ? node9298 : node9269;
												assign node9269 = (inp[2]) ? node9283 : node9270;
													assign node9270 = (inp[3]) ? node9276 : node9271;
														assign node9271 = (inp[0]) ? node9273 : 4'b0100;
															assign node9273 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node9276 = (inp[0]) ? node9280 : node9277;
															assign node9277 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node9280 = (inp[5]) ? 4'b0100 : 4'b0100;
													assign node9283 = (inp[3]) ? node9291 : node9284;
														assign node9284 = (inp[0]) ? node9288 : node9285;
															assign node9285 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node9288 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node9291 = (inp[0]) ? node9295 : node9292;
															assign node9292 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node9295 = (inp[5]) ? 4'b1001 : 4'b1001;
												assign node9298 = (inp[0]) ? node9310 : node9299;
													assign node9299 = (inp[15]) ? node9305 : node9300;
														assign node9300 = (inp[5]) ? node9302 : 4'b1011;
															assign node9302 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node9305 = (inp[3]) ? node9307 : 4'b1001;
															assign node9307 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node9310 = (inp[15]) ? node9316 : node9311;
														assign node9311 = (inp[3]) ? node9313 : 4'b1001;
															assign node9313 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node9316 = (inp[5]) ? node9318 : 4'b1011;
															assign node9318 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node9321 = (inp[7]) ? node9379 : node9322;
											assign node9322 = (inp[2]) ? node9350 : node9323;
												assign node9323 = (inp[14]) ? node9337 : node9324;
													assign node9324 = (inp[0]) ? node9330 : node9325;
														assign node9325 = (inp[3]) ? node9327 : 4'b0110;
															assign node9327 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node9330 = (inp[15]) ? node9334 : node9331;
															assign node9331 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node9334 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node9337 = (inp[5]) ? node9343 : node9338;
														assign node9338 = (inp[15]) ? 4'b1001 : node9339;
															assign node9339 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node9343 = (inp[15]) ? node9347 : node9344;
															assign node9344 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node9347 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node9350 = (inp[5]) ? node9366 : node9351;
													assign node9351 = (inp[14]) ? node9359 : node9352;
														assign node9352 = (inp[0]) ? node9356 : node9353;
															assign node9353 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node9356 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node9359 = (inp[15]) ? node9363 : node9360;
															assign node9360 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node9363 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node9366 = (inp[14]) ? node9374 : node9367;
														assign node9367 = (inp[3]) ? node9371 : node9368;
															assign node9368 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node9371 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node9374 = (inp[0]) ? 4'b1001 : node9375;
															assign node9375 = (inp[3]) ? 4'b1001 : 4'b1001;
											assign node9379 = (inp[14]) ? node9409 : node9380;
												assign node9380 = (inp[2]) ? node9396 : node9381;
													assign node9381 = (inp[0]) ? node9389 : node9382;
														assign node9382 = (inp[15]) ? node9386 : node9383;
															assign node9383 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node9386 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node9389 = (inp[15]) ? node9393 : node9390;
															assign node9390 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node9393 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node9396 = (inp[5]) ? node9402 : node9397;
														assign node9397 = (inp[3]) ? 4'b1000 : node9398;
															assign node9398 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node9402 = (inp[3]) ? node9406 : node9403;
															assign node9403 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node9406 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node9409 = (inp[3]) ? node9425 : node9410;
													assign node9410 = (inp[5]) ? node9418 : node9411;
														assign node9411 = (inp[15]) ? node9415 : node9412;
															assign node9412 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node9415 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node9418 = (inp[0]) ? node9422 : node9419;
															assign node9419 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node9422 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node9425 = (inp[5]) ? node9433 : node9426;
														assign node9426 = (inp[2]) ? node9430 : node9427;
															assign node9427 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node9430 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node9433 = (inp[15]) ? node9437 : node9434;
															assign node9434 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node9437 = (inp[0]) ? 4'b1000 : 4'b1010;
								assign node9440 = (inp[1]) ? node9672 : node9441;
									assign node9441 = (inp[7]) ? node9555 : node9442;
										assign node9442 = (inp[8]) ? node9498 : node9443;
											assign node9443 = (inp[14]) ? node9471 : node9444;
												assign node9444 = (inp[2]) ? node9458 : node9445;
													assign node9445 = (inp[15]) ? node9451 : node9446;
														assign node9446 = (inp[0]) ? node9448 : 4'b0111;
															assign node9448 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node9451 = (inp[0]) ? node9455 : node9452;
															assign node9452 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node9455 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node9458 = (inp[0]) ? node9464 : node9459;
														assign node9459 = (inp[15]) ? 4'b0100 : node9460;
															assign node9460 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node9464 = (inp[15]) ? node9468 : node9465;
															assign node9465 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node9468 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node9471 = (inp[2]) ? node9485 : node9472;
													assign node9472 = (inp[15]) ? node9478 : node9473;
														assign node9473 = (inp[0]) ? node9475 : 4'b0110;
															assign node9475 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node9478 = (inp[0]) ? node9482 : node9479;
															assign node9479 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node9482 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node9485 = (inp[0]) ? node9491 : node9486;
														assign node9486 = (inp[15]) ? 4'b0100 : node9487;
															assign node9487 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node9491 = (inp[15]) ? node9495 : node9492;
															assign node9492 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node9495 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node9498 = (inp[14]) ? node9530 : node9499;
												assign node9499 = (inp[2]) ? node9515 : node9500;
													assign node9500 = (inp[5]) ? node9508 : node9501;
														assign node9501 = (inp[0]) ? node9505 : node9502;
															assign node9502 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node9505 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node9508 = (inp[15]) ? node9512 : node9509;
															assign node9509 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node9512 = (inp[3]) ? 4'b0100 : 4'b0100;
													assign node9515 = (inp[0]) ? node9523 : node9516;
														assign node9516 = (inp[15]) ? node9520 : node9517;
															assign node9517 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node9520 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node9523 = (inp[15]) ? node9527 : node9524;
															assign node9524 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node9527 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node9530 = (inp[3]) ? node9546 : node9531;
													assign node9531 = (inp[5]) ? node9539 : node9532;
														assign node9532 = (inp[2]) ? node9536 : node9533;
															assign node9533 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node9536 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node9539 = (inp[15]) ? node9543 : node9540;
															assign node9540 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node9543 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node9546 = (inp[15]) ? 4'b1001 : node9547;
														assign node9547 = (inp[5]) ? node9551 : node9548;
															assign node9548 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node9551 = (inp[0]) ? 4'b1011 : 4'b1001;
										assign node9555 = (inp[8]) ? node9613 : node9556;
											assign node9556 = (inp[14]) ? node9582 : node9557;
												assign node9557 = (inp[2]) ? node9571 : node9558;
													assign node9558 = (inp[5]) ? node9566 : node9559;
														assign node9559 = (inp[0]) ? node9563 : node9560;
															assign node9560 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node9563 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node9566 = (inp[3]) ? 4'b0110 : node9567;
															assign node9567 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node9571 = (inp[0]) ? node9577 : node9572;
														assign node9572 = (inp[15]) ? node9574 : 4'b1011;
															assign node9574 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node9577 = (inp[15]) ? node9579 : 4'b1001;
															assign node9579 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node9582 = (inp[2]) ? node9598 : node9583;
													assign node9583 = (inp[3]) ? node9591 : node9584;
														assign node9584 = (inp[5]) ? node9588 : node9585;
															assign node9585 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node9588 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node9591 = (inp[15]) ? node9595 : node9592;
															assign node9592 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node9595 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node9598 = (inp[15]) ? node9606 : node9599;
														assign node9599 = (inp[0]) ? node9603 : node9600;
															assign node9600 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node9603 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node9606 = (inp[0]) ? node9610 : node9607;
															assign node9607 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node9610 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node9613 = (inp[14]) ? node9643 : node9614;
												assign node9614 = (inp[2]) ? node9630 : node9615;
													assign node9615 = (inp[3]) ? node9623 : node9616;
														assign node9616 = (inp[15]) ? node9620 : node9617;
															assign node9617 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node9620 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node9623 = (inp[5]) ? node9627 : node9624;
															assign node9624 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node9627 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node9630 = (inp[3]) ? node9638 : node9631;
														assign node9631 = (inp[15]) ? node9635 : node9632;
															assign node9632 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node9635 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node9638 = (inp[0]) ? node9640 : 4'b1010;
															assign node9640 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node9643 = (inp[2]) ? node9659 : node9644;
													assign node9644 = (inp[3]) ? node9652 : node9645;
														assign node9645 = (inp[5]) ? node9649 : node9646;
															assign node9646 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node9649 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node9652 = (inp[15]) ? node9656 : node9653;
															assign node9653 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node9656 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node9659 = (inp[0]) ? node9667 : node9660;
														assign node9660 = (inp[15]) ? node9664 : node9661;
															assign node9661 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node9664 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node9667 = (inp[15]) ? 4'b1010 : node9668;
															assign node9668 = (inp[3]) ? 4'b1010 : 4'b1000;
									assign node9672 = (inp[0]) ? node9776 : node9673;
										assign node9673 = (inp[15]) ? node9727 : node9674;
											assign node9674 = (inp[5]) ? node9698 : node9675;
												assign node9675 = (inp[8]) ? node9687 : node9676;
													assign node9676 = (inp[7]) ? node9682 : node9677;
														assign node9677 = (inp[14]) ? 4'b1010 : node9678;
															assign node9678 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node9682 = (inp[2]) ? 4'b1011 : node9683;
															assign node9683 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node9687 = (inp[7]) ? node9693 : node9688;
														assign node9688 = (inp[2]) ? 4'b1011 : node9689;
															assign node9689 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node9693 = (inp[14]) ? 4'b1010 : node9694;
															assign node9694 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node9698 = (inp[3]) ? node9714 : node9699;
													assign node9699 = (inp[8]) ? node9707 : node9700;
														assign node9700 = (inp[7]) ? node9704 : node9701;
															assign node9701 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node9704 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node9707 = (inp[7]) ? node9711 : node9708;
															assign node9708 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node9711 = (inp[14]) ? 4'b1010 : 4'b1010;
													assign node9714 = (inp[7]) ? node9722 : node9715;
														assign node9715 = (inp[8]) ? node9719 : node9716;
															assign node9716 = (inp[2]) ? 4'b1000 : 4'b1000;
															assign node9719 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node9722 = (inp[8]) ? node9724 : 4'b1001;
															assign node9724 = (inp[14]) ? 4'b1000 : 4'b1000;
											assign node9727 = (inp[5]) ? node9747 : node9728;
												assign node9728 = (inp[7]) ? node9740 : node9729;
													assign node9729 = (inp[8]) ? node9735 : node9730;
														assign node9730 = (inp[2]) ? 4'b1000 : node9731;
															assign node9731 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node9735 = (inp[2]) ? 4'b1001 : node9736;
															assign node9736 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node9740 = (inp[8]) ? node9742 : 4'b1001;
														assign node9742 = (inp[2]) ? 4'b1000 : node9743;
															assign node9743 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node9747 = (inp[3]) ? node9761 : node9748;
													assign node9748 = (inp[2]) ? node9754 : node9749;
														assign node9749 = (inp[14]) ? 4'b1001 : node9750;
															assign node9750 = (inp[7]) ? 4'b1000 : 4'b1000;
														assign node9754 = (inp[7]) ? node9758 : node9755;
															assign node9755 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node9758 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node9761 = (inp[14]) ? node9769 : node9762;
														assign node9762 = (inp[2]) ? node9766 : node9763;
															assign node9763 = (inp[8]) ? 4'b1010 : 4'b1010;
															assign node9766 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node9769 = (inp[2]) ? node9773 : node9770;
															assign node9770 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node9773 = (inp[7]) ? 4'b1010 : 4'b1010;
										assign node9776 = (inp[15]) ? node9838 : node9777;
											assign node9777 = (inp[5]) ? node9809 : node9778;
												assign node9778 = (inp[2]) ? node9794 : node9779;
													assign node9779 = (inp[8]) ? node9787 : node9780;
														assign node9780 = (inp[14]) ? node9784 : node9781;
															assign node9781 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node9784 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node9787 = (inp[3]) ? node9791 : node9788;
															assign node9788 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node9791 = (inp[14]) ? 4'b1000 : 4'b1000;
													assign node9794 = (inp[3]) ? node9802 : node9795;
														assign node9795 = (inp[14]) ? node9799 : node9796;
															assign node9796 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node9799 = (inp[7]) ? 4'b1000 : 4'b1000;
														assign node9802 = (inp[8]) ? node9806 : node9803;
															assign node9803 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node9806 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node9809 = (inp[3]) ? node9823 : node9810;
													assign node9810 = (inp[14]) ? node9816 : node9811;
														assign node9811 = (inp[8]) ? node9813 : 4'b1000;
															assign node9813 = (inp[2]) ? 4'b1000 : 4'b1000;
														assign node9816 = (inp[2]) ? node9820 : node9817;
															assign node9817 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node9820 = (inp[7]) ? 4'b1000 : 4'b1000;
													assign node9823 = (inp[14]) ? node9831 : node9824;
														assign node9824 = (inp[7]) ? node9828 : node9825;
															assign node9825 = (inp[2]) ? 4'b1010 : 4'b1010;
															assign node9828 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node9831 = (inp[7]) ? node9835 : node9832;
															assign node9832 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node9835 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node9838 = (inp[3]) ? node9862 : node9839;
												assign node9839 = (inp[7]) ? node9851 : node9840;
													assign node9840 = (inp[8]) ? node9846 : node9841;
														assign node9841 = (inp[14]) ? 4'b1010 : node9842;
															assign node9842 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node9846 = (inp[14]) ? 4'b1011 : node9847;
															assign node9847 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node9851 = (inp[8]) ? node9857 : node9852;
														assign node9852 = (inp[2]) ? 4'b1011 : node9853;
															assign node9853 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node9857 = (inp[2]) ? 4'b1010 : node9858;
															assign node9858 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node9862 = (inp[5]) ? node9876 : node9863;
													assign node9863 = (inp[14]) ? node9871 : node9864;
														assign node9864 = (inp[7]) ? node9868 : node9865;
															assign node9865 = (inp[2]) ? 4'b1010 : 4'b1010;
															assign node9868 = (inp[2]) ? 4'b1010 : 4'b1010;
														assign node9871 = (inp[8]) ? 4'b1010 : node9872;
															assign node9872 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node9876 = (inp[2]) ? node9884 : node9877;
														assign node9877 = (inp[8]) ? node9881 : node9878;
															assign node9878 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node9881 = (inp[14]) ? 4'b1000 : 4'b1000;
														assign node9884 = (inp[14]) ? node9888 : node9885;
															assign node9885 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node9888 = (inp[7]) ? 4'b1000 : 4'b1000;
							assign node9891 = (inp[13]) ? node10345 : node9892;
								assign node9892 = (inp[1]) ? node10124 : node9893;
									assign node9893 = (inp[7]) ? node10011 : node9894;
										assign node9894 = (inp[8]) ? node9948 : node9895;
											assign node9895 = (inp[2]) ? node9925 : node9896;
												assign node9896 = (inp[14]) ? node9910 : node9897;
													assign node9897 = (inp[3]) ? node9903 : node9898;
														assign node9898 = (inp[15]) ? node9900 : 4'b1011;
															assign node9900 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node9903 = (inp[0]) ? node9907 : node9904;
															assign node9904 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node9907 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node9910 = (inp[5]) ? node9918 : node9911;
														assign node9911 = (inp[0]) ? node9915 : node9912;
															assign node9912 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node9915 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node9918 = (inp[0]) ? node9922 : node9919;
															assign node9919 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node9922 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node9925 = (inp[0]) ? node9937 : node9926;
													assign node9926 = (inp[15]) ? node9932 : node9927;
														assign node9927 = (inp[5]) ? node9929 : 4'b1010;
															assign node9929 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node9932 = (inp[3]) ? node9934 : 4'b1000;
															assign node9934 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node9937 = (inp[15]) ? node9943 : node9938;
														assign node9938 = (inp[3]) ? node9940 : 4'b1000;
															assign node9940 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node9943 = (inp[3]) ? node9945 : 4'b1010;
															assign node9945 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node9948 = (inp[14]) ? node9980 : node9949;
												assign node9949 = (inp[2]) ? node9965 : node9950;
													assign node9950 = (inp[3]) ? node9958 : node9951;
														assign node9951 = (inp[5]) ? node9955 : node9952;
															assign node9952 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node9955 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node9958 = (inp[0]) ? node9962 : node9959;
															assign node9959 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node9962 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node9965 = (inp[0]) ? node9973 : node9966;
														assign node9966 = (inp[15]) ? node9970 : node9967;
															assign node9967 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node9970 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node9973 = (inp[15]) ? node9977 : node9974;
															assign node9974 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node9977 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node9980 = (inp[5]) ? node9996 : node9981;
													assign node9981 = (inp[3]) ? node9989 : node9982;
														assign node9982 = (inp[0]) ? node9986 : node9983;
															assign node9983 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node9986 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node9989 = (inp[2]) ? node9993 : node9990;
															assign node9990 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node9993 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node9996 = (inp[0]) ? node10004 : node9997;
														assign node9997 = (inp[2]) ? node10001 : node9998;
															assign node9998 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node10001 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node10004 = (inp[2]) ? node10008 : node10005;
															assign node10005 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node10008 = (inp[3]) ? 4'b1011 : 4'b1001;
										assign node10011 = (inp[8]) ? node10067 : node10012;
											assign node10012 = (inp[14]) ? node10044 : node10013;
												assign node10013 = (inp[2]) ? node10029 : node10014;
													assign node10014 = (inp[0]) ? node10022 : node10015;
														assign node10015 = (inp[15]) ? node10019 : node10016;
															assign node10016 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node10019 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node10022 = (inp[15]) ? node10026 : node10023;
															assign node10023 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node10026 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node10029 = (inp[5]) ? node10037 : node10030;
														assign node10030 = (inp[3]) ? node10034 : node10031;
															assign node10031 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node10034 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node10037 = (inp[3]) ? node10041 : node10038;
															assign node10038 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node10041 = (inp[15]) ? 4'b1001 : 4'b1001;
												assign node10044 = (inp[3]) ? node10052 : node10045;
													assign node10045 = (inp[0]) ? node10049 : node10046;
														assign node10046 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node10049 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node10052 = (inp[5]) ? node10060 : node10053;
														assign node10053 = (inp[2]) ? node10057 : node10054;
															assign node10054 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node10057 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node10060 = (inp[15]) ? node10064 : node10061;
															assign node10061 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node10064 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node10067 = (inp[14]) ? node10095 : node10068;
												assign node10068 = (inp[2]) ? node10082 : node10069;
													assign node10069 = (inp[3]) ? node10077 : node10070;
														assign node10070 = (inp[15]) ? node10074 : node10071;
															assign node10071 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node10074 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node10077 = (inp[0]) ? node10079 : 4'b1011;
															assign node10079 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node10082 = (inp[3]) ? node10088 : node10083;
														assign node10083 = (inp[5]) ? node10085 : 4'b1000;
															assign node10085 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node10088 = (inp[0]) ? node10092 : node10089;
															assign node10089 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node10092 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node10095 = (inp[2]) ? node10111 : node10096;
													assign node10096 = (inp[0]) ? node10104 : node10097;
														assign node10097 = (inp[15]) ? node10101 : node10098;
															assign node10098 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node10101 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node10104 = (inp[15]) ? node10108 : node10105;
															assign node10105 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node10108 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node10111 = (inp[5]) ? node10119 : node10112;
														assign node10112 = (inp[3]) ? node10116 : node10113;
															assign node10113 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node10116 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node10119 = (inp[3]) ? node10121 : 4'b1000;
															assign node10121 = (inp[15]) ? 4'b1000 : 4'b1000;
									assign node10124 = (inp[7]) ? node10230 : node10125;
										assign node10125 = (inp[8]) ? node10179 : node10126;
											assign node10126 = (inp[2]) ? node10156 : node10127;
												assign node10127 = (inp[14]) ? node10143 : node10128;
													assign node10128 = (inp[5]) ? node10136 : node10129;
														assign node10129 = (inp[0]) ? node10133 : node10130;
															assign node10130 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node10133 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node10136 = (inp[15]) ? node10140 : node10137;
															assign node10137 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node10140 = (inp[3]) ? 4'b1001 : 4'b1001;
													assign node10143 = (inp[15]) ? node10149 : node10144;
														assign node10144 = (inp[3]) ? node10146 : 4'b1000;
															assign node10146 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node10149 = (inp[0]) ? node10153 : node10150;
															assign node10150 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node10153 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node10156 = (inp[0]) ? node10168 : node10157;
													assign node10157 = (inp[15]) ? node10163 : node10158;
														assign node10158 = (inp[5]) ? node10160 : 4'b1010;
															assign node10160 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node10163 = (inp[5]) ? node10165 : 4'b1000;
															assign node10165 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node10168 = (inp[15]) ? node10174 : node10169;
														assign node10169 = (inp[5]) ? node10171 : 4'b1000;
															assign node10171 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node10174 = (inp[5]) ? node10176 : 4'b1010;
															assign node10176 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node10179 = (inp[14]) ? node10209 : node10180;
												assign node10180 = (inp[2]) ? node10194 : node10181;
													assign node10181 = (inp[0]) ? node10187 : node10182;
														assign node10182 = (inp[3]) ? node10184 : 4'b1000;
															assign node10184 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node10187 = (inp[15]) ? node10191 : node10188;
															assign node10188 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node10191 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node10194 = (inp[5]) ? node10202 : node10195;
														assign node10195 = (inp[15]) ? node10199 : node10196;
															assign node10196 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node10199 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node10202 = (inp[3]) ? node10206 : node10203;
															assign node10203 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node10206 = (inp[0]) ? 4'b0001 : 4'b0001;
												assign node10209 = (inp[5]) ? node10217 : node10210;
													assign node10210 = (inp[0]) ? node10214 : node10211;
														assign node10211 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node10214 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node10217 = (inp[3]) ? node10225 : node10218;
														assign node10218 = (inp[15]) ? node10222 : node10219;
															assign node10219 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node10222 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node10225 = (inp[2]) ? 4'b0001 : node10226;
															assign node10226 = (inp[0]) ? 4'b0001 : 4'b0001;
										assign node10230 = (inp[8]) ? node10288 : node10231;
											assign node10231 = (inp[14]) ? node10259 : node10232;
												assign node10232 = (inp[2]) ? node10246 : node10233;
													assign node10233 = (inp[3]) ? node10241 : node10234;
														assign node10234 = (inp[0]) ? node10238 : node10235;
															assign node10235 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node10238 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node10241 = (inp[0]) ? node10243 : 4'b1000;
															assign node10243 = (inp[5]) ? 4'b1000 : 4'b1000;
													assign node10246 = (inp[5]) ? node10252 : node10247;
														assign node10247 = (inp[3]) ? 4'b0011 : node10248;
															assign node10248 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node10252 = (inp[15]) ? node10256 : node10253;
															assign node10253 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node10256 = (inp[0]) ? 4'b0001 : 4'b0001;
												assign node10259 = (inp[2]) ? node10275 : node10260;
													assign node10260 = (inp[0]) ? node10268 : node10261;
														assign node10261 = (inp[15]) ? node10265 : node10262;
															assign node10262 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node10265 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node10268 = (inp[15]) ? node10272 : node10269;
															assign node10269 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node10272 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node10275 = (inp[0]) ? node10281 : node10276;
														assign node10276 = (inp[15]) ? node10278 : 4'b0011;
															assign node10278 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node10281 = (inp[15]) ? node10285 : node10282;
															assign node10282 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node10285 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node10288 = (inp[14]) ? node10316 : node10289;
												assign node10289 = (inp[2]) ? node10303 : node10290;
													assign node10290 = (inp[0]) ? node10298 : node10291;
														assign node10291 = (inp[15]) ? node10295 : node10292;
															assign node10292 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node10295 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node10298 = (inp[15]) ? 4'b0011 : node10299;
															assign node10299 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node10303 = (inp[3]) ? node10309 : node10304;
														assign node10304 = (inp[5]) ? 4'b0000 : node10305;
															assign node10305 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node10309 = (inp[0]) ? node10313 : node10310;
															assign node10310 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node10313 = (inp[15]) ? 4'b0000 : 4'b0000;
												assign node10316 = (inp[3]) ? node10332 : node10317;
													assign node10317 = (inp[5]) ? node10325 : node10318;
														assign node10318 = (inp[2]) ? node10322 : node10319;
															assign node10319 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node10322 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node10325 = (inp[0]) ? node10329 : node10326;
															assign node10326 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node10329 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node10332 = (inp[5]) ? node10340 : node10333;
														assign node10333 = (inp[15]) ? node10337 : node10334;
															assign node10334 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node10337 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node10340 = (inp[2]) ? 4'b0010 : node10341;
															assign node10341 = (inp[0]) ? 4'b0000 : 4'b0000;
								assign node10345 = (inp[1]) ? node10559 : node10346;
									assign node10346 = (inp[8]) ? node10452 : node10347;
										assign node10347 = (inp[7]) ? node10391 : node10348;
											assign node10348 = (inp[2]) ? node10372 : node10349;
												assign node10349 = (inp[14]) ? node10361 : node10350;
													assign node10350 = (inp[5]) ? node10356 : node10351;
														assign node10351 = (inp[3]) ? 4'b1001 : node10352;
															assign node10352 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node10356 = (inp[3]) ? 4'b1011 : node10357;
															assign node10357 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node10361 = (inp[0]) ? node10367 : node10362;
														assign node10362 = (inp[15]) ? node10364 : 4'b1010;
															assign node10364 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node10367 = (inp[15]) ? node10369 : 4'b1000;
															assign node10369 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node10372 = (inp[15]) ? node10380 : node10373;
													assign node10373 = (inp[0]) ? node10375 : 4'b1010;
														assign node10375 = (inp[5]) ? node10377 : 4'b1000;
															assign node10377 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node10380 = (inp[0]) ? node10386 : node10381;
														assign node10381 = (inp[3]) ? node10383 : 4'b1000;
															assign node10383 = (inp[14]) ? 4'b1010 : 4'b1000;
														assign node10386 = (inp[3]) ? node10388 : 4'b1010;
															assign node10388 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node10391 = (inp[2]) ? node10423 : node10392;
												assign node10392 = (inp[14]) ? node10408 : node10393;
													assign node10393 = (inp[15]) ? node10401 : node10394;
														assign node10394 = (inp[0]) ? node10398 : node10395;
															assign node10395 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node10398 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node10401 = (inp[0]) ? node10405 : node10402;
															assign node10402 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node10405 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node10408 = (inp[5]) ? node10416 : node10409;
														assign node10409 = (inp[3]) ? node10413 : node10410;
															assign node10410 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node10413 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node10416 = (inp[15]) ? node10420 : node10417;
															assign node10417 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node10420 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node10423 = (inp[5]) ? node10439 : node10424;
													assign node10424 = (inp[3]) ? node10432 : node10425;
														assign node10425 = (inp[15]) ? node10429 : node10426;
															assign node10426 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node10429 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node10432 = (inp[15]) ? node10436 : node10433;
															assign node10433 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node10436 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node10439 = (inp[14]) ? node10447 : node10440;
														assign node10440 = (inp[3]) ? node10444 : node10441;
															assign node10441 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node10444 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node10447 = (inp[15]) ? node10449 : 4'b0011;
															assign node10449 = (inp[3]) ? 4'b0001 : 4'b0001;
										assign node10452 = (inp[7]) ? node10504 : node10453;
											assign node10453 = (inp[2]) ? node10481 : node10454;
												assign node10454 = (inp[14]) ? node10470 : node10455;
													assign node10455 = (inp[3]) ? node10463 : node10456;
														assign node10456 = (inp[5]) ? node10460 : node10457;
															assign node10457 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node10460 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node10463 = (inp[15]) ? node10467 : node10464;
															assign node10464 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node10467 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node10470 = (inp[0]) ? node10476 : node10471;
														assign node10471 = (inp[15]) ? 4'b0001 : node10472;
															assign node10472 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node10476 = (inp[15]) ? 4'b0011 : node10477;
															assign node10477 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node10481 = (inp[0]) ? node10493 : node10482;
													assign node10482 = (inp[15]) ? node10488 : node10483;
														assign node10483 = (inp[5]) ? node10485 : 4'b0011;
															assign node10485 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node10488 = (inp[5]) ? node10490 : 4'b0001;
															assign node10490 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node10493 = (inp[15]) ? node10499 : node10494;
														assign node10494 = (inp[5]) ? node10496 : 4'b0001;
															assign node10496 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node10499 = (inp[5]) ? node10501 : 4'b0011;
															assign node10501 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node10504 = (inp[2]) ? node10532 : node10505;
												assign node10505 = (inp[14]) ? node10521 : node10506;
													assign node10506 = (inp[3]) ? node10514 : node10507;
														assign node10507 = (inp[15]) ? node10511 : node10508;
															assign node10508 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node10511 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node10514 = (inp[0]) ? node10518 : node10515;
															assign node10515 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node10518 = (inp[5]) ? 4'b0001 : 4'b0001;
													assign node10521 = (inp[0]) ? node10527 : node10522;
														assign node10522 = (inp[15]) ? 4'b0000 : node10523;
															assign node10523 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node10527 = (inp[15]) ? 4'b0010 : node10528;
															assign node10528 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node10532 = (inp[14]) ? node10546 : node10533;
													assign node10533 = (inp[0]) ? node10539 : node10534;
														assign node10534 = (inp[15]) ? 4'b0000 : node10535;
															assign node10535 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node10539 = (inp[15]) ? node10543 : node10540;
															assign node10540 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node10543 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node10546 = (inp[0]) ? node10554 : node10547;
														assign node10547 = (inp[15]) ? node10551 : node10548;
															assign node10548 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node10551 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node10554 = (inp[15]) ? node10556 : 4'b0000;
															assign node10556 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node10559 = (inp[2]) ? node10687 : node10560;
										assign node10560 = (inp[0]) ? node10624 : node10561;
											assign node10561 = (inp[15]) ? node10593 : node10562;
												assign node10562 = (inp[5]) ? node10578 : node10563;
													assign node10563 = (inp[3]) ? node10571 : node10564;
														assign node10564 = (inp[7]) ? node10568 : node10565;
															assign node10565 = (inp[14]) ? 4'b0010 : 4'b0010;
															assign node10568 = (inp[14]) ? 4'b0010 : 4'b0010;
														assign node10571 = (inp[8]) ? node10575 : node10572;
															assign node10572 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node10575 = (inp[7]) ? 4'b0010 : 4'b0010;
													assign node10578 = (inp[3]) ? node10586 : node10579;
														assign node10579 = (inp[14]) ? node10583 : node10580;
															assign node10580 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node10583 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node10586 = (inp[14]) ? node10590 : node10587;
															assign node10587 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node10590 = (inp[7]) ? 4'b0000 : 4'b0000;
												assign node10593 = (inp[5]) ? node10609 : node10594;
													assign node10594 = (inp[3]) ? node10602 : node10595;
														assign node10595 = (inp[14]) ? node10599 : node10596;
															assign node10596 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node10599 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node10602 = (inp[14]) ? node10606 : node10603;
															assign node10603 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node10606 = (inp[8]) ? 4'b0000 : 4'b0000;
													assign node10609 = (inp[3]) ? node10617 : node10610;
														assign node10610 = (inp[8]) ? node10614 : node10611;
															assign node10611 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node10614 = (inp[14]) ? 4'b0000 : 4'b0000;
														assign node10617 = (inp[14]) ? node10621 : node10618;
															assign node10618 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node10621 = (inp[8]) ? 4'b0010 : 4'b0010;
											assign node10624 = (inp[15]) ? node10656 : node10625;
												assign node10625 = (inp[5]) ? node10641 : node10626;
													assign node10626 = (inp[14]) ? node10634 : node10627;
														assign node10627 = (inp[7]) ? node10631 : node10628;
															assign node10628 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node10631 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node10634 = (inp[7]) ? node10638 : node10635;
															assign node10635 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node10638 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node10641 = (inp[3]) ? node10649 : node10642;
														assign node10642 = (inp[7]) ? node10646 : node10643;
															assign node10643 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node10646 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node10649 = (inp[7]) ? node10653 : node10650;
															assign node10650 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node10653 = (inp[14]) ? 4'b0010 : 4'b0010;
												assign node10656 = (inp[3]) ? node10672 : node10657;
													assign node10657 = (inp[14]) ? node10665 : node10658;
														assign node10658 = (inp[8]) ? node10662 : node10659;
															assign node10659 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node10662 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node10665 = (inp[7]) ? node10669 : node10666;
															assign node10666 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node10669 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node10672 = (inp[5]) ? node10680 : node10673;
														assign node10673 = (inp[7]) ? node10677 : node10674;
															assign node10674 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node10677 = (inp[14]) ? 4'b0010 : 4'b0010;
														assign node10680 = (inp[14]) ? node10684 : node10681;
															assign node10681 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node10684 = (inp[7]) ? 4'b0000 : 4'b0000;
										assign node10687 = (inp[15]) ? node10731 : node10688;
											assign node10688 = (inp[0]) ? node10710 : node10689;
												assign node10689 = (inp[5]) ? node10697 : node10690;
													assign node10690 = (inp[8]) ? node10694 : node10691;
														assign node10691 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node10694 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node10697 = (inp[3]) ? node10703 : node10698;
														assign node10698 = (inp[14]) ? node10700 : 4'b0010;
															assign node10700 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node10703 = (inp[7]) ? node10707 : node10704;
															assign node10704 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node10707 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node10710 = (inp[3]) ? node10718 : node10711;
													assign node10711 = (inp[8]) ? node10715 : node10712;
														assign node10712 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node10715 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node10718 = (inp[5]) ? node10726 : node10719;
														assign node10719 = (inp[14]) ? node10723 : node10720;
															assign node10720 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node10723 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node10726 = (inp[14]) ? node10728 : 4'b0011;
															assign node10728 = (inp[7]) ? 4'b0010 : 4'b0010;
											assign node10731 = (inp[0]) ? node10755 : node10732;
												assign node10732 = (inp[5]) ? node10740 : node10733;
													assign node10733 = (inp[8]) ? node10737 : node10734;
														assign node10734 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node10737 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node10740 = (inp[3]) ? node10748 : node10741;
														assign node10741 = (inp[7]) ? node10745 : node10742;
															assign node10742 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node10745 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node10748 = (inp[14]) ? node10752 : node10749;
															assign node10749 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node10752 = (inp[8]) ? 4'b0010 : 4'b0010;
												assign node10755 = (inp[3]) ? node10763 : node10756;
													assign node10756 = (inp[7]) ? node10760 : node10757;
														assign node10757 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node10760 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node10763 = (inp[5]) ? node10771 : node10764;
														assign node10764 = (inp[7]) ? node10768 : node10765;
															assign node10765 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node10768 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node10771 = (inp[7]) ? node10775 : node10772;
															assign node10772 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node10775 = (inp[8]) ? 4'b0000 : 4'b0001;
					assign node10778 = (inp[3]) ? node12338 : node10779;
						assign node10779 = (inp[2]) ? node11717 : node10780;
							assign node10780 = (inp[1]) ? node11222 : node10781;
								assign node10781 = (inp[7]) ? node10979 : node10782;
									assign node10782 = (inp[11]) ? node10888 : node10783;
										assign node10783 = (inp[6]) ? node10845 : node10784;
											assign node10784 = (inp[13]) ? node10816 : node10785;
												assign node10785 = (inp[14]) ? node10801 : node10786;
													assign node10786 = (inp[8]) ? node10794 : node10787;
														assign node10787 = (inp[5]) ? node10791 : node10788;
															assign node10788 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node10791 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node10794 = (inp[15]) ? node10798 : node10795;
															assign node10795 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node10798 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node10801 = (inp[8]) ? node10809 : node10802;
														assign node10802 = (inp[15]) ? node10806 : node10803;
															assign node10803 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node10806 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node10809 = (inp[0]) ? node10813 : node10810;
															assign node10810 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node10813 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node10816 = (inp[14]) ? node10832 : node10817;
													assign node10817 = (inp[8]) ? node10825 : node10818;
														assign node10818 = (inp[5]) ? node10822 : node10819;
															assign node10819 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node10822 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node10825 = (inp[0]) ? node10829 : node10826;
															assign node10826 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node10829 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node10832 = (inp[8]) ? node10838 : node10833;
														assign node10833 = (inp[0]) ? node10835 : 4'b1000;
															assign node10835 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node10838 = (inp[15]) ? node10842 : node10839;
															assign node10839 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node10842 = (inp[0]) ? 4'b0011 : 4'b0001;
											assign node10845 = (inp[14]) ? node10865 : node10846;
												assign node10846 = (inp[8]) ? node10858 : node10847;
													assign node10847 = (inp[5]) ? node10853 : node10848;
														assign node10848 = (inp[13]) ? node10850 : 4'b0001;
															assign node10850 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node10853 = (inp[13]) ? node10855 : 4'b0011;
															assign node10855 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node10858 = (inp[0]) ? node10862 : node10859;
														assign node10859 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node10862 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node10865 = (inp[8]) ? node10873 : node10866;
													assign node10866 = (inp[0]) ? node10870 : node10867;
														assign node10867 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node10870 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node10873 = (inp[13]) ? node10881 : node10874;
														assign node10874 = (inp[0]) ? node10878 : node10875;
															assign node10875 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node10878 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node10881 = (inp[5]) ? node10885 : node10882;
															assign node10882 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node10885 = (inp[15]) ? 4'b1001 : 4'b1001;
										assign node10888 = (inp[6]) ? node10926 : node10889;
											assign node10889 = (inp[14]) ? node10905 : node10890;
												assign node10890 = (inp[8]) ? node10898 : node10891;
													assign node10891 = (inp[15]) ? node10895 : node10892;
														assign node10892 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node10895 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node10898 = (inp[0]) ? node10902 : node10899;
														assign node10899 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node10902 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node10905 = (inp[8]) ? node10913 : node10906;
													assign node10906 = (inp[15]) ? node10910 : node10907;
														assign node10907 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node10910 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node10913 = (inp[13]) ? node10921 : node10914;
														assign node10914 = (inp[15]) ? node10918 : node10915;
															assign node10915 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node10918 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node10921 = (inp[5]) ? node10923 : 4'b1011;
															assign node10923 = (inp[0]) ? 4'b1001 : 4'b1001;
											assign node10926 = (inp[14]) ? node10956 : node10927;
												assign node10927 = (inp[8]) ? node10941 : node10928;
													assign node10928 = (inp[5]) ? node10936 : node10929;
														assign node10929 = (inp[15]) ? node10933 : node10930;
															assign node10930 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node10933 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node10936 = (inp[15]) ? node10938 : 4'b1001;
															assign node10938 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node10941 = (inp[5]) ? node10949 : node10942;
														assign node10942 = (inp[13]) ? node10946 : node10943;
															assign node10943 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node10946 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node10949 = (inp[13]) ? node10953 : node10950;
															assign node10950 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node10953 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node10956 = (inp[8]) ? node10964 : node10957;
													assign node10957 = (inp[0]) ? node10961 : node10958;
														assign node10958 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node10961 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node10964 = (inp[13]) ? node10972 : node10965;
														assign node10965 = (inp[0]) ? node10969 : node10966;
															assign node10966 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node10969 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node10972 = (inp[5]) ? node10976 : node10973;
															assign node10973 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node10976 = (inp[15]) ? 4'b0001 : 4'b0001;
									assign node10979 = (inp[5]) ? node11103 : node10980;
										assign node10980 = (inp[15]) ? node11044 : node10981;
											assign node10981 = (inp[0]) ? node11013 : node10982;
												assign node10982 = (inp[8]) ? node10998 : node10983;
													assign node10983 = (inp[14]) ? node10991 : node10984;
														assign node10984 = (inp[13]) ? node10988 : node10985;
															assign node10985 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node10988 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node10991 = (inp[6]) ? node10995 : node10992;
															assign node10992 = (inp[13]) ? 4'b0011 : 4'b0011;
															assign node10995 = (inp[11]) ? 4'b0011 : 4'b0011;
													assign node10998 = (inp[14]) ? node11006 : node10999;
														assign node10999 = (inp[13]) ? node11003 : node11000;
															assign node11000 = (inp[6]) ? 4'b0011 : 4'b1011;
															assign node11003 = (inp[11]) ? 4'b0011 : 4'b0011;
														assign node11006 = (inp[11]) ? node11010 : node11007;
															assign node11007 = (inp[13]) ? 4'b0010 : 4'b0010;
															assign node11010 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node11013 = (inp[6]) ? node11029 : node11014;
													assign node11014 = (inp[11]) ? node11022 : node11015;
														assign node11015 = (inp[13]) ? node11019 : node11016;
															assign node11016 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node11019 = (inp[14]) ? 4'b0000 : 4'b0000;
														assign node11022 = (inp[13]) ? node11026 : node11023;
															assign node11023 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node11026 = (inp[8]) ? 4'b1000 : 4'b0000;
													assign node11029 = (inp[11]) ? node11037 : node11030;
														assign node11030 = (inp[13]) ? node11034 : node11031;
															assign node11031 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node11034 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node11037 = (inp[13]) ? node11041 : node11038;
															assign node11038 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node11041 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node11044 = (inp[0]) ? node11074 : node11045;
												assign node11045 = (inp[8]) ? node11059 : node11046;
													assign node11046 = (inp[14]) ? node11054 : node11047;
														assign node11047 = (inp[13]) ? node11051 : node11048;
															assign node11048 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node11051 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node11054 = (inp[11]) ? 4'b0001 : node11055;
															assign node11055 = (inp[6]) ? 4'b0001 : 4'b0001;
													assign node11059 = (inp[14]) ? node11067 : node11060;
														assign node11060 = (inp[6]) ? node11064 : node11061;
															assign node11061 = (inp[11]) ? 4'b0001 : 4'b0001;
															assign node11064 = (inp[13]) ? 4'b0001 : 4'b0001;
														assign node11067 = (inp[6]) ? node11071 : node11068;
															assign node11068 = (inp[13]) ? 4'b0000 : 4'b0000;
															assign node11071 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node11074 = (inp[13]) ? node11090 : node11075;
													assign node11075 = (inp[6]) ? node11083 : node11076;
														assign node11076 = (inp[11]) ? node11080 : node11077;
															assign node11077 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node11080 = (inp[8]) ? 4'b0010 : 4'b0010;
														assign node11083 = (inp[11]) ? node11087 : node11084;
															assign node11084 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node11087 = (inp[8]) ? 4'b1010 : 4'b1010;
													assign node11090 = (inp[14]) ? node11098 : node11091;
														assign node11091 = (inp[8]) ? node11095 : node11092;
															assign node11092 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node11095 = (inp[11]) ? 4'b0011 : 4'b0011;
														assign node11098 = (inp[8]) ? node11100 : 4'b0011;
															assign node11100 = (inp[6]) ? 4'b0010 : 4'b0010;
										assign node11103 = (inp[11]) ? node11163 : node11104;
											assign node11104 = (inp[6]) ? node11132 : node11105;
												assign node11105 = (inp[13]) ? node11119 : node11106;
													assign node11106 = (inp[14]) ? node11112 : node11107;
														assign node11107 = (inp[8]) ? node11109 : 4'b1010;
															assign node11109 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node11112 = (inp[8]) ? node11116 : node11113;
															assign node11113 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node11116 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node11119 = (inp[8]) ? node11127 : node11120;
														assign node11120 = (inp[14]) ? node11124 : node11121;
															assign node11121 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node11124 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node11127 = (inp[14]) ? 4'b0010 : node11128;
															assign node11128 = (inp[15]) ? 4'b0001 : 4'b0001;
												assign node11132 = (inp[13]) ? node11148 : node11133;
													assign node11133 = (inp[0]) ? node11141 : node11134;
														assign node11134 = (inp[15]) ? node11138 : node11135;
															assign node11135 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node11138 = (inp[14]) ? 4'b0000 : 4'b0000;
														assign node11141 = (inp[15]) ? node11145 : node11142;
															assign node11142 = (inp[14]) ? 4'b0000 : 4'b0000;
															assign node11145 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node11148 = (inp[14]) ? node11156 : node11149;
														assign node11149 = (inp[8]) ? node11153 : node11150;
															assign node11150 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node11153 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node11156 = (inp[8]) ? node11160 : node11157;
															assign node11157 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node11160 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node11163 = (inp[6]) ? node11193 : node11164;
												assign node11164 = (inp[13]) ? node11180 : node11165;
													assign node11165 = (inp[8]) ? node11173 : node11166;
														assign node11166 = (inp[14]) ? node11170 : node11167;
															assign node11167 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node11170 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node11173 = (inp[14]) ? node11177 : node11174;
															assign node11174 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node11177 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node11180 = (inp[8]) ? node11188 : node11181;
														assign node11181 = (inp[14]) ? node11185 : node11182;
															assign node11182 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node11185 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node11188 = (inp[14]) ? 4'b1000 : node11189;
															assign node11189 = (inp[0]) ? 4'b1001 : 4'b1001;
												assign node11193 = (inp[13]) ? node11209 : node11194;
													assign node11194 = (inp[8]) ? node11202 : node11195;
														assign node11195 = (inp[14]) ? node11199 : node11196;
															assign node11196 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node11199 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node11202 = (inp[14]) ? node11206 : node11203;
															assign node11203 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node11206 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node11209 = (inp[8]) ? node11215 : node11210;
														assign node11210 = (inp[14]) ? node11212 : 4'b1010;
															assign node11212 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node11215 = (inp[14]) ? node11219 : node11216;
															assign node11216 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node11219 = (inp[15]) ? 4'b0000 : 4'b0000;
								assign node11222 = (inp[13]) ? node11472 : node11223;
									assign node11223 = (inp[0]) ? node11351 : node11224;
										assign node11224 = (inp[15]) ? node11288 : node11225;
											assign node11225 = (inp[7]) ? node11257 : node11226;
												assign node11226 = (inp[14]) ? node11242 : node11227;
													assign node11227 = (inp[8]) ? node11235 : node11228;
														assign node11228 = (inp[11]) ? node11232 : node11229;
															assign node11229 = (inp[6]) ? 4'b0011 : 4'b1011;
															assign node11232 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node11235 = (inp[6]) ? node11239 : node11236;
															assign node11236 = (inp[11]) ? 4'b0010 : 4'b1010;
															assign node11239 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node11242 = (inp[8]) ? node11250 : node11243;
														assign node11243 = (inp[11]) ? node11247 : node11244;
															assign node11244 = (inp[6]) ? 4'b0010 : 4'b1010;
															assign node11247 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node11250 = (inp[5]) ? node11254 : node11251;
															assign node11251 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node11254 = (inp[6]) ? 4'b0011 : 4'b0011;
												assign node11257 = (inp[14]) ? node11273 : node11258;
													assign node11258 = (inp[8]) ? node11266 : node11259;
														assign node11259 = (inp[5]) ? node11263 : node11260;
															assign node11260 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node11263 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node11266 = (inp[5]) ? node11270 : node11267;
															assign node11267 = (inp[11]) ? 4'b0011 : 4'b0011;
															assign node11270 = (inp[11]) ? 4'b0011 : 4'b0011;
													assign node11273 = (inp[8]) ? node11281 : node11274;
														assign node11274 = (inp[6]) ? node11278 : node11275;
															assign node11275 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node11278 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node11281 = (inp[11]) ? node11285 : node11282;
															assign node11282 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node11285 = (inp[6]) ? 4'b0010 : 4'b1010;
											assign node11288 = (inp[11]) ? node11320 : node11289;
												assign node11289 = (inp[8]) ? node11305 : node11290;
													assign node11290 = (inp[6]) ? node11298 : node11291;
														assign node11291 = (inp[14]) ? node11295 : node11292;
															assign node11292 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node11295 = (inp[7]) ? 4'b0001 : 4'b1000;
														assign node11298 = (inp[7]) ? node11302 : node11299;
															assign node11299 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node11302 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node11305 = (inp[6]) ? node11313 : node11306;
														assign node11306 = (inp[7]) ? node11310 : node11307;
															assign node11307 = (inp[14]) ? 4'b0001 : 4'b1000;
															assign node11310 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node11313 = (inp[7]) ? node11317 : node11314;
															assign node11314 = (inp[14]) ? 4'b1001 : 4'b0000;
															assign node11317 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node11320 = (inp[8]) ? node11336 : node11321;
													assign node11321 = (inp[6]) ? node11329 : node11322;
														assign node11322 = (inp[7]) ? node11326 : node11323;
															assign node11323 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node11326 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node11329 = (inp[14]) ? node11333 : node11330;
															assign node11330 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node11333 = (inp[7]) ? 4'b0001 : 4'b1000;
													assign node11336 = (inp[6]) ? node11344 : node11337;
														assign node11337 = (inp[5]) ? node11341 : node11338;
															assign node11338 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node11341 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node11344 = (inp[14]) ? node11348 : node11345;
															assign node11345 = (inp[7]) ? 4'b0001 : 4'b1000;
															assign node11348 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node11351 = (inp[15]) ? node11409 : node11352;
											assign node11352 = (inp[14]) ? node11378 : node11353;
												assign node11353 = (inp[11]) ? node11363 : node11354;
													assign node11354 = (inp[6]) ? 4'b0000 : node11355;
														assign node11355 = (inp[7]) ? node11359 : node11356;
															assign node11356 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node11359 = (inp[8]) ? 4'b0001 : 4'b1000;
													assign node11363 = (inp[6]) ? node11371 : node11364;
														assign node11364 = (inp[7]) ? node11368 : node11365;
															assign node11365 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node11368 = (inp[8]) ? 4'b1001 : 4'b0000;
														assign node11371 = (inp[7]) ? node11375 : node11372;
															assign node11372 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node11375 = (inp[8]) ? 4'b0001 : 4'b1000;
												assign node11378 = (inp[5]) ? node11394 : node11379;
													assign node11379 = (inp[6]) ? node11387 : node11380;
														assign node11380 = (inp[11]) ? node11384 : node11381;
															assign node11381 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node11384 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node11387 = (inp[11]) ? node11391 : node11388;
															assign node11388 = (inp[8]) ? 4'b1000 : 4'b0000;
															assign node11391 = (inp[7]) ? 4'b0000 : 4'b1000;
													assign node11394 = (inp[6]) ? node11402 : node11395;
														assign node11395 = (inp[11]) ? node11399 : node11396;
															assign node11396 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node11399 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node11402 = (inp[11]) ? node11406 : node11403;
															assign node11403 = (inp[8]) ? 4'b1000 : 4'b0000;
															assign node11406 = (inp[8]) ? 4'b0000 : 4'b0001;
											assign node11409 = (inp[7]) ? node11441 : node11410;
												assign node11410 = (inp[14]) ? node11426 : node11411;
													assign node11411 = (inp[8]) ? node11419 : node11412;
														assign node11412 = (inp[11]) ? node11416 : node11413;
															assign node11413 = (inp[6]) ? 4'b0011 : 4'b1011;
															assign node11416 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node11419 = (inp[5]) ? node11423 : node11420;
															assign node11420 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node11423 = (inp[11]) ? 4'b0010 : 4'b0010;
													assign node11426 = (inp[8]) ? node11434 : node11427;
														assign node11427 = (inp[5]) ? node11431 : node11428;
															assign node11428 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node11431 = (inp[11]) ? 4'b0010 : 4'b0010;
														assign node11434 = (inp[6]) ? node11438 : node11435;
															assign node11435 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node11438 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node11441 = (inp[6]) ? node11457 : node11442;
													assign node11442 = (inp[11]) ? node11450 : node11443;
														assign node11443 = (inp[14]) ? node11447 : node11444;
															assign node11444 = (inp[8]) ? 4'b0011 : 4'b1010;
															assign node11447 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node11450 = (inp[8]) ? node11454 : node11451;
															assign node11451 = (inp[14]) ? 4'b1011 : 4'b0010;
															assign node11454 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node11457 = (inp[11]) ? node11465 : node11458;
														assign node11458 = (inp[8]) ? node11462 : node11459;
															assign node11459 = (inp[14]) ? 4'b1011 : 4'b0010;
															assign node11462 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node11465 = (inp[8]) ? node11469 : node11466;
															assign node11466 = (inp[14]) ? 4'b0011 : 4'b1010;
															assign node11469 = (inp[14]) ? 4'b0010 : 4'b0011;
									assign node11472 = (inp[14]) ? node11596 : node11473;
										assign node11473 = (inp[7]) ? node11533 : node11474;
											assign node11474 = (inp[8]) ? node11504 : node11475;
												assign node11475 = (inp[5]) ? node11489 : node11476;
													assign node11476 = (inp[11]) ? node11484 : node11477;
														assign node11477 = (inp[6]) ? node11481 : node11478;
															assign node11478 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node11481 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node11484 = (inp[6]) ? node11486 : 4'b1001;
															assign node11486 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node11489 = (inp[0]) ? node11497 : node11490;
														assign node11490 = (inp[15]) ? node11494 : node11491;
															assign node11491 = (inp[11]) ? 4'b0011 : 4'b0011;
															assign node11494 = (inp[11]) ? 4'b0001 : 4'b0001;
														assign node11497 = (inp[15]) ? node11501 : node11498;
															assign node11498 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node11501 = (inp[6]) ? 4'b0011 : 4'b0011;
												assign node11504 = (inp[6]) ? node11520 : node11505;
													assign node11505 = (inp[11]) ? node11513 : node11506;
														assign node11506 = (inp[15]) ? node11510 : node11507;
															assign node11507 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node11510 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node11513 = (inp[0]) ? node11517 : node11514;
															assign node11514 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node11517 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node11520 = (inp[11]) ? node11526 : node11521;
														assign node11521 = (inp[0]) ? 4'b1000 : node11522;
															assign node11522 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node11526 = (inp[15]) ? node11530 : node11527;
															assign node11527 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node11530 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node11533 = (inp[8]) ? node11565 : node11534;
												assign node11534 = (inp[15]) ? node11550 : node11535;
													assign node11535 = (inp[0]) ? node11543 : node11536;
														assign node11536 = (inp[6]) ? node11540 : node11537;
															assign node11537 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node11540 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node11543 = (inp[11]) ? node11547 : node11544;
															assign node11544 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node11547 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node11550 = (inp[0]) ? node11558 : node11551;
														assign node11551 = (inp[6]) ? node11555 : node11552;
															assign node11552 = (inp[11]) ? 4'b1000 : 4'b0000;
															assign node11555 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node11558 = (inp[6]) ? node11562 : node11559;
															assign node11559 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node11562 = (inp[11]) ? 4'b0010 : 4'b1010;
												assign node11565 = (inp[6]) ? node11581 : node11566;
													assign node11566 = (inp[11]) ? node11574 : node11567;
														assign node11567 = (inp[15]) ? node11571 : node11568;
															assign node11568 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node11571 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node11574 = (inp[0]) ? node11578 : node11575;
															assign node11575 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node11578 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node11581 = (inp[11]) ? node11589 : node11582;
														assign node11582 = (inp[5]) ? node11586 : node11583;
															assign node11583 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node11586 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node11589 = (inp[0]) ? node11593 : node11590;
															assign node11590 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node11593 = (inp[15]) ? 4'b0011 : 4'b0001;
										assign node11596 = (inp[0]) ? node11656 : node11597;
											assign node11597 = (inp[15]) ? node11625 : node11598;
												assign node11598 = (inp[5]) ? node11612 : node11599;
													assign node11599 = (inp[7]) ? node11607 : node11600;
														assign node11600 = (inp[8]) ? node11604 : node11601;
															assign node11601 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node11604 = (inp[11]) ? 4'b0011 : 4'b0011;
														assign node11607 = (inp[8]) ? 4'b0010 : node11608;
															assign node11608 = (inp[6]) ? 4'b0011 : 4'b0011;
													assign node11612 = (inp[11]) ? node11620 : node11613;
														assign node11613 = (inp[6]) ? node11617 : node11614;
															assign node11614 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node11617 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node11620 = (inp[6]) ? node11622 : 4'b1010;
															assign node11622 = (inp[8]) ? 4'b0010 : 4'b0010;
												assign node11625 = (inp[6]) ? node11641 : node11626;
													assign node11626 = (inp[11]) ? node11634 : node11627;
														assign node11627 = (inp[8]) ? node11631 : node11628;
															assign node11628 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node11631 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node11634 = (inp[7]) ? node11638 : node11635;
															assign node11635 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node11638 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node11641 = (inp[11]) ? node11649 : node11642;
														assign node11642 = (inp[8]) ? node11646 : node11643;
															assign node11643 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node11646 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node11649 = (inp[5]) ? node11653 : node11650;
															assign node11650 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node11653 = (inp[7]) ? 4'b0000 : 4'b0000;
											assign node11656 = (inp[15]) ? node11688 : node11657;
												assign node11657 = (inp[6]) ? node11673 : node11658;
													assign node11658 = (inp[11]) ? node11666 : node11659;
														assign node11659 = (inp[8]) ? node11663 : node11660;
															assign node11660 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node11663 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node11666 = (inp[7]) ? node11670 : node11667;
															assign node11667 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node11670 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node11673 = (inp[11]) ? node11681 : node11674;
														assign node11674 = (inp[5]) ? node11678 : node11675;
															assign node11675 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node11678 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node11681 = (inp[5]) ? node11685 : node11682;
															assign node11682 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node11685 = (inp[7]) ? 4'b0000 : 4'b0000;
												assign node11688 = (inp[8]) ? node11702 : node11689;
													assign node11689 = (inp[7]) ? node11697 : node11690;
														assign node11690 = (inp[5]) ? node11694 : node11691;
															assign node11691 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node11694 = (inp[11]) ? 4'b0010 : 4'b0010;
														assign node11697 = (inp[5]) ? node11699 : 4'b1011;
															assign node11699 = (inp[6]) ? 4'b0011 : 4'b0011;
													assign node11702 = (inp[7]) ? node11710 : node11703;
														assign node11703 = (inp[6]) ? node11707 : node11704;
															assign node11704 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node11707 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node11710 = (inp[11]) ? node11714 : node11711;
															assign node11711 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node11714 = (inp[6]) ? 4'b0010 : 4'b1010;
							assign node11717 = (inp[15]) ? node12097 : node11718;
								assign node11718 = (inp[0]) ? node11870 : node11719;
									assign node11719 = (inp[7]) ? node11799 : node11720;
										assign node11720 = (inp[8]) ? node11760 : node11721;
											assign node11721 = (inp[1]) ? node11729 : node11722;
												assign node11722 = (inp[11]) ? node11726 : node11723;
													assign node11723 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node11726 = (inp[6]) ? 4'b1010 : 4'b0010;
												assign node11729 = (inp[11]) ? node11745 : node11730;
													assign node11730 = (inp[14]) ? node11738 : node11731;
														assign node11731 = (inp[5]) ? node11735 : node11732;
															assign node11732 = (inp[13]) ? 4'b0010 : 4'b0010;
															assign node11735 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node11738 = (inp[5]) ? node11742 : node11739;
															assign node11739 = (inp[13]) ? 4'b0010 : 4'b0010;
															assign node11742 = (inp[13]) ? 4'b0010 : 4'b0010;
													assign node11745 = (inp[14]) ? node11753 : node11746;
														assign node11746 = (inp[13]) ? node11750 : node11747;
															assign node11747 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node11750 = (inp[6]) ? 4'b0010 : 4'b1010;
														assign node11753 = (inp[6]) ? node11757 : node11754;
															assign node11754 = (inp[13]) ? 4'b1010 : 4'b0010;
															assign node11757 = (inp[13]) ? 4'b0010 : 4'b1010;
											assign node11760 = (inp[13]) ? node11776 : node11761;
												assign node11761 = (inp[11]) ? node11769 : node11762;
													assign node11762 = (inp[6]) ? node11766 : node11763;
														assign node11763 = (inp[1]) ? 4'b0011 : 4'b1011;
														assign node11766 = (inp[1]) ? 4'b1011 : 4'b0011;
													assign node11769 = (inp[1]) ? node11773 : node11770;
														assign node11770 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node11773 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node11776 = (inp[1]) ? node11784 : node11777;
													assign node11777 = (inp[11]) ? node11781 : node11778;
														assign node11778 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node11781 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node11784 = (inp[5]) ? node11792 : node11785;
														assign node11785 = (inp[11]) ? node11789 : node11786;
															assign node11786 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node11789 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node11792 = (inp[6]) ? node11796 : node11793;
															assign node11793 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node11796 = (inp[11]) ? 4'b0011 : 4'b1011;
										assign node11799 = (inp[8]) ? node11847 : node11800;
											assign node11800 = (inp[5]) ? node11824 : node11801;
												assign node11801 = (inp[11]) ? node11813 : node11802;
													assign node11802 = (inp[6]) ? node11808 : node11803;
														assign node11803 = (inp[1]) ? 4'b0011 : node11804;
															assign node11804 = (inp[13]) ? 4'b0011 : 4'b1011;
														assign node11808 = (inp[1]) ? 4'b1011 : node11809;
															assign node11809 = (inp[13]) ? 4'b1011 : 4'b0011;
													assign node11813 = (inp[6]) ? node11819 : node11814;
														assign node11814 = (inp[13]) ? 4'b1011 : node11815;
															assign node11815 = (inp[1]) ? 4'b1011 : 4'b0011;
														assign node11819 = (inp[13]) ? 4'b0011 : node11820;
															assign node11820 = (inp[1]) ? 4'b0011 : 4'b1011;
												assign node11824 = (inp[11]) ? node11836 : node11825;
													assign node11825 = (inp[6]) ? node11831 : node11826;
														assign node11826 = (inp[13]) ? 4'b0011 : node11827;
															assign node11827 = (inp[1]) ? 4'b0011 : 4'b1011;
														assign node11831 = (inp[1]) ? 4'b1011 : node11832;
															assign node11832 = (inp[13]) ? 4'b1011 : 4'b0011;
													assign node11836 = (inp[6]) ? node11842 : node11837;
														assign node11837 = (inp[1]) ? 4'b1011 : node11838;
															assign node11838 = (inp[13]) ? 4'b1011 : 4'b0011;
														assign node11842 = (inp[13]) ? 4'b0011 : node11843;
															assign node11843 = (inp[1]) ? 4'b0011 : 4'b1011;
											assign node11847 = (inp[11]) ? node11859 : node11848;
												assign node11848 = (inp[6]) ? node11854 : node11849;
													assign node11849 = (inp[1]) ? 4'b0010 : node11850;
														assign node11850 = (inp[13]) ? 4'b0010 : 4'b1010;
													assign node11854 = (inp[1]) ? 4'b1010 : node11855;
														assign node11855 = (inp[13]) ? 4'b1010 : 4'b0010;
												assign node11859 = (inp[6]) ? node11865 : node11860;
													assign node11860 = (inp[13]) ? 4'b1010 : node11861;
														assign node11861 = (inp[1]) ? 4'b1010 : 4'b0010;
													assign node11865 = (inp[1]) ? 4'b0010 : node11866;
														assign node11866 = (inp[13]) ? 4'b0010 : 4'b1010;
									assign node11870 = (inp[14]) ? node11994 : node11871;
										assign node11871 = (inp[5]) ? node11931 : node11872;
											assign node11872 = (inp[13]) ? node11904 : node11873;
												assign node11873 = (inp[7]) ? node11889 : node11874;
													assign node11874 = (inp[8]) ? node11882 : node11875;
														assign node11875 = (inp[11]) ? node11879 : node11876;
															assign node11876 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node11879 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node11882 = (inp[1]) ? node11886 : node11883;
															assign node11883 = (inp[11]) ? 4'b0001 : 4'b0001;
															assign node11886 = (inp[6]) ? 4'b0001 : 4'b0001;
													assign node11889 = (inp[8]) ? node11897 : node11890;
														assign node11890 = (inp[11]) ? node11894 : node11891;
															assign node11891 = (inp[1]) ? 4'b0001 : 4'b0001;
															assign node11894 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node11897 = (inp[6]) ? node11901 : node11898;
															assign node11898 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node11901 = (inp[11]) ? 4'b1000 : 4'b0000;
												assign node11904 = (inp[11]) ? node11920 : node11905;
													assign node11905 = (inp[6]) ? node11913 : node11906;
														assign node11906 = (inp[7]) ? node11910 : node11907;
															assign node11907 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node11910 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node11913 = (inp[8]) ? node11917 : node11914;
															assign node11914 = (inp[7]) ? 4'b1001 : 4'b0000;
															assign node11917 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node11920 = (inp[6]) ? node11926 : node11921;
														assign node11921 = (inp[1]) ? node11923 : 4'b1001;
															assign node11923 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node11926 = (inp[8]) ? node11928 : 4'b0001;
															assign node11928 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node11931 = (inp[11]) ? node11963 : node11932;
												assign node11932 = (inp[6]) ? node11948 : node11933;
													assign node11933 = (inp[1]) ? node11941 : node11934;
														assign node11934 = (inp[13]) ? node11938 : node11935;
															assign node11935 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node11938 = (inp[8]) ? 4'b0000 : 4'b1000;
														assign node11941 = (inp[8]) ? node11945 : node11942;
															assign node11942 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node11945 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node11948 = (inp[1]) ? node11956 : node11949;
														assign node11949 = (inp[13]) ? node11953 : node11950;
															assign node11950 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node11953 = (inp[8]) ? 4'b1000 : 4'b0000;
														assign node11956 = (inp[13]) ? node11960 : node11957;
															assign node11957 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node11960 = (inp[8]) ? 4'b1000 : 4'b1000;
												assign node11963 = (inp[6]) ? node11979 : node11964;
													assign node11964 = (inp[1]) ? node11972 : node11965;
														assign node11965 = (inp[13]) ? node11969 : node11966;
															assign node11966 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node11969 = (inp[8]) ? 4'b1001 : 4'b0000;
														assign node11972 = (inp[13]) ? node11976 : node11973;
															assign node11973 = (inp[7]) ? 4'b1000 : 4'b0000;
															assign node11976 = (inp[8]) ? 4'b1000 : 4'b1000;
													assign node11979 = (inp[13]) ? node11987 : node11980;
														assign node11980 = (inp[1]) ? node11984 : node11981;
															assign node11981 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node11984 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node11987 = (inp[7]) ? node11991 : node11988;
															assign node11988 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node11991 = (inp[8]) ? 4'b0000 : 4'b0001;
										assign node11994 = (inp[6]) ? node12046 : node11995;
											assign node11995 = (inp[11]) ? node12021 : node11996;
												assign node11996 = (inp[13]) ? node12012 : node11997;
													assign node11997 = (inp[1]) ? node12005 : node11998;
														assign node11998 = (inp[5]) ? node12002 : node11999;
															assign node11999 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node12002 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node12005 = (inp[8]) ? node12009 : node12006;
															assign node12006 = (inp[7]) ? 4'b0001 : 4'b1000;
															assign node12009 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node12012 = (inp[8]) ? node12018 : node12013;
														assign node12013 = (inp[7]) ? 4'b0001 : node12014;
															assign node12014 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node12018 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node12021 = (inp[1]) ? node12037 : node12022;
													assign node12022 = (inp[13]) ? node12030 : node12023;
														assign node12023 = (inp[8]) ? node12027 : node12024;
															assign node12024 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node12027 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node12030 = (inp[8]) ? node12034 : node12031;
															assign node12031 = (inp[7]) ? 4'b1001 : 4'b0000;
															assign node12034 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node12037 = (inp[7]) ? node12043 : node12038;
														assign node12038 = (inp[8]) ? 4'b1001 : node12039;
															assign node12039 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node12043 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node12046 = (inp[11]) ? node12072 : node12047;
												assign node12047 = (inp[1]) ? node12063 : node12048;
													assign node12048 = (inp[13]) ? node12056 : node12049;
														assign node12049 = (inp[7]) ? node12053 : node12050;
															assign node12050 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node12053 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node12056 = (inp[7]) ? node12060 : node12057;
															assign node12057 = (inp[8]) ? 4'b1001 : 4'b0000;
															assign node12060 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node12063 = (inp[8]) ? node12069 : node12064;
														assign node12064 = (inp[7]) ? 4'b1001 : node12065;
															assign node12065 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node12069 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node12072 = (inp[13]) ? node12088 : node12073;
													assign node12073 = (inp[1]) ? node12081 : node12074;
														assign node12074 = (inp[7]) ? node12078 : node12075;
															assign node12075 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node12078 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node12081 = (inp[8]) ? node12085 : node12082;
															assign node12082 = (inp[7]) ? 4'b0001 : 4'b1000;
															assign node12085 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node12088 = (inp[7]) ? node12094 : node12089;
														assign node12089 = (inp[8]) ? 4'b0001 : node12090;
															assign node12090 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node12094 = (inp[8]) ? 4'b0000 : 4'b0001;
								assign node12097 = (inp[0]) ? node12219 : node12098;
									assign node12098 = (inp[1]) ? node12168 : node12099;
										assign node12099 = (inp[6]) ? node12137 : node12100;
											assign node12100 = (inp[11]) ? node12116 : node12101;
												assign node12101 = (inp[13]) ? node12109 : node12102;
													assign node12102 = (inp[8]) ? node12106 : node12103;
														assign node12103 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node12106 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node12109 = (inp[8]) ? node12113 : node12110;
														assign node12110 = (inp[7]) ? 4'b0001 : 4'b1000;
														assign node12113 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node12116 = (inp[13]) ? node12130 : node12117;
													assign node12117 = (inp[14]) ? node12123 : node12118;
														assign node12118 = (inp[5]) ? 4'b0000 : node12119;
															assign node12119 = (inp[7]) ? 4'b0000 : 4'b0000;
														assign node12123 = (inp[5]) ? node12127 : node12124;
															assign node12124 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node12127 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node12130 = (inp[7]) ? node12134 : node12131;
														assign node12131 = (inp[8]) ? 4'b1001 : 4'b0000;
														assign node12134 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node12137 = (inp[11]) ? node12153 : node12138;
												assign node12138 = (inp[13]) ? node12146 : node12139;
													assign node12139 = (inp[7]) ? node12143 : node12140;
														assign node12140 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node12143 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node12146 = (inp[7]) ? node12150 : node12147;
														assign node12147 = (inp[8]) ? 4'b1001 : 4'b0000;
														assign node12150 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node12153 = (inp[13]) ? node12161 : node12154;
													assign node12154 = (inp[8]) ? node12158 : node12155;
														assign node12155 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node12158 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node12161 = (inp[7]) ? node12165 : node12162;
														assign node12162 = (inp[8]) ? 4'b0001 : 4'b1000;
														assign node12165 = (inp[8]) ? 4'b0000 : 4'b0001;
										assign node12168 = (inp[11]) ? node12200 : node12169;
											assign node12169 = (inp[6]) ? node12179 : node12170;
												assign node12170 = (inp[7]) ? node12176 : node12171;
													assign node12171 = (inp[8]) ? 4'b0001 : node12172;
														assign node12172 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node12176 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node12179 = (inp[13]) ? node12187 : node12180;
													assign node12180 = (inp[8]) ? node12184 : node12181;
														assign node12181 = (inp[7]) ? 4'b1001 : 4'b0000;
														assign node12184 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node12187 = (inp[5]) ? node12193 : node12188;
														assign node12188 = (inp[14]) ? 4'b1001 : node12189;
															assign node12189 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node12193 = (inp[14]) ? node12197 : node12194;
															assign node12194 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node12197 = (inp[7]) ? 4'b1000 : 4'b1000;
											assign node12200 = (inp[6]) ? node12210 : node12201;
												assign node12201 = (inp[7]) ? node12207 : node12202;
													assign node12202 = (inp[8]) ? 4'b1001 : node12203;
														assign node12203 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node12207 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node12210 = (inp[8]) ? node12216 : node12211;
													assign node12211 = (inp[7]) ? 4'b0001 : node12212;
														assign node12212 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node12216 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node12219 = (inp[11]) ? node12279 : node12220;
										assign node12220 = (inp[6]) ? node12254 : node12221;
											assign node12221 = (inp[1]) ? node12245 : node12222;
												assign node12222 = (inp[13]) ? node12238 : node12223;
													assign node12223 = (inp[14]) ? node12231 : node12224;
														assign node12224 = (inp[7]) ? node12228 : node12225;
															assign node12225 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node12228 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node12231 = (inp[5]) ? node12235 : node12232;
															assign node12232 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node12235 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node12238 = (inp[8]) ? node12242 : node12239;
														assign node12239 = (inp[7]) ? 4'b0011 : 4'b1010;
														assign node12242 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node12245 = (inp[7]) ? node12251 : node12246;
													assign node12246 = (inp[8]) ? 4'b0011 : node12247;
														assign node12247 = (inp[13]) ? 4'b0010 : 4'b1010;
													assign node12251 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node12254 = (inp[13]) ? node12270 : node12255;
												assign node12255 = (inp[1]) ? node12263 : node12256;
													assign node12256 = (inp[7]) ? node12260 : node12257;
														assign node12257 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node12260 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node12263 = (inp[7]) ? node12267 : node12264;
														assign node12264 = (inp[8]) ? 4'b1011 : 4'b0010;
														assign node12267 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node12270 = (inp[7]) ? node12276 : node12271;
													assign node12271 = (inp[8]) ? 4'b1011 : node12272;
														assign node12272 = (inp[1]) ? 4'b1010 : 4'b0010;
													assign node12276 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node12279 = (inp[6]) ? node12313 : node12280;
											assign node12280 = (inp[13]) ? node12304 : node12281;
												assign node12281 = (inp[1]) ? node12297 : node12282;
													assign node12282 = (inp[5]) ? node12290 : node12283;
														assign node12283 = (inp[14]) ? node12287 : node12284;
															assign node12284 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node12287 = (inp[8]) ? 4'b0010 : 4'b0010;
														assign node12290 = (inp[7]) ? node12294 : node12291;
															assign node12291 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node12294 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node12297 = (inp[7]) ? node12301 : node12298;
														assign node12298 = (inp[8]) ? 4'b1011 : 4'b0010;
														assign node12301 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node12304 = (inp[8]) ? node12310 : node12305;
													assign node12305 = (inp[7]) ? 4'b1011 : node12306;
														assign node12306 = (inp[1]) ? 4'b1010 : 4'b0010;
													assign node12310 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node12313 = (inp[13]) ? node12329 : node12314;
												assign node12314 = (inp[1]) ? node12322 : node12315;
													assign node12315 = (inp[8]) ? node12319 : node12316;
														assign node12316 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node12319 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node12322 = (inp[8]) ? node12326 : node12323;
														assign node12323 = (inp[7]) ? 4'b0011 : 4'b1010;
														assign node12326 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node12329 = (inp[7]) ? node12335 : node12330;
													assign node12330 = (inp[8]) ? 4'b0011 : node12331;
														assign node12331 = (inp[1]) ? 4'b0010 : 4'b1010;
													assign node12335 = (inp[8]) ? 4'b0010 : 4'b0011;
						assign node12338 = (inp[7]) ? node13300 : node12339;
							assign node12339 = (inp[8]) ? node12819 : node12340;
								assign node12340 = (inp[14]) ? node12586 : node12341;
									assign node12341 = (inp[2]) ? node12467 : node12342;
										assign node12342 = (inp[15]) ? node12404 : node12343;
											assign node12343 = (inp[1]) ? node12373 : node12344;
												assign node12344 = (inp[13]) ? node12358 : node12345;
													assign node12345 = (inp[0]) ? node12353 : node12346;
														assign node12346 = (inp[5]) ? node12350 : node12347;
															assign node12347 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node12350 = (inp[11]) ? 4'b0001 : 4'b0001;
														assign node12353 = (inp[5]) ? 4'b1011 : node12354;
															assign node12354 = (inp[6]) ? 4'b0001 : 4'b0001;
													assign node12358 = (inp[6]) ? node12366 : node12359;
														assign node12359 = (inp[11]) ? node12363 : node12360;
															assign node12360 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node12363 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node12366 = (inp[11]) ? node12370 : node12367;
															assign node12367 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node12370 = (inp[5]) ? 4'b1001 : 4'b1001;
												assign node12373 = (inp[5]) ? node12389 : node12374;
													assign node12374 = (inp[0]) ? node12382 : node12375;
														assign node12375 = (inp[11]) ? node12379 : node12376;
															assign node12376 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node12379 = (inp[13]) ? 4'b1011 : 4'b0011;
														assign node12382 = (inp[11]) ? node12386 : node12383;
															assign node12383 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node12386 = (inp[6]) ? 4'b0001 : 4'b0001;
													assign node12389 = (inp[0]) ? node12397 : node12390;
														assign node12390 = (inp[6]) ? node12394 : node12391;
															assign node12391 = (inp[11]) ? 4'b0001 : 4'b0001;
															assign node12394 = (inp[13]) ? 4'b0001 : 4'b0001;
														assign node12397 = (inp[11]) ? node12401 : node12398;
															assign node12398 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node12401 = (inp[13]) ? 4'b0011 : 4'b0011;
											assign node12404 = (inp[5]) ? node12436 : node12405;
												assign node12405 = (inp[0]) ? node12421 : node12406;
													assign node12406 = (inp[11]) ? node12414 : node12407;
														assign node12407 = (inp[6]) ? node12411 : node12408;
															assign node12408 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node12411 = (inp[1]) ? 4'b0001 : 4'b0001;
														assign node12414 = (inp[6]) ? node12418 : node12415;
															assign node12415 = (inp[1]) ? 4'b0001 : 4'b0001;
															assign node12418 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node12421 = (inp[1]) ? node12429 : node12422;
														assign node12422 = (inp[6]) ? node12426 : node12423;
															assign node12423 = (inp[13]) ? 4'b1011 : 4'b0011;
															assign node12426 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node12429 = (inp[11]) ? node12433 : node12430;
															assign node12430 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node12433 = (inp[6]) ? 4'b0011 : 4'b0011;
												assign node12436 = (inp[0]) ? node12452 : node12437;
													assign node12437 = (inp[11]) ? node12445 : node12438;
														assign node12438 = (inp[6]) ? node12442 : node12439;
															assign node12439 = (inp[1]) ? 4'b0011 : 4'b1011;
															assign node12442 = (inp[13]) ? 4'b0011 : 4'b0011;
														assign node12445 = (inp[6]) ? node12449 : node12446;
															assign node12446 = (inp[1]) ? 4'b0011 : 4'b0011;
															assign node12449 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node12452 = (inp[6]) ? node12460 : node12453;
														assign node12453 = (inp[11]) ? node12457 : node12454;
															assign node12454 = (inp[1]) ? 4'b0001 : 4'b1001;
															assign node12457 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node12460 = (inp[11]) ? node12464 : node12461;
															assign node12461 = (inp[13]) ? 4'b0001 : 4'b0001;
															assign node12464 = (inp[13]) ? 4'b0001 : 4'b1001;
										assign node12467 = (inp[15]) ? node12529 : node12468;
											assign node12468 = (inp[11]) ? node12498 : node12469;
												assign node12469 = (inp[6]) ? node12485 : node12470;
													assign node12470 = (inp[13]) ? node12478 : node12471;
														assign node12471 = (inp[1]) ? node12475 : node12472;
															assign node12472 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node12475 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node12478 = (inp[1]) ? node12482 : node12479;
															assign node12479 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node12482 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node12485 = (inp[13]) ? node12493 : node12486;
														assign node12486 = (inp[5]) ? node12490 : node12487;
															assign node12487 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node12490 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node12493 = (inp[1]) ? 4'b1000 : node12494;
															assign node12494 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node12498 = (inp[6]) ? node12514 : node12499;
													assign node12499 = (inp[13]) ? node12507 : node12500;
														assign node12500 = (inp[1]) ? node12504 : node12501;
															assign node12501 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node12504 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node12507 = (inp[1]) ? node12511 : node12508;
															assign node12508 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node12511 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node12514 = (inp[1]) ? node12522 : node12515;
														assign node12515 = (inp[13]) ? node12519 : node12516;
															assign node12516 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node12519 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node12522 = (inp[13]) ? node12526 : node12523;
															assign node12523 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node12526 = (inp[5]) ? 4'b0000 : 4'b0000;
											assign node12529 = (inp[6]) ? node12557 : node12530;
												assign node12530 = (inp[11]) ? node12546 : node12531;
													assign node12531 = (inp[13]) ? node12539 : node12532;
														assign node12532 = (inp[0]) ? node12536 : node12533;
															assign node12533 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node12536 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node12539 = (inp[1]) ? node12543 : node12540;
															assign node12540 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node12543 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node12546 = (inp[1]) ? node12552 : node12547;
														assign node12547 = (inp[5]) ? node12549 : 4'b0000;
															assign node12549 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node12552 = (inp[13]) ? node12554 : 4'b0000;
															assign node12554 = (inp[5]) ? 4'b1000 : 4'b1000;
												assign node12557 = (inp[11]) ? node12571 : node12558;
													assign node12558 = (inp[1]) ? node12564 : node12559;
														assign node12559 = (inp[13]) ? 4'b0010 : node12560;
															assign node12560 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node12564 = (inp[13]) ? node12568 : node12565;
															assign node12565 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node12568 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node12571 = (inp[13]) ? node12579 : node12572;
														assign node12572 = (inp[1]) ? node12576 : node12573;
															assign node12573 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node12576 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node12579 = (inp[1]) ? node12583 : node12580;
															assign node12580 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node12583 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node12586 = (inp[1]) ? node12702 : node12587;
										assign node12587 = (inp[5]) ? node12643 : node12588;
											assign node12588 = (inp[0]) ? node12612 : node12589;
												assign node12589 = (inp[15]) ? node12597 : node12590;
													assign node12590 = (inp[11]) ? node12594 : node12591;
														assign node12591 = (inp[6]) ? 4'b0010 : 4'b1010;
														assign node12594 = (inp[6]) ? 4'b1010 : 4'b0010;
													assign node12597 = (inp[2]) ? node12605 : node12598;
														assign node12598 = (inp[11]) ? node12602 : node12599;
															assign node12599 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node12602 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node12605 = (inp[6]) ? node12609 : node12606;
															assign node12606 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node12609 = (inp[11]) ? 4'b1000 : 4'b0000;
												assign node12612 = (inp[15]) ? node12628 : node12613;
													assign node12613 = (inp[13]) ? node12621 : node12614;
														assign node12614 = (inp[2]) ? node12618 : node12615;
															assign node12615 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node12618 = (inp[11]) ? 4'b0000 : 4'b0000;
														assign node12621 = (inp[6]) ? node12625 : node12622;
															assign node12622 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node12625 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node12628 = (inp[2]) ? node12636 : node12629;
														assign node12629 = (inp[11]) ? node12633 : node12630;
															assign node12630 = (inp[6]) ? 4'b0010 : 4'b1010;
															assign node12633 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node12636 = (inp[11]) ? node12640 : node12637;
															assign node12637 = (inp[6]) ? 4'b0010 : 4'b1010;
															assign node12640 = (inp[6]) ? 4'b1010 : 4'b0010;
											assign node12643 = (inp[0]) ? node12671 : node12644;
												assign node12644 = (inp[15]) ? node12658 : node12645;
													assign node12645 = (inp[2]) ? node12653 : node12646;
														assign node12646 = (inp[13]) ? node12650 : node12647;
															assign node12647 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node12650 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node12653 = (inp[13]) ? 4'b0000 : node12654;
															assign node12654 = (inp[11]) ? 4'b0000 : 4'b0000;
													assign node12658 = (inp[2]) ? node12666 : node12659;
														assign node12659 = (inp[13]) ? node12663 : node12660;
															assign node12660 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node12663 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node12666 = (inp[13]) ? 4'b1010 : node12667;
															assign node12667 = (inp[11]) ? 4'b0010 : 4'b0010;
												assign node12671 = (inp[15]) ? node12687 : node12672;
													assign node12672 = (inp[13]) ? node12680 : node12673;
														assign node12673 = (inp[6]) ? node12677 : node12674;
															assign node12674 = (inp[11]) ? 4'b0010 : 4'b1010;
															assign node12677 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node12680 = (inp[2]) ? node12684 : node12681;
															assign node12681 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node12684 = (inp[6]) ? 4'b0010 : 4'b0010;
													assign node12687 = (inp[2]) ? node12695 : node12688;
														assign node12688 = (inp[13]) ? node12692 : node12689;
															assign node12689 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node12692 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node12695 = (inp[11]) ? node12699 : node12696;
															assign node12696 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node12699 = (inp[6]) ? 4'b1000 : 4'b0000;
										assign node12702 = (inp[13]) ? node12760 : node12703;
											assign node12703 = (inp[11]) ? node12733 : node12704;
												assign node12704 = (inp[6]) ? node12720 : node12705;
													assign node12705 = (inp[2]) ? node12713 : node12706;
														assign node12706 = (inp[5]) ? node12710 : node12707;
															assign node12707 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node12710 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node12713 = (inp[0]) ? node12717 : node12714;
															assign node12714 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node12717 = (inp[5]) ? 4'b1000 : 4'b1000;
													assign node12720 = (inp[2]) ? node12726 : node12721;
														assign node12721 = (inp[15]) ? 4'b0000 : node12722;
															assign node12722 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node12726 = (inp[0]) ? node12730 : node12727;
															assign node12727 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node12730 = (inp[15]) ? 4'b0000 : 4'b0000;
												assign node12733 = (inp[6]) ? node12747 : node12734;
													assign node12734 = (inp[2]) ? node12742 : node12735;
														assign node12735 = (inp[15]) ? node12739 : node12736;
															assign node12736 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node12739 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node12742 = (inp[5]) ? node12744 : 4'b0000;
															assign node12744 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node12747 = (inp[15]) ? node12755 : node12748;
														assign node12748 = (inp[2]) ? node12752 : node12749;
															assign node12749 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node12752 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node12755 = (inp[5]) ? node12757 : 4'b1010;
															assign node12757 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node12760 = (inp[11]) ? node12792 : node12761;
												assign node12761 = (inp[6]) ? node12777 : node12762;
													assign node12762 = (inp[15]) ? node12770 : node12763;
														assign node12763 = (inp[5]) ? node12767 : node12764;
															assign node12764 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node12767 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node12770 = (inp[5]) ? node12774 : node12771;
															assign node12771 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node12774 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node12777 = (inp[15]) ? node12785 : node12778;
														assign node12778 = (inp[0]) ? node12782 : node12779;
															assign node12779 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node12782 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node12785 = (inp[0]) ? node12789 : node12786;
															assign node12786 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node12789 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node12792 = (inp[6]) ? node12808 : node12793;
													assign node12793 = (inp[5]) ? node12801 : node12794;
														assign node12794 = (inp[2]) ? node12798 : node12795;
															assign node12795 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node12798 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node12801 = (inp[2]) ? node12805 : node12802;
															assign node12802 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node12805 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node12808 = (inp[2]) ? node12814 : node12809;
														assign node12809 = (inp[5]) ? 4'b0000 : node12810;
															assign node12810 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node12814 = (inp[5]) ? node12816 : 4'b0000;
															assign node12816 = (inp[0]) ? 4'b0000 : 4'b0000;
								assign node12819 = (inp[14]) ? node13065 : node12820;
									assign node12820 = (inp[2]) ? node12942 : node12821;
										assign node12821 = (inp[5]) ? node12885 : node12822;
											assign node12822 = (inp[13]) ? node12854 : node12823;
												assign node12823 = (inp[6]) ? node12839 : node12824;
													assign node12824 = (inp[11]) ? node12832 : node12825;
														assign node12825 = (inp[1]) ? node12829 : node12826;
															assign node12826 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node12829 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node12832 = (inp[15]) ? node12836 : node12833;
															assign node12833 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node12836 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node12839 = (inp[11]) ? node12847 : node12840;
														assign node12840 = (inp[0]) ? node12844 : node12841;
															assign node12841 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node12844 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node12847 = (inp[1]) ? node12851 : node12848;
															assign node12848 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node12851 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node12854 = (inp[1]) ? node12870 : node12855;
													assign node12855 = (inp[0]) ? node12863 : node12856;
														assign node12856 = (inp[15]) ? node12860 : node12857;
															assign node12857 = (inp[11]) ? 4'b0010 : 4'b1010;
															assign node12860 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node12863 = (inp[15]) ? node12867 : node12864;
															assign node12864 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node12867 = (inp[11]) ? 4'b0010 : 4'b0010;
													assign node12870 = (inp[0]) ? node12878 : node12871;
														assign node12871 = (inp[15]) ? node12875 : node12872;
															assign node12872 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node12875 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node12878 = (inp[15]) ? node12882 : node12879;
															assign node12879 = (inp[11]) ? 4'b1000 : 4'b0000;
															assign node12882 = (inp[6]) ? 4'b0010 : 4'b1010;
											assign node12885 = (inp[15]) ? node12913 : node12886;
												assign node12886 = (inp[0]) ? node12900 : node12887;
													assign node12887 = (inp[11]) ? node12895 : node12888;
														assign node12888 = (inp[6]) ? node12892 : node12889;
															assign node12889 = (inp[1]) ? 4'b0000 : 4'b1000;
															assign node12892 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node12895 = (inp[6]) ? node12897 : 4'b0000;
															assign node12897 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node12900 = (inp[6]) ? node12906 : node12901;
														assign node12901 = (inp[11]) ? node12903 : 4'b1010;
															assign node12903 = (inp[1]) ? 4'b0010 : 4'b0010;
														assign node12906 = (inp[11]) ? node12910 : node12907;
															assign node12907 = (inp[1]) ? 4'b0010 : 4'b0010;
															assign node12910 = (inp[1]) ? 4'b0010 : 4'b1010;
												assign node12913 = (inp[0]) ? node12927 : node12914;
													assign node12914 = (inp[11]) ? node12920 : node12915;
														assign node12915 = (inp[6]) ? 4'b0010 : node12916;
															assign node12916 = (inp[13]) ? 4'b0010 : 4'b1010;
														assign node12920 = (inp[6]) ? node12924 : node12921;
															assign node12921 = (inp[1]) ? 4'b1010 : 4'b0010;
															assign node12924 = (inp[13]) ? 4'b0010 : 4'b1010;
													assign node12927 = (inp[13]) ? node12935 : node12928;
														assign node12928 = (inp[1]) ? node12932 : node12929;
															assign node12929 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node12932 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node12935 = (inp[6]) ? node12939 : node12936;
															assign node12936 = (inp[1]) ? 4'b0000 : 4'b0000;
															assign node12939 = (inp[11]) ? 4'b0000 : 4'b0000;
										assign node12942 = (inp[13]) ? node13006 : node12943;
											assign node12943 = (inp[15]) ? node12975 : node12944;
												assign node12944 = (inp[6]) ? node12960 : node12945;
													assign node12945 = (inp[11]) ? node12953 : node12946;
														assign node12946 = (inp[1]) ? node12950 : node12947;
															assign node12947 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node12950 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node12953 = (inp[1]) ? node12957 : node12954;
															assign node12954 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node12957 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node12960 = (inp[11]) ? node12968 : node12961;
														assign node12961 = (inp[1]) ? node12965 : node12962;
															assign node12962 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node12965 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node12968 = (inp[1]) ? node12972 : node12969;
															assign node12969 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node12972 = (inp[5]) ? 4'b0001 : 4'b0001;
												assign node12975 = (inp[6]) ? node12991 : node12976;
													assign node12976 = (inp[11]) ? node12984 : node12977;
														assign node12977 = (inp[1]) ? node12981 : node12978;
															assign node12978 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node12981 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node12984 = (inp[1]) ? node12988 : node12985;
															assign node12985 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node12988 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node12991 = (inp[1]) ? node12999 : node12992;
														assign node12992 = (inp[11]) ? node12996 : node12993;
															assign node12993 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node12996 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node12999 = (inp[11]) ? node13003 : node13000;
															assign node13000 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node13003 = (inp[5]) ? 4'b0001 : 4'b0001;
											assign node13006 = (inp[6]) ? node13036 : node13007;
												assign node13007 = (inp[11]) ? node13021 : node13008;
													assign node13008 = (inp[0]) ? node13014 : node13009;
														assign node13009 = (inp[1]) ? node13011 : 4'b0011;
															assign node13011 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node13014 = (inp[1]) ? node13018 : node13015;
															assign node13015 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node13018 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node13021 = (inp[0]) ? node13029 : node13022;
														assign node13022 = (inp[15]) ? node13026 : node13023;
															assign node13023 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node13026 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node13029 = (inp[5]) ? node13033 : node13030;
															assign node13030 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node13033 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node13036 = (inp[11]) ? node13050 : node13037;
													assign node13037 = (inp[15]) ? node13043 : node13038;
														assign node13038 = (inp[0]) ? node13040 : 4'b1001;
															assign node13040 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node13043 = (inp[0]) ? node13047 : node13044;
															assign node13044 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node13047 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node13050 = (inp[5]) ? node13058 : node13051;
														assign node13051 = (inp[15]) ? node13055 : node13052;
															assign node13052 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node13055 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node13058 = (inp[0]) ? node13062 : node13059;
															assign node13059 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node13062 = (inp[15]) ? 4'b0001 : 4'b0011;
									assign node13065 = (inp[15]) ? node13185 : node13066;
										assign node13066 = (inp[1]) ? node13126 : node13067;
											assign node13067 = (inp[6]) ? node13097 : node13068;
												assign node13068 = (inp[5]) ? node13082 : node13069;
													assign node13069 = (inp[0]) ? node13075 : node13070;
														assign node13070 = (inp[2]) ? node13072 : 4'b0011;
															assign node13072 = (inp[13]) ? 4'b0011 : 4'b0011;
														assign node13075 = (inp[11]) ? node13079 : node13076;
															assign node13076 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node13079 = (inp[13]) ? 4'b1001 : 4'b0001;
													assign node13082 = (inp[0]) ? node13090 : node13083;
														assign node13083 = (inp[13]) ? node13087 : node13084;
															assign node13084 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node13087 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node13090 = (inp[11]) ? node13094 : node13091;
															assign node13091 = (inp[13]) ? 4'b0011 : 4'b1011;
															assign node13094 = (inp[13]) ? 4'b1011 : 4'b0011;
												assign node13097 = (inp[13]) ? node13111 : node13098;
													assign node13098 = (inp[11]) ? node13104 : node13099;
														assign node13099 = (inp[2]) ? 4'b0001 : node13100;
															assign node13100 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node13104 = (inp[0]) ? node13108 : node13105;
															assign node13105 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node13108 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node13111 = (inp[11]) ? node13119 : node13112;
														assign node13112 = (inp[5]) ? node13116 : node13113;
															assign node13113 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node13116 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node13119 = (inp[5]) ? node13123 : node13120;
															assign node13120 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node13123 = (inp[0]) ? 4'b0011 : 4'b0001;
											assign node13126 = (inp[2]) ? node13158 : node13127;
												assign node13127 = (inp[13]) ? node13143 : node13128;
													assign node13128 = (inp[6]) ? node13136 : node13129;
														assign node13129 = (inp[11]) ? node13133 : node13130;
															assign node13130 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node13133 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node13136 = (inp[11]) ? node13140 : node13137;
															assign node13137 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node13140 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node13143 = (inp[5]) ? node13151 : node13144;
														assign node13144 = (inp[0]) ? node13148 : node13145;
															assign node13145 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node13148 = (inp[6]) ? 4'b0001 : 4'b0001;
														assign node13151 = (inp[0]) ? node13155 : node13152;
															assign node13152 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node13155 = (inp[11]) ? 4'b0011 : 4'b0011;
												assign node13158 = (inp[0]) ? node13174 : node13159;
													assign node13159 = (inp[5]) ? node13167 : node13160;
														assign node13160 = (inp[11]) ? node13164 : node13161;
															assign node13161 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node13164 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node13167 = (inp[11]) ? node13171 : node13168;
															assign node13168 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node13171 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node13174 = (inp[5]) ? node13180 : node13175;
														assign node13175 = (inp[11]) ? node13177 : 4'b0001;
															assign node13177 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node13180 = (inp[6]) ? 4'b0011 : node13181;
															assign node13181 = (inp[11]) ? 4'b1011 : 4'b0011;
										assign node13185 = (inp[2]) ? node13243 : node13186;
											assign node13186 = (inp[5]) ? node13214 : node13187;
												assign node13187 = (inp[0]) ? node13201 : node13188;
													assign node13188 = (inp[13]) ? node13194 : node13189;
														assign node13189 = (inp[11]) ? node13191 : 4'b0001;
															assign node13191 = (inp[1]) ? 4'b0001 : 4'b0001;
														assign node13194 = (inp[6]) ? node13198 : node13195;
															assign node13195 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node13198 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node13201 = (inp[6]) ? node13207 : node13202;
														assign node13202 = (inp[11]) ? node13204 : 4'b0011;
															assign node13204 = (inp[1]) ? 4'b1011 : 4'b0011;
														assign node13207 = (inp[11]) ? node13211 : node13208;
															assign node13208 = (inp[1]) ? 4'b1011 : 4'b0011;
															assign node13211 = (inp[1]) ? 4'b0011 : 4'b0011;
												assign node13214 = (inp[0]) ? node13228 : node13215;
													assign node13215 = (inp[11]) ? node13221 : node13216;
														assign node13216 = (inp[6]) ? 4'b1011 : node13217;
															assign node13217 = (inp[1]) ? 4'b0011 : 4'b0011;
														assign node13221 = (inp[6]) ? node13225 : node13222;
															assign node13222 = (inp[1]) ? 4'b1011 : 4'b0011;
															assign node13225 = (inp[1]) ? 4'b0011 : 4'b0011;
													assign node13228 = (inp[13]) ? node13236 : node13229;
														assign node13229 = (inp[11]) ? node13233 : node13230;
															assign node13230 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node13233 = (inp[1]) ? 4'b0001 : 4'b0001;
														assign node13236 = (inp[1]) ? node13240 : node13237;
															assign node13237 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node13240 = (inp[6]) ? 4'b0001 : 4'b0001;
											assign node13243 = (inp[0]) ? node13275 : node13244;
												assign node13244 = (inp[5]) ? node13260 : node13245;
													assign node13245 = (inp[13]) ? node13253 : node13246;
														assign node13246 = (inp[6]) ? node13250 : node13247;
															assign node13247 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node13250 = (inp[11]) ? 4'b0001 : 4'b0001;
														assign node13253 = (inp[6]) ? node13257 : node13254;
															assign node13254 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node13257 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node13260 = (inp[11]) ? node13268 : node13261;
														assign node13261 = (inp[6]) ? node13265 : node13262;
															assign node13262 = (inp[13]) ? 4'b0011 : 4'b0011;
															assign node13265 = (inp[1]) ? 4'b1011 : 4'b0011;
														assign node13268 = (inp[6]) ? node13272 : node13269;
															assign node13269 = (inp[13]) ? 4'b1011 : 4'b0011;
															assign node13272 = (inp[1]) ? 4'b0011 : 4'b1011;
												assign node13275 = (inp[5]) ? node13289 : node13276;
													assign node13276 = (inp[11]) ? node13284 : node13277;
														assign node13277 = (inp[6]) ? node13281 : node13278;
															assign node13278 = (inp[13]) ? 4'b0011 : 4'b0011;
															assign node13281 = (inp[1]) ? 4'b1011 : 4'b0011;
														assign node13284 = (inp[6]) ? node13286 : 4'b1011;
															assign node13286 = (inp[13]) ? 4'b0011 : 4'b1011;
													assign node13289 = (inp[11]) ? node13297 : node13290;
														assign node13290 = (inp[6]) ? node13294 : node13291;
															assign node13291 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node13294 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node13297 = (inp[6]) ? 4'b0001 : 4'b1001;
							assign node13300 = (inp[8]) ? node13784 : node13301;
								assign node13301 = (inp[14]) ? node13549 : node13302;
									assign node13302 = (inp[2]) ? node13428 : node13303;
										assign node13303 = (inp[6]) ? node13365 : node13304;
											assign node13304 = (inp[11]) ? node13336 : node13305;
												assign node13305 = (inp[1]) ? node13321 : node13306;
													assign node13306 = (inp[5]) ? node13314 : node13307;
														assign node13307 = (inp[15]) ? node13311 : node13308;
															assign node13308 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node13311 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node13314 = (inp[15]) ? node13318 : node13315;
															assign node13315 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node13318 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node13321 = (inp[13]) ? node13329 : node13322;
														assign node13322 = (inp[0]) ? node13326 : node13323;
															assign node13323 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node13326 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node13329 = (inp[5]) ? node13333 : node13330;
															assign node13330 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node13333 = (inp[15]) ? 4'b0000 : 4'b0000;
												assign node13336 = (inp[1]) ? node13352 : node13337;
													assign node13337 = (inp[0]) ? node13345 : node13338;
														assign node13338 = (inp[15]) ? node13342 : node13339;
															assign node13339 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node13342 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node13345 = (inp[5]) ? node13349 : node13346;
															assign node13346 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node13349 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node13352 = (inp[13]) ? node13360 : node13353;
														assign node13353 = (inp[15]) ? node13357 : node13354;
															assign node13354 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node13357 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node13360 = (inp[0]) ? node13362 : 4'b1000;
															assign node13362 = (inp[5]) ? 4'b1000 : 4'b1000;
											assign node13365 = (inp[11]) ? node13397 : node13366;
												assign node13366 = (inp[13]) ? node13382 : node13367;
													assign node13367 = (inp[0]) ? node13375 : node13368;
														assign node13368 = (inp[5]) ? node13372 : node13369;
															assign node13369 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node13372 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node13375 = (inp[5]) ? node13379 : node13376;
															assign node13376 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node13379 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node13382 = (inp[1]) ? node13390 : node13383;
														assign node13383 = (inp[5]) ? node13387 : node13384;
															assign node13384 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node13387 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node13390 = (inp[0]) ? node13394 : node13391;
															assign node13391 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node13394 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node13397 = (inp[1]) ? node13413 : node13398;
													assign node13398 = (inp[13]) ? node13406 : node13399;
														assign node13399 = (inp[0]) ? node13403 : node13400;
															assign node13400 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node13403 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node13406 = (inp[15]) ? node13410 : node13407;
															assign node13407 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node13410 = (inp[5]) ? 4'b1000 : 4'b1000;
													assign node13413 = (inp[13]) ? node13421 : node13414;
														assign node13414 = (inp[15]) ? node13418 : node13415;
															assign node13415 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node13418 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node13421 = (inp[15]) ? node13425 : node13422;
															assign node13422 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node13425 = (inp[0]) ? 4'b0010 : 4'b0000;
										assign node13428 = (inp[15]) ? node13488 : node13429;
											assign node13429 = (inp[6]) ? node13459 : node13430;
												assign node13430 = (inp[11]) ? node13444 : node13431;
													assign node13431 = (inp[1]) ? node13437 : node13432;
														assign node13432 = (inp[13]) ? node13434 : 4'b1011;
															assign node13434 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node13437 = (inp[0]) ? node13441 : node13438;
															assign node13438 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node13441 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node13444 = (inp[13]) ? node13452 : node13445;
														assign node13445 = (inp[1]) ? node13449 : node13446;
															assign node13446 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node13449 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node13452 = (inp[1]) ? node13456 : node13453;
															assign node13453 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node13456 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node13459 = (inp[11]) ? node13475 : node13460;
													assign node13460 = (inp[1]) ? node13468 : node13461;
														assign node13461 = (inp[13]) ? node13465 : node13462;
															assign node13462 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node13465 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node13468 = (inp[5]) ? node13472 : node13469;
															assign node13469 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node13472 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node13475 = (inp[13]) ? node13483 : node13476;
														assign node13476 = (inp[1]) ? node13480 : node13477;
															assign node13477 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node13480 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node13483 = (inp[0]) ? node13485 : 4'b0001;
															assign node13485 = (inp[5]) ? 4'b0011 : 4'b0001;
											assign node13488 = (inp[13]) ? node13520 : node13489;
												assign node13489 = (inp[11]) ? node13505 : node13490;
													assign node13490 = (inp[1]) ? node13498 : node13491;
														assign node13491 = (inp[6]) ? node13495 : node13492;
															assign node13492 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node13495 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node13498 = (inp[6]) ? node13502 : node13499;
															assign node13499 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node13502 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node13505 = (inp[6]) ? node13513 : node13506;
														assign node13506 = (inp[1]) ? node13510 : node13507;
															assign node13507 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node13510 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node13513 = (inp[1]) ? node13517 : node13514;
															assign node13514 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node13517 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node13520 = (inp[0]) ? node13536 : node13521;
													assign node13521 = (inp[5]) ? node13529 : node13522;
														assign node13522 = (inp[11]) ? node13526 : node13523;
															assign node13523 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node13526 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node13529 = (inp[6]) ? node13533 : node13530;
															assign node13530 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node13533 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node13536 = (inp[5]) ? node13542 : node13537;
														assign node13537 = (inp[11]) ? node13539 : 4'b0011;
															assign node13539 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node13542 = (inp[11]) ? node13546 : node13543;
															assign node13543 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node13546 = (inp[6]) ? 4'b0001 : 4'b1001;
									assign node13549 = (inp[15]) ? node13673 : node13550;
										assign node13550 = (inp[13]) ? node13610 : node13551;
											assign node13551 = (inp[5]) ? node13579 : node13552;
												assign node13552 = (inp[0]) ? node13564 : node13553;
													assign node13553 = (inp[6]) ? node13559 : node13554;
														assign node13554 = (inp[2]) ? 4'b1011 : node13555;
															assign node13555 = (inp[1]) ? 4'b0011 : 4'b0011;
														assign node13559 = (inp[2]) ? 4'b0011 : node13560;
															assign node13560 = (inp[11]) ? 4'b0011 : 4'b0011;
													assign node13564 = (inp[2]) ? node13572 : node13565;
														assign node13565 = (inp[11]) ? node13569 : node13566;
															assign node13566 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node13569 = (inp[1]) ? 4'b0001 : 4'b0001;
														assign node13572 = (inp[6]) ? node13576 : node13573;
															assign node13573 = (inp[11]) ? 4'b0001 : 4'b0001;
															assign node13576 = (inp[1]) ? 4'b0001 : 4'b0001;
												assign node13579 = (inp[0]) ? node13595 : node13580;
													assign node13580 = (inp[6]) ? node13588 : node13581;
														assign node13581 = (inp[2]) ? node13585 : node13582;
															assign node13582 = (inp[1]) ? 4'b0001 : 4'b0001;
															assign node13585 = (inp[1]) ? 4'b0001 : 4'b0001;
														assign node13588 = (inp[1]) ? node13592 : node13589;
															assign node13589 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node13592 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node13595 = (inp[1]) ? node13603 : node13596;
														assign node13596 = (inp[11]) ? node13600 : node13597;
															assign node13597 = (inp[6]) ? 4'b0011 : 4'b1011;
															assign node13600 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node13603 = (inp[2]) ? node13607 : node13604;
															assign node13604 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node13607 = (inp[11]) ? 4'b0011 : 4'b0011;
											assign node13610 = (inp[1]) ? node13642 : node13611;
												assign node13611 = (inp[11]) ? node13627 : node13612;
													assign node13612 = (inp[6]) ? node13620 : node13613;
														assign node13613 = (inp[5]) ? node13617 : node13614;
															assign node13614 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node13617 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node13620 = (inp[2]) ? node13624 : node13621;
															assign node13621 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node13624 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node13627 = (inp[6]) ? node13635 : node13628;
														assign node13628 = (inp[5]) ? node13632 : node13629;
															assign node13629 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node13632 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node13635 = (inp[2]) ? node13639 : node13636;
															assign node13636 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node13639 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node13642 = (inp[11]) ? node13658 : node13643;
													assign node13643 = (inp[6]) ? node13651 : node13644;
														assign node13644 = (inp[5]) ? node13648 : node13645;
															assign node13645 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node13648 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node13651 = (inp[2]) ? node13655 : node13652;
															assign node13652 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node13655 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node13658 = (inp[6]) ? node13666 : node13659;
														assign node13659 = (inp[5]) ? node13663 : node13660;
															assign node13660 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node13663 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node13666 = (inp[2]) ? node13670 : node13667;
															assign node13667 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node13670 = (inp[0]) ? 4'b0001 : 4'b0001;
										assign node13673 = (inp[11]) ? node13729 : node13674;
											assign node13674 = (inp[6]) ? node13706 : node13675;
												assign node13675 = (inp[1]) ? node13691 : node13676;
													assign node13676 = (inp[13]) ? node13684 : node13677;
														assign node13677 = (inp[0]) ? node13681 : node13678;
															assign node13678 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node13681 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node13684 = (inp[5]) ? node13688 : node13685;
															assign node13685 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node13688 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node13691 = (inp[13]) ? node13699 : node13692;
														assign node13692 = (inp[2]) ? node13696 : node13693;
															assign node13693 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node13696 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node13699 = (inp[5]) ? node13703 : node13700;
															assign node13700 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node13703 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node13706 = (inp[13]) ? node13722 : node13707;
													assign node13707 = (inp[1]) ? node13715 : node13708;
														assign node13708 = (inp[2]) ? node13712 : node13709;
															assign node13709 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node13712 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node13715 = (inp[2]) ? node13719 : node13716;
															assign node13716 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node13719 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node13722 = (inp[0]) ? node13726 : node13723;
														assign node13723 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node13726 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node13729 = (inp[6]) ? node13753 : node13730;
												assign node13730 = (inp[13]) ? node13746 : node13731;
													assign node13731 = (inp[1]) ? node13739 : node13732;
														assign node13732 = (inp[5]) ? node13736 : node13733;
															assign node13733 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node13736 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node13739 = (inp[2]) ? node13743 : node13740;
															assign node13740 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node13743 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node13746 = (inp[0]) ? node13750 : node13747;
														assign node13747 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node13750 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node13753 = (inp[13]) ? node13769 : node13754;
													assign node13754 = (inp[1]) ? node13762 : node13755;
														assign node13755 = (inp[0]) ? node13759 : node13756;
															assign node13756 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node13759 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node13762 = (inp[5]) ? node13766 : node13763;
															assign node13763 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node13766 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node13769 = (inp[2]) ? node13777 : node13770;
														assign node13770 = (inp[5]) ? node13774 : node13771;
															assign node13771 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node13774 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node13777 = (inp[0]) ? node13781 : node13778;
															assign node13778 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node13781 = (inp[5]) ? 4'b0001 : 4'b0011;
								assign node13784 = (inp[2]) ? node14022 : node13785;
									assign node13785 = (inp[14]) ? node13901 : node13786;
										assign node13786 = (inp[5]) ? node13844 : node13787;
											assign node13787 = (inp[1]) ? node13815 : node13788;
												assign node13788 = (inp[13]) ? node13804 : node13789;
													assign node13789 = (inp[15]) ? node13797 : node13790;
														assign node13790 = (inp[0]) ? node13794 : node13791;
															assign node13791 = (inp[11]) ? 4'b0011 : 4'b0011;
															assign node13794 = (inp[6]) ? 4'b0001 : 4'b0001;
														assign node13797 = (inp[0]) ? node13801 : node13798;
															assign node13798 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node13801 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node13804 = (inp[11]) ? node13810 : node13805;
														assign node13805 = (inp[6]) ? node13807 : 4'b0001;
															assign node13807 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node13810 = (inp[6]) ? 4'b0001 : node13811;
															assign node13811 = (inp[0]) ? 4'b1001 : 4'b1001;
												assign node13815 = (inp[0]) ? node13831 : node13816;
													assign node13816 = (inp[15]) ? node13824 : node13817;
														assign node13817 = (inp[6]) ? node13821 : node13818;
															assign node13818 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node13821 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node13824 = (inp[11]) ? node13828 : node13825;
															assign node13825 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node13828 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node13831 = (inp[15]) ? node13839 : node13832;
														assign node13832 = (inp[11]) ? node13836 : node13833;
															assign node13833 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node13836 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node13839 = (inp[11]) ? 4'b0011 : node13840;
															assign node13840 = (inp[6]) ? 4'b1011 : 4'b0011;
											assign node13844 = (inp[15]) ? node13874 : node13845;
												assign node13845 = (inp[0]) ? node13861 : node13846;
													assign node13846 = (inp[11]) ? node13854 : node13847;
														assign node13847 = (inp[6]) ? node13851 : node13848;
															assign node13848 = (inp[13]) ? 4'b0001 : 4'b0001;
															assign node13851 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node13854 = (inp[6]) ? node13858 : node13855;
															assign node13855 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node13858 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node13861 = (inp[11]) ? node13867 : node13862;
														assign node13862 = (inp[6]) ? node13864 : 4'b0011;
															assign node13864 = (inp[1]) ? 4'b1011 : 4'b0011;
														assign node13867 = (inp[6]) ? node13871 : node13868;
															assign node13868 = (inp[1]) ? 4'b1011 : 4'b0011;
															assign node13871 = (inp[1]) ? 4'b0011 : 4'b0011;
												assign node13874 = (inp[0]) ? node13890 : node13875;
													assign node13875 = (inp[11]) ? node13883 : node13876;
														assign node13876 = (inp[6]) ? node13880 : node13877;
															assign node13877 = (inp[1]) ? 4'b0011 : 4'b0011;
															assign node13880 = (inp[1]) ? 4'b1011 : 4'b0011;
														assign node13883 = (inp[6]) ? node13887 : node13884;
															assign node13884 = (inp[1]) ? 4'b1011 : 4'b0011;
															assign node13887 = (inp[1]) ? 4'b0011 : 4'b0011;
													assign node13890 = (inp[13]) ? node13896 : node13891;
														assign node13891 = (inp[1]) ? node13893 : 4'b0001;
															assign node13893 = (inp[6]) ? 4'b0001 : 4'b0001;
														assign node13896 = (inp[1]) ? 4'b0001 : node13897;
															assign node13897 = (inp[6]) ? 4'b1001 : 4'b0001;
										assign node13901 = (inp[1]) ? node13959 : node13902;
											assign node13902 = (inp[11]) ? node13930 : node13903;
												assign node13903 = (inp[13]) ? node13917 : node13904;
													assign node13904 = (inp[6]) ? node13912 : node13905;
														assign node13905 = (inp[5]) ? node13909 : node13906;
															assign node13906 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node13909 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node13912 = (inp[15]) ? node13914 : 4'b0000;
															assign node13914 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node13917 = (inp[6]) ? node13923 : node13918;
														assign node13918 = (inp[0]) ? 4'b0010 : node13919;
															assign node13919 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node13923 = (inp[15]) ? node13927 : node13924;
															assign node13924 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node13927 = (inp[5]) ? 4'b1000 : 4'b1000;
												assign node13930 = (inp[13]) ? node13944 : node13931;
													assign node13931 = (inp[6]) ? node13939 : node13932;
														assign node13932 = (inp[5]) ? node13936 : node13933;
															assign node13933 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node13936 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node13939 = (inp[15]) ? node13941 : 4'b1010;
															assign node13941 = (inp[5]) ? 4'b1000 : 4'b1000;
													assign node13944 = (inp[6]) ? node13952 : node13945;
														assign node13945 = (inp[15]) ? node13949 : node13946;
															assign node13946 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node13949 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node13952 = (inp[0]) ? node13956 : node13953;
															assign node13953 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node13956 = (inp[5]) ? 4'b0000 : 4'b0000;
											assign node13959 = (inp[0]) ? node13991 : node13960;
												assign node13960 = (inp[6]) ? node13976 : node13961;
													assign node13961 = (inp[11]) ? node13969 : node13962;
														assign node13962 = (inp[5]) ? node13966 : node13963;
															assign node13963 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node13966 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node13969 = (inp[15]) ? node13973 : node13970;
															assign node13970 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node13973 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node13976 = (inp[11]) ? node13984 : node13977;
														assign node13977 = (inp[15]) ? node13981 : node13978;
															assign node13978 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node13981 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node13984 = (inp[15]) ? node13988 : node13985;
															assign node13985 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node13988 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node13991 = (inp[11]) ? node14007 : node13992;
													assign node13992 = (inp[6]) ? node14000 : node13993;
														assign node13993 = (inp[5]) ? node13997 : node13994;
															assign node13994 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node13997 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node14000 = (inp[13]) ? node14004 : node14001;
															assign node14001 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node14004 = (inp[5]) ? 4'b1000 : 4'b1000;
													assign node14007 = (inp[6]) ? node14015 : node14008;
														assign node14008 = (inp[5]) ? node14012 : node14009;
															assign node14009 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node14012 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node14015 = (inp[5]) ? node14019 : node14016;
															assign node14016 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node14019 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node14022 = (inp[13]) ? node14142 : node14023;
										assign node14023 = (inp[11]) ? node14083 : node14024;
											assign node14024 = (inp[1]) ? node14052 : node14025;
												assign node14025 = (inp[6]) ? node14039 : node14026;
													assign node14026 = (inp[14]) ? node14032 : node14027;
														assign node14027 = (inp[5]) ? node14029 : 4'b1010;
															assign node14029 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node14032 = (inp[5]) ? node14036 : node14033;
															assign node14033 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node14036 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node14039 = (inp[15]) ? node14047 : node14040;
														assign node14040 = (inp[0]) ? node14044 : node14041;
															assign node14041 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node14044 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node14047 = (inp[14]) ? 4'b0010 : node14048;
															assign node14048 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node14052 = (inp[6]) ? node14068 : node14053;
													assign node14053 = (inp[15]) ? node14061 : node14054;
														assign node14054 = (inp[14]) ? node14058 : node14055;
															assign node14055 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node14058 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node14061 = (inp[5]) ? node14065 : node14062;
															assign node14062 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node14065 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node14068 = (inp[15]) ? node14076 : node14069;
														assign node14069 = (inp[14]) ? node14073 : node14070;
															assign node14070 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node14073 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node14076 = (inp[14]) ? node14080 : node14077;
															assign node14077 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node14080 = (inp[5]) ? 4'b1000 : 4'b1000;
											assign node14083 = (inp[1]) ? node14111 : node14084;
												assign node14084 = (inp[6]) ? node14100 : node14085;
													assign node14085 = (inp[0]) ? node14093 : node14086;
														assign node14086 = (inp[15]) ? node14090 : node14087;
															assign node14087 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node14090 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node14093 = (inp[15]) ? node14097 : node14094;
															assign node14094 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node14097 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node14100 = (inp[14]) ? node14106 : node14101;
														assign node14101 = (inp[0]) ? node14103 : 4'b1010;
															assign node14103 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node14106 = (inp[5]) ? 4'b1000 : node14107;
															assign node14107 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node14111 = (inp[6]) ? node14127 : node14112;
													assign node14112 = (inp[0]) ? node14120 : node14113;
														assign node14113 = (inp[14]) ? node14117 : node14114;
															assign node14114 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node14117 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node14120 = (inp[15]) ? node14124 : node14121;
															assign node14121 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node14124 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node14127 = (inp[0]) ? node14135 : node14128;
														assign node14128 = (inp[15]) ? node14132 : node14129;
															assign node14129 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node14132 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node14135 = (inp[14]) ? node14139 : node14136;
															assign node14136 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node14139 = (inp[15]) ? 4'b0000 : 4'b0000;
										assign node14142 = (inp[5]) ? node14204 : node14143;
											assign node14143 = (inp[15]) ? node14173 : node14144;
												assign node14144 = (inp[0]) ? node14158 : node14145;
													assign node14145 = (inp[14]) ? node14153 : node14146;
														assign node14146 = (inp[6]) ? node14150 : node14147;
															assign node14147 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node14150 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node14153 = (inp[1]) ? 4'b0010 : node14154;
															assign node14154 = (inp[6]) ? 4'b0010 : 4'b0010;
													assign node14158 = (inp[14]) ? node14166 : node14159;
														assign node14159 = (inp[6]) ? node14163 : node14160;
															assign node14160 = (inp[11]) ? 4'b1000 : 4'b0000;
															assign node14163 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node14166 = (inp[11]) ? node14170 : node14167;
															assign node14167 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node14170 = (inp[6]) ? 4'b0000 : 4'b1000;
												assign node14173 = (inp[0]) ? node14189 : node14174;
													assign node14174 = (inp[14]) ? node14182 : node14175;
														assign node14175 = (inp[6]) ? node14179 : node14176;
															assign node14176 = (inp[11]) ? 4'b1000 : 4'b0000;
															assign node14179 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node14182 = (inp[11]) ? node14186 : node14183;
															assign node14183 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node14186 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node14189 = (inp[14]) ? node14197 : node14190;
														assign node14190 = (inp[1]) ? node14194 : node14191;
															assign node14191 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node14194 = (inp[11]) ? 4'b0010 : 4'b0010;
														assign node14197 = (inp[1]) ? node14201 : node14198;
															assign node14198 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node14201 = (inp[6]) ? 4'b0010 : 4'b0010;
											assign node14204 = (inp[15]) ? node14236 : node14205;
												assign node14205 = (inp[0]) ? node14221 : node14206;
													assign node14206 = (inp[14]) ? node14214 : node14207;
														assign node14207 = (inp[11]) ? node14211 : node14208;
															assign node14208 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node14211 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node14214 = (inp[1]) ? node14218 : node14215;
															assign node14215 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node14218 = (inp[6]) ? 4'b0000 : 4'b0000;
													assign node14221 = (inp[1]) ? node14229 : node14222;
														assign node14222 = (inp[6]) ? node14226 : node14223;
															assign node14223 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node14226 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node14229 = (inp[6]) ? node14233 : node14230;
															assign node14230 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node14233 = (inp[11]) ? 4'b0010 : 4'b1010;
												assign node14236 = (inp[0]) ? node14244 : node14237;
													assign node14237 = (inp[11]) ? node14241 : node14238;
														assign node14238 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node14241 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node14244 = (inp[1]) ? node14252 : node14245;
														assign node14245 = (inp[6]) ? node14249 : node14246;
															assign node14246 = (inp[11]) ? 4'b1000 : 4'b0000;
															assign node14249 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node14252 = (inp[14]) ? node14256 : node14253;
															assign node14253 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node14256 = (inp[6]) ? 4'b0000 : 4'b0000;
			assign node14259 = (inp[10]) ? node21487 : node14260;
				assign node14260 = (inp[12]) ? node17882 : node14261;
					assign node14261 = (inp[6]) ? node16067 : node14262;
						assign node14262 = (inp[11]) ? node15182 : node14263;
							assign node14263 = (inp[1]) ? node14729 : node14264;
								assign node14264 = (inp[13]) ? node14514 : node14265;
									assign node14265 = (inp[5]) ? node14393 : node14266;
										assign node14266 = (inp[2]) ? node14330 : node14267;
											assign node14267 = (inp[3]) ? node14299 : node14268;
												assign node14268 = (inp[14]) ? node14284 : node14269;
													assign node14269 = (inp[0]) ? node14277 : node14270;
														assign node14270 = (inp[15]) ? node14274 : node14271;
															assign node14271 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node14274 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node14277 = (inp[15]) ? node14281 : node14278;
															assign node14278 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node14281 = (inp[8]) ? 4'b1010 : 4'b1010;
													assign node14284 = (inp[7]) ? node14292 : node14285;
														assign node14285 = (inp[8]) ? node14289 : node14286;
															assign node14286 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node14289 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node14292 = (inp[8]) ? node14296 : node14293;
															assign node14293 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node14296 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node14299 = (inp[14]) ? node14315 : node14300;
													assign node14300 = (inp[7]) ? node14308 : node14301;
														assign node14301 = (inp[8]) ? node14305 : node14302;
															assign node14302 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node14305 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node14308 = (inp[8]) ? node14312 : node14309;
															assign node14309 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node14312 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node14315 = (inp[8]) ? node14323 : node14316;
														assign node14316 = (inp[7]) ? node14320 : node14317;
															assign node14317 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node14320 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node14323 = (inp[7]) ? node14327 : node14324;
															assign node14324 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node14327 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node14330 = (inp[14]) ? node14362 : node14331;
												assign node14331 = (inp[7]) ? node14347 : node14332;
													assign node14332 = (inp[8]) ? node14340 : node14333;
														assign node14333 = (inp[15]) ? node14337 : node14334;
															assign node14334 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node14337 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node14340 = (inp[0]) ? node14344 : node14341;
															assign node14341 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node14344 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node14347 = (inp[8]) ? node14355 : node14348;
														assign node14348 = (inp[15]) ? node14352 : node14349;
															assign node14349 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node14352 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node14355 = (inp[3]) ? node14359 : node14356;
															assign node14356 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node14359 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node14362 = (inp[15]) ? node14378 : node14363;
													assign node14363 = (inp[0]) ? node14371 : node14364;
														assign node14364 = (inp[7]) ? node14368 : node14365;
															assign node14365 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node14368 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node14371 = (inp[8]) ? node14375 : node14372;
															assign node14372 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node14375 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node14378 = (inp[0]) ? node14386 : node14379;
														assign node14379 = (inp[8]) ? node14383 : node14380;
															assign node14380 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node14383 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node14386 = (inp[7]) ? node14390 : node14387;
															assign node14387 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node14390 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node14393 = (inp[0]) ? node14453 : node14394;
											assign node14394 = (inp[14]) ? node14426 : node14395;
												assign node14395 = (inp[15]) ? node14411 : node14396;
													assign node14396 = (inp[3]) ? node14404 : node14397;
														assign node14397 = (inp[8]) ? node14401 : node14398;
															assign node14398 = (inp[2]) ? 4'b1010 : 4'b1010;
															assign node14401 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node14404 = (inp[2]) ? node14408 : node14405;
															assign node14405 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node14408 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node14411 = (inp[3]) ? node14419 : node14412;
														assign node14412 = (inp[2]) ? node14416 : node14413;
															assign node14413 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node14416 = (inp[7]) ? 4'b1000 : 4'b1000;
														assign node14419 = (inp[2]) ? node14423 : node14420;
															assign node14420 = (inp[8]) ? 4'b1010 : 4'b1010;
															assign node14423 = (inp[7]) ? 4'b1010 : 4'b1010;
												assign node14426 = (inp[15]) ? node14440 : node14427;
													assign node14427 = (inp[3]) ? node14433 : node14428;
														assign node14428 = (inp[8]) ? 4'b1010 : node14429;
															assign node14429 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node14433 = (inp[8]) ? node14437 : node14434;
															assign node14434 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node14437 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node14440 = (inp[3]) ? node14448 : node14441;
														assign node14441 = (inp[8]) ? node14445 : node14442;
															assign node14442 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node14445 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node14448 = (inp[8]) ? node14450 : 4'b1010;
															assign node14450 = (inp[7]) ? 4'b1010 : 4'b1011;
											assign node14453 = (inp[8]) ? node14485 : node14454;
												assign node14454 = (inp[7]) ? node14470 : node14455;
													assign node14455 = (inp[2]) ? node14463 : node14456;
														assign node14456 = (inp[14]) ? node14460 : node14457;
															assign node14457 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node14460 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node14463 = (inp[3]) ? node14467 : node14464;
															assign node14464 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node14467 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node14470 = (inp[2]) ? node14478 : node14471;
														assign node14471 = (inp[14]) ? node14475 : node14472;
															assign node14472 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node14475 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node14478 = (inp[3]) ? node14482 : node14479;
															assign node14479 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node14482 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node14485 = (inp[7]) ? node14501 : node14486;
													assign node14486 = (inp[2]) ? node14494 : node14487;
														assign node14487 = (inp[14]) ? node14491 : node14488;
															assign node14488 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node14491 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node14494 = (inp[3]) ? node14498 : node14495;
															assign node14495 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node14498 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node14501 = (inp[2]) ? node14507 : node14502;
														assign node14502 = (inp[14]) ? 4'b1000 : node14503;
															assign node14503 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node14507 = (inp[3]) ? node14511 : node14508;
															assign node14508 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node14511 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node14514 = (inp[8]) ? node14620 : node14515;
										assign node14515 = (inp[7]) ? node14569 : node14516;
											assign node14516 = (inp[2]) ? node14546 : node14517;
												assign node14517 = (inp[14]) ? node14533 : node14518;
													assign node14518 = (inp[3]) ? node14526 : node14519;
														assign node14519 = (inp[0]) ? node14523 : node14520;
															assign node14520 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node14523 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node14526 = (inp[5]) ? node14530 : node14527;
															assign node14527 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node14530 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node14533 = (inp[5]) ? node14539 : node14534;
														assign node14534 = (inp[15]) ? 4'b1010 : node14535;
															assign node14535 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node14539 = (inp[15]) ? node14543 : node14540;
															assign node14540 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node14543 = (inp[3]) ? 4'b1000 : 4'b1000;
												assign node14546 = (inp[15]) ? node14558 : node14547;
													assign node14547 = (inp[0]) ? node14553 : node14548;
														assign node14548 = (inp[5]) ? node14550 : 4'b1010;
															assign node14550 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node14553 = (inp[3]) ? node14555 : 4'b1000;
															assign node14555 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node14558 = (inp[0]) ? node14564 : node14559;
														assign node14559 = (inp[5]) ? node14561 : 4'b1000;
															assign node14561 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node14564 = (inp[5]) ? node14566 : 4'b1010;
															assign node14566 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node14569 = (inp[2]) ? node14597 : node14570;
												assign node14570 = (inp[14]) ? node14584 : node14571;
													assign node14571 = (inp[15]) ? node14577 : node14572;
														assign node14572 = (inp[5]) ? node14574 : 4'b1010;
															assign node14574 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node14577 = (inp[0]) ? node14581 : node14578;
															assign node14578 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node14581 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node14584 = (inp[3]) ? node14592 : node14585;
														assign node14585 = (inp[0]) ? node14589 : node14586;
															assign node14586 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node14589 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node14592 = (inp[15]) ? 4'b0011 : node14593;
															assign node14593 = (inp[0]) ? 4'b0001 : 4'b0001;
												assign node14597 = (inp[15]) ? node14609 : node14598;
													assign node14598 = (inp[0]) ? node14604 : node14599;
														assign node14599 = (inp[3]) ? node14601 : 4'b0011;
															assign node14601 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node14604 = (inp[3]) ? node14606 : 4'b0001;
															assign node14606 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node14609 = (inp[0]) ? node14615 : node14610;
														assign node14610 = (inp[5]) ? node14612 : 4'b0001;
															assign node14612 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node14615 = (inp[5]) ? node14617 : 4'b0011;
															assign node14617 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node14620 = (inp[7]) ? node14676 : node14621;
											assign node14621 = (inp[14]) ? node14653 : node14622;
												assign node14622 = (inp[2]) ? node14638 : node14623;
													assign node14623 = (inp[5]) ? node14631 : node14624;
														assign node14624 = (inp[15]) ? node14628 : node14625;
															assign node14625 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node14628 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node14631 = (inp[3]) ? node14635 : node14632;
															assign node14632 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node14635 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node14638 = (inp[0]) ? node14646 : node14639;
														assign node14639 = (inp[15]) ? node14643 : node14640;
															assign node14640 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node14643 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node14646 = (inp[15]) ? node14650 : node14647;
															assign node14647 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node14650 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node14653 = (inp[5]) ? node14661 : node14654;
													assign node14654 = (inp[0]) ? node14658 : node14655;
														assign node14655 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node14658 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node14661 = (inp[15]) ? node14669 : node14662;
														assign node14662 = (inp[0]) ? node14666 : node14663;
															assign node14663 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node14666 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node14669 = (inp[0]) ? node14673 : node14670;
															assign node14670 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node14673 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node14676 = (inp[14]) ? node14706 : node14677;
												assign node14677 = (inp[2]) ? node14693 : node14678;
													assign node14678 = (inp[0]) ? node14686 : node14679;
														assign node14679 = (inp[15]) ? node14683 : node14680;
															assign node14680 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node14683 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node14686 = (inp[15]) ? node14690 : node14687;
															assign node14687 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node14690 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node14693 = (inp[5]) ? node14701 : node14694;
														assign node14694 = (inp[0]) ? node14698 : node14695;
															assign node14695 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node14698 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node14701 = (inp[0]) ? node14703 : 4'b0010;
															assign node14703 = (inp[15]) ? 4'b0000 : 4'b0000;
												assign node14706 = (inp[0]) ? node14718 : node14707;
													assign node14707 = (inp[15]) ? node14713 : node14708;
														assign node14708 = (inp[3]) ? node14710 : 4'b0010;
															assign node14710 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node14713 = (inp[5]) ? node14715 : 4'b0000;
															assign node14715 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node14718 = (inp[15]) ? node14724 : node14719;
														assign node14719 = (inp[3]) ? node14721 : 4'b0000;
															assign node14721 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node14724 = (inp[5]) ? node14726 : 4'b0010;
															assign node14726 = (inp[3]) ? 4'b0000 : 4'b0010;
								assign node14729 = (inp[13]) ? node14951 : node14730;
									assign node14730 = (inp[7]) ? node14844 : node14731;
										assign node14731 = (inp[8]) ? node14791 : node14732;
											assign node14732 = (inp[14]) ? node14760 : node14733;
												assign node14733 = (inp[2]) ? node14747 : node14734;
													assign node14734 = (inp[0]) ? node14740 : node14735;
														assign node14735 = (inp[15]) ? node14737 : 4'b1011;
															assign node14737 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node14740 = (inp[15]) ? node14744 : node14741;
															assign node14741 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node14744 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node14747 = (inp[3]) ? node14753 : node14748;
														assign node14748 = (inp[15]) ? 4'b1000 : node14749;
															assign node14749 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node14753 = (inp[0]) ? node14757 : node14754;
															assign node14754 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node14757 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node14760 = (inp[2]) ? node14776 : node14761;
													assign node14761 = (inp[5]) ? node14769 : node14762;
														assign node14762 = (inp[3]) ? node14766 : node14763;
															assign node14763 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node14766 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node14769 = (inp[15]) ? node14773 : node14770;
															assign node14770 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node14773 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node14776 = (inp[3]) ? node14784 : node14777;
														assign node14777 = (inp[0]) ? node14781 : node14778;
															assign node14778 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node14781 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node14784 = (inp[15]) ? node14788 : node14785;
															assign node14785 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node14788 = (inp[5]) ? 4'b1000 : 4'b1000;
											assign node14791 = (inp[14]) ? node14819 : node14792;
												assign node14792 = (inp[2]) ? node14806 : node14793;
													assign node14793 = (inp[15]) ? node14799 : node14794;
														assign node14794 = (inp[0]) ? node14796 : 4'b1010;
															assign node14796 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node14799 = (inp[0]) ? node14803 : node14800;
															assign node14800 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node14803 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node14806 = (inp[5]) ? node14814 : node14807;
														assign node14807 = (inp[3]) ? node14811 : node14808;
															assign node14808 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node14811 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node14814 = (inp[3]) ? node14816 : 4'b0001;
															assign node14816 = (inp[0]) ? 4'b0001 : 4'b0001;
												assign node14819 = (inp[2]) ? node14831 : node14820;
													assign node14820 = (inp[0]) ? node14826 : node14821;
														assign node14821 = (inp[15]) ? 4'b0001 : node14822;
															assign node14822 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node14826 = (inp[15]) ? 4'b0011 : node14827;
															assign node14827 = (inp[3]) ? 4'b0001 : 4'b0001;
													assign node14831 = (inp[5]) ? node14839 : node14832;
														assign node14832 = (inp[15]) ? node14836 : node14833;
															assign node14833 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node14836 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node14839 = (inp[15]) ? node14841 : 4'b0011;
															assign node14841 = (inp[0]) ? 4'b0011 : 4'b0001;
										assign node14844 = (inp[8]) ? node14896 : node14845;
											assign node14845 = (inp[14]) ? node14873 : node14846;
												assign node14846 = (inp[2]) ? node14860 : node14847;
													assign node14847 = (inp[15]) ? node14853 : node14848;
														assign node14848 = (inp[0]) ? node14850 : 4'b1010;
															assign node14850 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node14853 = (inp[0]) ? node14857 : node14854;
															assign node14854 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node14857 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node14860 = (inp[3]) ? node14868 : node14861;
														assign node14861 = (inp[15]) ? node14865 : node14862;
															assign node14862 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node14865 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node14868 = (inp[15]) ? node14870 : 4'b0011;
															assign node14870 = (inp[5]) ? 4'b0001 : 4'b0001;
												assign node14873 = (inp[0]) ? node14885 : node14874;
													assign node14874 = (inp[15]) ? node14880 : node14875;
														assign node14875 = (inp[5]) ? node14877 : 4'b0011;
															assign node14877 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node14880 = (inp[3]) ? node14882 : 4'b0001;
															assign node14882 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node14885 = (inp[15]) ? node14891 : node14886;
														assign node14886 = (inp[5]) ? node14888 : 4'b0001;
															assign node14888 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node14891 = (inp[3]) ? node14893 : 4'b0011;
															assign node14893 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node14896 = (inp[14]) ? node14928 : node14897;
												assign node14897 = (inp[2]) ? node14913 : node14898;
													assign node14898 = (inp[5]) ? node14906 : node14899;
														assign node14899 = (inp[15]) ? node14903 : node14900;
															assign node14900 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node14903 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node14906 = (inp[3]) ? node14910 : node14907;
															assign node14907 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node14910 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node14913 = (inp[3]) ? node14921 : node14914;
														assign node14914 = (inp[0]) ? node14918 : node14915;
															assign node14915 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node14918 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node14921 = (inp[15]) ? node14925 : node14922;
															assign node14922 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node14925 = (inp[5]) ? 4'b0000 : 4'b0000;
												assign node14928 = (inp[15]) ? node14940 : node14929;
													assign node14929 = (inp[0]) ? node14935 : node14930;
														assign node14930 = (inp[3]) ? node14932 : 4'b0010;
															assign node14932 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node14935 = (inp[5]) ? node14937 : 4'b0000;
															assign node14937 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node14940 = (inp[0]) ? node14946 : node14941;
														assign node14941 = (inp[3]) ? node14943 : 4'b0000;
															assign node14943 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node14946 = (inp[3]) ? node14948 : 4'b0010;
															assign node14948 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node14951 = (inp[0]) ? node15069 : node14952;
										assign node14952 = (inp[15]) ? node15016 : node14953;
											assign node14953 = (inp[5]) ? node14985 : node14954;
												assign node14954 = (inp[14]) ? node14970 : node14955;
													assign node14955 = (inp[7]) ? node14963 : node14956;
														assign node14956 = (inp[8]) ? node14960 : node14957;
															assign node14957 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node14960 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node14963 = (inp[2]) ? node14967 : node14964;
															assign node14964 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node14967 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node14970 = (inp[3]) ? node14978 : node14971;
														assign node14971 = (inp[8]) ? node14975 : node14972;
															assign node14972 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node14975 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node14978 = (inp[2]) ? node14982 : node14979;
															assign node14979 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node14982 = (inp[8]) ? 4'b0010 : 4'b0010;
												assign node14985 = (inp[3]) ? node15001 : node14986;
													assign node14986 = (inp[2]) ? node14994 : node14987;
														assign node14987 = (inp[14]) ? node14991 : node14988;
															assign node14988 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node14991 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node14994 = (inp[7]) ? node14998 : node14995;
															assign node14995 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node14998 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node15001 = (inp[8]) ? node15009 : node15002;
														assign node15002 = (inp[7]) ? node15006 : node15003;
															assign node15003 = (inp[14]) ? 4'b0000 : 4'b0000;
															assign node15006 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node15009 = (inp[7]) ? node15013 : node15010;
															assign node15010 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node15013 = (inp[2]) ? 4'b0000 : 4'b0000;
											assign node15016 = (inp[3]) ? node15040 : node15017;
												assign node15017 = (inp[7]) ? node15029 : node15018;
													assign node15018 = (inp[8]) ? node15024 : node15019;
														assign node15019 = (inp[14]) ? 4'b0000 : node15020;
															assign node15020 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node15024 = (inp[14]) ? 4'b0001 : node15025;
															assign node15025 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node15029 = (inp[8]) ? node15035 : node15030;
														assign node15030 = (inp[2]) ? 4'b0001 : node15031;
															assign node15031 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node15035 = (inp[14]) ? 4'b0000 : node15036;
															assign node15036 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node15040 = (inp[5]) ? node15056 : node15041;
													assign node15041 = (inp[14]) ? node15049 : node15042;
														assign node15042 = (inp[7]) ? node15046 : node15043;
															assign node15043 = (inp[2]) ? 4'b0000 : 4'b0000;
															assign node15046 = (inp[2]) ? 4'b0000 : 4'b0000;
														assign node15049 = (inp[2]) ? node15053 : node15050;
															assign node15050 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node15053 = (inp[7]) ? 4'b0000 : 4'b0000;
													assign node15056 = (inp[7]) ? node15064 : node15057;
														assign node15057 = (inp[8]) ? node15061 : node15058;
															assign node15058 = (inp[14]) ? 4'b0010 : 4'b0010;
															assign node15061 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node15064 = (inp[8]) ? node15066 : 4'b0011;
															assign node15066 = (inp[2]) ? 4'b0010 : 4'b0010;
										assign node15069 = (inp[15]) ? node15129 : node15070;
											assign node15070 = (inp[3]) ? node15100 : node15071;
												assign node15071 = (inp[5]) ? node15085 : node15072;
													assign node15072 = (inp[7]) ? node15078 : node15073;
														assign node15073 = (inp[8]) ? 4'b0001 : node15074;
															assign node15074 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node15078 = (inp[2]) ? node15082 : node15079;
															assign node15079 = (inp[14]) ? 4'b0000 : 4'b0000;
															assign node15082 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node15085 = (inp[8]) ? node15093 : node15086;
														assign node15086 = (inp[7]) ? node15090 : node15087;
															assign node15087 = (inp[2]) ? 4'b0000 : 4'b0000;
															assign node15090 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node15093 = (inp[7]) ? node15097 : node15094;
															assign node15094 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node15097 = (inp[2]) ? 4'b0000 : 4'b0000;
												assign node15100 = (inp[5]) ? node15116 : node15101;
													assign node15101 = (inp[2]) ? node15109 : node15102;
														assign node15102 = (inp[7]) ? node15106 : node15103;
															assign node15103 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node15106 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node15109 = (inp[8]) ? node15113 : node15110;
															assign node15110 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node15113 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node15116 = (inp[2]) ? node15122 : node15117;
														assign node15117 = (inp[14]) ? node15119 : 4'b0011;
															assign node15119 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node15122 = (inp[8]) ? node15126 : node15123;
															assign node15123 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node15126 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node15129 = (inp[5]) ? node15153 : node15130;
												assign node15130 = (inp[8]) ? node15142 : node15131;
													assign node15131 = (inp[7]) ? node15137 : node15132;
														assign node15132 = (inp[14]) ? 4'b0010 : node15133;
															assign node15133 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node15137 = (inp[14]) ? 4'b0011 : node15138;
															assign node15138 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node15142 = (inp[7]) ? node15148 : node15143;
														assign node15143 = (inp[2]) ? 4'b0011 : node15144;
															assign node15144 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node15148 = (inp[2]) ? 4'b0010 : node15149;
															assign node15149 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node15153 = (inp[3]) ? node15169 : node15154;
													assign node15154 = (inp[2]) ? node15162 : node15155;
														assign node15155 = (inp[8]) ? node15159 : node15156;
															assign node15156 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node15159 = (inp[14]) ? 4'b0010 : 4'b0010;
														assign node15162 = (inp[14]) ? node15166 : node15163;
															assign node15163 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node15166 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node15169 = (inp[8]) ? node15177 : node15170;
														assign node15170 = (inp[7]) ? node15174 : node15171;
															assign node15171 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node15174 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node15177 = (inp[7]) ? node15179 : 4'b0001;
															assign node15179 = (inp[14]) ? 4'b0000 : 4'b0001;
							assign node15182 = (inp[1]) ? node15630 : node15183;
								assign node15183 = (inp[13]) ? node15409 : node15184;
									assign node15184 = (inp[8]) ? node15302 : node15185;
										assign node15185 = (inp[7]) ? node15243 : node15186;
											assign node15186 = (inp[14]) ? node15214 : node15187;
												assign node15187 = (inp[2]) ? node15201 : node15188;
													assign node15188 = (inp[15]) ? node15196 : node15189;
														assign node15189 = (inp[0]) ? node15193 : node15190;
															assign node15190 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node15193 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node15196 = (inp[0]) ? node15198 : 4'b0001;
															assign node15198 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node15201 = (inp[15]) ? node15209 : node15202;
														assign node15202 = (inp[0]) ? node15206 : node15203;
															assign node15203 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node15206 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node15209 = (inp[0]) ? 4'b0010 : node15210;
															assign node15210 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node15214 = (inp[5]) ? node15228 : node15215;
													assign node15215 = (inp[2]) ? node15221 : node15216;
														assign node15216 = (inp[15]) ? 4'b0010 : node15217;
															assign node15217 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node15221 = (inp[15]) ? node15225 : node15222;
															assign node15222 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node15225 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node15228 = (inp[15]) ? node15236 : node15229;
														assign node15229 = (inp[3]) ? node15233 : node15230;
															assign node15230 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node15233 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node15236 = (inp[3]) ? node15240 : node15237;
															assign node15237 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node15240 = (inp[0]) ? 4'b0000 : 4'b0010;
											assign node15243 = (inp[2]) ? node15273 : node15244;
												assign node15244 = (inp[14]) ? node15260 : node15245;
													assign node15245 = (inp[15]) ? node15253 : node15246;
														assign node15246 = (inp[0]) ? node15250 : node15247;
															assign node15247 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node15250 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node15253 = (inp[0]) ? node15257 : node15254;
															assign node15254 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node15257 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node15260 = (inp[0]) ? node15266 : node15261;
														assign node15261 = (inp[5]) ? node15263 : 4'b0011;
															assign node15263 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node15266 = (inp[15]) ? node15270 : node15267;
															assign node15267 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node15270 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node15273 = (inp[14]) ? node15287 : node15274;
													assign node15274 = (inp[15]) ? node15280 : node15275;
														assign node15275 = (inp[0]) ? 4'b0001 : node15276;
															assign node15276 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node15280 = (inp[0]) ? node15284 : node15281;
															assign node15281 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node15284 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node15287 = (inp[5]) ? node15295 : node15288;
														assign node15288 = (inp[0]) ? node15292 : node15289;
															assign node15289 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node15292 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node15295 = (inp[3]) ? node15299 : node15296;
															assign node15296 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node15299 = (inp[0]) ? 4'b0001 : 4'b0011;
										assign node15302 = (inp[7]) ? node15358 : node15303;
											assign node15303 = (inp[14]) ? node15335 : node15304;
												assign node15304 = (inp[2]) ? node15320 : node15305;
													assign node15305 = (inp[5]) ? node15313 : node15306;
														assign node15306 = (inp[0]) ? node15310 : node15307;
															assign node15307 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node15310 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node15313 = (inp[3]) ? node15317 : node15314;
															assign node15314 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node15317 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node15320 = (inp[3]) ? node15328 : node15321;
														assign node15321 = (inp[5]) ? node15325 : node15322;
															assign node15322 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node15325 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node15328 = (inp[15]) ? node15332 : node15329;
															assign node15329 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node15332 = (inp[5]) ? 4'b0001 : 4'b0001;
												assign node15335 = (inp[0]) ? node15347 : node15336;
													assign node15336 = (inp[15]) ? node15342 : node15337;
														assign node15337 = (inp[3]) ? node15339 : 4'b0011;
															assign node15339 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node15342 = (inp[5]) ? node15344 : 4'b0001;
															assign node15344 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node15347 = (inp[15]) ? node15353 : node15348;
														assign node15348 = (inp[5]) ? node15350 : 4'b0001;
															assign node15350 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node15353 = (inp[5]) ? node15355 : 4'b0011;
															assign node15355 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node15358 = (inp[2]) ? node15388 : node15359;
												assign node15359 = (inp[14]) ? node15375 : node15360;
													assign node15360 = (inp[5]) ? node15368 : node15361;
														assign node15361 = (inp[3]) ? node15365 : node15362;
															assign node15362 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node15365 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node15368 = (inp[0]) ? node15372 : node15369;
															assign node15369 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node15372 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node15375 = (inp[15]) ? node15381 : node15376;
														assign node15376 = (inp[3]) ? node15378 : 4'b0000;
															assign node15378 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node15381 = (inp[0]) ? node15385 : node15382;
															assign node15382 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node15385 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node15388 = (inp[15]) ? node15398 : node15389;
													assign node15389 = (inp[0]) ? node15393 : node15390;
														assign node15390 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node15393 = (inp[3]) ? node15395 : 4'b0000;
															assign node15395 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node15398 = (inp[0]) ? node15404 : node15399;
														assign node15399 = (inp[3]) ? node15401 : 4'b0000;
															assign node15401 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node15404 = (inp[5]) ? node15406 : 4'b0010;
															assign node15406 = (inp[3]) ? 4'b0000 : 4'b0010;
									assign node15409 = (inp[7]) ? node15515 : node15410;
										assign node15410 = (inp[8]) ? node15462 : node15411;
											assign node15411 = (inp[2]) ? node15441 : node15412;
												assign node15412 = (inp[14]) ? node15428 : node15413;
													assign node15413 = (inp[0]) ? node15421 : node15414;
														assign node15414 = (inp[15]) ? node15418 : node15415;
															assign node15415 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node15418 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node15421 = (inp[15]) ? node15425 : node15422;
															assign node15422 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node15425 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node15428 = (inp[0]) ? node15434 : node15429;
														assign node15429 = (inp[15]) ? 4'b0000 : node15430;
															assign node15430 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node15434 = (inp[15]) ? node15438 : node15435;
															assign node15435 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node15438 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node15441 = (inp[5]) ? node15449 : node15442;
													assign node15442 = (inp[15]) ? node15446 : node15443;
														assign node15443 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node15446 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node15449 = (inp[14]) ? node15455 : node15450;
														assign node15450 = (inp[3]) ? node15452 : 4'b0010;
															assign node15452 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node15455 = (inp[3]) ? node15459 : node15456;
															assign node15456 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node15459 = (inp[15]) ? 4'b0000 : 4'b0000;
											assign node15462 = (inp[2]) ? node15492 : node15463;
												assign node15463 = (inp[14]) ? node15479 : node15464;
													assign node15464 = (inp[0]) ? node15472 : node15465;
														assign node15465 = (inp[15]) ? node15469 : node15466;
															assign node15466 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node15469 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node15472 = (inp[15]) ? node15476 : node15473;
															assign node15473 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node15476 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node15479 = (inp[3]) ? node15485 : node15480;
														assign node15480 = (inp[15]) ? 4'b1011 : node15481;
															assign node15481 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node15485 = (inp[15]) ? node15489 : node15486;
															assign node15486 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node15489 = (inp[0]) ? 4'b1001 : 4'b1001;
												assign node15492 = (inp[3]) ? node15500 : node15493;
													assign node15493 = (inp[15]) ? node15497 : node15494;
														assign node15494 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node15497 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node15500 = (inp[15]) ? node15508 : node15501;
														assign node15501 = (inp[14]) ? node15505 : node15502;
															assign node15502 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node15505 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node15508 = (inp[0]) ? node15512 : node15509;
															assign node15509 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node15512 = (inp[5]) ? 4'b1001 : 4'b1011;
										assign node15515 = (inp[8]) ? node15577 : node15516;
											assign node15516 = (inp[2]) ? node15546 : node15517;
												assign node15517 = (inp[14]) ? node15533 : node15518;
													assign node15518 = (inp[5]) ? node15526 : node15519;
														assign node15519 = (inp[0]) ? node15523 : node15520;
															assign node15520 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node15523 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node15526 = (inp[15]) ? node15530 : node15527;
															assign node15527 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node15530 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node15533 = (inp[15]) ? node15539 : node15534;
														assign node15534 = (inp[0]) ? 4'b1001 : node15535;
															assign node15535 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node15539 = (inp[0]) ? node15543 : node15540;
															assign node15540 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node15543 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node15546 = (inp[14]) ? node15562 : node15547;
													assign node15547 = (inp[15]) ? node15555 : node15548;
														assign node15548 = (inp[0]) ? node15552 : node15549;
															assign node15549 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node15552 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node15555 = (inp[0]) ? node15559 : node15556;
															assign node15556 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node15559 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node15562 = (inp[15]) ? node15570 : node15563;
														assign node15563 = (inp[0]) ? node15567 : node15564;
															assign node15564 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node15567 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node15570 = (inp[0]) ? node15574 : node15571;
															assign node15571 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node15574 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node15577 = (inp[14]) ? node15607 : node15578;
												assign node15578 = (inp[2]) ? node15594 : node15579;
													assign node15579 = (inp[0]) ? node15587 : node15580;
														assign node15580 = (inp[15]) ? node15584 : node15581;
															assign node15581 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node15584 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node15587 = (inp[15]) ? node15591 : node15588;
															assign node15588 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node15591 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node15594 = (inp[5]) ? node15602 : node15595;
														assign node15595 = (inp[15]) ? node15599 : node15596;
															assign node15596 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node15599 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node15602 = (inp[3]) ? 4'b1000 : node15603;
															assign node15603 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node15607 = (inp[15]) ? node15619 : node15608;
													assign node15608 = (inp[0]) ? node15614 : node15609;
														assign node15609 = (inp[5]) ? node15611 : 4'b1010;
															assign node15611 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node15614 = (inp[3]) ? node15616 : 4'b1000;
															assign node15616 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node15619 = (inp[0]) ? node15625 : node15620;
														assign node15620 = (inp[5]) ? node15622 : 4'b1000;
															assign node15622 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node15625 = (inp[5]) ? node15627 : 4'b1010;
															assign node15627 = (inp[3]) ? 4'b1000 : 4'b1010;
								assign node15630 = (inp[13]) ? node15854 : node15631;
									assign node15631 = (inp[7]) ? node15733 : node15632;
										assign node15632 = (inp[8]) ? node15682 : node15633;
											assign node15633 = (inp[14]) ? node15659 : node15634;
												assign node15634 = (inp[2]) ? node15648 : node15635;
													assign node15635 = (inp[0]) ? node15641 : node15636;
														assign node15636 = (inp[15]) ? node15638 : 4'b0011;
															assign node15638 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node15641 = (inp[15]) ? node15645 : node15642;
															assign node15642 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node15645 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node15648 = (inp[0]) ? node15654 : node15649;
														assign node15649 = (inp[15]) ? 4'b0000 : node15650;
															assign node15650 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node15654 = (inp[15]) ? 4'b0010 : node15655;
															assign node15655 = (inp[5]) ? 4'b0000 : 4'b0000;
												assign node15659 = (inp[15]) ? node15671 : node15660;
													assign node15660 = (inp[0]) ? node15666 : node15661;
														assign node15661 = (inp[5]) ? node15663 : 4'b0010;
															assign node15663 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node15666 = (inp[5]) ? node15668 : 4'b0000;
															assign node15668 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node15671 = (inp[0]) ? node15677 : node15672;
														assign node15672 = (inp[3]) ? node15674 : 4'b0000;
															assign node15674 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node15677 = (inp[3]) ? node15679 : 4'b0010;
															assign node15679 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node15682 = (inp[2]) ? node15710 : node15683;
												assign node15683 = (inp[14]) ? node15697 : node15684;
													assign node15684 = (inp[0]) ? node15692 : node15685;
														assign node15685 = (inp[15]) ? node15689 : node15686;
															assign node15686 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node15689 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node15692 = (inp[15]) ? 4'b0010 : node15693;
															assign node15693 = (inp[5]) ? 4'b0000 : 4'b0000;
													assign node15697 = (inp[0]) ? node15703 : node15698;
														assign node15698 = (inp[15]) ? 4'b1001 : node15699;
															assign node15699 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node15703 = (inp[15]) ? node15707 : node15704;
															assign node15704 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node15707 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node15710 = (inp[15]) ? node15722 : node15711;
													assign node15711 = (inp[0]) ? node15717 : node15712;
														assign node15712 = (inp[5]) ? node15714 : 4'b1011;
															assign node15714 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node15717 = (inp[3]) ? node15719 : 4'b1001;
															assign node15719 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node15722 = (inp[0]) ? node15728 : node15723;
														assign node15723 = (inp[5]) ? node15725 : 4'b1001;
															assign node15725 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node15728 = (inp[3]) ? node15730 : 4'b1011;
															assign node15730 = (inp[5]) ? 4'b1001 : 4'b1011;
										assign node15733 = (inp[8]) ? node15795 : node15734;
											assign node15734 = (inp[14]) ? node15764 : node15735;
												assign node15735 = (inp[2]) ? node15751 : node15736;
													assign node15736 = (inp[5]) ? node15744 : node15737;
														assign node15737 = (inp[15]) ? node15741 : node15738;
															assign node15738 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node15741 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node15744 = (inp[15]) ? node15748 : node15745;
															assign node15745 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node15748 = (inp[3]) ? 4'b0000 : 4'b0000;
													assign node15751 = (inp[0]) ? node15757 : node15752;
														assign node15752 = (inp[15]) ? node15754 : 4'b1011;
															assign node15754 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node15757 = (inp[15]) ? node15761 : node15758;
															assign node15758 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node15761 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node15764 = (inp[2]) ? node15780 : node15765;
													assign node15765 = (inp[15]) ? node15773 : node15766;
														assign node15766 = (inp[0]) ? node15770 : node15767;
															assign node15767 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node15770 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node15773 = (inp[0]) ? node15777 : node15774;
															assign node15774 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node15777 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node15780 = (inp[3]) ? node15788 : node15781;
														assign node15781 = (inp[0]) ? node15785 : node15782;
															assign node15782 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node15785 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node15788 = (inp[0]) ? node15792 : node15789;
															assign node15789 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node15792 = (inp[5]) ? 4'b1001 : 4'b1001;
											assign node15795 = (inp[14]) ? node15827 : node15796;
												assign node15796 = (inp[2]) ? node15812 : node15797;
													assign node15797 = (inp[3]) ? node15805 : node15798;
														assign node15798 = (inp[0]) ? node15802 : node15799;
															assign node15799 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node15802 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node15805 = (inp[5]) ? node15809 : node15806;
															assign node15806 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node15809 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node15812 = (inp[15]) ? node15820 : node15813;
														assign node15813 = (inp[0]) ? node15817 : node15814;
															assign node15814 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node15817 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node15820 = (inp[0]) ? node15824 : node15821;
															assign node15821 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node15824 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node15827 = (inp[3]) ? node15841 : node15828;
													assign node15828 = (inp[2]) ? node15836 : node15829;
														assign node15829 = (inp[5]) ? node15833 : node15830;
															assign node15830 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node15833 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node15836 = (inp[0]) ? 4'b1010 : node15837;
															assign node15837 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node15841 = (inp[0]) ? node15849 : node15842;
														assign node15842 = (inp[5]) ? node15846 : node15843;
															assign node15843 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node15846 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node15849 = (inp[2]) ? 4'b1000 : node15850;
															assign node15850 = (inp[5]) ? 4'b1000 : 4'b1000;
									assign node15854 = (inp[5]) ? node15950 : node15855;
										assign node15855 = (inp[15]) ? node15903 : node15856;
											assign node15856 = (inp[0]) ? node15880 : node15857;
												assign node15857 = (inp[7]) ? node15869 : node15858;
													assign node15858 = (inp[8]) ? node15864 : node15859;
														assign node15859 = (inp[14]) ? 4'b1010 : node15860;
															assign node15860 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node15864 = (inp[2]) ? 4'b1011 : node15865;
															assign node15865 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node15869 = (inp[8]) ? node15875 : node15870;
														assign node15870 = (inp[2]) ? 4'b1011 : node15871;
															assign node15871 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node15875 = (inp[14]) ? 4'b1010 : node15876;
															assign node15876 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node15880 = (inp[8]) ? node15892 : node15881;
													assign node15881 = (inp[7]) ? node15887 : node15882;
														assign node15882 = (inp[14]) ? 4'b1000 : node15883;
															assign node15883 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node15887 = (inp[2]) ? 4'b1001 : node15888;
															assign node15888 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node15892 = (inp[7]) ? node15898 : node15893;
														assign node15893 = (inp[2]) ? 4'b1001 : node15894;
															assign node15894 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node15898 = (inp[2]) ? 4'b1000 : node15899;
															assign node15899 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node15903 = (inp[0]) ? node15927 : node15904;
												assign node15904 = (inp[7]) ? node15916 : node15905;
													assign node15905 = (inp[8]) ? node15911 : node15906;
														assign node15906 = (inp[2]) ? 4'b1000 : node15907;
															assign node15907 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node15911 = (inp[2]) ? 4'b1001 : node15912;
															assign node15912 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node15916 = (inp[8]) ? node15922 : node15917;
														assign node15917 = (inp[14]) ? 4'b1001 : node15918;
															assign node15918 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node15922 = (inp[14]) ? 4'b1000 : node15923;
															assign node15923 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node15927 = (inp[7]) ? node15939 : node15928;
													assign node15928 = (inp[8]) ? node15934 : node15929;
														assign node15929 = (inp[14]) ? 4'b1010 : node15930;
															assign node15930 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node15934 = (inp[14]) ? 4'b1011 : node15935;
															assign node15935 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node15939 = (inp[8]) ? node15945 : node15940;
														assign node15940 = (inp[2]) ? 4'b1011 : node15941;
															assign node15941 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node15945 = (inp[2]) ? 4'b1010 : node15946;
															assign node15946 = (inp[14]) ? 4'b1010 : 4'b1011;
										assign node15950 = (inp[0]) ? node16006 : node15951;
											assign node15951 = (inp[15]) ? node15979 : node15952;
												assign node15952 = (inp[3]) ? node15966 : node15953;
													assign node15953 = (inp[7]) ? node15961 : node15954;
														assign node15954 = (inp[8]) ? node15958 : node15955;
															assign node15955 = (inp[2]) ? 4'b1010 : 4'b1010;
															assign node15958 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node15961 = (inp[8]) ? node15963 : 4'b1011;
															assign node15963 = (inp[14]) ? 4'b1010 : 4'b1010;
													assign node15966 = (inp[14]) ? node15972 : node15967;
														assign node15967 = (inp[8]) ? node15969 : 4'b1000;
															assign node15969 = (inp[2]) ? 4'b1000 : 4'b1000;
														assign node15972 = (inp[7]) ? node15976 : node15973;
															assign node15973 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node15976 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node15979 = (inp[3]) ? node15991 : node15980;
													assign node15980 = (inp[7]) ? node15986 : node15981;
														assign node15981 = (inp[8]) ? 4'b1001 : node15982;
															assign node15982 = (inp[2]) ? 4'b1000 : 4'b1000;
														assign node15986 = (inp[8]) ? 4'b1000 : node15987;
															assign node15987 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node15991 = (inp[7]) ? node15999 : node15992;
														assign node15992 = (inp[8]) ? node15996 : node15993;
															assign node15993 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node15996 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node15999 = (inp[8]) ? node16003 : node16000;
															assign node16000 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node16003 = (inp[14]) ? 4'b1010 : 4'b1011;
											assign node16006 = (inp[3]) ? node16038 : node16007;
												assign node16007 = (inp[15]) ? node16023 : node16008;
													assign node16008 = (inp[2]) ? node16016 : node16009;
														assign node16009 = (inp[8]) ? node16013 : node16010;
															assign node16010 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node16013 = (inp[7]) ? 4'b1000 : 4'b1000;
														assign node16016 = (inp[14]) ? node16020 : node16017;
															assign node16017 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node16020 = (inp[7]) ? 4'b1000 : 4'b1000;
													assign node16023 = (inp[7]) ? node16031 : node16024;
														assign node16024 = (inp[8]) ? node16028 : node16025;
															assign node16025 = (inp[2]) ? 4'b1010 : 4'b1010;
															assign node16028 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node16031 = (inp[8]) ? node16035 : node16032;
															assign node16032 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node16035 = (inp[14]) ? 4'b1010 : 4'b1010;
												assign node16038 = (inp[15]) ? node16052 : node16039;
													assign node16039 = (inp[7]) ? node16047 : node16040;
														assign node16040 = (inp[8]) ? node16044 : node16041;
															assign node16041 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node16044 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node16047 = (inp[8]) ? node16049 : 4'b1011;
															assign node16049 = (inp[14]) ? 4'b1010 : 4'b1010;
													assign node16052 = (inp[8]) ? node16060 : node16053;
														assign node16053 = (inp[7]) ? node16057 : node16054;
															assign node16054 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node16057 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node16060 = (inp[7]) ? node16064 : node16061;
															assign node16061 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node16064 = (inp[2]) ? 4'b1000 : 4'b1001;
						assign node16067 = (inp[11]) ? node16971 : node16068;
							assign node16068 = (inp[13]) ? node16518 : node16069;
								assign node16069 = (inp[1]) ? node16293 : node16070;
									assign node16070 = (inp[3]) ? node16172 : node16071;
										assign node16071 = (inp[14]) ? node16133 : node16072;
											assign node16072 = (inp[7]) ? node16102 : node16073;
												assign node16073 = (inp[15]) ? node16087 : node16074;
													assign node16074 = (inp[0]) ? node16082 : node16075;
														assign node16075 = (inp[8]) ? node16079 : node16076;
															assign node16076 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node16079 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node16082 = (inp[8]) ? node16084 : 4'b0001;
															assign node16084 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node16087 = (inp[0]) ? node16095 : node16088;
														assign node16088 = (inp[2]) ? node16092 : node16089;
															assign node16089 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node16092 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node16095 = (inp[2]) ? node16099 : node16096;
															assign node16096 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node16099 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node16102 = (inp[0]) ? node16118 : node16103;
													assign node16103 = (inp[15]) ? node16111 : node16104;
														assign node16104 = (inp[8]) ? node16108 : node16105;
															assign node16105 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node16108 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node16111 = (inp[5]) ? node16115 : node16112;
															assign node16112 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node16115 = (inp[2]) ? 4'b0000 : 4'b0000;
													assign node16118 = (inp[15]) ? node16126 : node16119;
														assign node16119 = (inp[5]) ? node16123 : node16120;
															assign node16120 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node16123 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node16126 = (inp[2]) ? node16130 : node16127;
															assign node16127 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node16130 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node16133 = (inp[7]) ? node16149 : node16134;
												assign node16134 = (inp[8]) ? node16142 : node16135;
													assign node16135 = (inp[15]) ? node16139 : node16136;
														assign node16136 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node16139 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node16142 = (inp[15]) ? node16146 : node16143;
														assign node16143 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node16146 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node16149 = (inp[8]) ? node16157 : node16150;
													assign node16150 = (inp[0]) ? node16154 : node16151;
														assign node16151 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node16154 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node16157 = (inp[2]) ? node16165 : node16158;
														assign node16158 = (inp[5]) ? node16162 : node16159;
															assign node16159 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node16162 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node16165 = (inp[5]) ? node16169 : node16166;
															assign node16166 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node16169 = (inp[0]) ? 4'b0000 : 4'b0000;
										assign node16172 = (inp[2]) ? node16234 : node16173;
											assign node16173 = (inp[0]) ? node16203 : node16174;
												assign node16174 = (inp[14]) ? node16188 : node16175;
													assign node16175 = (inp[5]) ? node16183 : node16176;
														assign node16176 = (inp[15]) ? node16180 : node16177;
															assign node16177 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node16180 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node16183 = (inp[15]) ? node16185 : 4'b0001;
															assign node16185 = (inp[7]) ? 4'b0010 : 4'b0010;
													assign node16188 = (inp[8]) ? node16196 : node16189;
														assign node16189 = (inp[7]) ? node16193 : node16190;
															assign node16190 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node16193 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node16196 = (inp[7]) ? node16200 : node16197;
															assign node16197 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node16200 = (inp[15]) ? 4'b0000 : 4'b0000;
												assign node16203 = (inp[7]) ? node16219 : node16204;
													assign node16204 = (inp[15]) ? node16212 : node16205;
														assign node16205 = (inp[5]) ? node16209 : node16206;
															assign node16206 = (inp[14]) ? 4'b0000 : 4'b0000;
															assign node16209 = (inp[8]) ? 4'b0010 : 4'b0010;
														assign node16212 = (inp[5]) ? node16216 : node16213;
															assign node16213 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node16216 = (inp[8]) ? 4'b0000 : 4'b0000;
													assign node16219 = (inp[15]) ? node16227 : node16220;
														assign node16220 = (inp[5]) ? node16224 : node16221;
															assign node16221 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node16224 = (inp[8]) ? 4'b0010 : 4'b0010;
														assign node16227 = (inp[5]) ? node16231 : node16228;
															assign node16228 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node16231 = (inp[8]) ? 4'b0000 : 4'b0000;
											assign node16234 = (inp[5]) ? node16264 : node16235;
												assign node16235 = (inp[0]) ? node16249 : node16236;
													assign node16236 = (inp[15]) ? node16242 : node16237;
														assign node16237 = (inp[14]) ? 4'b0010 : node16238;
															assign node16238 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node16242 = (inp[8]) ? node16246 : node16243;
															assign node16243 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node16246 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node16249 = (inp[15]) ? node16257 : node16250;
														assign node16250 = (inp[7]) ? node16254 : node16251;
															assign node16251 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node16254 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node16257 = (inp[14]) ? node16261 : node16258;
															assign node16258 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node16261 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node16264 = (inp[7]) ? node16278 : node16265;
													assign node16265 = (inp[8]) ? node16273 : node16266;
														assign node16266 = (inp[14]) ? node16270 : node16267;
															assign node16267 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node16270 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node16273 = (inp[14]) ? node16275 : 4'b0011;
															assign node16275 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node16278 = (inp[8]) ? node16286 : node16279;
														assign node16279 = (inp[0]) ? node16283 : node16280;
															assign node16280 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node16283 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node16286 = (inp[14]) ? node16290 : node16287;
															assign node16287 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node16290 = (inp[15]) ? 4'b0000 : 4'b0000;
									assign node16293 = (inp[7]) ? node16407 : node16294;
										assign node16294 = (inp[8]) ? node16356 : node16295;
											assign node16295 = (inp[2]) ? node16325 : node16296;
												assign node16296 = (inp[14]) ? node16310 : node16297;
													assign node16297 = (inp[3]) ? node16305 : node16298;
														assign node16298 = (inp[5]) ? node16302 : node16299;
															assign node16299 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node16302 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node16305 = (inp[15]) ? 4'b0001 : node16306;
															assign node16306 = (inp[5]) ? 4'b0001 : 4'b0001;
													assign node16310 = (inp[15]) ? node16318 : node16311;
														assign node16311 = (inp[0]) ? node16315 : node16312;
															assign node16312 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node16315 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node16318 = (inp[0]) ? node16322 : node16319;
															assign node16319 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node16322 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node16325 = (inp[5]) ? node16341 : node16326;
													assign node16326 = (inp[14]) ? node16334 : node16327;
														assign node16327 = (inp[0]) ? node16331 : node16328;
															assign node16328 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node16331 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node16334 = (inp[0]) ? node16338 : node16335;
															assign node16335 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node16338 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node16341 = (inp[0]) ? node16349 : node16342;
														assign node16342 = (inp[15]) ? node16346 : node16343;
															assign node16343 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node16346 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node16349 = (inp[3]) ? node16353 : node16350;
															assign node16350 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node16353 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node16356 = (inp[14]) ? node16384 : node16357;
												assign node16357 = (inp[2]) ? node16373 : node16358;
													assign node16358 = (inp[5]) ? node16366 : node16359;
														assign node16359 = (inp[3]) ? node16363 : node16360;
															assign node16360 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node16363 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node16366 = (inp[0]) ? node16370 : node16367;
															assign node16367 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node16370 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node16373 = (inp[5]) ? node16379 : node16374;
														assign node16374 = (inp[3]) ? 4'b1011 : node16375;
															assign node16375 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node16379 = (inp[3]) ? 4'b1001 : node16380;
															assign node16380 = (inp[0]) ? 4'b1001 : 4'b1001;
												assign node16384 = (inp[3]) ? node16392 : node16385;
													assign node16385 = (inp[0]) ? node16389 : node16386;
														assign node16386 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node16389 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node16392 = (inp[5]) ? node16400 : node16393;
														assign node16393 = (inp[15]) ? node16397 : node16394;
															assign node16394 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node16397 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node16400 = (inp[0]) ? node16404 : node16401;
															assign node16401 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node16404 = (inp[15]) ? 4'b1001 : 4'b1011;
										assign node16407 = (inp[8]) ? node16457 : node16408;
											assign node16408 = (inp[14]) ? node16434 : node16409;
												assign node16409 = (inp[2]) ? node16425 : node16410;
													assign node16410 = (inp[0]) ? node16418 : node16411;
														assign node16411 = (inp[15]) ? node16415 : node16412;
															assign node16412 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node16415 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node16418 = (inp[15]) ? node16422 : node16419;
															assign node16419 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node16422 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node16425 = (inp[5]) ? 4'b1001 : node16426;
														assign node16426 = (inp[15]) ? node16430 : node16427;
															assign node16427 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node16430 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node16434 = (inp[15]) ? node16446 : node16435;
													assign node16435 = (inp[0]) ? node16441 : node16436;
														assign node16436 = (inp[3]) ? node16438 : 4'b1011;
															assign node16438 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node16441 = (inp[5]) ? node16443 : 4'b1001;
															assign node16443 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node16446 = (inp[0]) ? node16452 : node16447;
														assign node16447 = (inp[3]) ? node16449 : 4'b1001;
															assign node16449 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node16452 = (inp[5]) ? node16454 : 4'b1011;
															assign node16454 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node16457 = (inp[14]) ? node16487 : node16458;
												assign node16458 = (inp[2]) ? node16472 : node16459;
													assign node16459 = (inp[3]) ? node16467 : node16460;
														assign node16460 = (inp[5]) ? node16464 : node16461;
															assign node16461 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node16464 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node16467 = (inp[0]) ? node16469 : 4'b1001;
															assign node16469 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node16472 = (inp[3]) ? node16480 : node16473;
														assign node16473 = (inp[5]) ? node16477 : node16474;
															assign node16474 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node16477 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node16480 = (inp[0]) ? node16484 : node16481;
															assign node16481 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node16484 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node16487 = (inp[5]) ? node16503 : node16488;
													assign node16488 = (inp[2]) ? node16496 : node16489;
														assign node16489 = (inp[3]) ? node16493 : node16490;
															assign node16490 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node16493 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node16496 = (inp[15]) ? node16500 : node16497;
															assign node16497 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node16500 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node16503 = (inp[15]) ? node16511 : node16504;
														assign node16504 = (inp[3]) ? node16508 : node16505;
															assign node16505 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node16508 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node16511 = (inp[2]) ? node16515 : node16512;
															assign node16512 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node16515 = (inp[3]) ? 4'b1000 : 4'b1000;
								assign node16518 = (inp[1]) ? node16744 : node16519;
									assign node16519 = (inp[7]) ? node16637 : node16520;
										assign node16520 = (inp[8]) ? node16578 : node16521;
											assign node16521 = (inp[14]) ? node16549 : node16522;
												assign node16522 = (inp[2]) ? node16536 : node16523;
													assign node16523 = (inp[15]) ? node16529 : node16524;
														assign node16524 = (inp[0]) ? 4'b0001 : node16525;
															assign node16525 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node16529 = (inp[0]) ? node16533 : node16530;
															assign node16530 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node16533 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node16536 = (inp[0]) ? node16544 : node16537;
														assign node16537 = (inp[15]) ? node16541 : node16538;
															assign node16538 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node16541 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node16544 = (inp[15]) ? 4'b0010 : node16545;
															assign node16545 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node16549 = (inp[3]) ? node16565 : node16550;
													assign node16550 = (inp[2]) ? node16558 : node16551;
														assign node16551 = (inp[0]) ? node16555 : node16552;
															assign node16552 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node16555 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node16558 = (inp[15]) ? node16562 : node16559;
															assign node16559 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node16562 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node16565 = (inp[2]) ? node16573 : node16566;
														assign node16566 = (inp[5]) ? node16570 : node16567;
															assign node16567 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node16570 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node16573 = (inp[0]) ? node16575 : 4'b0000;
															assign node16575 = (inp[5]) ? 4'b0000 : 4'b0000;
											assign node16578 = (inp[14]) ? node16608 : node16579;
												assign node16579 = (inp[2]) ? node16595 : node16580;
													assign node16580 = (inp[5]) ? node16588 : node16581;
														assign node16581 = (inp[0]) ? node16585 : node16582;
															assign node16582 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node16585 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node16588 = (inp[15]) ? node16592 : node16589;
															assign node16589 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node16592 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node16595 = (inp[3]) ? node16601 : node16596;
														assign node16596 = (inp[5]) ? 4'b1011 : node16597;
															assign node16597 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node16601 = (inp[5]) ? node16605 : node16602;
															assign node16602 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node16605 = (inp[15]) ? 4'b1001 : 4'b1001;
												assign node16608 = (inp[3]) ? node16622 : node16609;
													assign node16609 = (inp[2]) ? node16617 : node16610;
														assign node16610 = (inp[5]) ? node16614 : node16611;
															assign node16611 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node16614 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node16617 = (inp[5]) ? node16619 : 4'b1001;
															assign node16619 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node16622 = (inp[2]) ? node16630 : node16623;
														assign node16623 = (inp[5]) ? node16627 : node16624;
															assign node16624 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node16627 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node16630 = (inp[15]) ? node16634 : node16631;
															assign node16631 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node16634 = (inp[0]) ? 4'b1001 : 4'b1001;
										assign node16637 = (inp[8]) ? node16691 : node16638;
											assign node16638 = (inp[14]) ? node16668 : node16639;
												assign node16639 = (inp[2]) ? node16653 : node16640;
													assign node16640 = (inp[15]) ? node16646 : node16641;
														assign node16641 = (inp[0]) ? node16643 : 4'b0010;
															assign node16643 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node16646 = (inp[0]) ? node16650 : node16647;
															assign node16647 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node16650 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node16653 = (inp[15]) ? node16661 : node16654;
														assign node16654 = (inp[0]) ? node16658 : node16655;
															assign node16655 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node16658 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node16661 = (inp[0]) ? node16665 : node16662;
															assign node16662 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node16665 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node16668 = (inp[0]) ? node16680 : node16669;
													assign node16669 = (inp[15]) ? node16675 : node16670;
														assign node16670 = (inp[5]) ? node16672 : 4'b1011;
															assign node16672 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node16675 = (inp[5]) ? node16677 : 4'b1001;
															assign node16677 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node16680 = (inp[15]) ? node16686 : node16681;
														assign node16681 = (inp[5]) ? node16683 : 4'b1001;
															assign node16683 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node16686 = (inp[3]) ? node16688 : 4'b1011;
															assign node16688 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node16691 = (inp[14]) ? node16721 : node16692;
												assign node16692 = (inp[2]) ? node16708 : node16693;
													assign node16693 = (inp[5]) ? node16701 : node16694;
														assign node16694 = (inp[3]) ? node16698 : node16695;
															assign node16695 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node16698 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node16701 = (inp[3]) ? node16705 : node16702;
															assign node16702 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node16705 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node16708 = (inp[0]) ? node16716 : node16709;
														assign node16709 = (inp[15]) ? node16713 : node16710;
															assign node16710 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node16713 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node16716 = (inp[3]) ? node16718 : 4'b1010;
															assign node16718 = (inp[5]) ? 4'b1000 : 4'b1000;
												assign node16721 = (inp[15]) ? node16733 : node16722;
													assign node16722 = (inp[0]) ? node16728 : node16723;
														assign node16723 = (inp[3]) ? node16725 : 4'b1010;
															assign node16725 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node16728 = (inp[5]) ? node16730 : 4'b1000;
															assign node16730 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node16733 = (inp[0]) ? node16739 : node16734;
														assign node16734 = (inp[3]) ? node16736 : 4'b1000;
															assign node16736 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node16739 = (inp[3]) ? node16741 : 4'b1010;
															assign node16741 = (inp[5]) ? 4'b1000 : 4'b1010;
									assign node16744 = (inp[0]) ? node16862 : node16745;
										assign node16745 = (inp[15]) ? node16805 : node16746;
											assign node16746 = (inp[3]) ? node16778 : node16747;
												assign node16747 = (inp[5]) ? node16763 : node16748;
													assign node16748 = (inp[14]) ? node16756 : node16749;
														assign node16749 = (inp[7]) ? node16753 : node16750;
															assign node16750 = (inp[8]) ? 4'b1010 : 4'b1010;
															assign node16753 = (inp[2]) ? 4'b1010 : 4'b1010;
														assign node16756 = (inp[7]) ? node16760 : node16757;
															assign node16757 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node16760 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node16763 = (inp[2]) ? node16771 : node16764;
														assign node16764 = (inp[14]) ? node16768 : node16765;
															assign node16765 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node16768 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node16771 = (inp[8]) ? node16775 : node16772;
															assign node16772 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node16775 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node16778 = (inp[5]) ? node16792 : node16779;
													assign node16779 = (inp[7]) ? node16787 : node16780;
														assign node16780 = (inp[8]) ? node16784 : node16781;
															assign node16781 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node16784 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node16787 = (inp[14]) ? 4'b1010 : node16788;
															assign node16788 = (inp[2]) ? 4'b1010 : 4'b1010;
													assign node16792 = (inp[7]) ? node16800 : node16793;
														assign node16793 = (inp[8]) ? node16797 : node16794;
															assign node16794 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node16797 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node16800 = (inp[14]) ? 4'b1001 : node16801;
															assign node16801 = (inp[2]) ? 4'b1000 : 4'b1000;
											assign node16805 = (inp[3]) ? node16835 : node16806;
												assign node16806 = (inp[2]) ? node16820 : node16807;
													assign node16807 = (inp[14]) ? node16815 : node16808;
														assign node16808 = (inp[5]) ? node16812 : node16809;
															assign node16809 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node16812 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node16815 = (inp[8]) ? node16817 : 4'b1001;
															assign node16817 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node16820 = (inp[5]) ? node16828 : node16821;
														assign node16821 = (inp[7]) ? node16825 : node16822;
															assign node16822 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node16825 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node16828 = (inp[7]) ? node16832 : node16829;
															assign node16829 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node16832 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node16835 = (inp[5]) ? node16849 : node16836;
													assign node16836 = (inp[8]) ? node16842 : node16837;
														assign node16837 = (inp[7]) ? 4'b1001 : node16838;
															assign node16838 = (inp[2]) ? 4'b1000 : 4'b1000;
														assign node16842 = (inp[7]) ? node16846 : node16843;
															assign node16843 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node16846 = (inp[2]) ? 4'b1000 : 4'b1000;
													assign node16849 = (inp[2]) ? node16855 : node16850;
														assign node16850 = (inp[7]) ? node16852 : 4'b1011;
															assign node16852 = (inp[14]) ? 4'b1010 : 4'b1010;
														assign node16855 = (inp[14]) ? node16859 : node16856;
															assign node16856 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node16859 = (inp[8]) ? 4'b1010 : 4'b1010;
										assign node16862 = (inp[15]) ? node16916 : node16863;
											assign node16863 = (inp[3]) ? node16887 : node16864;
												assign node16864 = (inp[7]) ? node16876 : node16865;
													assign node16865 = (inp[8]) ? node16871 : node16866;
														assign node16866 = (inp[14]) ? 4'b1000 : node16867;
															assign node16867 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node16871 = (inp[2]) ? 4'b1001 : node16872;
															assign node16872 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node16876 = (inp[8]) ? node16882 : node16877;
														assign node16877 = (inp[14]) ? 4'b1001 : node16878;
															assign node16878 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node16882 = (inp[2]) ? 4'b1000 : node16883;
															assign node16883 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node16887 = (inp[5]) ? node16903 : node16888;
													assign node16888 = (inp[14]) ? node16896 : node16889;
														assign node16889 = (inp[2]) ? node16893 : node16890;
															assign node16890 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node16893 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node16896 = (inp[2]) ? node16900 : node16897;
															assign node16897 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node16900 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node16903 = (inp[2]) ? node16909 : node16904;
														assign node16904 = (inp[7]) ? 4'b1010 : node16905;
															assign node16905 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node16909 = (inp[14]) ? node16913 : node16910;
															assign node16910 = (inp[8]) ? 4'b1010 : 4'b1010;
															assign node16913 = (inp[7]) ? 4'b1010 : 4'b1010;
											assign node16916 = (inp[5]) ? node16944 : node16917;
												assign node16917 = (inp[3]) ? node16931 : node16918;
													assign node16918 = (inp[2]) ? node16926 : node16919;
														assign node16919 = (inp[7]) ? node16923 : node16920;
															assign node16920 = (inp[8]) ? 4'b1010 : 4'b1010;
															assign node16923 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node16926 = (inp[7]) ? node16928 : 4'b1011;
															assign node16928 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node16931 = (inp[7]) ? node16937 : node16932;
														assign node16932 = (inp[8]) ? 4'b1011 : node16933;
															assign node16933 = (inp[14]) ? 4'b1010 : 4'b1010;
														assign node16937 = (inp[8]) ? node16941 : node16938;
															assign node16938 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node16941 = (inp[14]) ? 4'b1010 : 4'b1010;
												assign node16944 = (inp[3]) ? node16958 : node16945;
													assign node16945 = (inp[8]) ? node16951 : node16946;
														assign node16946 = (inp[7]) ? 4'b1011 : node16947;
															assign node16947 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node16951 = (inp[7]) ? node16955 : node16952;
															assign node16952 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node16955 = (inp[14]) ? 4'b1010 : 4'b1010;
													assign node16958 = (inp[8]) ? node16966 : node16959;
														assign node16959 = (inp[7]) ? node16963 : node16960;
															assign node16960 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node16963 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node16966 = (inp[7]) ? 4'b1000 : node16967;
															assign node16967 = (inp[2]) ? 4'b1001 : 4'b1000;
							assign node16971 = (inp[13]) ? node17427 : node16972;
								assign node16972 = (inp[1]) ? node17200 : node16973;
									assign node16973 = (inp[3]) ? node17081 : node16974;
										assign node16974 = (inp[2]) ? node17036 : node16975;
											assign node16975 = (inp[8]) ? node17005 : node16976;
												assign node16976 = (inp[5]) ? node16992 : node16977;
													assign node16977 = (inp[7]) ? node16985 : node16978;
														assign node16978 = (inp[14]) ? node16982 : node16979;
															assign node16979 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node16982 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node16985 = (inp[14]) ? node16989 : node16986;
															assign node16986 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node16989 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node16992 = (inp[7]) ? node16998 : node16993;
														assign node16993 = (inp[14]) ? node16995 : 4'b1001;
															assign node16995 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node16998 = (inp[14]) ? node17002 : node16999;
															assign node16999 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node17002 = (inp[15]) ? 4'b1001 : 4'b1001;
												assign node17005 = (inp[7]) ? node17021 : node17006;
													assign node17006 = (inp[14]) ? node17014 : node17007;
														assign node17007 = (inp[0]) ? node17011 : node17008;
															assign node17008 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node17011 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node17014 = (inp[15]) ? node17018 : node17015;
															assign node17015 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node17018 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node17021 = (inp[14]) ? node17029 : node17022;
														assign node17022 = (inp[5]) ? node17026 : node17023;
															assign node17023 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node17026 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node17029 = (inp[15]) ? node17033 : node17030;
															assign node17030 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node17033 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node17036 = (inp[8]) ? node17052 : node17037;
												assign node17037 = (inp[7]) ? node17045 : node17038;
													assign node17038 = (inp[15]) ? node17042 : node17039;
														assign node17039 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node17042 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node17045 = (inp[0]) ? node17049 : node17046;
														assign node17046 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node17049 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node17052 = (inp[7]) ? node17066 : node17053;
													assign node17053 = (inp[14]) ? node17059 : node17054;
														assign node17054 = (inp[0]) ? node17056 : 4'b1001;
															assign node17056 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node17059 = (inp[5]) ? node17063 : node17060;
															assign node17060 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node17063 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node17066 = (inp[14]) ? node17074 : node17067;
														assign node17067 = (inp[15]) ? node17071 : node17068;
															assign node17068 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node17071 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node17074 = (inp[0]) ? node17078 : node17075;
															assign node17075 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node17078 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node17081 = (inp[2]) ? node17143 : node17082;
											assign node17082 = (inp[5]) ? node17114 : node17083;
												assign node17083 = (inp[8]) ? node17099 : node17084;
													assign node17084 = (inp[15]) ? node17092 : node17085;
														assign node17085 = (inp[0]) ? node17089 : node17086;
															assign node17086 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node17089 = (inp[14]) ? 4'b1000 : 4'b1000;
														assign node17092 = (inp[0]) ? node17096 : node17093;
															assign node17093 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node17096 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node17099 = (inp[15]) ? node17107 : node17100;
														assign node17100 = (inp[0]) ? node17104 : node17101;
															assign node17101 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node17104 = (inp[7]) ? 4'b1000 : 4'b1000;
														assign node17107 = (inp[0]) ? node17111 : node17108;
															assign node17108 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node17111 = (inp[7]) ? 4'b1010 : 4'b1010;
												assign node17114 = (inp[15]) ? node17128 : node17115;
													assign node17115 = (inp[0]) ? node17121 : node17116;
														assign node17116 = (inp[7]) ? 4'b1000 : node17117;
															assign node17117 = (inp[14]) ? 4'b1000 : 4'b1000;
														assign node17121 = (inp[14]) ? node17125 : node17122;
															assign node17122 = (inp[8]) ? 4'b1010 : 4'b1010;
															assign node17125 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node17128 = (inp[0]) ? node17136 : node17129;
														assign node17129 = (inp[8]) ? node17133 : node17130;
															assign node17130 = (inp[14]) ? 4'b1010 : 4'b1011;
															assign node17133 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node17136 = (inp[8]) ? node17140 : node17137;
															assign node17137 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node17140 = (inp[7]) ? 4'b1001 : 4'b1000;
											assign node17143 = (inp[14]) ? node17173 : node17144;
												assign node17144 = (inp[5]) ? node17160 : node17145;
													assign node17145 = (inp[15]) ? node17153 : node17146;
														assign node17146 = (inp[0]) ? node17150 : node17147;
															assign node17147 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node17150 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node17153 = (inp[0]) ? node17157 : node17154;
															assign node17154 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node17157 = (inp[8]) ? 4'b1010 : 4'b1010;
													assign node17160 = (inp[0]) ? node17168 : node17161;
														assign node17161 = (inp[15]) ? node17165 : node17162;
															assign node17162 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node17165 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node17168 = (inp[15]) ? node17170 : 4'b1011;
															assign node17170 = (inp[8]) ? 4'b1000 : 4'b1000;
												assign node17173 = (inp[7]) ? node17187 : node17174;
													assign node17174 = (inp[8]) ? node17180 : node17175;
														assign node17175 = (inp[5]) ? node17177 : 4'b1010;
															assign node17177 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node17180 = (inp[15]) ? node17184 : node17181;
															assign node17181 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node17184 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node17187 = (inp[8]) ? node17193 : node17188;
														assign node17188 = (inp[5]) ? 4'b1011 : node17189;
															assign node17189 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node17193 = (inp[15]) ? node17197 : node17194;
															assign node17194 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node17197 = (inp[5]) ? 4'b1000 : 4'b1000;
									assign node17200 = (inp[8]) ? node17310 : node17201;
										assign node17201 = (inp[7]) ? node17257 : node17202;
											assign node17202 = (inp[2]) ? node17234 : node17203;
												assign node17203 = (inp[14]) ? node17219 : node17204;
													assign node17204 = (inp[0]) ? node17212 : node17205;
														assign node17205 = (inp[15]) ? node17209 : node17206;
															assign node17206 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node17209 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node17212 = (inp[15]) ? node17216 : node17213;
															assign node17213 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node17216 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node17219 = (inp[5]) ? node17227 : node17220;
														assign node17220 = (inp[3]) ? node17224 : node17221;
															assign node17221 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node17224 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node17227 = (inp[0]) ? node17231 : node17228;
															assign node17228 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node17231 = (inp[3]) ? 4'b1000 : 4'b1000;
												assign node17234 = (inp[3]) ? node17242 : node17235;
													assign node17235 = (inp[15]) ? node17239 : node17236;
														assign node17236 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node17239 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node17242 = (inp[5]) ? node17250 : node17243;
														assign node17243 = (inp[14]) ? node17247 : node17244;
															assign node17244 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node17247 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node17250 = (inp[15]) ? node17254 : node17251;
															assign node17251 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node17254 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node17257 = (inp[14]) ? node17287 : node17258;
												assign node17258 = (inp[2]) ? node17274 : node17259;
													assign node17259 = (inp[3]) ? node17267 : node17260;
														assign node17260 = (inp[5]) ? node17264 : node17261;
															assign node17261 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node17264 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node17267 = (inp[15]) ? node17271 : node17268;
															assign node17268 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node17271 = (inp[5]) ? 4'b1000 : 4'b1000;
													assign node17274 = (inp[5]) ? node17280 : node17275;
														assign node17275 = (inp[3]) ? node17277 : 4'b0001;
															assign node17277 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node17280 = (inp[0]) ? node17284 : node17281;
															assign node17281 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node17284 = (inp[3]) ? 4'b0001 : 4'b0001;
												assign node17287 = (inp[0]) ? node17299 : node17288;
													assign node17288 = (inp[15]) ? node17294 : node17289;
														assign node17289 = (inp[3]) ? node17291 : 4'b0011;
															assign node17291 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node17294 = (inp[5]) ? node17296 : 4'b0001;
															assign node17296 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node17299 = (inp[15]) ? node17305 : node17300;
														assign node17300 = (inp[5]) ? node17302 : 4'b0001;
															assign node17302 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node17305 = (inp[5]) ? node17307 : 4'b0011;
															assign node17307 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node17310 = (inp[7]) ? node17366 : node17311;
											assign node17311 = (inp[2]) ? node17343 : node17312;
												assign node17312 = (inp[14]) ? node17328 : node17313;
													assign node17313 = (inp[5]) ? node17321 : node17314;
														assign node17314 = (inp[3]) ? node17318 : node17315;
															assign node17315 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node17318 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node17321 = (inp[3]) ? node17325 : node17322;
															assign node17322 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node17325 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node17328 = (inp[5]) ? node17336 : node17329;
														assign node17329 = (inp[0]) ? node17333 : node17330;
															assign node17330 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node17333 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node17336 = (inp[3]) ? node17340 : node17337;
															assign node17337 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node17340 = (inp[15]) ? 4'b0001 : 4'b0001;
												assign node17343 = (inp[0]) ? node17355 : node17344;
													assign node17344 = (inp[15]) ? node17350 : node17345;
														assign node17345 = (inp[5]) ? node17347 : 4'b0011;
															assign node17347 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node17350 = (inp[3]) ? node17352 : 4'b0001;
															assign node17352 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node17355 = (inp[15]) ? node17361 : node17356;
														assign node17356 = (inp[3]) ? node17358 : 4'b0001;
															assign node17358 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node17361 = (inp[5]) ? node17363 : 4'b0011;
															assign node17363 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node17366 = (inp[2]) ? node17398 : node17367;
												assign node17367 = (inp[14]) ? node17383 : node17368;
													assign node17368 = (inp[0]) ? node17376 : node17369;
														assign node17369 = (inp[15]) ? node17373 : node17370;
															assign node17370 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node17373 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node17376 = (inp[15]) ? node17380 : node17377;
															assign node17377 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node17380 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node17383 = (inp[5]) ? node17391 : node17384;
														assign node17384 = (inp[15]) ? node17388 : node17385;
															assign node17385 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node17388 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node17391 = (inp[0]) ? node17395 : node17392;
															assign node17392 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node17395 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node17398 = (inp[14]) ? node17414 : node17399;
													assign node17399 = (inp[3]) ? node17407 : node17400;
														assign node17400 = (inp[15]) ? node17404 : node17401;
															assign node17401 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node17404 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node17407 = (inp[0]) ? node17411 : node17408;
															assign node17408 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node17411 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node17414 = (inp[15]) ? node17420 : node17415;
														assign node17415 = (inp[0]) ? 4'b0000 : node17416;
															assign node17416 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node17420 = (inp[0]) ? node17424 : node17421;
															assign node17421 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node17424 = (inp[3]) ? 4'b0000 : 4'b0010;
								assign node17427 = (inp[1]) ? node17657 : node17428;
									assign node17428 = (inp[7]) ? node17550 : node17429;
										assign node17429 = (inp[8]) ? node17491 : node17430;
											assign node17430 = (inp[2]) ? node17460 : node17431;
												assign node17431 = (inp[14]) ? node17447 : node17432;
													assign node17432 = (inp[3]) ? node17440 : node17433;
														assign node17433 = (inp[5]) ? node17437 : node17434;
															assign node17434 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node17437 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node17440 = (inp[5]) ? node17444 : node17441;
															assign node17441 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node17444 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node17447 = (inp[0]) ? node17453 : node17448;
														assign node17448 = (inp[15]) ? 4'b1000 : node17449;
															assign node17449 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node17453 = (inp[15]) ? node17457 : node17454;
															assign node17454 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node17457 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node17460 = (inp[3]) ? node17476 : node17461;
													assign node17461 = (inp[14]) ? node17469 : node17462;
														assign node17462 = (inp[0]) ? node17466 : node17463;
															assign node17463 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node17466 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node17469 = (inp[0]) ? node17473 : node17470;
															assign node17470 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node17473 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node17476 = (inp[5]) ? node17484 : node17477;
														assign node17477 = (inp[0]) ? node17481 : node17478;
															assign node17478 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node17481 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node17484 = (inp[14]) ? node17488 : node17485;
															assign node17485 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node17488 = (inp[0]) ? 4'b1000 : 4'b1000;
											assign node17491 = (inp[14]) ? node17521 : node17492;
												assign node17492 = (inp[2]) ? node17506 : node17493;
													assign node17493 = (inp[5]) ? node17501 : node17494;
														assign node17494 = (inp[3]) ? node17498 : node17495;
															assign node17495 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node17498 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node17501 = (inp[0]) ? 4'b1010 : node17502;
															assign node17502 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node17506 = (inp[5]) ? node17514 : node17507;
														assign node17507 = (inp[3]) ? node17511 : node17508;
															assign node17508 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node17511 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node17514 = (inp[0]) ? node17518 : node17515;
															assign node17515 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node17518 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node17521 = (inp[3]) ? node17535 : node17522;
													assign node17522 = (inp[2]) ? node17530 : node17523;
														assign node17523 = (inp[15]) ? node17527 : node17524;
															assign node17524 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node17527 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node17530 = (inp[5]) ? 4'b0011 : node17531;
															assign node17531 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node17535 = (inp[0]) ? node17543 : node17536;
														assign node17536 = (inp[5]) ? node17540 : node17537;
															assign node17537 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node17540 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node17543 = (inp[5]) ? node17547 : node17544;
															assign node17544 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node17547 = (inp[15]) ? 4'b0001 : 4'b0011;
										assign node17550 = (inp[8]) ? node17604 : node17551;
											assign node17551 = (inp[2]) ? node17581 : node17552;
												assign node17552 = (inp[14]) ? node17568 : node17553;
													assign node17553 = (inp[15]) ? node17561 : node17554;
														assign node17554 = (inp[0]) ? node17558 : node17555;
															assign node17555 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node17558 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node17561 = (inp[0]) ? node17565 : node17562;
															assign node17562 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node17565 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node17568 = (inp[3]) ? node17574 : node17569;
														assign node17569 = (inp[5]) ? 4'b0011 : node17570;
															assign node17570 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node17574 = (inp[15]) ? node17578 : node17575;
															assign node17575 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node17578 = (inp[5]) ? 4'b0001 : 4'b0001;
												assign node17581 = (inp[15]) ? node17593 : node17582;
													assign node17582 = (inp[0]) ? node17588 : node17583;
														assign node17583 = (inp[5]) ? node17585 : 4'b0011;
															assign node17585 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node17588 = (inp[3]) ? node17590 : 4'b0001;
															assign node17590 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node17593 = (inp[0]) ? node17599 : node17594;
														assign node17594 = (inp[3]) ? node17596 : 4'b0001;
															assign node17596 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node17599 = (inp[5]) ? node17601 : 4'b0011;
															assign node17601 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node17604 = (inp[14]) ? node17634 : node17605;
												assign node17605 = (inp[2]) ? node17621 : node17606;
													assign node17606 = (inp[3]) ? node17614 : node17607;
														assign node17607 = (inp[0]) ? node17611 : node17608;
															assign node17608 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node17611 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node17614 = (inp[15]) ? node17618 : node17615;
															assign node17615 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node17618 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node17621 = (inp[3]) ? node17627 : node17622;
														assign node17622 = (inp[5]) ? node17624 : 4'b0010;
															assign node17624 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node17627 = (inp[5]) ? node17631 : node17628;
															assign node17628 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node17631 = (inp[0]) ? 4'b0000 : 4'b0000;
												assign node17634 = (inp[15]) ? node17646 : node17635;
													assign node17635 = (inp[0]) ? node17641 : node17636;
														assign node17636 = (inp[3]) ? node17638 : 4'b0010;
															assign node17638 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node17641 = (inp[5]) ? node17643 : 4'b0000;
															assign node17643 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node17646 = (inp[0]) ? node17652 : node17647;
														assign node17647 = (inp[5]) ? node17649 : 4'b0000;
															assign node17649 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node17652 = (inp[5]) ? node17654 : 4'b0010;
															assign node17654 = (inp[3]) ? 4'b0000 : 4'b0010;
									assign node17657 = (inp[2]) ? node17775 : node17658;
										assign node17658 = (inp[14]) ? node17718 : node17659;
											assign node17659 = (inp[15]) ? node17691 : node17660;
												assign node17660 = (inp[0]) ? node17676 : node17661;
													assign node17661 = (inp[5]) ? node17669 : node17662;
														assign node17662 = (inp[8]) ? node17666 : node17663;
															assign node17663 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node17666 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node17669 = (inp[3]) ? node17673 : node17670;
															assign node17670 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node17673 = (inp[8]) ? 4'b0000 : 4'b0000;
													assign node17676 = (inp[3]) ? node17684 : node17677;
														assign node17677 = (inp[7]) ? node17681 : node17678;
															assign node17678 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node17681 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node17684 = (inp[5]) ? node17688 : node17685;
															assign node17685 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node17688 = (inp[8]) ? 4'b0010 : 4'b0010;
												assign node17691 = (inp[0]) ? node17705 : node17692;
													assign node17692 = (inp[3]) ? node17698 : node17693;
														assign node17693 = (inp[7]) ? 4'b0000 : node17694;
															assign node17694 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node17698 = (inp[5]) ? node17702 : node17699;
															assign node17699 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node17702 = (inp[7]) ? 4'b0010 : 4'b0010;
													assign node17705 = (inp[3]) ? node17713 : node17706;
														assign node17706 = (inp[7]) ? node17710 : node17707;
															assign node17707 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node17710 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node17713 = (inp[5]) ? node17715 : 4'b0010;
															assign node17715 = (inp[8]) ? 4'b0000 : 4'b0000;
											assign node17718 = (inp[7]) ? node17750 : node17719;
												assign node17719 = (inp[8]) ? node17735 : node17720;
													assign node17720 = (inp[0]) ? node17728 : node17721;
														assign node17721 = (inp[15]) ? node17725 : node17722;
															assign node17722 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node17725 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node17728 = (inp[15]) ? node17732 : node17729;
															assign node17729 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node17732 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node17735 = (inp[5]) ? node17743 : node17736;
														assign node17736 = (inp[0]) ? node17740 : node17737;
															assign node17737 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node17740 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node17743 = (inp[0]) ? node17747 : node17744;
															assign node17744 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node17747 = (inp[3]) ? 4'b0001 : 4'b0001;
												assign node17750 = (inp[8]) ? node17764 : node17751;
													assign node17751 = (inp[3]) ? node17757 : node17752;
														assign node17752 = (inp[5]) ? 4'b0001 : node17753;
															assign node17753 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node17757 = (inp[15]) ? node17761 : node17758;
															assign node17758 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node17761 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node17764 = (inp[3]) ? node17770 : node17765;
														assign node17765 = (inp[5]) ? 4'b0000 : node17766;
															assign node17766 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node17770 = (inp[5]) ? node17772 : 4'b0000;
															assign node17772 = (inp[15]) ? 4'b0000 : 4'b0000;
										assign node17775 = (inp[0]) ? node17821 : node17776;
											assign node17776 = (inp[15]) ? node17798 : node17777;
												assign node17777 = (inp[5]) ? node17785 : node17778;
													assign node17778 = (inp[7]) ? node17782 : node17779;
														assign node17779 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node17782 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node17785 = (inp[3]) ? node17791 : node17786;
														assign node17786 = (inp[8]) ? node17788 : 4'b0011;
															assign node17788 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node17791 = (inp[14]) ? node17795 : node17792;
															assign node17792 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node17795 = (inp[8]) ? 4'b0000 : 4'b0000;
												assign node17798 = (inp[5]) ? node17806 : node17799;
													assign node17799 = (inp[7]) ? node17803 : node17800;
														assign node17800 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node17803 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node17806 = (inp[3]) ? node17814 : node17807;
														assign node17807 = (inp[14]) ? node17811 : node17808;
															assign node17808 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node17811 = (inp[7]) ? 4'b0000 : 4'b0000;
														assign node17814 = (inp[14]) ? node17818 : node17815;
															assign node17815 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node17818 = (inp[8]) ? 4'b0010 : 4'b0010;
											assign node17821 = (inp[15]) ? node17851 : node17822;
												assign node17822 = (inp[3]) ? node17838 : node17823;
													assign node17823 = (inp[5]) ? node17831 : node17824;
														assign node17824 = (inp[8]) ? node17828 : node17825;
															assign node17825 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node17828 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node17831 = (inp[8]) ? node17835 : node17832;
															assign node17832 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node17835 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node17838 = (inp[5]) ? node17844 : node17839;
														assign node17839 = (inp[7]) ? 4'b0000 : node17840;
															assign node17840 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node17844 = (inp[7]) ? node17848 : node17845;
															assign node17845 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node17848 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node17851 = (inp[5]) ? node17867 : node17852;
													assign node17852 = (inp[3]) ? node17860 : node17853;
														assign node17853 = (inp[7]) ? node17857 : node17854;
															assign node17854 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node17857 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node17860 = (inp[8]) ? node17864 : node17861;
															assign node17861 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node17864 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node17867 = (inp[3]) ? node17875 : node17868;
														assign node17868 = (inp[14]) ? node17872 : node17869;
															assign node17869 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node17872 = (inp[8]) ? 4'b0010 : 4'b0010;
														assign node17875 = (inp[7]) ? node17879 : node17876;
															assign node17876 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node17879 = (inp[8]) ? 4'b0000 : 4'b0001;
					assign node17882 = (inp[11]) ? node19676 : node17883;
						assign node17883 = (inp[6]) ? node18759 : node17884;
							assign node17884 = (inp[1]) ? node18326 : node17885;
								assign node17885 = (inp[13]) ? node18107 : node17886;
									assign node17886 = (inp[0]) ? node17990 : node17887;
										assign node17887 = (inp[15]) ? node17937 : node17888;
											assign node17888 = (inp[5]) ? node17912 : node17889;
												assign node17889 = (inp[2]) ? node17905 : node17890;
													assign node17890 = (inp[14]) ? node17898 : node17891;
														assign node17891 = (inp[7]) ? node17895 : node17892;
															assign node17892 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node17895 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node17898 = (inp[3]) ? node17902 : node17899;
															assign node17899 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node17902 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node17905 = (inp[8]) ? node17909 : node17906;
														assign node17906 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node17909 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node17912 = (inp[3]) ? node17926 : node17913;
													assign node17913 = (inp[7]) ? node17919 : node17914;
														assign node17914 = (inp[2]) ? 4'b1011 : node17915;
															assign node17915 = (inp[14]) ? 4'b1010 : 4'b1010;
														assign node17919 = (inp[8]) ? node17923 : node17920;
															assign node17920 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node17923 = (inp[14]) ? 4'b1010 : 4'b1010;
													assign node17926 = (inp[8]) ? node17932 : node17927;
														assign node17927 = (inp[7]) ? node17929 : 4'b1000;
															assign node17929 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node17932 = (inp[7]) ? 4'b1000 : node17933;
															assign node17933 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node17937 = (inp[5]) ? node17961 : node17938;
												assign node17938 = (inp[2]) ? node17954 : node17939;
													assign node17939 = (inp[8]) ? node17947 : node17940;
														assign node17940 = (inp[14]) ? node17944 : node17941;
															assign node17941 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node17944 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node17947 = (inp[7]) ? node17951 : node17948;
															assign node17948 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node17951 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node17954 = (inp[7]) ? node17958 : node17955;
														assign node17955 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node17958 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node17961 = (inp[3]) ? node17975 : node17962;
													assign node17962 = (inp[14]) ? node17970 : node17963;
														assign node17963 = (inp[7]) ? node17967 : node17964;
															assign node17964 = (inp[2]) ? 4'b1000 : 4'b1000;
															assign node17967 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node17970 = (inp[8]) ? node17972 : 4'b1000;
															assign node17972 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node17975 = (inp[8]) ? node17983 : node17976;
														assign node17976 = (inp[7]) ? node17980 : node17977;
															assign node17977 = (inp[2]) ? 4'b1010 : 4'b1010;
															assign node17980 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node17983 = (inp[7]) ? node17987 : node17984;
															assign node17984 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node17987 = (inp[14]) ? 4'b1010 : 4'b1010;
										assign node17990 = (inp[15]) ? node18046 : node17991;
											assign node17991 = (inp[3]) ? node18015 : node17992;
												assign node17992 = (inp[14]) ? node18008 : node17993;
													assign node17993 = (inp[8]) ? node18001 : node17994;
														assign node17994 = (inp[2]) ? node17998 : node17995;
															assign node17995 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node17998 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node18001 = (inp[2]) ? node18005 : node18002;
															assign node18002 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node18005 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node18008 = (inp[8]) ? node18012 : node18009;
														assign node18009 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node18012 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node18015 = (inp[5]) ? node18031 : node18016;
													assign node18016 = (inp[2]) ? node18024 : node18017;
														assign node18017 = (inp[14]) ? node18021 : node18018;
															assign node18018 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node18021 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node18024 = (inp[8]) ? node18028 : node18025;
															assign node18025 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node18028 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node18031 = (inp[7]) ? node18039 : node18032;
														assign node18032 = (inp[8]) ? node18036 : node18033;
															assign node18033 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node18036 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node18039 = (inp[8]) ? node18043 : node18040;
															assign node18040 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node18043 = (inp[2]) ? 4'b1010 : 4'b1010;
											assign node18046 = (inp[5]) ? node18078 : node18047;
												assign node18047 = (inp[14]) ? node18063 : node18048;
													assign node18048 = (inp[7]) ? node18056 : node18049;
														assign node18049 = (inp[3]) ? node18053 : node18050;
															assign node18050 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node18053 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node18056 = (inp[8]) ? node18060 : node18057;
															assign node18057 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node18060 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node18063 = (inp[2]) ? node18071 : node18064;
														assign node18064 = (inp[7]) ? node18068 : node18065;
															assign node18065 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node18068 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node18071 = (inp[3]) ? node18075 : node18072;
															assign node18072 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node18075 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node18078 = (inp[3]) ? node18092 : node18079;
													assign node18079 = (inp[7]) ? node18085 : node18080;
														assign node18080 = (inp[8]) ? node18082 : 4'b1010;
															assign node18082 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node18085 = (inp[8]) ? node18089 : node18086;
															assign node18086 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node18089 = (inp[2]) ? 4'b1010 : 4'b1010;
													assign node18092 = (inp[7]) ? node18100 : node18093;
														assign node18093 = (inp[8]) ? node18097 : node18094;
															assign node18094 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node18097 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node18100 = (inp[8]) ? node18104 : node18101;
															assign node18101 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node18104 = (inp[14]) ? 4'b1000 : 4'b1000;
									assign node18107 = (inp[8]) ? node18227 : node18108;
										assign node18108 = (inp[7]) ? node18172 : node18109;
											assign node18109 = (inp[2]) ? node18141 : node18110;
												assign node18110 = (inp[14]) ? node18126 : node18111;
													assign node18111 = (inp[3]) ? node18119 : node18112;
														assign node18112 = (inp[15]) ? node18116 : node18113;
															assign node18113 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node18116 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node18119 = (inp[0]) ? node18123 : node18120;
															assign node18120 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node18123 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node18126 = (inp[5]) ? node18134 : node18127;
														assign node18127 = (inp[3]) ? node18131 : node18128;
															assign node18128 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node18131 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node18134 = (inp[0]) ? node18138 : node18135;
															assign node18135 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node18138 = (inp[3]) ? 4'b1000 : 4'b1000;
												assign node18141 = (inp[14]) ? node18157 : node18142;
													assign node18142 = (inp[15]) ? node18150 : node18143;
														assign node18143 = (inp[0]) ? node18147 : node18144;
															assign node18144 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node18147 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node18150 = (inp[0]) ? node18154 : node18151;
															assign node18151 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node18154 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node18157 = (inp[15]) ? node18165 : node18158;
														assign node18158 = (inp[0]) ? node18162 : node18159;
															assign node18159 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node18162 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node18165 = (inp[0]) ? node18169 : node18166;
															assign node18166 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node18169 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node18172 = (inp[2]) ? node18204 : node18173;
												assign node18173 = (inp[14]) ? node18189 : node18174;
													assign node18174 = (inp[3]) ? node18182 : node18175;
														assign node18175 = (inp[5]) ? node18179 : node18176;
															assign node18176 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node18179 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node18182 = (inp[5]) ? node18186 : node18183;
															assign node18183 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node18186 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node18189 = (inp[0]) ? node18197 : node18190;
														assign node18190 = (inp[15]) ? node18194 : node18191;
															assign node18191 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node18194 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node18197 = (inp[15]) ? node18201 : node18198;
															assign node18198 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node18201 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node18204 = (inp[0]) ? node18216 : node18205;
													assign node18205 = (inp[15]) ? node18211 : node18206;
														assign node18206 = (inp[5]) ? node18208 : 4'b0011;
															assign node18208 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node18211 = (inp[3]) ? node18213 : 4'b0001;
															assign node18213 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node18216 = (inp[15]) ? node18222 : node18217;
														assign node18217 = (inp[5]) ? node18219 : 4'b0001;
															assign node18219 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node18222 = (inp[3]) ? node18224 : 4'b0011;
															assign node18224 = (inp[5]) ? 4'b0001 : 4'b0011;
										assign node18227 = (inp[7]) ? node18277 : node18228;
											assign node18228 = (inp[14]) ? node18254 : node18229;
												assign node18229 = (inp[2]) ? node18243 : node18230;
													assign node18230 = (inp[5]) ? node18238 : node18231;
														assign node18231 = (inp[0]) ? node18235 : node18232;
															assign node18232 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node18235 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node18238 = (inp[0]) ? node18240 : 4'b1000;
															assign node18240 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node18243 = (inp[0]) ? node18247 : node18244;
														assign node18244 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node18247 = (inp[15]) ? node18251 : node18248;
															assign node18248 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node18251 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node18254 = (inp[3]) ? node18262 : node18255;
													assign node18255 = (inp[15]) ? node18259 : node18256;
														assign node18256 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node18259 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node18262 = (inp[15]) ? node18270 : node18263;
														assign node18263 = (inp[0]) ? node18267 : node18264;
															assign node18264 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node18267 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node18270 = (inp[0]) ? node18274 : node18271;
															assign node18271 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node18274 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node18277 = (inp[14]) ? node18303 : node18278;
												assign node18278 = (inp[2]) ? node18292 : node18279;
													assign node18279 = (inp[15]) ? node18287 : node18280;
														assign node18280 = (inp[0]) ? node18284 : node18281;
															assign node18281 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node18284 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node18287 = (inp[5]) ? node18289 : 4'b0001;
															assign node18289 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node18292 = (inp[3]) ? node18298 : node18293;
														assign node18293 = (inp[15]) ? 4'b0000 : node18294;
															assign node18294 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node18298 = (inp[5]) ? node18300 : 4'b0010;
															assign node18300 = (inp[15]) ? 4'b0000 : 4'b0000;
												assign node18303 = (inp[15]) ? node18315 : node18304;
													assign node18304 = (inp[0]) ? node18310 : node18305;
														assign node18305 = (inp[3]) ? node18307 : 4'b0010;
															assign node18307 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node18310 = (inp[3]) ? node18312 : 4'b0000;
															assign node18312 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node18315 = (inp[0]) ? node18321 : node18316;
														assign node18316 = (inp[3]) ? node18318 : 4'b0000;
															assign node18318 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node18321 = (inp[5]) ? node18323 : 4'b0010;
															assign node18323 = (inp[3]) ? 4'b0000 : 4'b0010;
								assign node18326 = (inp[13]) ? node18538 : node18327;
									assign node18327 = (inp[8]) ? node18439 : node18328;
										assign node18328 = (inp[7]) ? node18386 : node18329;
											assign node18329 = (inp[2]) ? node18359 : node18330;
												assign node18330 = (inp[14]) ? node18346 : node18331;
													assign node18331 = (inp[5]) ? node18339 : node18332;
														assign node18332 = (inp[0]) ? node18336 : node18333;
															assign node18333 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node18336 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node18339 = (inp[3]) ? node18343 : node18340;
															assign node18340 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node18343 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node18346 = (inp[3]) ? node18354 : node18347;
														assign node18347 = (inp[0]) ? node18351 : node18348;
															assign node18348 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node18351 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node18354 = (inp[0]) ? node18356 : 4'b1010;
															assign node18356 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node18359 = (inp[14]) ? node18375 : node18360;
													assign node18360 = (inp[3]) ? node18368 : node18361;
														assign node18361 = (inp[5]) ? node18365 : node18362;
															assign node18362 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node18365 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node18368 = (inp[0]) ? node18372 : node18369;
															assign node18369 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node18372 = (inp[5]) ? 4'b1000 : 4'b1000;
													assign node18375 = (inp[15]) ? node18381 : node18376;
														assign node18376 = (inp[0]) ? node18378 : 4'b1010;
															assign node18378 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node18381 = (inp[0]) ? 4'b1010 : node18382;
															assign node18382 = (inp[5]) ? 4'b1000 : 4'b1000;
											assign node18386 = (inp[2]) ? node18416 : node18387;
												assign node18387 = (inp[14]) ? node18403 : node18388;
													assign node18388 = (inp[3]) ? node18396 : node18389;
														assign node18389 = (inp[0]) ? node18393 : node18390;
															assign node18390 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node18393 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node18396 = (inp[0]) ? node18400 : node18397;
															assign node18397 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node18400 = (inp[5]) ? 4'b1000 : 4'b1000;
													assign node18403 = (inp[3]) ? node18409 : node18404;
														assign node18404 = (inp[5]) ? node18406 : 4'b0011;
															assign node18406 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node18409 = (inp[15]) ? node18413 : node18410;
															assign node18410 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node18413 = (inp[5]) ? 4'b0001 : 4'b0001;
												assign node18416 = (inp[0]) ? node18428 : node18417;
													assign node18417 = (inp[15]) ? node18423 : node18418;
														assign node18418 = (inp[3]) ? node18420 : 4'b0011;
															assign node18420 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node18423 = (inp[5]) ? node18425 : 4'b0001;
															assign node18425 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node18428 = (inp[15]) ? node18434 : node18429;
														assign node18429 = (inp[5]) ? node18431 : 4'b0001;
															assign node18431 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node18434 = (inp[3]) ? node18436 : 4'b0011;
															assign node18436 = (inp[5]) ? 4'b0001 : 4'b0011;
										assign node18439 = (inp[7]) ? node18491 : node18440;
											assign node18440 = (inp[2]) ? node18468 : node18441;
												assign node18441 = (inp[14]) ? node18457 : node18442;
													assign node18442 = (inp[0]) ? node18450 : node18443;
														assign node18443 = (inp[15]) ? node18447 : node18444;
															assign node18444 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node18447 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node18450 = (inp[15]) ? node18454 : node18451;
															assign node18451 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node18454 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node18457 = (inp[15]) ? node18463 : node18458;
														assign node18458 = (inp[0]) ? node18460 : 4'b0011;
															assign node18460 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node18463 = (inp[0]) ? 4'b0011 : node18464;
															assign node18464 = (inp[3]) ? 4'b0001 : 4'b0001;
												assign node18468 = (inp[5]) ? node18476 : node18469;
													assign node18469 = (inp[0]) ? node18473 : node18470;
														assign node18470 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node18473 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node18476 = (inp[15]) ? node18484 : node18477;
														assign node18477 = (inp[3]) ? node18481 : node18478;
															assign node18478 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node18481 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node18484 = (inp[0]) ? node18488 : node18485;
															assign node18485 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node18488 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node18491 = (inp[2]) ? node18519 : node18492;
												assign node18492 = (inp[14]) ? node18506 : node18493;
													assign node18493 = (inp[3]) ? node18501 : node18494;
														assign node18494 = (inp[15]) ? node18498 : node18495;
															assign node18495 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node18498 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node18501 = (inp[15]) ? node18503 : 4'b0001;
															assign node18503 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node18506 = (inp[3]) ? node18514 : node18507;
														assign node18507 = (inp[0]) ? node18511 : node18508;
															assign node18508 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node18511 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node18514 = (inp[15]) ? 4'b0010 : node18515;
															assign node18515 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node18519 = (inp[0]) ? node18531 : node18520;
													assign node18520 = (inp[15]) ? node18526 : node18521;
														assign node18521 = (inp[5]) ? node18523 : 4'b0010;
															assign node18523 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node18526 = (inp[5]) ? node18528 : 4'b0000;
															assign node18528 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node18531 = (inp[15]) ? 4'b0010 : node18532;
														assign node18532 = (inp[5]) ? node18534 : 4'b0000;
															assign node18534 = (inp[3]) ? 4'b0010 : 4'b0000;
									assign node18538 = (inp[8]) ? node18646 : node18539;
										assign node18539 = (inp[7]) ? node18593 : node18540;
											assign node18540 = (inp[14]) ? node18570 : node18541;
												assign node18541 = (inp[2]) ? node18557 : node18542;
													assign node18542 = (inp[3]) ? node18550 : node18543;
														assign node18543 = (inp[15]) ? node18547 : node18544;
															assign node18544 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node18547 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node18550 = (inp[15]) ? node18554 : node18551;
															assign node18551 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node18554 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node18557 = (inp[0]) ? node18565 : node18558;
														assign node18558 = (inp[15]) ? node18562 : node18559;
															assign node18559 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node18562 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node18565 = (inp[3]) ? node18567 : 4'b0010;
															assign node18567 = (inp[15]) ? 4'b0000 : 4'b0000;
												assign node18570 = (inp[0]) ? node18582 : node18571;
													assign node18571 = (inp[15]) ? node18577 : node18572;
														assign node18572 = (inp[3]) ? node18574 : 4'b0010;
															assign node18574 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node18577 = (inp[5]) ? node18579 : 4'b0000;
															assign node18579 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node18582 = (inp[15]) ? node18588 : node18583;
														assign node18583 = (inp[2]) ? 4'b0000 : node18584;
															assign node18584 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node18588 = (inp[3]) ? node18590 : 4'b0010;
															assign node18590 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node18593 = (inp[14]) ? node18625 : node18594;
												assign node18594 = (inp[2]) ? node18610 : node18595;
													assign node18595 = (inp[3]) ? node18603 : node18596;
														assign node18596 = (inp[5]) ? node18600 : node18597;
															assign node18597 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node18600 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node18603 = (inp[0]) ? node18607 : node18604;
															assign node18604 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node18607 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node18610 = (inp[3]) ? node18618 : node18611;
														assign node18611 = (inp[15]) ? node18615 : node18612;
															assign node18612 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node18615 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node18618 = (inp[0]) ? node18622 : node18619;
															assign node18619 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node18622 = (inp[5]) ? 4'b0001 : 4'b0001;
												assign node18625 = (inp[3]) ? node18633 : node18626;
													assign node18626 = (inp[15]) ? node18630 : node18627;
														assign node18627 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node18630 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node18633 = (inp[2]) ? node18641 : node18634;
														assign node18634 = (inp[5]) ? node18638 : node18635;
															assign node18635 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node18638 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node18641 = (inp[5]) ? node18643 : 4'b0011;
															assign node18643 = (inp[15]) ? 4'b0001 : 4'b0001;
										assign node18646 = (inp[7]) ? node18698 : node18647;
											assign node18647 = (inp[14]) ? node18675 : node18648;
												assign node18648 = (inp[2]) ? node18662 : node18649;
													assign node18649 = (inp[0]) ? node18657 : node18650;
														assign node18650 = (inp[15]) ? node18654 : node18651;
															assign node18651 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node18654 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node18657 = (inp[5]) ? node18659 : 4'b0010;
															assign node18659 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node18662 = (inp[3]) ? node18668 : node18663;
														assign node18663 = (inp[5]) ? node18665 : 4'b0001;
															assign node18665 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node18668 = (inp[0]) ? node18672 : node18669;
															assign node18669 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node18672 = (inp[15]) ? 4'b0001 : 4'b0001;
												assign node18675 = (inp[15]) ? node18687 : node18676;
													assign node18676 = (inp[0]) ? node18682 : node18677;
														assign node18677 = (inp[3]) ? node18679 : 4'b0011;
															assign node18679 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node18682 = (inp[5]) ? node18684 : 4'b0001;
															assign node18684 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node18687 = (inp[0]) ? node18693 : node18688;
														assign node18688 = (inp[3]) ? node18690 : 4'b0001;
															assign node18690 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node18693 = (inp[3]) ? node18695 : 4'b0011;
															assign node18695 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node18698 = (inp[14]) ? node18728 : node18699;
												assign node18699 = (inp[2]) ? node18715 : node18700;
													assign node18700 = (inp[3]) ? node18708 : node18701;
														assign node18701 = (inp[5]) ? node18705 : node18702;
															assign node18702 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node18705 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node18708 = (inp[15]) ? node18712 : node18709;
															assign node18709 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node18712 = (inp[5]) ? 4'b0001 : 4'b0001;
													assign node18715 = (inp[3]) ? node18721 : node18716;
														assign node18716 = (inp[0]) ? node18718 : 4'b0000;
															assign node18718 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node18721 = (inp[5]) ? node18725 : node18722;
															assign node18722 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node18725 = (inp[0]) ? 4'b0000 : 4'b0000;
												assign node18728 = (inp[2]) ? node18744 : node18729;
													assign node18729 = (inp[3]) ? node18737 : node18730;
														assign node18730 = (inp[0]) ? node18734 : node18731;
															assign node18731 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node18734 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node18737 = (inp[15]) ? node18741 : node18738;
															assign node18738 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node18741 = (inp[5]) ? 4'b0000 : 4'b0000;
													assign node18744 = (inp[3]) ? node18752 : node18745;
														assign node18745 = (inp[0]) ? node18749 : node18746;
															assign node18746 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node18749 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node18752 = (inp[5]) ? node18756 : node18753;
															assign node18753 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node18756 = (inp[15]) ? 4'b0000 : 4'b0000;
							assign node18759 = (inp[1]) ? node19203 : node18760;
								assign node18760 = (inp[13]) ? node18982 : node18761;
									assign node18761 = (inp[0]) ? node18869 : node18762;
										assign node18762 = (inp[15]) ? node18814 : node18763;
											assign node18763 = (inp[5]) ? node18787 : node18764;
												assign node18764 = (inp[7]) ? node18776 : node18765;
													assign node18765 = (inp[8]) ? node18771 : node18766;
														assign node18766 = (inp[2]) ? 4'b0010 : node18767;
															assign node18767 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node18771 = (inp[14]) ? 4'b0011 : node18772;
															assign node18772 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node18776 = (inp[8]) ? node18782 : node18777;
														assign node18777 = (inp[2]) ? 4'b0011 : node18778;
															assign node18778 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node18782 = (inp[2]) ? 4'b0010 : node18783;
															assign node18783 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node18787 = (inp[3]) ? node18803 : node18788;
													assign node18788 = (inp[2]) ? node18796 : node18789;
														assign node18789 = (inp[8]) ? node18793 : node18790;
															assign node18790 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node18793 = (inp[14]) ? 4'b0010 : 4'b0010;
														assign node18796 = (inp[7]) ? node18800 : node18797;
															assign node18797 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node18800 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node18803 = (inp[7]) ? node18807 : node18804;
														assign node18804 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node18807 = (inp[8]) ? node18811 : node18808;
															assign node18808 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node18811 = (inp[2]) ? 4'b0000 : 4'b0000;
											assign node18814 = (inp[5]) ? node18838 : node18815;
												assign node18815 = (inp[14]) ? node18831 : node18816;
													assign node18816 = (inp[3]) ? node18824 : node18817;
														assign node18817 = (inp[7]) ? node18821 : node18818;
															assign node18818 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node18821 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node18824 = (inp[8]) ? node18828 : node18825;
															assign node18825 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node18828 = (inp[7]) ? 4'b0000 : 4'b0000;
													assign node18831 = (inp[8]) ? node18835 : node18832;
														assign node18832 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node18835 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node18838 = (inp[3]) ? node18854 : node18839;
													assign node18839 = (inp[7]) ? node18847 : node18840;
														assign node18840 = (inp[8]) ? node18844 : node18841;
															assign node18841 = (inp[2]) ? 4'b0000 : 4'b0000;
															assign node18844 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node18847 = (inp[8]) ? node18851 : node18848;
															assign node18848 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node18851 = (inp[14]) ? 4'b0000 : 4'b0001;
													assign node18854 = (inp[8]) ? node18862 : node18855;
														assign node18855 = (inp[7]) ? node18859 : node18856;
															assign node18856 = (inp[14]) ? 4'b0010 : 4'b0010;
															assign node18859 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node18862 = (inp[7]) ? node18866 : node18863;
															assign node18863 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node18866 = (inp[2]) ? 4'b0010 : 4'b0010;
										assign node18869 = (inp[15]) ? node18925 : node18870;
											assign node18870 = (inp[3]) ? node18894 : node18871;
												assign node18871 = (inp[8]) ? node18883 : node18872;
													assign node18872 = (inp[7]) ? node18878 : node18873;
														assign node18873 = (inp[2]) ? 4'b0000 : node18874;
															assign node18874 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node18878 = (inp[2]) ? 4'b0001 : node18879;
															assign node18879 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node18883 = (inp[7]) ? node18889 : node18884;
														assign node18884 = (inp[14]) ? 4'b0001 : node18885;
															assign node18885 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node18889 = (inp[14]) ? 4'b0000 : node18890;
															assign node18890 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node18894 = (inp[5]) ? node18910 : node18895;
													assign node18895 = (inp[14]) ? node18903 : node18896;
														assign node18896 = (inp[2]) ? node18900 : node18897;
															assign node18897 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node18900 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node18903 = (inp[2]) ? node18907 : node18904;
															assign node18904 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node18907 = (inp[7]) ? 4'b0000 : 4'b0000;
													assign node18910 = (inp[14]) ? node18918 : node18911;
														assign node18911 = (inp[8]) ? node18915 : node18912;
															assign node18912 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node18915 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node18918 = (inp[7]) ? node18922 : node18919;
															assign node18919 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node18922 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node18925 = (inp[3]) ? node18955 : node18926;
												assign node18926 = (inp[5]) ? node18942 : node18927;
													assign node18927 = (inp[14]) ? node18935 : node18928;
														assign node18928 = (inp[7]) ? node18932 : node18929;
															assign node18929 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node18932 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node18935 = (inp[2]) ? node18939 : node18936;
															assign node18936 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node18939 = (inp[7]) ? 4'b0010 : 4'b0010;
													assign node18942 = (inp[14]) ? node18948 : node18943;
														assign node18943 = (inp[2]) ? node18945 : 4'b0010;
															assign node18945 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node18948 = (inp[7]) ? node18952 : node18949;
															assign node18949 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node18952 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node18955 = (inp[5]) ? node18967 : node18956;
													assign node18956 = (inp[2]) ? node18962 : node18957;
														assign node18957 = (inp[7]) ? node18959 : 4'b0011;
															assign node18959 = (inp[14]) ? 4'b0010 : 4'b0010;
														assign node18962 = (inp[7]) ? 4'b0010 : node18963;
															assign node18963 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node18967 = (inp[2]) ? node18975 : node18968;
														assign node18968 = (inp[8]) ? node18972 : node18969;
															assign node18969 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node18972 = (inp[7]) ? 4'b0000 : 4'b0000;
														assign node18975 = (inp[7]) ? node18979 : node18976;
															assign node18976 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node18979 = (inp[8]) ? 4'b0000 : 4'b0001;
									assign node18982 = (inp[8]) ? node19088 : node18983;
										assign node18983 = (inp[7]) ? node19035 : node18984;
											assign node18984 = (inp[2]) ? node19012 : node18985;
												assign node18985 = (inp[14]) ? node18999 : node18986;
													assign node18986 = (inp[0]) ? node18992 : node18987;
														assign node18987 = (inp[15]) ? node18989 : 4'b0011;
															assign node18989 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node18992 = (inp[15]) ? node18996 : node18993;
															assign node18993 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node18996 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node18999 = (inp[5]) ? node19007 : node19000;
														assign node19000 = (inp[3]) ? node19004 : node19001;
															assign node19001 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node19004 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node19007 = (inp[3]) ? 4'b0000 : node19008;
															assign node19008 = (inp[15]) ? 4'b0000 : 4'b0000;
												assign node19012 = (inp[3]) ? node19020 : node19013;
													assign node19013 = (inp[0]) ? node19017 : node19014;
														assign node19014 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node19017 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node19020 = (inp[0]) ? node19028 : node19021;
														assign node19021 = (inp[14]) ? node19025 : node19022;
															assign node19022 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node19025 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node19028 = (inp[5]) ? node19032 : node19029;
															assign node19029 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node19032 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node19035 = (inp[2]) ? node19065 : node19036;
												assign node19036 = (inp[14]) ? node19052 : node19037;
													assign node19037 = (inp[15]) ? node19045 : node19038;
														assign node19038 = (inp[0]) ? node19042 : node19039;
															assign node19039 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node19042 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node19045 = (inp[0]) ? node19049 : node19046;
															assign node19046 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node19049 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node19052 = (inp[0]) ? node19060 : node19053;
														assign node19053 = (inp[15]) ? node19057 : node19054;
															assign node19054 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node19057 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node19060 = (inp[15]) ? 4'b1101 : node19061;
															assign node19061 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node19065 = (inp[0]) ? node19077 : node19066;
													assign node19066 = (inp[15]) ? node19072 : node19067;
														assign node19067 = (inp[5]) ? 4'b1101 : node19068;
															assign node19068 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node19072 = (inp[5]) ? 4'b1111 : node19073;
															assign node19073 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node19077 = (inp[15]) ? node19083 : node19078;
														assign node19078 = (inp[5]) ? 4'b1111 : node19079;
															assign node19079 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node19083 = (inp[5]) ? 4'b1101 : node19084;
															assign node19084 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node19088 = (inp[7]) ? node19144 : node19089;
											assign node19089 = (inp[2]) ? node19121 : node19090;
												assign node19090 = (inp[14]) ? node19106 : node19091;
													assign node19091 = (inp[3]) ? node19099 : node19092;
														assign node19092 = (inp[0]) ? node19096 : node19093;
															assign node19093 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node19096 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node19099 = (inp[0]) ? node19103 : node19100;
															assign node19100 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node19103 = (inp[5]) ? 4'b0000 : 4'b0000;
													assign node19106 = (inp[5]) ? node19114 : node19107;
														assign node19107 = (inp[3]) ? node19111 : node19108;
															assign node19108 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node19111 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node19114 = (inp[3]) ? node19118 : node19115;
															assign node19115 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node19118 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node19121 = (inp[5]) ? node19137 : node19122;
													assign node19122 = (inp[14]) ? node19130 : node19123;
														assign node19123 = (inp[3]) ? node19127 : node19124;
															assign node19124 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node19127 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node19130 = (inp[0]) ? node19134 : node19131;
															assign node19131 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node19134 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node19137 = (inp[15]) ? node19141 : node19138;
														assign node19138 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node19141 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node19144 = (inp[14]) ? node19174 : node19145;
												assign node19145 = (inp[2]) ? node19161 : node19146;
													assign node19146 = (inp[5]) ? node19154 : node19147;
														assign node19147 = (inp[0]) ? node19151 : node19148;
															assign node19148 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node19151 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node19154 = (inp[0]) ? node19158 : node19155;
															assign node19155 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node19158 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node19161 = (inp[15]) ? node19167 : node19162;
														assign node19162 = (inp[0]) ? node19164 : 4'b1100;
															assign node19164 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node19167 = (inp[0]) ? node19171 : node19168;
															assign node19168 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node19171 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node19174 = (inp[2]) ? node19190 : node19175;
													assign node19175 = (inp[5]) ? node19183 : node19176;
														assign node19176 = (inp[3]) ? node19180 : node19177;
															assign node19177 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node19180 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node19183 = (inp[15]) ? node19187 : node19184;
															assign node19184 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node19187 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node19190 = (inp[0]) ? node19196 : node19191;
														assign node19191 = (inp[15]) ? node19193 : 4'b1100;
															assign node19193 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node19196 = (inp[15]) ? node19200 : node19197;
															assign node19197 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node19200 = (inp[3]) ? 4'b1100 : 4'b1100;
								assign node19203 = (inp[13]) ? node19441 : node19204;
									assign node19204 = (inp[8]) ? node19322 : node19205;
										assign node19205 = (inp[7]) ? node19263 : node19206;
											assign node19206 = (inp[14]) ? node19232 : node19207;
												assign node19207 = (inp[2]) ? node19223 : node19208;
													assign node19208 = (inp[15]) ? node19216 : node19209;
														assign node19209 = (inp[0]) ? node19213 : node19210;
															assign node19210 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node19213 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node19216 = (inp[0]) ? node19220 : node19217;
															assign node19217 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node19220 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node19223 = (inp[5]) ? node19225 : 4'b0010;
														assign node19225 = (inp[15]) ? node19229 : node19226;
															assign node19226 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node19229 = (inp[3]) ? 4'b0000 : 4'b0000;
												assign node19232 = (inp[3]) ? node19248 : node19233;
													assign node19233 = (inp[5]) ? node19241 : node19234;
														assign node19234 = (inp[2]) ? node19238 : node19235;
															assign node19235 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node19238 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node19241 = (inp[0]) ? node19245 : node19242;
															assign node19242 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node19245 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node19248 = (inp[5]) ? node19256 : node19249;
														assign node19249 = (inp[2]) ? node19253 : node19250;
															assign node19250 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node19253 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node19256 = (inp[2]) ? node19260 : node19257;
															assign node19257 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node19260 = (inp[0]) ? 4'b0000 : 4'b0000;
											assign node19263 = (inp[2]) ? node19293 : node19264;
												assign node19264 = (inp[14]) ? node19280 : node19265;
													assign node19265 = (inp[5]) ? node19273 : node19266;
														assign node19266 = (inp[3]) ? node19270 : node19267;
															assign node19267 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node19270 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node19273 = (inp[3]) ? node19277 : node19274;
															assign node19274 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node19277 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node19280 = (inp[5]) ? node19286 : node19281;
														assign node19281 = (inp[15]) ? node19283 : 4'b1101;
															assign node19283 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node19286 = (inp[15]) ? node19290 : node19287;
															assign node19287 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node19290 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node19293 = (inp[14]) ? node19309 : node19294;
													assign node19294 = (inp[0]) ? node19302 : node19295;
														assign node19295 = (inp[15]) ? node19299 : node19296;
															assign node19296 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node19299 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node19302 = (inp[15]) ? node19306 : node19303;
															assign node19303 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node19306 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node19309 = (inp[0]) ? node19315 : node19310;
														assign node19310 = (inp[15]) ? 4'b1111 : node19311;
															assign node19311 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node19315 = (inp[15]) ? node19319 : node19316;
															assign node19316 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node19319 = (inp[5]) ? 4'b1101 : 4'b1101;
										assign node19322 = (inp[7]) ? node19384 : node19323;
											assign node19323 = (inp[14]) ? node19353 : node19324;
												assign node19324 = (inp[2]) ? node19340 : node19325;
													assign node19325 = (inp[5]) ? node19333 : node19326;
														assign node19326 = (inp[0]) ? node19330 : node19327;
															assign node19327 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node19330 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node19333 = (inp[15]) ? node19337 : node19334;
															assign node19334 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node19337 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node19340 = (inp[5]) ? node19346 : node19341;
														assign node19341 = (inp[15]) ? node19343 : 4'b1101;
															assign node19343 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node19346 = (inp[3]) ? node19350 : node19347;
															assign node19347 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node19350 = (inp[15]) ? 4'b1101 : 4'b1101;
												assign node19353 = (inp[2]) ? node19369 : node19354;
													assign node19354 = (inp[15]) ? node19362 : node19355;
														assign node19355 = (inp[0]) ? node19359 : node19356;
															assign node19356 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node19359 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node19362 = (inp[0]) ? node19366 : node19363;
															assign node19363 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node19366 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node19369 = (inp[5]) ? node19377 : node19370;
														assign node19370 = (inp[0]) ? node19374 : node19371;
															assign node19371 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node19374 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node19377 = (inp[15]) ? node19381 : node19378;
															assign node19378 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node19381 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node19384 = (inp[14]) ? node19416 : node19385;
												assign node19385 = (inp[2]) ? node19401 : node19386;
													assign node19386 = (inp[0]) ? node19394 : node19387;
														assign node19387 = (inp[15]) ? node19391 : node19388;
															assign node19388 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node19391 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node19394 = (inp[15]) ? node19398 : node19395;
															assign node19395 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node19398 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node19401 = (inp[3]) ? node19409 : node19402;
														assign node19402 = (inp[5]) ? node19406 : node19403;
															assign node19403 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node19406 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node19409 = (inp[15]) ? node19413 : node19410;
															assign node19410 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node19413 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node19416 = (inp[2]) ? node19432 : node19417;
													assign node19417 = (inp[0]) ? node19425 : node19418;
														assign node19418 = (inp[15]) ? node19422 : node19419;
															assign node19419 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node19422 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node19425 = (inp[15]) ? node19429 : node19426;
															assign node19426 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node19429 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node19432 = (inp[15]) ? node19438 : node19433;
														assign node19433 = (inp[0]) ? 4'b1110 : node19434;
															assign node19434 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node19438 = (inp[0]) ? 4'b1100 : 4'b1110;
									assign node19441 = (inp[15]) ? node19557 : node19442;
										assign node19442 = (inp[0]) ? node19496 : node19443;
											assign node19443 = (inp[5]) ? node19473 : node19444;
												assign node19444 = (inp[3]) ? node19458 : node19445;
													assign node19445 = (inp[8]) ? node19451 : node19446;
														assign node19446 = (inp[7]) ? 4'b1111 : node19447;
															assign node19447 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node19451 = (inp[7]) ? node19455 : node19452;
															assign node19452 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node19455 = (inp[2]) ? 4'b1110 : 4'b1110;
													assign node19458 = (inp[8]) ? node19466 : node19459;
														assign node19459 = (inp[7]) ? node19463 : node19460;
															assign node19460 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node19463 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node19466 = (inp[7]) ? node19470 : node19467;
															assign node19467 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node19470 = (inp[14]) ? 4'b1100 : 4'b1100;
												assign node19473 = (inp[14]) ? node19489 : node19474;
													assign node19474 = (inp[8]) ? node19482 : node19475;
														assign node19475 = (inp[3]) ? node19479 : node19476;
															assign node19476 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node19479 = (inp[2]) ? 4'b1100 : 4'b1100;
														assign node19482 = (inp[3]) ? node19486 : node19483;
															assign node19483 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node19486 = (inp[7]) ? 4'b1100 : 4'b1100;
													assign node19489 = (inp[7]) ? node19493 : node19490;
														assign node19490 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node19493 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node19496 = (inp[3]) ? node19526 : node19497;
												assign node19497 = (inp[5]) ? node19513 : node19498;
													assign node19498 = (inp[8]) ? node19506 : node19499;
														assign node19499 = (inp[7]) ? node19503 : node19500;
															assign node19500 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node19503 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node19506 = (inp[7]) ? node19510 : node19507;
															assign node19507 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node19510 = (inp[14]) ? 4'b1100 : 4'b1100;
													assign node19513 = (inp[7]) ? node19521 : node19514;
														assign node19514 = (inp[8]) ? node19518 : node19515;
															assign node19515 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node19518 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node19521 = (inp[8]) ? 4'b1110 : node19522;
															assign node19522 = (inp[14]) ? 4'b1111 : 4'b1110;
												assign node19526 = (inp[2]) ? node19542 : node19527;
													assign node19527 = (inp[8]) ? node19535 : node19528;
														assign node19528 = (inp[7]) ? node19532 : node19529;
															assign node19529 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node19532 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node19535 = (inp[14]) ? node19539 : node19536;
															assign node19536 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node19539 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node19542 = (inp[5]) ? node19550 : node19543;
														assign node19543 = (inp[14]) ? node19547 : node19544;
															assign node19544 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node19547 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node19550 = (inp[8]) ? node19554 : node19551;
															assign node19551 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node19554 = (inp[7]) ? 4'b1110 : 4'b1111;
										assign node19557 = (inp[0]) ? node19617 : node19558;
											assign node19558 = (inp[3]) ? node19586 : node19559;
												assign node19559 = (inp[5]) ? node19573 : node19560;
													assign node19560 = (inp[7]) ? node19566 : node19561;
														assign node19561 = (inp[8]) ? node19563 : 4'b1100;
															assign node19563 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node19566 = (inp[8]) ? node19570 : node19567;
															assign node19567 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node19570 = (inp[2]) ? 4'b1100 : 4'b1100;
													assign node19573 = (inp[2]) ? node19579 : node19574;
														assign node19574 = (inp[7]) ? 4'b1111 : node19575;
															assign node19575 = (inp[14]) ? 4'b1110 : 4'b1110;
														assign node19579 = (inp[7]) ? node19583 : node19580;
															assign node19580 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node19583 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node19586 = (inp[14]) ? node19602 : node19587;
													assign node19587 = (inp[7]) ? node19595 : node19588;
														assign node19588 = (inp[2]) ? node19592 : node19589;
															assign node19589 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node19592 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node19595 = (inp[2]) ? node19599 : node19596;
															assign node19596 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node19599 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node19602 = (inp[2]) ? node19610 : node19603;
														assign node19603 = (inp[5]) ? node19607 : node19604;
															assign node19604 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node19607 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node19610 = (inp[7]) ? node19614 : node19611;
															assign node19611 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node19614 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node19617 = (inp[3]) ? node19645 : node19618;
												assign node19618 = (inp[5]) ? node19634 : node19619;
													assign node19619 = (inp[2]) ? node19627 : node19620;
														assign node19620 = (inp[14]) ? node19624 : node19621;
															assign node19621 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node19624 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node19627 = (inp[14]) ? node19631 : node19628;
															assign node19628 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node19631 = (inp[7]) ? 4'b1110 : 4'b1110;
													assign node19634 = (inp[8]) ? node19638 : node19635;
														assign node19635 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node19638 = (inp[7]) ? node19642 : node19639;
															assign node19639 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node19642 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node19645 = (inp[2]) ? node19661 : node19646;
													assign node19646 = (inp[8]) ? node19654 : node19647;
														assign node19647 = (inp[7]) ? node19651 : node19648;
															assign node19648 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node19651 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node19654 = (inp[5]) ? node19658 : node19655;
															assign node19655 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node19658 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node19661 = (inp[14]) ? node19669 : node19662;
														assign node19662 = (inp[8]) ? node19666 : node19663;
															assign node19663 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node19666 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node19669 = (inp[5]) ? node19673 : node19670;
															assign node19670 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node19673 = (inp[8]) ? 4'b1100 : 4'b1100;
						assign node19676 = (inp[6]) ? node20584 : node19677;
							assign node19677 = (inp[1]) ? node20141 : node19678;
								assign node19678 = (inp[13]) ? node19924 : node19679;
									assign node19679 = (inp[5]) ? node19803 : node19680;
										assign node19680 = (inp[8]) ? node19742 : node19681;
											assign node19681 = (inp[7]) ? node19711 : node19682;
												assign node19682 = (inp[2]) ? node19696 : node19683;
													assign node19683 = (inp[14]) ? node19691 : node19684;
														assign node19684 = (inp[0]) ? node19688 : node19685;
															assign node19685 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node19688 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node19691 = (inp[3]) ? node19693 : 4'b0010;
															assign node19693 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node19696 = (inp[14]) ? node19704 : node19697;
														assign node19697 = (inp[3]) ? node19701 : node19698;
															assign node19698 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node19701 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node19704 = (inp[0]) ? node19708 : node19705;
															assign node19705 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node19708 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node19711 = (inp[2]) ? node19727 : node19712;
													assign node19712 = (inp[14]) ? node19720 : node19713;
														assign node19713 = (inp[0]) ? node19717 : node19714;
															assign node19714 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node19717 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node19720 = (inp[3]) ? node19724 : node19721;
															assign node19721 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node19724 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node19727 = (inp[14]) ? node19735 : node19728;
														assign node19728 = (inp[0]) ? node19732 : node19729;
															assign node19729 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node19732 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node19735 = (inp[3]) ? node19739 : node19736;
															assign node19736 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node19739 = (inp[15]) ? 4'b0001 : 4'b0001;
											assign node19742 = (inp[7]) ? node19774 : node19743;
												assign node19743 = (inp[14]) ? node19759 : node19744;
													assign node19744 = (inp[2]) ? node19752 : node19745;
														assign node19745 = (inp[3]) ? node19749 : node19746;
															assign node19746 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node19749 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node19752 = (inp[0]) ? node19756 : node19753;
															assign node19753 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node19756 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node19759 = (inp[3]) ? node19767 : node19760;
														assign node19760 = (inp[0]) ? node19764 : node19761;
															assign node19761 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node19764 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node19767 = (inp[2]) ? node19771 : node19768;
															assign node19768 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node19771 = (inp[0]) ? 4'b0001 : 4'b0001;
												assign node19774 = (inp[2]) ? node19788 : node19775;
													assign node19775 = (inp[14]) ? node19783 : node19776;
														assign node19776 = (inp[15]) ? node19780 : node19777;
															assign node19777 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node19780 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node19783 = (inp[3]) ? 4'b0000 : node19784;
															assign node19784 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node19788 = (inp[3]) ? node19796 : node19789;
														assign node19789 = (inp[0]) ? node19793 : node19790;
															assign node19790 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node19793 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node19796 = (inp[15]) ? node19800 : node19797;
															assign node19797 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node19800 = (inp[0]) ? 4'b0010 : 4'b0000;
										assign node19803 = (inp[15]) ? node19863 : node19804;
											assign node19804 = (inp[2]) ? node19832 : node19805;
												assign node19805 = (inp[7]) ? node19819 : node19806;
													assign node19806 = (inp[14]) ? node19812 : node19807;
														assign node19807 = (inp[8]) ? 4'b0010 : node19808;
															assign node19808 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node19812 = (inp[8]) ? node19816 : node19813;
															assign node19813 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node19816 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node19819 = (inp[3]) ? node19827 : node19820;
														assign node19820 = (inp[0]) ? node19824 : node19821;
															assign node19821 = (inp[14]) ? 4'b0010 : 4'b0010;
															assign node19824 = (inp[14]) ? 4'b0000 : 4'b0000;
														assign node19827 = (inp[0]) ? node19829 : 4'b0000;
															assign node19829 = (inp[8]) ? 4'b0010 : 4'b0010;
												assign node19832 = (inp[3]) ? node19848 : node19833;
													assign node19833 = (inp[0]) ? node19841 : node19834;
														assign node19834 = (inp[8]) ? node19838 : node19835;
															assign node19835 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node19838 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node19841 = (inp[7]) ? node19845 : node19842;
															assign node19842 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node19845 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node19848 = (inp[0]) ? node19856 : node19849;
														assign node19849 = (inp[7]) ? node19853 : node19850;
															assign node19850 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node19853 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node19856 = (inp[14]) ? node19860 : node19857;
															assign node19857 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node19860 = (inp[8]) ? 4'b0010 : 4'b0010;
											assign node19863 = (inp[14]) ? node19895 : node19864;
												assign node19864 = (inp[0]) ? node19880 : node19865;
													assign node19865 = (inp[3]) ? node19873 : node19866;
														assign node19866 = (inp[8]) ? node19870 : node19867;
															assign node19867 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node19870 = (inp[2]) ? 4'b0000 : 4'b0000;
														assign node19873 = (inp[2]) ? node19877 : node19874;
															assign node19874 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node19877 = (inp[7]) ? 4'b0010 : 4'b0010;
													assign node19880 = (inp[3]) ? node19888 : node19881;
														assign node19881 = (inp[7]) ? node19885 : node19882;
															assign node19882 = (inp[2]) ? 4'b0010 : 4'b0010;
															assign node19885 = (inp[2]) ? 4'b0010 : 4'b0010;
														assign node19888 = (inp[7]) ? node19892 : node19889;
															assign node19889 = (inp[2]) ? 4'b0000 : 4'b0000;
															assign node19892 = (inp[2]) ? 4'b0000 : 4'b0000;
												assign node19895 = (inp[8]) ? node19909 : node19896;
													assign node19896 = (inp[7]) ? node19904 : node19897;
														assign node19897 = (inp[0]) ? node19901 : node19898;
															assign node19898 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node19901 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node19904 = (inp[3]) ? 4'b0001 : node19905;
															assign node19905 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node19909 = (inp[7]) ? node19917 : node19910;
														assign node19910 = (inp[3]) ? node19914 : node19911;
															assign node19911 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node19914 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node19917 = (inp[3]) ? node19921 : node19918;
															assign node19918 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node19921 = (inp[0]) ? 4'b0000 : 4'b0010;
									assign node19924 = (inp[8]) ? node20034 : node19925;
										assign node19925 = (inp[7]) ? node19977 : node19926;
											assign node19926 = (inp[14]) ? node19956 : node19927;
												assign node19927 = (inp[2]) ? node19943 : node19928;
													assign node19928 = (inp[0]) ? node19936 : node19929;
														assign node19929 = (inp[15]) ? node19933 : node19930;
															assign node19930 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node19933 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node19936 = (inp[15]) ? node19940 : node19937;
															assign node19937 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node19940 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node19943 = (inp[15]) ? node19951 : node19944;
														assign node19944 = (inp[0]) ? node19948 : node19945;
															assign node19945 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node19948 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node19951 = (inp[0]) ? node19953 : 4'b0000;
															assign node19953 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node19956 = (inp[15]) ? node19968 : node19957;
													assign node19957 = (inp[0]) ? node19963 : node19958;
														assign node19958 = (inp[3]) ? node19960 : 4'b0010;
															assign node19960 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node19963 = (inp[3]) ? node19965 : 4'b0000;
															assign node19965 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node19968 = (inp[0]) ? node19974 : node19969;
														assign node19969 = (inp[5]) ? node19971 : 4'b0000;
															assign node19971 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node19974 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node19977 = (inp[14]) ? node20005 : node19978;
												assign node19978 = (inp[2]) ? node19992 : node19979;
													assign node19979 = (inp[3]) ? node19985 : node19980;
														assign node19980 = (inp[5]) ? node19982 : 4'b0000;
															assign node19982 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node19985 = (inp[15]) ? node19989 : node19986;
															assign node19986 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node19989 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node19992 = (inp[5]) ? node19998 : node19993;
														assign node19993 = (inp[0]) ? node19995 : 4'b1111;
															assign node19995 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node19998 = (inp[15]) ? node20002 : node19999;
															assign node19999 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node20002 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node20005 = (inp[3]) ? node20021 : node20006;
													assign node20006 = (inp[15]) ? node20014 : node20007;
														assign node20007 = (inp[5]) ? node20011 : node20008;
															assign node20008 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node20011 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node20014 = (inp[2]) ? node20018 : node20015;
															assign node20015 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node20018 = (inp[0]) ? 4'b1101 : 4'b1101;
													assign node20021 = (inp[5]) ? node20027 : node20022;
														assign node20022 = (inp[0]) ? node20024 : 4'b1111;
															assign node20024 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node20027 = (inp[2]) ? node20031 : node20028;
															assign node20028 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node20031 = (inp[15]) ? 4'b1101 : 4'b1101;
										assign node20034 = (inp[7]) ? node20090 : node20035;
											assign node20035 = (inp[14]) ? node20061 : node20036;
												assign node20036 = (inp[2]) ? node20048 : node20037;
													assign node20037 = (inp[0]) ? node20043 : node20038;
														assign node20038 = (inp[15]) ? 4'b0000 : node20039;
															assign node20039 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node20043 = (inp[15]) ? 4'b0010 : node20044;
															assign node20044 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node20048 = (inp[15]) ? node20056 : node20049;
														assign node20049 = (inp[0]) ? node20053 : node20050;
															assign node20050 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node20053 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node20056 = (inp[3]) ? 4'b1101 : node20057;
															assign node20057 = (inp[0]) ? 4'b1101 : 4'b1101;
												assign node20061 = (inp[2]) ? node20075 : node20062;
													assign node20062 = (inp[5]) ? node20070 : node20063;
														assign node20063 = (inp[0]) ? node20067 : node20064;
															assign node20064 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node20067 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node20070 = (inp[3]) ? 4'b1111 : node20071;
															assign node20071 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node20075 = (inp[15]) ? node20083 : node20076;
														assign node20076 = (inp[0]) ? node20080 : node20077;
															assign node20077 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node20080 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node20083 = (inp[0]) ? node20087 : node20084;
															assign node20084 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node20087 = (inp[5]) ? 4'b1101 : 4'b1101;
											assign node20090 = (inp[2]) ? node20118 : node20091;
												assign node20091 = (inp[14]) ? node20105 : node20092;
													assign node20092 = (inp[5]) ? node20098 : node20093;
														assign node20093 = (inp[0]) ? node20095 : 4'b1111;
															assign node20095 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node20098 = (inp[15]) ? node20102 : node20099;
															assign node20099 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node20102 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node20105 = (inp[5]) ? node20113 : node20106;
														assign node20106 = (inp[3]) ? node20110 : node20107;
															assign node20107 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node20110 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node20113 = (inp[3]) ? 4'b1100 : node20114;
															assign node20114 = (inp[15]) ? 4'b1100 : 4'b1100;
												assign node20118 = (inp[0]) ? node20130 : node20119;
													assign node20119 = (inp[15]) ? node20125 : node20120;
														assign node20120 = (inp[3]) ? 4'b1100 : node20121;
															assign node20121 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node20125 = (inp[3]) ? 4'b1110 : node20126;
															assign node20126 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node20130 = (inp[15]) ? node20136 : node20131;
														assign node20131 = (inp[3]) ? 4'b1110 : node20132;
															assign node20132 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node20136 = (inp[5]) ? 4'b1100 : node20137;
															assign node20137 = (inp[3]) ? 4'b1100 : 4'b1110;
								assign node20141 = (inp[13]) ? node20361 : node20142;
									assign node20142 = (inp[8]) ? node20254 : node20143;
										assign node20143 = (inp[7]) ? node20197 : node20144;
											assign node20144 = (inp[14]) ? node20174 : node20145;
												assign node20145 = (inp[2]) ? node20161 : node20146;
													assign node20146 = (inp[5]) ? node20154 : node20147;
														assign node20147 = (inp[3]) ? node20151 : node20148;
															assign node20148 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node20151 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node20154 = (inp[3]) ? node20158 : node20155;
															assign node20155 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node20158 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node20161 = (inp[5]) ? node20169 : node20162;
														assign node20162 = (inp[3]) ? node20166 : node20163;
															assign node20163 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node20166 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node20169 = (inp[3]) ? node20171 : 4'b0010;
															assign node20171 = (inp[15]) ? 4'b0000 : 4'b0000;
												assign node20174 = (inp[0]) ? node20186 : node20175;
													assign node20175 = (inp[15]) ? node20181 : node20176;
														assign node20176 = (inp[3]) ? node20178 : 4'b0010;
															assign node20178 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node20181 = (inp[5]) ? node20183 : 4'b0000;
															assign node20183 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node20186 = (inp[15]) ? node20192 : node20187;
														assign node20187 = (inp[5]) ? node20189 : 4'b0000;
															assign node20189 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node20192 = (inp[5]) ? node20194 : 4'b0010;
															assign node20194 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node20197 = (inp[2]) ? node20223 : node20198;
												assign node20198 = (inp[14]) ? node20214 : node20199;
													assign node20199 = (inp[3]) ? node20207 : node20200;
														assign node20200 = (inp[15]) ? node20204 : node20201;
															assign node20201 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node20204 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node20207 = (inp[15]) ? node20211 : node20208;
															assign node20208 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node20211 = (inp[5]) ? 4'b0000 : 4'b0000;
													assign node20214 = (inp[15]) ? node20218 : node20215;
														assign node20215 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node20218 = (inp[0]) ? node20220 : 4'b1111;
															assign node20220 = (inp[5]) ? 4'b1101 : 4'b1101;
												assign node20223 = (inp[14]) ? node20239 : node20224;
													assign node20224 = (inp[5]) ? node20232 : node20225;
														assign node20225 = (inp[15]) ? node20229 : node20226;
															assign node20226 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node20229 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node20232 = (inp[0]) ? node20236 : node20233;
															assign node20233 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node20236 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node20239 = (inp[15]) ? node20247 : node20240;
														assign node20240 = (inp[0]) ? node20244 : node20241;
															assign node20241 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node20244 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node20247 = (inp[0]) ? node20251 : node20248;
															assign node20248 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node20251 = (inp[5]) ? 4'b1101 : 4'b1101;
										assign node20254 = (inp[7]) ? node20308 : node20255;
											assign node20255 = (inp[14]) ? node20285 : node20256;
												assign node20256 = (inp[2]) ? node20272 : node20257;
													assign node20257 = (inp[5]) ? node20265 : node20258;
														assign node20258 = (inp[15]) ? node20262 : node20259;
															assign node20259 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node20262 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node20265 = (inp[0]) ? node20269 : node20266;
															assign node20266 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node20269 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node20272 = (inp[15]) ? node20280 : node20273;
														assign node20273 = (inp[0]) ? node20277 : node20274;
															assign node20274 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node20277 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node20280 = (inp[0]) ? 4'b1101 : node20281;
															assign node20281 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node20285 = (inp[15]) ? node20297 : node20286;
													assign node20286 = (inp[0]) ? node20292 : node20287;
														assign node20287 = (inp[3]) ? 4'b1101 : node20288;
															assign node20288 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node20292 = (inp[5]) ? 4'b1111 : node20293;
															assign node20293 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node20297 = (inp[0]) ? node20303 : node20298;
														assign node20298 = (inp[5]) ? 4'b1111 : node20299;
															assign node20299 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node20303 = (inp[5]) ? 4'b1101 : node20304;
															assign node20304 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node20308 = (inp[2]) ? node20338 : node20309;
												assign node20309 = (inp[14]) ? node20323 : node20310;
													assign node20310 = (inp[15]) ? node20316 : node20311;
														assign node20311 = (inp[0]) ? 4'b1111 : node20312;
															assign node20312 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node20316 = (inp[0]) ? node20320 : node20317;
															assign node20317 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node20320 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node20323 = (inp[0]) ? node20331 : node20324;
														assign node20324 = (inp[15]) ? node20328 : node20325;
															assign node20325 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node20328 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node20331 = (inp[15]) ? node20335 : node20332;
															assign node20332 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node20335 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node20338 = (inp[15]) ? node20350 : node20339;
													assign node20339 = (inp[0]) ? node20345 : node20340;
														assign node20340 = (inp[3]) ? 4'b1100 : node20341;
															assign node20341 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node20345 = (inp[5]) ? 4'b1110 : node20346;
															assign node20346 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node20350 = (inp[0]) ? node20356 : node20351;
														assign node20351 = (inp[5]) ? 4'b1110 : node20352;
															assign node20352 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node20356 = (inp[3]) ? 4'b1100 : node20357;
															assign node20357 = (inp[5]) ? 4'b1100 : 4'b1110;
									assign node20361 = (inp[0]) ? node20463 : node20362;
										assign node20362 = (inp[15]) ? node20414 : node20363;
											assign node20363 = (inp[3]) ? node20391 : node20364;
												assign node20364 = (inp[5]) ? node20378 : node20365;
													assign node20365 = (inp[7]) ? node20373 : node20366;
														assign node20366 = (inp[8]) ? node20370 : node20367;
															assign node20367 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node20370 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node20373 = (inp[8]) ? 4'b1110 : node20374;
															assign node20374 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node20378 = (inp[7]) ? node20386 : node20379;
														assign node20379 = (inp[8]) ? node20383 : node20380;
															assign node20380 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node20383 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node20386 = (inp[2]) ? 4'b1101 : node20387;
															assign node20387 = (inp[14]) ? 4'b1100 : 4'b1100;
												assign node20391 = (inp[8]) ? node20403 : node20392;
													assign node20392 = (inp[7]) ? node20398 : node20393;
														assign node20393 = (inp[2]) ? 4'b1100 : node20394;
															assign node20394 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node20398 = (inp[2]) ? 4'b1101 : node20399;
															assign node20399 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node20403 = (inp[7]) ? node20409 : node20404;
														assign node20404 = (inp[14]) ? 4'b1101 : node20405;
															assign node20405 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node20409 = (inp[2]) ? 4'b1100 : node20410;
															assign node20410 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node20414 = (inp[5]) ? node20440 : node20415;
												assign node20415 = (inp[3]) ? node20429 : node20416;
													assign node20416 = (inp[14]) ? node20422 : node20417;
														assign node20417 = (inp[2]) ? 4'b1100 : node20418;
															assign node20418 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node20422 = (inp[2]) ? node20426 : node20423;
															assign node20423 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node20426 = (inp[7]) ? 4'b1100 : 4'b1100;
													assign node20429 = (inp[8]) ? node20435 : node20430;
														assign node20430 = (inp[14]) ? 4'b1110 : node20431;
															assign node20431 = (inp[2]) ? 4'b1110 : 4'b1110;
														assign node20435 = (inp[7]) ? node20437 : 4'b1111;
															assign node20437 = (inp[14]) ? 4'b1110 : 4'b1110;
												assign node20440 = (inp[8]) ? node20452 : node20441;
													assign node20441 = (inp[7]) ? node20447 : node20442;
														assign node20442 = (inp[14]) ? 4'b1110 : node20443;
															assign node20443 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node20447 = (inp[14]) ? 4'b1111 : node20448;
															assign node20448 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node20452 = (inp[7]) ? node20458 : node20453;
														assign node20453 = (inp[14]) ? 4'b1111 : node20454;
															assign node20454 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node20458 = (inp[2]) ? 4'b1110 : node20459;
															assign node20459 = (inp[14]) ? 4'b1110 : 4'b1111;
										assign node20463 = (inp[15]) ? node20525 : node20464;
											assign node20464 = (inp[5]) ? node20494 : node20465;
												assign node20465 = (inp[3]) ? node20479 : node20466;
													assign node20466 = (inp[2]) ? node20472 : node20467;
														assign node20467 = (inp[7]) ? 4'b1101 : node20468;
															assign node20468 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node20472 = (inp[8]) ? node20476 : node20473;
															assign node20473 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node20476 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node20479 = (inp[14]) ? node20487 : node20480;
														assign node20480 = (inp[2]) ? node20484 : node20481;
															assign node20481 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node20484 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node20487 = (inp[7]) ? node20491 : node20488;
															assign node20488 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node20491 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node20494 = (inp[2]) ? node20510 : node20495;
													assign node20495 = (inp[14]) ? node20503 : node20496;
														assign node20496 = (inp[3]) ? node20500 : node20497;
															assign node20497 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node20500 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node20503 = (inp[3]) ? node20507 : node20504;
															assign node20504 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node20507 = (inp[7]) ? 4'b1110 : 4'b1110;
													assign node20510 = (inp[3]) ? node20518 : node20511;
														assign node20511 = (inp[7]) ? node20515 : node20512;
															assign node20512 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node20515 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node20518 = (inp[8]) ? node20522 : node20519;
															assign node20519 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node20522 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node20525 = (inp[5]) ? node20555 : node20526;
												assign node20526 = (inp[3]) ? node20542 : node20527;
													assign node20527 = (inp[7]) ? node20535 : node20528;
														assign node20528 = (inp[8]) ? node20532 : node20529;
															assign node20529 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node20532 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node20535 = (inp[8]) ? node20539 : node20536;
															assign node20536 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node20539 = (inp[2]) ? 4'b1110 : 4'b1110;
													assign node20542 = (inp[8]) ? node20550 : node20543;
														assign node20543 = (inp[7]) ? node20547 : node20544;
															assign node20544 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node20547 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node20550 = (inp[14]) ? 4'b1101 : node20551;
															assign node20551 = (inp[2]) ? 4'b1100 : 4'b1100;
												assign node20555 = (inp[3]) ? node20571 : node20556;
													assign node20556 = (inp[8]) ? node20564 : node20557;
														assign node20557 = (inp[7]) ? node20561 : node20558;
															assign node20558 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node20561 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node20564 = (inp[7]) ? node20568 : node20565;
															assign node20565 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node20568 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node20571 = (inp[2]) ? node20579 : node20572;
														assign node20572 = (inp[14]) ? node20576 : node20573;
															assign node20573 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node20576 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node20579 = (inp[14]) ? 4'b1100 : node20580;
															assign node20580 = (inp[7]) ? 4'b1100 : 4'b1100;
							assign node20584 = (inp[13]) ? node21040 : node20585;
								assign node20585 = (inp[1]) ? node20821 : node20586;
									assign node20586 = (inp[14]) ? node20712 : node20587;
										assign node20587 = (inp[8]) ? node20651 : node20588;
											assign node20588 = (inp[3]) ? node20620 : node20589;
												assign node20589 = (inp[7]) ? node20605 : node20590;
													assign node20590 = (inp[2]) ? node20598 : node20591;
														assign node20591 = (inp[15]) ? node20595 : node20592;
															assign node20592 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node20595 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node20598 = (inp[0]) ? node20602 : node20599;
															assign node20599 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node20602 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node20605 = (inp[2]) ? node20613 : node20606;
														assign node20606 = (inp[5]) ? node20610 : node20607;
															assign node20607 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node20610 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node20613 = (inp[0]) ? node20617 : node20614;
															assign node20614 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node20617 = (inp[15]) ? 4'b1101 : 4'b1101;
												assign node20620 = (inp[2]) ? node20636 : node20621;
													assign node20621 = (inp[7]) ? node20629 : node20622;
														assign node20622 = (inp[5]) ? node20626 : node20623;
															assign node20623 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node20626 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node20629 = (inp[5]) ? node20633 : node20630;
															assign node20630 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node20633 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node20636 = (inp[7]) ? node20644 : node20637;
														assign node20637 = (inp[5]) ? node20641 : node20638;
															assign node20638 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node20641 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node20644 = (inp[5]) ? node20648 : node20645;
															assign node20645 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node20648 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node20651 = (inp[15]) ? node20683 : node20652;
												assign node20652 = (inp[0]) ? node20668 : node20653;
													assign node20653 = (inp[3]) ? node20661 : node20654;
														assign node20654 = (inp[5]) ? node20658 : node20655;
															assign node20655 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node20658 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node20661 = (inp[2]) ? node20665 : node20662;
															assign node20662 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node20665 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node20668 = (inp[5]) ? node20676 : node20669;
														assign node20669 = (inp[3]) ? node20673 : node20670;
															assign node20670 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node20673 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node20676 = (inp[7]) ? node20680 : node20677;
															assign node20677 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node20680 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node20683 = (inp[0]) ? node20699 : node20684;
													assign node20684 = (inp[5]) ? node20692 : node20685;
														assign node20685 = (inp[3]) ? node20689 : node20686;
															assign node20686 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node20689 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node20692 = (inp[2]) ? node20696 : node20693;
															assign node20693 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node20696 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node20699 = (inp[3]) ? node20705 : node20700;
														assign node20700 = (inp[5]) ? node20702 : 4'b1110;
															assign node20702 = (inp[2]) ? 4'b1100 : 4'b1100;
														assign node20705 = (inp[5]) ? node20709 : node20706;
															assign node20706 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node20709 = (inp[7]) ? 4'b1100 : 4'b1100;
										assign node20712 = (inp[8]) ? node20766 : node20713;
											assign node20713 = (inp[7]) ? node20735 : node20714;
												assign node20714 = (inp[3]) ? node20728 : node20715;
													assign node20715 = (inp[5]) ? node20723 : node20716;
														assign node20716 = (inp[2]) ? node20720 : node20717;
															assign node20717 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node20720 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node20723 = (inp[0]) ? 4'b1110 : node20724;
															assign node20724 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node20728 = (inp[0]) ? node20732 : node20729;
														assign node20729 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node20732 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node20735 = (inp[5]) ? node20751 : node20736;
													assign node20736 = (inp[0]) ? node20744 : node20737;
														assign node20737 = (inp[2]) ? node20741 : node20738;
															assign node20738 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node20741 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node20744 = (inp[15]) ? node20748 : node20745;
															assign node20745 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node20748 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node20751 = (inp[3]) ? node20759 : node20752;
														assign node20752 = (inp[15]) ? node20756 : node20753;
															assign node20753 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node20756 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node20759 = (inp[2]) ? node20763 : node20760;
															assign node20760 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node20763 = (inp[15]) ? 4'b1101 : 4'b1101;
											assign node20766 = (inp[7]) ? node20790 : node20767;
												assign node20767 = (inp[0]) ? node20779 : node20768;
													assign node20768 = (inp[15]) ? node20774 : node20769;
														assign node20769 = (inp[5]) ? 4'b1101 : node20770;
															assign node20770 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node20774 = (inp[3]) ? 4'b1111 : node20775;
															assign node20775 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node20779 = (inp[15]) ? node20785 : node20780;
														assign node20780 = (inp[3]) ? 4'b1111 : node20781;
															assign node20781 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node20785 = (inp[3]) ? 4'b1101 : node20786;
															assign node20786 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node20790 = (inp[2]) ? node20806 : node20791;
													assign node20791 = (inp[3]) ? node20799 : node20792;
														assign node20792 = (inp[0]) ? node20796 : node20793;
															assign node20793 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node20796 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node20799 = (inp[5]) ? node20803 : node20800;
															assign node20800 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node20803 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node20806 = (inp[5]) ? node20814 : node20807;
														assign node20807 = (inp[15]) ? node20811 : node20808;
															assign node20808 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node20811 = (inp[3]) ? 4'b1100 : 4'b1100;
														assign node20814 = (inp[15]) ? node20818 : node20815;
															assign node20815 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node20818 = (inp[0]) ? 4'b1100 : 4'b1110;
									assign node20821 = (inp[8]) ? node20939 : node20822;
										assign node20822 = (inp[7]) ? node20880 : node20823;
											assign node20823 = (inp[14]) ? node20851 : node20824;
												assign node20824 = (inp[2]) ? node20838 : node20825;
													assign node20825 = (inp[0]) ? node20833 : node20826;
														assign node20826 = (inp[15]) ? node20830 : node20827;
															assign node20827 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node20830 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node20833 = (inp[15]) ? node20835 : 4'b1111;
															assign node20835 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node20838 = (inp[5]) ? node20844 : node20839;
														assign node20839 = (inp[0]) ? 4'b1100 : node20840;
															assign node20840 = (inp[3]) ? 4'b1100 : 4'b1100;
														assign node20844 = (inp[3]) ? node20848 : node20845;
															assign node20845 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node20848 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node20851 = (inp[5]) ? node20865 : node20852;
													assign node20852 = (inp[2]) ? node20860 : node20853;
														assign node20853 = (inp[3]) ? node20857 : node20854;
															assign node20854 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node20857 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node20860 = (inp[15]) ? node20862 : 4'b1100;
															assign node20862 = (inp[0]) ? 4'b1100 : 4'b1100;
													assign node20865 = (inp[3]) ? node20873 : node20866;
														assign node20866 = (inp[15]) ? node20870 : node20867;
															assign node20867 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node20870 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node20873 = (inp[0]) ? node20877 : node20874;
															assign node20874 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node20877 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node20880 = (inp[14]) ? node20910 : node20881;
												assign node20881 = (inp[2]) ? node20897 : node20882;
													assign node20882 = (inp[15]) ? node20890 : node20883;
														assign node20883 = (inp[0]) ? node20887 : node20884;
															assign node20884 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node20887 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node20890 = (inp[0]) ? node20894 : node20891;
															assign node20891 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node20894 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node20897 = (inp[0]) ? node20905 : node20898;
														assign node20898 = (inp[15]) ? node20902 : node20899;
															assign node20899 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node20902 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node20905 = (inp[5]) ? 4'b0111 : node20906;
															assign node20906 = (inp[3]) ? 4'b0101 : 4'b0101;
												assign node20910 = (inp[3]) ? node20924 : node20911;
													assign node20911 = (inp[5]) ? node20919 : node20912;
														assign node20912 = (inp[15]) ? node20916 : node20913;
															assign node20913 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node20916 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node20919 = (inp[2]) ? 4'b0101 : node20920;
															assign node20920 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node20924 = (inp[2]) ? node20932 : node20925;
														assign node20925 = (inp[15]) ? node20929 : node20926;
															assign node20926 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node20929 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node20932 = (inp[15]) ? node20936 : node20933;
															assign node20933 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node20936 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node20939 = (inp[7]) ? node20991 : node20940;
											assign node20940 = (inp[14]) ? node20970 : node20941;
												assign node20941 = (inp[2]) ? node20957 : node20942;
													assign node20942 = (inp[0]) ? node20950 : node20943;
														assign node20943 = (inp[15]) ? node20947 : node20944;
															assign node20944 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node20947 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node20950 = (inp[15]) ? node20954 : node20951;
															assign node20951 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node20954 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node20957 = (inp[15]) ? node20963 : node20958;
														assign node20958 = (inp[3]) ? 4'b0101 : node20959;
															assign node20959 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node20963 = (inp[0]) ? node20967 : node20964;
															assign node20964 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node20967 = (inp[3]) ? 4'b0101 : 4'b0101;
												assign node20970 = (inp[5]) ? node20984 : node20971;
													assign node20971 = (inp[2]) ? node20979 : node20972;
														assign node20972 = (inp[0]) ? node20976 : node20973;
															assign node20973 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node20976 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node20979 = (inp[3]) ? 4'b0111 : node20980;
															assign node20980 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node20984 = (inp[15]) ? node20988 : node20985;
														assign node20985 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node20988 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node20991 = (inp[14]) ? node21019 : node20992;
												assign node20992 = (inp[2]) ? node21006 : node20993;
													assign node20993 = (inp[5]) ? node21001 : node20994;
														assign node20994 = (inp[0]) ? node20998 : node20995;
															assign node20995 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node20998 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node21001 = (inp[15]) ? node21003 : 4'b0101;
															assign node21003 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node21006 = (inp[0]) ? node21012 : node21007;
														assign node21007 = (inp[15]) ? node21009 : 4'b0100;
															assign node21009 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node21012 = (inp[15]) ? node21016 : node21013;
															assign node21013 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node21016 = (inp[3]) ? 4'b0100 : 4'b0100;
												assign node21019 = (inp[5]) ? node21033 : node21020;
													assign node21020 = (inp[2]) ? node21028 : node21021;
														assign node21021 = (inp[15]) ? node21025 : node21022;
															assign node21022 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node21025 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node21028 = (inp[3]) ? node21030 : 4'b0100;
															assign node21030 = (inp[0]) ? 4'b0100 : 4'b0100;
													assign node21033 = (inp[0]) ? node21037 : node21034;
														assign node21034 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node21037 = (inp[15]) ? 4'b0100 : 4'b0110;
								assign node21040 = (inp[1]) ? node21264 : node21041;
									assign node21041 = (inp[8]) ? node21153 : node21042;
										assign node21042 = (inp[7]) ? node21100 : node21043;
											assign node21043 = (inp[14]) ? node21069 : node21044;
												assign node21044 = (inp[2]) ? node21058 : node21045;
													assign node21045 = (inp[3]) ? node21053 : node21046;
														assign node21046 = (inp[0]) ? node21050 : node21047;
															assign node21047 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node21050 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node21053 = (inp[5]) ? 4'b1101 : node21054;
															assign node21054 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node21058 = (inp[5]) ? node21064 : node21059;
														assign node21059 = (inp[0]) ? 4'b1100 : node21060;
															assign node21060 = (inp[3]) ? 4'b1100 : 4'b1100;
														assign node21064 = (inp[3]) ? 4'b1110 : node21065;
															assign node21065 = (inp[15]) ? 4'b1100 : 4'b1100;
												assign node21069 = (inp[3]) ? node21085 : node21070;
													assign node21070 = (inp[15]) ? node21078 : node21071;
														assign node21071 = (inp[2]) ? node21075 : node21072;
															assign node21072 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node21075 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node21078 = (inp[5]) ? node21082 : node21079;
															assign node21079 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node21082 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node21085 = (inp[2]) ? node21093 : node21086;
														assign node21086 = (inp[0]) ? node21090 : node21087;
															assign node21087 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node21090 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node21093 = (inp[15]) ? node21097 : node21094;
															assign node21094 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node21097 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node21100 = (inp[14]) ? node21130 : node21101;
												assign node21101 = (inp[2]) ? node21117 : node21102;
													assign node21102 = (inp[3]) ? node21110 : node21103;
														assign node21103 = (inp[5]) ? node21107 : node21104;
															assign node21104 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node21107 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node21110 = (inp[0]) ? node21114 : node21111;
															assign node21111 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node21114 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node21117 = (inp[3]) ? node21123 : node21118;
														assign node21118 = (inp[15]) ? node21120 : 4'b0111;
															assign node21120 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node21123 = (inp[15]) ? node21127 : node21124;
															assign node21124 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node21127 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node21130 = (inp[0]) ? node21142 : node21131;
													assign node21131 = (inp[15]) ? node21137 : node21132;
														assign node21132 = (inp[5]) ? 4'b0101 : node21133;
															assign node21133 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node21137 = (inp[5]) ? 4'b0111 : node21138;
															assign node21138 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node21142 = (inp[15]) ? node21148 : node21143;
														assign node21143 = (inp[5]) ? 4'b0111 : node21144;
															assign node21144 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node21148 = (inp[5]) ? 4'b0101 : node21149;
															assign node21149 = (inp[3]) ? 4'b0101 : 4'b0111;
										assign node21153 = (inp[7]) ? node21205 : node21154;
											assign node21154 = (inp[2]) ? node21182 : node21155;
												assign node21155 = (inp[14]) ? node21169 : node21156;
													assign node21156 = (inp[5]) ? node21164 : node21157;
														assign node21157 = (inp[0]) ? node21161 : node21158;
															assign node21158 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node21161 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node21164 = (inp[3]) ? node21166 : 4'b1100;
															assign node21166 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node21169 = (inp[3]) ? node21175 : node21170;
														assign node21170 = (inp[5]) ? 4'b0101 : node21171;
															assign node21171 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node21175 = (inp[0]) ? node21179 : node21176;
															assign node21176 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node21179 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node21182 = (inp[5]) ? node21198 : node21183;
													assign node21183 = (inp[0]) ? node21191 : node21184;
														assign node21184 = (inp[15]) ? node21188 : node21185;
															assign node21185 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node21188 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node21191 = (inp[14]) ? node21195 : node21192;
															assign node21192 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node21195 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node21198 = (inp[15]) ? node21202 : node21199;
														assign node21199 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node21202 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node21205 = (inp[14]) ? node21233 : node21206;
												assign node21206 = (inp[2]) ? node21220 : node21207;
													assign node21207 = (inp[5]) ? node21213 : node21208;
														assign node21208 = (inp[15]) ? 4'b0111 : node21209;
															assign node21209 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node21213 = (inp[15]) ? node21217 : node21214;
															assign node21214 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node21217 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node21220 = (inp[15]) ? node21228 : node21221;
														assign node21221 = (inp[0]) ? node21225 : node21222;
															assign node21222 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node21225 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node21228 = (inp[0]) ? node21230 : 4'b0110;
															assign node21230 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node21233 = (inp[2]) ? node21249 : node21234;
													assign node21234 = (inp[3]) ? node21242 : node21235;
														assign node21235 = (inp[0]) ? node21239 : node21236;
															assign node21236 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node21239 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node21242 = (inp[0]) ? node21246 : node21243;
															assign node21243 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node21246 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node21249 = (inp[3]) ? node21257 : node21250;
														assign node21250 = (inp[0]) ? node21254 : node21251;
															assign node21251 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node21254 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node21257 = (inp[5]) ? node21261 : node21258;
															assign node21258 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node21261 = (inp[0]) ? 4'b0100 : 4'b0100;
									assign node21264 = (inp[0]) ? node21374 : node21265;
										assign node21265 = (inp[15]) ? node21321 : node21266;
											assign node21266 = (inp[5]) ? node21298 : node21267;
												assign node21267 = (inp[3]) ? node21283 : node21268;
													assign node21268 = (inp[7]) ? node21276 : node21269;
														assign node21269 = (inp[8]) ? node21273 : node21270;
															assign node21270 = (inp[2]) ? 4'b0110 : 4'b0110;
															assign node21273 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node21276 = (inp[8]) ? node21280 : node21277;
															assign node21277 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node21280 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node21283 = (inp[7]) ? node21291 : node21284;
														assign node21284 = (inp[8]) ? node21288 : node21285;
															assign node21285 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node21288 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node21291 = (inp[8]) ? node21295 : node21292;
															assign node21292 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node21295 = (inp[2]) ? 4'b0100 : 4'b0100;
												assign node21298 = (inp[8]) ? node21310 : node21299;
													assign node21299 = (inp[7]) ? node21305 : node21300;
														assign node21300 = (inp[14]) ? 4'b0100 : node21301;
															assign node21301 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node21305 = (inp[2]) ? 4'b0101 : node21306;
															assign node21306 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node21310 = (inp[7]) ? node21316 : node21311;
														assign node21311 = (inp[2]) ? 4'b0101 : node21312;
															assign node21312 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node21316 = (inp[14]) ? 4'b0100 : node21317;
															assign node21317 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node21321 = (inp[3]) ? node21351 : node21322;
												assign node21322 = (inp[5]) ? node21338 : node21323;
													assign node21323 = (inp[2]) ? node21331 : node21324;
														assign node21324 = (inp[7]) ? node21328 : node21325;
															assign node21325 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node21328 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node21331 = (inp[14]) ? node21335 : node21332;
															assign node21332 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node21335 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node21338 = (inp[7]) ? node21344 : node21339;
														assign node21339 = (inp[14]) ? 4'b0111 : node21340;
															assign node21340 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node21344 = (inp[8]) ? node21348 : node21345;
															assign node21345 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node21348 = (inp[14]) ? 4'b0110 : 4'b0110;
												assign node21351 = (inp[8]) ? node21363 : node21352;
													assign node21352 = (inp[7]) ? node21358 : node21353;
														assign node21353 = (inp[14]) ? 4'b0110 : node21354;
															assign node21354 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node21358 = (inp[2]) ? 4'b0111 : node21359;
															assign node21359 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node21363 = (inp[7]) ? node21369 : node21364;
														assign node21364 = (inp[2]) ? 4'b0111 : node21365;
															assign node21365 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node21369 = (inp[2]) ? 4'b0110 : node21370;
															assign node21370 = (inp[14]) ? 4'b0110 : 4'b0111;
										assign node21374 = (inp[15]) ? node21436 : node21375;
											assign node21375 = (inp[5]) ? node21405 : node21376;
												assign node21376 = (inp[3]) ? node21390 : node21377;
													assign node21377 = (inp[2]) ? node21385 : node21378;
														assign node21378 = (inp[8]) ? node21382 : node21379;
															assign node21379 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node21382 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node21385 = (inp[14]) ? 4'b0100 : node21386;
															assign node21386 = (inp[8]) ? 4'b0100 : 4'b0100;
													assign node21390 = (inp[7]) ? node21398 : node21391;
														assign node21391 = (inp[8]) ? node21395 : node21392;
															assign node21392 = (inp[2]) ? 4'b0110 : 4'b0110;
															assign node21395 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node21398 = (inp[8]) ? node21402 : node21399;
															assign node21399 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node21402 = (inp[2]) ? 4'b0110 : 4'b0110;
												assign node21405 = (inp[14]) ? node21421 : node21406;
													assign node21406 = (inp[7]) ? node21414 : node21407;
														assign node21407 = (inp[8]) ? node21411 : node21408;
															assign node21408 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node21411 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node21414 = (inp[3]) ? node21418 : node21415;
															assign node21415 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node21418 = (inp[8]) ? 4'b0110 : 4'b0110;
													assign node21421 = (inp[3]) ? node21429 : node21422;
														assign node21422 = (inp[8]) ? node21426 : node21423;
															assign node21423 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node21426 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node21429 = (inp[7]) ? node21433 : node21430;
															assign node21430 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node21433 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node21436 = (inp[5]) ? node21468 : node21437;
												assign node21437 = (inp[3]) ? node21453 : node21438;
													assign node21438 = (inp[2]) ? node21446 : node21439;
														assign node21439 = (inp[8]) ? node21443 : node21440;
															assign node21440 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node21443 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node21446 = (inp[7]) ? node21450 : node21447;
															assign node21447 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node21450 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node21453 = (inp[14]) ? node21461 : node21454;
														assign node21454 = (inp[7]) ? node21458 : node21455;
															assign node21455 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node21458 = (inp[2]) ? 4'b0100 : 4'b0100;
														assign node21461 = (inp[2]) ? node21465 : node21462;
															assign node21462 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node21465 = (inp[7]) ? 4'b0100 : 4'b0100;
												assign node21468 = (inp[8]) ? node21480 : node21469;
													assign node21469 = (inp[7]) ? node21475 : node21470;
														assign node21470 = (inp[14]) ? 4'b0100 : node21471;
															assign node21471 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node21475 = (inp[14]) ? 4'b0101 : node21476;
															assign node21476 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node21480 = (inp[7]) ? node21482 : 4'b0101;
														assign node21482 = (inp[2]) ? 4'b0100 : node21483;
															assign node21483 = (inp[14]) ? 4'b0100 : 4'b0101;
				assign node21487 = (inp[12]) ? node25083 : node21488;
					assign node21488 = (inp[6]) ? node23278 : node21489;
						assign node21489 = (inp[11]) ? node22355 : node21490;
							assign node21490 = (inp[13]) ? node21928 : node21491;
								assign node21491 = (inp[1]) ? node21699 : node21492;
									assign node21492 = (inp[0]) ? node21596 : node21493;
										assign node21493 = (inp[15]) ? node21547 : node21494;
											assign node21494 = (inp[5]) ? node21518 : node21495;
												assign node21495 = (inp[7]) ? node21507 : node21496;
													assign node21496 = (inp[8]) ? node21502 : node21497;
														assign node21497 = (inp[14]) ? 4'b1010 : node21498;
															assign node21498 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node21502 = (inp[2]) ? 4'b1011 : node21503;
															assign node21503 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node21507 = (inp[8]) ? node21513 : node21508;
														assign node21508 = (inp[14]) ? 4'b1011 : node21509;
															assign node21509 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node21513 = (inp[14]) ? 4'b1010 : node21514;
															assign node21514 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node21518 = (inp[3]) ? node21532 : node21519;
													assign node21519 = (inp[2]) ? node21525 : node21520;
														assign node21520 = (inp[14]) ? node21522 : 4'b1010;
															assign node21522 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node21525 = (inp[8]) ? node21529 : node21526;
															assign node21526 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node21529 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node21532 = (inp[8]) ? node21540 : node21533;
														assign node21533 = (inp[7]) ? node21537 : node21534;
															assign node21534 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node21537 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node21540 = (inp[7]) ? node21544 : node21541;
															assign node21541 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node21544 = (inp[2]) ? 4'b1000 : 4'b1000;
											assign node21547 = (inp[3]) ? node21569 : node21548;
												assign node21548 = (inp[14]) ? node21562 : node21549;
													assign node21549 = (inp[8]) ? node21555 : node21550;
														assign node21550 = (inp[2]) ? node21552 : 4'b1000;
															assign node21552 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node21555 = (inp[5]) ? node21559 : node21556;
															assign node21556 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node21559 = (inp[7]) ? 4'b1000 : 4'b1000;
													assign node21562 = (inp[7]) ? node21566 : node21563;
														assign node21563 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node21566 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node21569 = (inp[5]) ? node21583 : node21570;
													assign node21570 = (inp[7]) ? node21576 : node21571;
														assign node21571 = (inp[8]) ? node21573 : 4'b1000;
															assign node21573 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node21576 = (inp[8]) ? node21580 : node21577;
															assign node21577 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node21580 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node21583 = (inp[2]) ? node21589 : node21584;
														assign node21584 = (inp[8]) ? node21586 : 4'b1010;
															assign node21586 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node21589 = (inp[8]) ? node21593 : node21590;
															assign node21590 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node21593 = (inp[7]) ? 4'b1010 : 4'b1011;
										assign node21596 = (inp[15]) ? node21646 : node21597;
											assign node21597 = (inp[5]) ? node21621 : node21598;
												assign node21598 = (inp[8]) ? node21610 : node21599;
													assign node21599 = (inp[7]) ? node21605 : node21600;
														assign node21600 = (inp[14]) ? 4'b1000 : node21601;
															assign node21601 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node21605 = (inp[14]) ? 4'b1001 : node21606;
															assign node21606 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node21610 = (inp[7]) ? node21616 : node21611;
														assign node21611 = (inp[2]) ? 4'b1001 : node21612;
															assign node21612 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node21616 = (inp[14]) ? 4'b1000 : node21617;
															assign node21617 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node21621 = (inp[3]) ? node21635 : node21622;
													assign node21622 = (inp[14]) ? node21628 : node21623;
														assign node21623 = (inp[2]) ? 4'b1000 : node21624;
															assign node21624 = (inp[7]) ? 4'b1000 : 4'b1000;
														assign node21628 = (inp[2]) ? node21632 : node21629;
															assign node21629 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node21632 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node21635 = (inp[7]) ? node21641 : node21636;
														assign node21636 = (inp[8]) ? 4'b1011 : node21637;
															assign node21637 = (inp[2]) ? 4'b1010 : 4'b1010;
														assign node21641 = (inp[8]) ? 4'b1010 : node21642;
															assign node21642 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node21646 = (inp[3]) ? node21670 : node21647;
												assign node21647 = (inp[8]) ? node21659 : node21648;
													assign node21648 = (inp[7]) ? node21654 : node21649;
														assign node21649 = (inp[2]) ? 4'b1010 : node21650;
															assign node21650 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node21654 = (inp[2]) ? 4'b1011 : node21655;
															assign node21655 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node21659 = (inp[7]) ? node21665 : node21660;
														assign node21660 = (inp[14]) ? 4'b1011 : node21661;
															assign node21661 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node21665 = (inp[2]) ? 4'b1010 : node21666;
															assign node21666 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node21670 = (inp[5]) ? node21686 : node21671;
													assign node21671 = (inp[7]) ? node21679 : node21672;
														assign node21672 = (inp[8]) ? node21676 : node21673;
															assign node21673 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node21676 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node21679 = (inp[8]) ? node21683 : node21680;
															assign node21680 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node21683 = (inp[2]) ? 4'b1010 : 4'b1010;
													assign node21686 = (inp[2]) ? node21692 : node21687;
														assign node21687 = (inp[14]) ? node21689 : 4'b1001;
															assign node21689 = (inp[7]) ? 4'b1000 : 4'b1000;
														assign node21692 = (inp[7]) ? node21696 : node21693;
															assign node21693 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node21696 = (inp[8]) ? 4'b1000 : 4'b1001;
									assign node21699 = (inp[8]) ? node21813 : node21700;
										assign node21700 = (inp[7]) ? node21758 : node21701;
											assign node21701 = (inp[14]) ? node21729 : node21702;
												assign node21702 = (inp[2]) ? node21718 : node21703;
													assign node21703 = (inp[5]) ? node21711 : node21704;
														assign node21704 = (inp[0]) ? node21708 : node21705;
															assign node21705 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node21708 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node21711 = (inp[15]) ? node21715 : node21712;
															assign node21712 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node21715 = (inp[3]) ? 4'b1001 : 4'b1001;
													assign node21718 = (inp[0]) ? node21724 : node21719;
														assign node21719 = (inp[5]) ? node21721 : 4'b1000;
															assign node21721 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node21724 = (inp[3]) ? node21726 : 4'b1010;
															assign node21726 = (inp[5]) ? 4'b1000 : 4'b1000;
												assign node21729 = (inp[5]) ? node21743 : node21730;
													assign node21730 = (inp[3]) ? node21738 : node21731;
														assign node21731 = (inp[15]) ? node21735 : node21732;
															assign node21732 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node21735 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node21738 = (inp[2]) ? 4'b1000 : node21739;
															assign node21739 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node21743 = (inp[0]) ? node21751 : node21744;
														assign node21744 = (inp[3]) ? node21748 : node21745;
															assign node21745 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node21748 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node21751 = (inp[2]) ? node21755 : node21752;
															assign node21752 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node21755 = (inp[15]) ? 4'b1000 : 4'b1000;
											assign node21758 = (inp[2]) ? node21790 : node21759;
												assign node21759 = (inp[14]) ? node21775 : node21760;
													assign node21760 = (inp[5]) ? node21768 : node21761;
														assign node21761 = (inp[15]) ? node21765 : node21762;
															assign node21762 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node21765 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node21768 = (inp[3]) ? node21772 : node21769;
															assign node21769 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node21772 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node21775 = (inp[5]) ? node21783 : node21776;
														assign node21776 = (inp[0]) ? node21780 : node21777;
															assign node21777 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node21780 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node21783 = (inp[15]) ? node21787 : node21784;
															assign node21784 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node21787 = (inp[3]) ? 4'b0001 : 4'b0001;
												assign node21790 = (inp[15]) ? node21802 : node21791;
													assign node21791 = (inp[0]) ? node21797 : node21792;
														assign node21792 = (inp[3]) ? node21794 : 4'b0011;
															assign node21794 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node21797 = (inp[5]) ? node21799 : 4'b0001;
															assign node21799 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node21802 = (inp[0]) ? node21808 : node21803;
														assign node21803 = (inp[3]) ? node21805 : 4'b0001;
															assign node21805 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node21808 = (inp[5]) ? node21810 : 4'b0011;
															assign node21810 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node21813 = (inp[7]) ? node21875 : node21814;
											assign node21814 = (inp[2]) ? node21844 : node21815;
												assign node21815 = (inp[14]) ? node21831 : node21816;
													assign node21816 = (inp[5]) ? node21824 : node21817;
														assign node21817 = (inp[0]) ? node21821 : node21818;
															assign node21818 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node21821 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node21824 = (inp[3]) ? node21828 : node21825;
															assign node21825 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node21828 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node21831 = (inp[15]) ? node21839 : node21832;
														assign node21832 = (inp[0]) ? node21836 : node21833;
															assign node21833 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node21836 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node21839 = (inp[0]) ? node21841 : 4'b0001;
															assign node21841 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node21844 = (inp[14]) ? node21860 : node21845;
													assign node21845 = (inp[5]) ? node21853 : node21846;
														assign node21846 = (inp[3]) ? node21850 : node21847;
															assign node21847 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node21850 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node21853 = (inp[15]) ? node21857 : node21854;
															assign node21854 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node21857 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node21860 = (inp[3]) ? node21868 : node21861;
														assign node21861 = (inp[15]) ? node21865 : node21862;
															assign node21862 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node21865 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node21868 = (inp[5]) ? node21872 : node21869;
															assign node21869 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node21872 = (inp[15]) ? 4'b0001 : 4'b0001;
											assign node21875 = (inp[2]) ? node21905 : node21876;
												assign node21876 = (inp[14]) ? node21892 : node21877;
													assign node21877 = (inp[3]) ? node21885 : node21878;
														assign node21878 = (inp[0]) ? node21882 : node21879;
															assign node21879 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node21882 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node21885 = (inp[15]) ? node21889 : node21886;
															assign node21886 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node21889 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node21892 = (inp[3]) ? node21900 : node21893;
														assign node21893 = (inp[15]) ? node21897 : node21894;
															assign node21894 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node21897 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node21900 = (inp[0]) ? 4'b0010 : node21901;
															assign node21901 = (inp[5]) ? 4'b0000 : 4'b0000;
												assign node21905 = (inp[15]) ? node21917 : node21906;
													assign node21906 = (inp[0]) ? node21912 : node21907;
														assign node21907 = (inp[3]) ? node21909 : 4'b0010;
															assign node21909 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node21912 = (inp[3]) ? node21914 : 4'b0000;
															assign node21914 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node21917 = (inp[0]) ? node21923 : node21918;
														assign node21918 = (inp[3]) ? node21920 : 4'b0000;
															assign node21920 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node21923 = (inp[3]) ? node21925 : 4'b0010;
															assign node21925 = (inp[5]) ? 4'b0000 : 4'b0010;
								assign node21928 = (inp[1]) ? node22148 : node21929;
									assign node21929 = (inp[7]) ? node22035 : node21930;
										assign node21930 = (inp[8]) ? node21984 : node21931;
											assign node21931 = (inp[14]) ? node21961 : node21932;
												assign node21932 = (inp[2]) ? node21948 : node21933;
													assign node21933 = (inp[5]) ? node21941 : node21934;
														assign node21934 = (inp[0]) ? node21938 : node21935;
															assign node21935 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node21938 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node21941 = (inp[15]) ? node21945 : node21942;
															assign node21942 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node21945 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node21948 = (inp[0]) ? node21956 : node21949;
														assign node21949 = (inp[15]) ? node21953 : node21950;
															assign node21950 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node21953 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node21956 = (inp[3]) ? node21958 : 4'b1010;
															assign node21958 = (inp[5]) ? 4'b1000 : 4'b1000;
												assign node21961 = (inp[0]) ? node21973 : node21962;
													assign node21962 = (inp[15]) ? node21968 : node21963;
														assign node21963 = (inp[5]) ? node21965 : 4'b1010;
															assign node21965 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node21968 = (inp[5]) ? node21970 : 4'b1000;
															assign node21970 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node21973 = (inp[15]) ? node21979 : node21974;
														assign node21974 = (inp[5]) ? node21976 : 4'b1000;
															assign node21976 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node21979 = (inp[5]) ? node21981 : 4'b1010;
															assign node21981 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node21984 = (inp[2]) ? node22014 : node21985;
												assign node21985 = (inp[14]) ? node21999 : node21986;
													assign node21986 = (inp[3]) ? node21992 : node21987;
														assign node21987 = (inp[5]) ? 4'b1000 : node21988;
															assign node21988 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node21992 = (inp[5]) ? node21996 : node21993;
															assign node21993 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node21996 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node21999 = (inp[5]) ? node22007 : node22000;
														assign node22000 = (inp[15]) ? node22004 : node22001;
															assign node22001 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node22004 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node22007 = (inp[0]) ? node22011 : node22008;
															assign node22008 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node22011 = (inp[3]) ? 4'b0001 : 4'b0001;
												assign node22014 = (inp[0]) ? node22026 : node22015;
													assign node22015 = (inp[15]) ? node22021 : node22016;
														assign node22016 = (inp[5]) ? node22018 : 4'b0011;
															assign node22018 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node22021 = (inp[5]) ? node22023 : 4'b0001;
															assign node22023 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node22026 = (inp[15]) ? node22032 : node22027;
														assign node22027 = (inp[5]) ? node22029 : 4'b0001;
															assign node22029 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node22032 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node22035 = (inp[8]) ? node22093 : node22036;
											assign node22036 = (inp[14]) ? node22064 : node22037;
												assign node22037 = (inp[2]) ? node22053 : node22038;
													assign node22038 = (inp[15]) ? node22046 : node22039;
														assign node22039 = (inp[0]) ? node22043 : node22040;
															assign node22040 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node22043 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node22046 = (inp[3]) ? node22050 : node22047;
															assign node22047 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node22050 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node22053 = (inp[15]) ? node22059 : node22054;
														assign node22054 = (inp[0]) ? 4'b0001 : node22055;
															assign node22055 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node22059 = (inp[3]) ? node22061 : 4'b0011;
															assign node22061 = (inp[0]) ? 4'b0001 : 4'b0001;
												assign node22064 = (inp[2]) ? node22078 : node22065;
													assign node22065 = (inp[3]) ? node22073 : node22066;
														assign node22066 = (inp[5]) ? node22070 : node22067;
															assign node22067 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node22070 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node22073 = (inp[0]) ? node22075 : 4'b0011;
															assign node22075 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node22078 = (inp[5]) ? node22086 : node22079;
														assign node22079 = (inp[15]) ? node22083 : node22080;
															assign node22080 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node22083 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node22086 = (inp[15]) ? node22090 : node22087;
															assign node22087 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node22090 = (inp[3]) ? 4'b0001 : 4'b0001;
											assign node22093 = (inp[2]) ? node22125 : node22094;
												assign node22094 = (inp[14]) ? node22110 : node22095;
													assign node22095 = (inp[3]) ? node22103 : node22096;
														assign node22096 = (inp[15]) ? node22100 : node22097;
															assign node22097 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node22100 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node22103 = (inp[15]) ? node22107 : node22104;
															assign node22104 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node22107 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node22110 = (inp[15]) ? node22118 : node22111;
														assign node22111 = (inp[0]) ? node22115 : node22112;
															assign node22112 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node22115 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node22118 = (inp[0]) ? node22122 : node22119;
															assign node22119 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node22122 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node22125 = (inp[0]) ? node22137 : node22126;
													assign node22126 = (inp[15]) ? node22132 : node22127;
														assign node22127 = (inp[5]) ? node22129 : 4'b0010;
															assign node22129 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node22132 = (inp[5]) ? node22134 : 4'b0000;
															assign node22134 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node22137 = (inp[15]) ? node22143 : node22138;
														assign node22138 = (inp[3]) ? node22140 : 4'b0000;
															assign node22140 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node22143 = (inp[3]) ? node22145 : 4'b0010;
															assign node22145 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node22148 = (inp[7]) ? node22254 : node22149;
										assign node22149 = (inp[8]) ? node22203 : node22150;
											assign node22150 = (inp[14]) ? node22180 : node22151;
												assign node22151 = (inp[2]) ? node22167 : node22152;
													assign node22152 = (inp[3]) ? node22160 : node22153;
														assign node22153 = (inp[0]) ? node22157 : node22154;
															assign node22154 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node22157 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node22160 = (inp[5]) ? node22164 : node22161;
															assign node22161 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node22164 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node22167 = (inp[0]) ? node22173 : node22168;
														assign node22168 = (inp[15]) ? node22170 : 4'b0010;
															assign node22170 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node22173 = (inp[15]) ? node22177 : node22174;
															assign node22174 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node22177 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node22180 = (inp[0]) ? node22192 : node22181;
													assign node22181 = (inp[15]) ? node22187 : node22182;
														assign node22182 = (inp[5]) ? node22184 : 4'b0010;
															assign node22184 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node22187 = (inp[5]) ? node22189 : 4'b0000;
															assign node22189 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node22192 = (inp[15]) ? node22198 : node22193;
														assign node22193 = (inp[5]) ? node22195 : 4'b0000;
															assign node22195 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node22198 = (inp[5]) ? node22200 : 4'b0010;
															assign node22200 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node22203 = (inp[2]) ? node22231 : node22204;
												assign node22204 = (inp[14]) ? node22218 : node22205;
													assign node22205 = (inp[3]) ? node22211 : node22206;
														assign node22206 = (inp[5]) ? node22208 : 4'b0010;
															assign node22208 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node22211 = (inp[5]) ? node22215 : node22212;
															assign node22212 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node22215 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node22218 = (inp[0]) ? node22224 : node22219;
														assign node22219 = (inp[3]) ? node22221 : 4'b0011;
															assign node22221 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node22224 = (inp[15]) ? node22228 : node22225;
															assign node22225 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node22228 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node22231 = (inp[15]) ? node22243 : node22232;
													assign node22232 = (inp[0]) ? node22238 : node22233;
														assign node22233 = (inp[3]) ? node22235 : 4'b0011;
															assign node22235 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node22238 = (inp[3]) ? node22240 : 4'b0001;
															assign node22240 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node22243 = (inp[0]) ? node22249 : node22244;
														assign node22244 = (inp[5]) ? node22246 : 4'b0001;
															assign node22246 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node22249 = (inp[3]) ? node22251 : 4'b0011;
															assign node22251 = (inp[14]) ? 4'b0011 : 4'b0001;
										assign node22254 = (inp[8]) ? node22304 : node22255;
											assign node22255 = (inp[2]) ? node22281 : node22256;
												assign node22256 = (inp[14]) ? node22270 : node22257;
													assign node22257 = (inp[15]) ? node22265 : node22258;
														assign node22258 = (inp[0]) ? node22262 : node22259;
															assign node22259 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node22262 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node22265 = (inp[0]) ? node22267 : 4'b0000;
															assign node22267 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node22270 = (inp[15]) ? node22276 : node22271;
														assign node22271 = (inp[0]) ? 4'b0001 : node22272;
															assign node22272 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node22276 = (inp[0]) ? 4'b0011 : node22277;
															assign node22277 = (inp[3]) ? 4'b0001 : 4'b0001;
												assign node22281 = (inp[0]) ? node22293 : node22282;
													assign node22282 = (inp[15]) ? node22288 : node22283;
														assign node22283 = (inp[3]) ? node22285 : 4'b0011;
															assign node22285 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node22288 = (inp[5]) ? node22290 : 4'b0001;
															assign node22290 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node22293 = (inp[15]) ? node22299 : node22294;
														assign node22294 = (inp[3]) ? node22296 : 4'b0001;
															assign node22296 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node22299 = (inp[3]) ? node22301 : 4'b0011;
															assign node22301 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node22304 = (inp[2]) ? node22332 : node22305;
												assign node22305 = (inp[14]) ? node22319 : node22306;
													assign node22306 = (inp[15]) ? node22312 : node22307;
														assign node22307 = (inp[0]) ? 4'b0001 : node22308;
															assign node22308 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node22312 = (inp[0]) ? node22316 : node22313;
															assign node22313 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node22316 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node22319 = (inp[0]) ? node22325 : node22320;
														assign node22320 = (inp[15]) ? 4'b0000 : node22321;
															assign node22321 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node22325 = (inp[15]) ? node22329 : node22326;
															assign node22326 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node22329 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node22332 = (inp[3]) ? node22340 : node22333;
													assign node22333 = (inp[15]) ? node22337 : node22334;
														assign node22334 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node22337 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node22340 = (inp[14]) ? node22348 : node22341;
														assign node22341 = (inp[5]) ? node22345 : node22342;
															assign node22342 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node22345 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node22348 = (inp[0]) ? node22352 : node22349;
															assign node22349 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node22352 = (inp[5]) ? 4'b0000 : 4'b0000;
							assign node22355 = (inp[1]) ? node22823 : node22356;
								assign node22356 = (inp[13]) ? node22606 : node22357;
									assign node22357 = (inp[5]) ? node22481 : node22358;
										assign node22358 = (inp[2]) ? node22420 : node22359;
											assign node22359 = (inp[15]) ? node22391 : node22360;
												assign node22360 = (inp[0]) ? node22376 : node22361;
													assign node22361 = (inp[3]) ? node22369 : node22362;
														assign node22362 = (inp[7]) ? node22366 : node22363;
															assign node22363 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node22366 = (inp[8]) ? 4'b0010 : 4'b0010;
														assign node22369 = (inp[14]) ? node22373 : node22370;
															assign node22370 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node22373 = (inp[7]) ? 4'b0010 : 4'b0010;
													assign node22376 = (inp[7]) ? node22384 : node22377;
														assign node22377 = (inp[3]) ? node22381 : node22378;
															assign node22378 = (inp[14]) ? 4'b0000 : 4'b0000;
															assign node22381 = (inp[14]) ? 4'b0000 : 4'b0000;
														assign node22384 = (inp[8]) ? node22388 : node22385;
															assign node22385 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node22388 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node22391 = (inp[0]) ? node22407 : node22392;
													assign node22392 = (inp[3]) ? node22400 : node22393;
														assign node22393 = (inp[14]) ? node22397 : node22394;
															assign node22394 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node22397 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node22400 = (inp[8]) ? node22404 : node22401;
															assign node22401 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node22404 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node22407 = (inp[8]) ? node22415 : node22408;
														assign node22408 = (inp[3]) ? node22412 : node22409;
															assign node22409 = (inp[14]) ? 4'b0010 : 4'b0010;
															assign node22412 = (inp[14]) ? 4'b0010 : 4'b0010;
														assign node22415 = (inp[7]) ? node22417 : 4'b0011;
															assign node22417 = (inp[14]) ? 4'b0010 : 4'b0011;
											assign node22420 = (inp[14]) ? node22452 : node22421;
												assign node22421 = (inp[7]) ? node22437 : node22422;
													assign node22422 = (inp[8]) ? node22430 : node22423;
														assign node22423 = (inp[0]) ? node22427 : node22424;
															assign node22424 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node22427 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node22430 = (inp[0]) ? node22434 : node22431;
															assign node22431 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node22434 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node22437 = (inp[8]) ? node22445 : node22438;
														assign node22438 = (inp[0]) ? node22442 : node22439;
															assign node22439 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node22442 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node22445 = (inp[0]) ? node22449 : node22446;
															assign node22446 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node22449 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node22452 = (inp[3]) ? node22466 : node22453;
													assign node22453 = (inp[8]) ? node22459 : node22454;
														assign node22454 = (inp[7]) ? 4'b0011 : node22455;
															assign node22455 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node22459 = (inp[7]) ? node22463 : node22460;
															assign node22460 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node22463 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node22466 = (inp[15]) ? node22474 : node22467;
														assign node22467 = (inp[0]) ? node22471 : node22468;
															assign node22468 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node22471 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node22474 = (inp[0]) ? node22478 : node22475;
															assign node22475 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node22478 = (inp[7]) ? 4'b0010 : 4'b0010;
										assign node22481 = (inp[0]) ? node22543 : node22482;
											assign node22482 = (inp[7]) ? node22514 : node22483;
												assign node22483 = (inp[8]) ? node22499 : node22484;
													assign node22484 = (inp[2]) ? node22492 : node22485;
														assign node22485 = (inp[14]) ? node22489 : node22486;
															assign node22486 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node22489 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node22492 = (inp[15]) ? node22496 : node22493;
															assign node22493 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node22496 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node22499 = (inp[2]) ? node22507 : node22500;
														assign node22500 = (inp[14]) ? node22504 : node22501;
															assign node22501 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node22504 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node22507 = (inp[14]) ? node22511 : node22508;
															assign node22508 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node22511 = (inp[15]) ? 4'b0001 : 4'b0001;
												assign node22514 = (inp[8]) ? node22530 : node22515;
													assign node22515 = (inp[14]) ? node22523 : node22516;
														assign node22516 = (inp[2]) ? node22520 : node22517;
															assign node22517 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node22520 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node22523 = (inp[3]) ? node22527 : node22524;
															assign node22524 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node22527 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node22530 = (inp[14]) ? node22538 : node22531;
														assign node22531 = (inp[2]) ? node22535 : node22532;
															assign node22532 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node22535 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node22538 = (inp[3]) ? 4'b0000 : node22539;
															assign node22539 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node22543 = (inp[8]) ? node22575 : node22544;
												assign node22544 = (inp[7]) ? node22560 : node22545;
													assign node22545 = (inp[14]) ? node22553 : node22546;
														assign node22546 = (inp[2]) ? node22550 : node22547;
															assign node22547 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node22550 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node22553 = (inp[3]) ? node22557 : node22554;
															assign node22554 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node22557 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node22560 = (inp[2]) ? node22568 : node22561;
														assign node22561 = (inp[14]) ? node22565 : node22562;
															assign node22562 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node22565 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node22568 = (inp[3]) ? node22572 : node22569;
															assign node22569 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node22572 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node22575 = (inp[7]) ? node22591 : node22576;
													assign node22576 = (inp[14]) ? node22584 : node22577;
														assign node22577 = (inp[2]) ? node22581 : node22578;
															assign node22578 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node22581 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node22584 = (inp[3]) ? node22588 : node22585;
															assign node22585 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node22588 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node22591 = (inp[14]) ? node22599 : node22592;
														assign node22592 = (inp[2]) ? node22596 : node22593;
															assign node22593 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node22596 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node22599 = (inp[15]) ? node22603 : node22600;
															assign node22600 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node22603 = (inp[3]) ? 4'b0000 : 4'b0010;
									assign node22606 = (inp[7]) ? node22718 : node22607;
										assign node22607 = (inp[8]) ? node22661 : node22608;
											assign node22608 = (inp[2]) ? node22638 : node22609;
												assign node22609 = (inp[14]) ? node22623 : node22610;
													assign node22610 = (inp[5]) ? node22618 : node22611;
														assign node22611 = (inp[0]) ? node22615 : node22612;
															assign node22612 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node22615 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node22618 = (inp[15]) ? 4'b0001 : node22619;
															assign node22619 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node22623 = (inp[5]) ? node22631 : node22624;
														assign node22624 = (inp[0]) ? node22628 : node22625;
															assign node22625 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node22628 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node22631 = (inp[3]) ? node22635 : node22632;
															assign node22632 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node22635 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node22638 = (inp[15]) ? node22650 : node22639;
													assign node22639 = (inp[0]) ? node22645 : node22640;
														assign node22640 = (inp[5]) ? node22642 : 4'b0010;
															assign node22642 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node22645 = (inp[3]) ? node22647 : 4'b0000;
															assign node22647 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node22650 = (inp[0]) ? node22656 : node22651;
														assign node22651 = (inp[3]) ? node22653 : 4'b0000;
															assign node22653 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node22656 = (inp[5]) ? node22658 : 4'b0010;
															assign node22658 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node22661 = (inp[14]) ? node22689 : node22662;
												assign node22662 = (inp[2]) ? node22678 : node22663;
													assign node22663 = (inp[0]) ? node22671 : node22664;
														assign node22664 = (inp[15]) ? node22668 : node22665;
															assign node22665 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node22668 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node22671 = (inp[15]) ? node22675 : node22672;
															assign node22672 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node22675 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node22678 = (inp[5]) ? node22684 : node22679;
														assign node22679 = (inp[3]) ? 4'b1101 : node22680;
															assign node22680 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node22684 = (inp[0]) ? node22686 : 4'b1111;
															assign node22686 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node22689 = (inp[2]) ? node22703 : node22690;
													assign node22690 = (inp[3]) ? node22698 : node22691;
														assign node22691 = (inp[15]) ? node22695 : node22692;
															assign node22692 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node22695 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node22698 = (inp[15]) ? 4'b1111 : node22699;
															assign node22699 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node22703 = (inp[3]) ? node22711 : node22704;
														assign node22704 = (inp[5]) ? node22708 : node22705;
															assign node22705 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node22708 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node22711 = (inp[5]) ? node22715 : node22712;
															assign node22712 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node22715 = (inp[15]) ? 4'b1101 : 4'b1101;
										assign node22718 = (inp[8]) ? node22772 : node22719;
											assign node22719 = (inp[14]) ? node22749 : node22720;
												assign node22720 = (inp[2]) ? node22736 : node22721;
													assign node22721 = (inp[0]) ? node22729 : node22722;
														assign node22722 = (inp[15]) ? node22726 : node22723;
															assign node22723 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node22726 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node22729 = (inp[15]) ? node22733 : node22730;
															assign node22730 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node22733 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node22736 = (inp[3]) ? node22744 : node22737;
														assign node22737 = (inp[15]) ? node22741 : node22738;
															assign node22738 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node22741 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node22744 = (inp[5]) ? node22746 : 4'b1111;
															assign node22746 = (inp[15]) ? 4'b1101 : 4'b1101;
												assign node22749 = (inp[5]) ? node22765 : node22750;
													assign node22750 = (inp[15]) ? node22758 : node22751;
														assign node22751 = (inp[0]) ? node22755 : node22752;
															assign node22752 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node22755 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node22758 = (inp[0]) ? node22762 : node22759;
															assign node22759 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node22762 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node22765 = (inp[0]) ? node22769 : node22766;
														assign node22766 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node22769 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node22772 = (inp[14]) ? node22800 : node22773;
												assign node22773 = (inp[2]) ? node22789 : node22774;
													assign node22774 = (inp[15]) ? node22782 : node22775;
														assign node22775 = (inp[0]) ? node22779 : node22776;
															assign node22776 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node22779 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node22782 = (inp[0]) ? node22786 : node22783;
															assign node22783 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node22786 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node22789 = (inp[5]) ? node22795 : node22790;
														assign node22790 = (inp[0]) ? 4'b1100 : node22791;
															assign node22791 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node22795 = (inp[0]) ? node22797 : 4'b1110;
															assign node22797 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node22800 = (inp[5]) ? node22816 : node22801;
													assign node22801 = (inp[15]) ? node22809 : node22802;
														assign node22802 = (inp[0]) ? node22806 : node22803;
															assign node22803 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node22806 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node22809 = (inp[0]) ? node22813 : node22810;
															assign node22810 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node22813 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node22816 = (inp[0]) ? node22820 : node22817;
														assign node22817 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node22820 = (inp[15]) ? 4'b1100 : 4'b1110;
								assign node22823 = (inp[13]) ? node23037 : node22824;
									assign node22824 = (inp[8]) ? node22930 : node22825;
										assign node22825 = (inp[7]) ? node22879 : node22826;
											assign node22826 = (inp[14]) ? node22858 : node22827;
												assign node22827 = (inp[2]) ? node22843 : node22828;
													assign node22828 = (inp[5]) ? node22836 : node22829;
														assign node22829 = (inp[3]) ? node22833 : node22830;
															assign node22830 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node22833 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node22836 = (inp[0]) ? node22840 : node22837;
															assign node22837 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node22840 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node22843 = (inp[3]) ? node22851 : node22844;
														assign node22844 = (inp[0]) ? node22848 : node22845;
															assign node22845 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node22848 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node22851 = (inp[5]) ? node22855 : node22852;
															assign node22852 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node22855 = (inp[0]) ? 4'b0000 : 4'b0000;
												assign node22858 = (inp[0]) ? node22868 : node22859;
													assign node22859 = (inp[15]) ? node22865 : node22860;
														assign node22860 = (inp[5]) ? node22862 : 4'b0010;
															assign node22862 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node22865 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node22868 = (inp[15]) ? node22874 : node22869;
														assign node22869 = (inp[3]) ? node22871 : 4'b0000;
															assign node22871 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node22874 = (inp[5]) ? node22876 : 4'b0010;
															assign node22876 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node22879 = (inp[2]) ? node22909 : node22880;
												assign node22880 = (inp[14]) ? node22896 : node22881;
													assign node22881 = (inp[5]) ? node22889 : node22882;
														assign node22882 = (inp[3]) ? node22886 : node22883;
															assign node22883 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node22886 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node22889 = (inp[0]) ? node22893 : node22890;
															assign node22890 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node22893 = (inp[3]) ? 4'b0000 : 4'b0000;
													assign node22896 = (inp[15]) ? node22902 : node22897;
														assign node22897 = (inp[0]) ? 4'b1111 : node22898;
															assign node22898 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node22902 = (inp[0]) ? node22906 : node22903;
															assign node22903 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node22906 = (inp[5]) ? 4'b1101 : 4'b1101;
												assign node22909 = (inp[0]) ? node22919 : node22910;
													assign node22910 = (inp[15]) ? node22916 : node22911;
														assign node22911 = (inp[3]) ? 4'b1101 : node22912;
															assign node22912 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node22916 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node22919 = (inp[15]) ? node22925 : node22920;
														assign node22920 = (inp[3]) ? 4'b1111 : node22921;
															assign node22921 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node22925 = (inp[3]) ? 4'b1101 : node22926;
															assign node22926 = (inp[5]) ? 4'b1101 : 4'b1111;
										assign node22930 = (inp[7]) ? node22990 : node22931;
											assign node22931 = (inp[2]) ? node22961 : node22932;
												assign node22932 = (inp[14]) ? node22948 : node22933;
													assign node22933 = (inp[3]) ? node22941 : node22934;
														assign node22934 = (inp[0]) ? node22938 : node22935;
															assign node22935 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node22938 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node22941 = (inp[5]) ? node22945 : node22942;
															assign node22942 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node22945 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node22948 = (inp[0]) ? node22954 : node22949;
														assign node22949 = (inp[3]) ? 4'b1111 : node22950;
															assign node22950 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node22954 = (inp[15]) ? node22958 : node22955;
															assign node22955 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node22958 = (inp[5]) ? 4'b1101 : 4'b1101;
												assign node22961 = (inp[14]) ? node22977 : node22962;
													assign node22962 = (inp[0]) ? node22970 : node22963;
														assign node22963 = (inp[15]) ? node22967 : node22964;
															assign node22964 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node22967 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node22970 = (inp[15]) ? node22974 : node22971;
															assign node22971 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node22974 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node22977 = (inp[5]) ? node22983 : node22978;
														assign node22978 = (inp[15]) ? node22980 : 4'b1111;
															assign node22980 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node22983 = (inp[0]) ? node22987 : node22984;
															assign node22984 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node22987 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node22990 = (inp[2]) ? node23014 : node22991;
												assign node22991 = (inp[14]) ? node23005 : node22992;
													assign node22992 = (inp[0]) ? node23000 : node22993;
														assign node22993 = (inp[15]) ? node22997 : node22994;
															assign node22994 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node22997 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node23000 = (inp[15]) ? 4'b1101 : node23001;
															assign node23001 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node23005 = (inp[0]) ? 4'b1110 : node23006;
														assign node23006 = (inp[15]) ? node23010 : node23007;
															assign node23007 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node23010 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node23014 = (inp[0]) ? node23026 : node23015;
													assign node23015 = (inp[15]) ? node23021 : node23016;
														assign node23016 = (inp[5]) ? 4'b1100 : node23017;
															assign node23017 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node23021 = (inp[5]) ? 4'b1110 : node23022;
															assign node23022 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node23026 = (inp[15]) ? node23032 : node23027;
														assign node23027 = (inp[3]) ? 4'b1110 : node23028;
															assign node23028 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node23032 = (inp[5]) ? 4'b1100 : node23033;
															assign node23033 = (inp[3]) ? 4'b1100 : 4'b1110;
									assign node23037 = (inp[14]) ? node23163 : node23038;
										assign node23038 = (inp[3]) ? node23102 : node23039;
											assign node23039 = (inp[8]) ? node23071 : node23040;
												assign node23040 = (inp[0]) ? node23056 : node23041;
													assign node23041 = (inp[7]) ? node23049 : node23042;
														assign node23042 = (inp[2]) ? node23046 : node23043;
															assign node23043 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node23046 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node23049 = (inp[2]) ? node23053 : node23050;
															assign node23050 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node23053 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node23056 = (inp[15]) ? node23064 : node23057;
														assign node23057 = (inp[5]) ? node23061 : node23058;
															assign node23058 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node23061 = (inp[7]) ? 4'b1110 : 4'b1110;
														assign node23064 = (inp[5]) ? node23068 : node23065;
															assign node23065 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node23068 = (inp[7]) ? 4'b1100 : 4'b1100;
												assign node23071 = (inp[2]) ? node23087 : node23072;
													assign node23072 = (inp[7]) ? node23080 : node23073;
														assign node23073 = (inp[15]) ? node23077 : node23074;
															assign node23074 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node23077 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node23080 = (inp[0]) ? node23084 : node23081;
															assign node23081 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node23084 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node23087 = (inp[7]) ? node23095 : node23088;
														assign node23088 = (inp[0]) ? node23092 : node23089;
															assign node23089 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node23092 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node23095 = (inp[15]) ? node23099 : node23096;
															assign node23096 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node23099 = (inp[0]) ? 4'b1100 : 4'b1100;
											assign node23102 = (inp[5]) ? node23132 : node23103;
												assign node23103 = (inp[0]) ? node23117 : node23104;
													assign node23104 = (inp[15]) ? node23110 : node23105;
														assign node23105 = (inp[7]) ? 4'b1101 : node23106;
															assign node23106 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node23110 = (inp[2]) ? node23114 : node23111;
															assign node23111 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node23114 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node23117 = (inp[15]) ? node23125 : node23118;
														assign node23118 = (inp[7]) ? node23122 : node23119;
															assign node23119 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node23122 = (inp[2]) ? 4'b1110 : 4'b1110;
														assign node23125 = (inp[8]) ? node23129 : node23126;
															assign node23126 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node23129 = (inp[2]) ? 4'b1100 : 4'b1100;
												assign node23132 = (inp[7]) ? node23148 : node23133;
													assign node23133 = (inp[0]) ? node23141 : node23134;
														assign node23134 = (inp[15]) ? node23138 : node23135;
															assign node23135 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node23138 = (inp[2]) ? 4'b1110 : 4'b1110;
														assign node23141 = (inp[15]) ? node23145 : node23142;
															assign node23142 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node23145 = (inp[8]) ? 4'b1100 : 4'b1100;
													assign node23148 = (inp[8]) ? node23156 : node23149;
														assign node23149 = (inp[2]) ? node23153 : node23150;
															assign node23150 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node23153 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node23156 = (inp[2]) ? node23160 : node23157;
															assign node23157 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node23160 = (inp[15]) ? 4'b1100 : 4'b1100;
										assign node23163 = (inp[2]) ? node23221 : node23164;
											assign node23164 = (inp[8]) ? node23194 : node23165;
												assign node23165 = (inp[7]) ? node23179 : node23166;
													assign node23166 = (inp[15]) ? node23174 : node23167;
														assign node23167 = (inp[0]) ? node23171 : node23168;
															assign node23168 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node23171 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node23174 = (inp[0]) ? 4'b1100 : node23175;
															assign node23175 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node23179 = (inp[5]) ? node23187 : node23180;
														assign node23180 = (inp[0]) ? node23184 : node23181;
															assign node23181 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node23184 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node23187 = (inp[3]) ? node23191 : node23188;
															assign node23188 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node23191 = (inp[15]) ? 4'b1101 : 4'b1101;
												assign node23194 = (inp[7]) ? node23206 : node23195;
													assign node23195 = (inp[0]) ? node23203 : node23196;
														assign node23196 = (inp[15]) ? node23200 : node23197;
															assign node23197 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node23200 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node23203 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node23206 = (inp[5]) ? node23214 : node23207;
														assign node23207 = (inp[15]) ? node23211 : node23208;
															assign node23208 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node23211 = (inp[3]) ? 4'b1100 : 4'b1100;
														assign node23214 = (inp[3]) ? node23218 : node23215;
															assign node23215 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node23218 = (inp[0]) ? 4'b1100 : 4'b1100;
											assign node23221 = (inp[3]) ? node23251 : node23222;
												assign node23222 = (inp[5]) ? node23238 : node23223;
													assign node23223 = (inp[0]) ? node23231 : node23224;
														assign node23224 = (inp[15]) ? node23228 : node23225;
															assign node23225 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node23228 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node23231 = (inp[15]) ? node23235 : node23232;
															assign node23232 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node23235 = (inp[7]) ? 4'b1110 : 4'b1110;
													assign node23238 = (inp[15]) ? node23244 : node23239;
														assign node23239 = (inp[0]) ? node23241 : 4'b1101;
															assign node23241 = (inp[7]) ? 4'b1110 : 4'b1110;
														assign node23244 = (inp[0]) ? node23248 : node23245;
															assign node23245 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node23248 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node23251 = (inp[5]) ? node23267 : node23252;
													assign node23252 = (inp[15]) ? node23260 : node23253;
														assign node23253 = (inp[0]) ? node23257 : node23254;
															assign node23254 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node23257 = (inp[7]) ? 4'b1110 : 4'b1110;
														assign node23260 = (inp[0]) ? node23264 : node23261;
															assign node23261 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node23264 = (inp[7]) ? 4'b1100 : 4'b1100;
													assign node23267 = (inp[7]) ? node23273 : node23268;
														assign node23268 = (inp[8]) ? 4'b1101 : node23269;
															assign node23269 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node23273 = (inp[8]) ? node23275 : 4'b1111;
															assign node23275 = (inp[15]) ? 4'b1110 : 4'b1100;
						assign node23278 = (inp[11]) ? node24192 : node23279;
							assign node23279 = (inp[1]) ? node23717 : node23280;
								assign node23280 = (inp[13]) ? node23498 : node23281;
									assign node23281 = (inp[15]) ? node23389 : node23282;
										assign node23282 = (inp[0]) ? node23336 : node23283;
											assign node23283 = (inp[5]) ? node23307 : node23284;
												assign node23284 = (inp[7]) ? node23296 : node23285;
													assign node23285 = (inp[8]) ? node23291 : node23286;
														assign node23286 = (inp[2]) ? 4'b0010 : node23287;
															assign node23287 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node23291 = (inp[2]) ? 4'b0011 : node23292;
															assign node23292 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node23296 = (inp[8]) ? node23302 : node23297;
														assign node23297 = (inp[14]) ? 4'b0011 : node23298;
															assign node23298 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node23302 = (inp[2]) ? 4'b0010 : node23303;
															assign node23303 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node23307 = (inp[3]) ? node23321 : node23308;
													assign node23308 = (inp[2]) ? node23314 : node23309;
														assign node23309 = (inp[7]) ? node23311 : 4'b0011;
															assign node23311 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node23314 = (inp[14]) ? node23318 : node23315;
															assign node23315 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node23318 = (inp[8]) ? 4'b0010 : 4'b0010;
													assign node23321 = (inp[7]) ? node23329 : node23322;
														assign node23322 = (inp[8]) ? node23326 : node23323;
															assign node23323 = (inp[14]) ? 4'b0000 : 4'b0000;
															assign node23326 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node23329 = (inp[8]) ? node23333 : node23330;
															assign node23330 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node23333 = (inp[14]) ? 4'b0000 : 4'b0000;
											assign node23336 = (inp[3]) ? node23360 : node23337;
												assign node23337 = (inp[14]) ? node23353 : node23338;
													assign node23338 = (inp[2]) ? node23346 : node23339;
														assign node23339 = (inp[5]) ? node23343 : node23340;
															assign node23340 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node23343 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node23346 = (inp[8]) ? node23350 : node23347;
															assign node23347 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node23350 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node23353 = (inp[7]) ? node23357 : node23354;
														assign node23354 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node23357 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node23360 = (inp[5]) ? node23374 : node23361;
													assign node23361 = (inp[8]) ? node23369 : node23362;
														assign node23362 = (inp[7]) ? node23366 : node23363;
															assign node23363 = (inp[2]) ? 4'b0000 : 4'b0000;
															assign node23366 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node23369 = (inp[7]) ? 4'b0000 : node23370;
															assign node23370 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node23374 = (inp[2]) ? node23382 : node23375;
														assign node23375 = (inp[8]) ? node23379 : node23376;
															assign node23376 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node23379 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node23382 = (inp[14]) ? node23386 : node23383;
															assign node23383 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node23386 = (inp[8]) ? 4'b0010 : 4'b0010;
										assign node23389 = (inp[0]) ? node23449 : node23390;
											assign node23390 = (inp[5]) ? node23422 : node23391;
												assign node23391 = (inp[3]) ? node23407 : node23392;
													assign node23392 = (inp[14]) ? node23400 : node23393;
														assign node23393 = (inp[8]) ? node23397 : node23394;
															assign node23394 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node23397 = (inp[2]) ? 4'b0000 : 4'b0000;
														assign node23400 = (inp[2]) ? node23404 : node23401;
															assign node23401 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node23404 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node23407 = (inp[8]) ? node23415 : node23408;
														assign node23408 = (inp[7]) ? node23412 : node23409;
															assign node23409 = (inp[2]) ? 4'b0000 : 4'b0000;
															assign node23412 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node23415 = (inp[7]) ? node23419 : node23416;
															assign node23416 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node23419 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node23422 = (inp[3]) ? node23436 : node23423;
													assign node23423 = (inp[7]) ? node23429 : node23424;
														assign node23424 = (inp[8]) ? node23426 : 4'b0000;
															assign node23426 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node23429 = (inp[8]) ? node23433 : node23430;
															assign node23430 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node23433 = (inp[2]) ? 4'b0000 : 4'b0000;
													assign node23436 = (inp[2]) ? node23444 : node23437;
														assign node23437 = (inp[7]) ? node23441 : node23438;
															assign node23438 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node23441 = (inp[8]) ? 4'b0010 : 4'b0010;
														assign node23444 = (inp[8]) ? node23446 : 4'b0010;
															assign node23446 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node23449 = (inp[3]) ? node23471 : node23450;
												assign node23450 = (inp[8]) ? node23462 : node23451;
													assign node23451 = (inp[7]) ? node23457 : node23452;
														assign node23452 = (inp[2]) ? 4'b0010 : node23453;
															assign node23453 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node23457 = (inp[14]) ? 4'b0011 : node23458;
															assign node23458 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node23462 = (inp[7]) ? node23466 : node23463;
														assign node23463 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node23466 = (inp[14]) ? 4'b0010 : node23467;
															assign node23467 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node23471 = (inp[5]) ? node23485 : node23472;
													assign node23472 = (inp[8]) ? node23478 : node23473;
														assign node23473 = (inp[7]) ? node23475 : 4'b0010;
															assign node23475 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node23478 = (inp[7]) ? node23482 : node23479;
															assign node23479 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node23482 = (inp[14]) ? 4'b0010 : 4'b0010;
													assign node23485 = (inp[2]) ? node23493 : node23486;
														assign node23486 = (inp[7]) ? node23490 : node23487;
															assign node23487 = (inp[14]) ? 4'b0000 : 4'b0000;
															assign node23490 = (inp[8]) ? 4'b0000 : 4'b0000;
														assign node23493 = (inp[14]) ? node23495 : 4'b0000;
															assign node23495 = (inp[7]) ? 4'b0000 : 4'b0000;
									assign node23498 = (inp[8]) ? node23614 : node23499;
										assign node23499 = (inp[7]) ? node23553 : node23500;
											assign node23500 = (inp[2]) ? node23530 : node23501;
												assign node23501 = (inp[14]) ? node23515 : node23502;
													assign node23502 = (inp[15]) ? node23510 : node23503;
														assign node23503 = (inp[0]) ? node23507 : node23504;
															assign node23504 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node23507 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node23510 = (inp[5]) ? node23512 : 4'b0011;
															assign node23512 = (inp[3]) ? 4'b0001 : 4'b0001;
													assign node23515 = (inp[3]) ? node23523 : node23516;
														assign node23516 = (inp[15]) ? node23520 : node23517;
															assign node23517 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node23520 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node23523 = (inp[5]) ? node23527 : node23524;
															assign node23524 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node23527 = (inp[0]) ? 4'b0000 : 4'b0000;
												assign node23530 = (inp[3]) ? node23538 : node23531;
													assign node23531 = (inp[0]) ? node23535 : node23532;
														assign node23532 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node23535 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node23538 = (inp[0]) ? node23546 : node23539;
														assign node23539 = (inp[15]) ? node23543 : node23540;
															assign node23540 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node23543 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node23546 = (inp[5]) ? node23550 : node23547;
															assign node23547 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node23550 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node23553 = (inp[2]) ? node23583 : node23554;
												assign node23554 = (inp[14]) ? node23570 : node23555;
													assign node23555 = (inp[3]) ? node23563 : node23556;
														assign node23556 = (inp[15]) ? node23560 : node23557;
															assign node23557 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node23560 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node23563 = (inp[15]) ? node23567 : node23564;
															assign node23564 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node23567 = (inp[5]) ? 4'b0000 : 4'b0000;
													assign node23570 = (inp[0]) ? node23578 : node23571;
														assign node23571 = (inp[15]) ? node23575 : node23572;
															assign node23572 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node23575 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node23578 = (inp[15]) ? 4'b1101 : node23579;
															assign node23579 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node23583 = (inp[14]) ? node23599 : node23584;
													assign node23584 = (inp[5]) ? node23592 : node23585;
														assign node23585 = (inp[3]) ? node23589 : node23586;
															assign node23586 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node23589 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node23592 = (inp[0]) ? node23596 : node23593;
															assign node23593 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node23596 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node23599 = (inp[15]) ? node23607 : node23600;
														assign node23600 = (inp[0]) ? node23604 : node23601;
															assign node23601 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node23604 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node23607 = (inp[0]) ? node23611 : node23608;
															assign node23608 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node23611 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node23614 = (inp[7]) ? node23668 : node23615;
											assign node23615 = (inp[2]) ? node23645 : node23616;
												assign node23616 = (inp[14]) ? node23630 : node23617;
													assign node23617 = (inp[0]) ? node23625 : node23618;
														assign node23618 = (inp[15]) ? node23622 : node23619;
															assign node23619 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node23622 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node23625 = (inp[15]) ? node23627 : 4'b0000;
															assign node23627 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node23630 = (inp[3]) ? node23638 : node23631;
														assign node23631 = (inp[0]) ? node23635 : node23632;
															assign node23632 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node23635 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node23638 = (inp[0]) ? node23642 : node23639;
															assign node23639 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node23642 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node23645 = (inp[3]) ? node23661 : node23646;
													assign node23646 = (inp[0]) ? node23654 : node23647;
														assign node23647 = (inp[15]) ? node23651 : node23648;
															assign node23648 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node23651 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node23654 = (inp[15]) ? node23658 : node23655;
															assign node23655 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node23658 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node23661 = (inp[15]) ? node23665 : node23662;
														assign node23662 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node23665 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node23668 = (inp[2]) ? node23694 : node23669;
												assign node23669 = (inp[14]) ? node23683 : node23670;
													assign node23670 = (inp[3]) ? node23676 : node23671;
														assign node23671 = (inp[5]) ? node23673 : 4'b1101;
															assign node23673 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node23676 = (inp[15]) ? node23680 : node23677;
															assign node23677 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node23680 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node23683 = (inp[0]) ? node23691 : node23684;
														assign node23684 = (inp[15]) ? node23688 : node23685;
															assign node23685 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node23688 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node23691 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node23694 = (inp[0]) ? node23706 : node23695;
													assign node23695 = (inp[15]) ? node23701 : node23696;
														assign node23696 = (inp[5]) ? 4'b1100 : node23697;
															assign node23697 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node23701 = (inp[3]) ? 4'b1110 : node23702;
															assign node23702 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node23706 = (inp[15]) ? node23712 : node23707;
														assign node23707 = (inp[5]) ? 4'b1110 : node23708;
															assign node23708 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node23712 = (inp[3]) ? 4'b1100 : node23713;
															assign node23713 = (inp[5]) ? 4'b1100 : 4'b1110;
								assign node23717 = (inp[13]) ? node23953 : node23718;
									assign node23718 = (inp[8]) ? node23834 : node23719;
										assign node23719 = (inp[7]) ? node23775 : node23720;
											assign node23720 = (inp[14]) ? node23746 : node23721;
												assign node23721 = (inp[2]) ? node23733 : node23722;
													assign node23722 = (inp[5]) ? node23728 : node23723;
														assign node23723 = (inp[15]) ? 4'b0011 : node23724;
															assign node23724 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node23728 = (inp[0]) ? node23730 : 4'b0001;
															assign node23730 = (inp[3]) ? 4'b0001 : 4'b0001;
													assign node23733 = (inp[0]) ? node23741 : node23734;
														assign node23734 = (inp[15]) ? node23738 : node23735;
															assign node23735 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node23738 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node23741 = (inp[15]) ? 4'b0010 : node23742;
															assign node23742 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node23746 = (inp[2]) ? node23760 : node23747;
													assign node23747 = (inp[5]) ? node23755 : node23748;
														assign node23748 = (inp[0]) ? node23752 : node23749;
															assign node23749 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node23752 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node23755 = (inp[3]) ? node23757 : 4'b0000;
															assign node23757 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node23760 = (inp[0]) ? node23768 : node23761;
														assign node23761 = (inp[15]) ? node23765 : node23762;
															assign node23762 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node23765 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node23768 = (inp[15]) ? node23772 : node23769;
															assign node23769 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node23772 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node23775 = (inp[14]) ? node23805 : node23776;
												assign node23776 = (inp[2]) ? node23792 : node23777;
													assign node23777 = (inp[15]) ? node23785 : node23778;
														assign node23778 = (inp[0]) ? node23782 : node23779;
															assign node23779 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node23782 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node23785 = (inp[0]) ? node23789 : node23786;
															assign node23786 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node23789 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node23792 = (inp[0]) ? node23798 : node23793;
														assign node23793 = (inp[5]) ? 4'b1111 : node23794;
															assign node23794 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node23798 = (inp[15]) ? node23802 : node23799;
															assign node23799 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node23802 = (inp[3]) ? 4'b1101 : 4'b1101;
												assign node23805 = (inp[2]) ? node23819 : node23806;
													assign node23806 = (inp[0]) ? node23812 : node23807;
														assign node23807 = (inp[15]) ? 4'b1111 : node23808;
															assign node23808 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node23812 = (inp[15]) ? node23816 : node23813;
															assign node23813 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node23816 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node23819 = (inp[5]) ? node23827 : node23820;
														assign node23820 = (inp[15]) ? node23824 : node23821;
															assign node23821 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node23824 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node23827 = (inp[0]) ? node23831 : node23828;
															assign node23828 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node23831 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node23834 = (inp[7]) ? node23892 : node23835;
											assign node23835 = (inp[14]) ? node23863 : node23836;
												assign node23836 = (inp[2]) ? node23850 : node23837;
													assign node23837 = (inp[15]) ? node23845 : node23838;
														assign node23838 = (inp[0]) ? node23842 : node23839;
															assign node23839 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node23842 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node23845 = (inp[0]) ? 4'b0010 : node23846;
															assign node23846 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node23850 = (inp[5]) ? node23858 : node23851;
														assign node23851 = (inp[15]) ? node23855 : node23852;
															assign node23852 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node23855 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node23858 = (inp[0]) ? 4'b1101 : node23859;
															assign node23859 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node23863 = (inp[2]) ? node23879 : node23864;
													assign node23864 = (inp[5]) ? node23872 : node23865;
														assign node23865 = (inp[3]) ? node23869 : node23866;
															assign node23866 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node23869 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node23872 = (inp[0]) ? node23876 : node23873;
															assign node23873 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node23876 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node23879 = (inp[5]) ? node23885 : node23880;
														assign node23880 = (inp[3]) ? node23882 : 4'b1111;
															assign node23882 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node23885 = (inp[3]) ? node23889 : node23886;
															assign node23886 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node23889 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node23892 = (inp[14]) ? node23922 : node23893;
												assign node23893 = (inp[2]) ? node23909 : node23894;
													assign node23894 = (inp[5]) ? node23902 : node23895;
														assign node23895 = (inp[3]) ? node23899 : node23896;
															assign node23896 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node23899 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node23902 = (inp[0]) ? node23906 : node23903;
															assign node23903 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node23906 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node23909 = (inp[5]) ? node23915 : node23910;
														assign node23910 = (inp[0]) ? 4'b1100 : node23911;
															assign node23911 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node23915 = (inp[0]) ? node23919 : node23916;
															assign node23916 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node23919 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node23922 = (inp[3]) ? node23938 : node23923;
													assign node23923 = (inp[5]) ? node23931 : node23924;
														assign node23924 = (inp[2]) ? node23928 : node23925;
															assign node23925 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node23928 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node23931 = (inp[15]) ? node23935 : node23932;
															assign node23932 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node23935 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node23938 = (inp[2]) ? node23946 : node23939;
														assign node23939 = (inp[0]) ? node23943 : node23940;
															assign node23940 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node23943 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node23946 = (inp[0]) ? node23950 : node23947;
															assign node23947 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node23950 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node23953 = (inp[5]) ? node24077 : node23954;
										assign node23954 = (inp[3]) ? node24016 : node23955;
											assign node23955 = (inp[2]) ? node23987 : node23956;
												assign node23956 = (inp[0]) ? node23972 : node23957;
													assign node23957 = (inp[15]) ? node23965 : node23958;
														assign node23958 = (inp[7]) ? node23962 : node23959;
															assign node23959 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node23962 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node23965 = (inp[14]) ? node23969 : node23966;
															assign node23966 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node23969 = (inp[7]) ? 4'b1100 : 4'b1100;
													assign node23972 = (inp[15]) ? node23980 : node23973;
														assign node23973 = (inp[14]) ? node23977 : node23974;
															assign node23974 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node23977 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node23980 = (inp[8]) ? node23984 : node23981;
															assign node23981 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node23984 = (inp[14]) ? 4'b1110 : 4'b1110;
												assign node23987 = (inp[7]) ? node24003 : node23988;
													assign node23988 = (inp[8]) ? node23996 : node23989;
														assign node23989 = (inp[14]) ? node23993 : node23990;
															assign node23990 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node23993 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node23996 = (inp[14]) ? node24000 : node23997;
															assign node23997 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node24000 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node24003 = (inp[8]) ? node24011 : node24004;
														assign node24004 = (inp[0]) ? node24008 : node24005;
															assign node24005 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node24008 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node24011 = (inp[14]) ? 4'b1100 : node24012;
															assign node24012 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node24016 = (inp[15]) ? node24046 : node24017;
												assign node24017 = (inp[0]) ? node24031 : node24018;
													assign node24018 = (inp[8]) ? node24026 : node24019;
														assign node24019 = (inp[7]) ? node24023 : node24020;
															assign node24020 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node24023 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node24026 = (inp[7]) ? 4'b1100 : node24027;
															assign node24027 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node24031 = (inp[2]) ? node24039 : node24032;
														assign node24032 = (inp[7]) ? node24036 : node24033;
															assign node24033 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node24036 = (inp[14]) ? 4'b1110 : 4'b1110;
														assign node24039 = (inp[7]) ? node24043 : node24040;
															assign node24040 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node24043 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node24046 = (inp[0]) ? node24062 : node24047;
													assign node24047 = (inp[2]) ? node24055 : node24048;
														assign node24048 = (inp[14]) ? node24052 : node24049;
															assign node24049 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node24052 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node24055 = (inp[7]) ? node24059 : node24056;
															assign node24056 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node24059 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node24062 = (inp[8]) ? node24070 : node24063;
														assign node24063 = (inp[7]) ? node24067 : node24064;
															assign node24064 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node24067 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node24070 = (inp[7]) ? node24074 : node24071;
															assign node24071 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node24074 = (inp[2]) ? 4'b1100 : 4'b1100;
										assign node24077 = (inp[8]) ? node24129 : node24078;
											assign node24078 = (inp[7]) ? node24100 : node24079;
												assign node24079 = (inp[2]) ? node24093 : node24080;
													assign node24080 = (inp[14]) ? node24088 : node24081;
														assign node24081 = (inp[3]) ? node24085 : node24082;
															assign node24082 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node24085 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node24088 = (inp[3]) ? 4'b1110 : node24089;
															assign node24089 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node24093 = (inp[15]) ? node24097 : node24094;
														assign node24094 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node24097 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node24100 = (inp[14]) ? node24114 : node24101;
													assign node24101 = (inp[2]) ? node24107 : node24102;
														assign node24102 = (inp[0]) ? 4'b1110 : node24103;
															assign node24103 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node24107 = (inp[15]) ? node24111 : node24108;
															assign node24108 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node24111 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node24114 = (inp[2]) ? node24122 : node24115;
														assign node24115 = (inp[0]) ? node24119 : node24116;
															assign node24116 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node24119 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node24122 = (inp[15]) ? node24126 : node24123;
															assign node24123 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node24126 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node24129 = (inp[7]) ? node24161 : node24130;
												assign node24130 = (inp[2]) ? node24146 : node24131;
													assign node24131 = (inp[14]) ? node24139 : node24132;
														assign node24132 = (inp[15]) ? node24136 : node24133;
															assign node24133 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node24136 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node24139 = (inp[0]) ? node24143 : node24140;
															assign node24140 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node24143 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node24146 = (inp[3]) ? node24154 : node24147;
														assign node24147 = (inp[15]) ? node24151 : node24148;
															assign node24148 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node24151 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node24154 = (inp[14]) ? node24158 : node24155;
															assign node24155 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node24158 = (inp[0]) ? 4'b1101 : 4'b1101;
												assign node24161 = (inp[14]) ? node24177 : node24162;
													assign node24162 = (inp[2]) ? node24170 : node24163;
														assign node24163 = (inp[3]) ? node24167 : node24164;
															assign node24164 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node24167 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node24170 = (inp[3]) ? node24174 : node24171;
															assign node24171 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node24174 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node24177 = (inp[3]) ? node24185 : node24178;
														assign node24178 = (inp[2]) ? node24182 : node24179;
															assign node24179 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node24182 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node24185 = (inp[0]) ? node24189 : node24186;
															assign node24186 = (inp[2]) ? 4'b1110 : 4'b1100;
															assign node24189 = (inp[15]) ? 4'b1100 : 4'b1110;
							assign node24192 = (inp[1]) ? node24644 : node24193;
								assign node24193 = (inp[13]) ? node24427 : node24194;
									assign node24194 = (inp[7]) ? node24302 : node24195;
										assign node24195 = (inp[8]) ? node24251 : node24196;
											assign node24196 = (inp[14]) ? node24228 : node24197;
												assign node24197 = (inp[2]) ? node24213 : node24198;
													assign node24198 = (inp[0]) ? node24206 : node24199;
														assign node24199 = (inp[15]) ? node24203 : node24200;
															assign node24200 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node24203 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node24206 = (inp[15]) ? node24210 : node24207;
															assign node24207 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node24210 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node24213 = (inp[15]) ? node24221 : node24214;
														assign node24214 = (inp[0]) ? node24218 : node24215;
															assign node24215 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node24218 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node24221 = (inp[0]) ? node24225 : node24222;
															assign node24222 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node24225 = (inp[3]) ? 4'b1100 : 4'b1100;
												assign node24228 = (inp[5]) ? node24244 : node24229;
													assign node24229 = (inp[3]) ? node24237 : node24230;
														assign node24230 = (inp[0]) ? node24234 : node24231;
															assign node24231 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node24234 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node24237 = (inp[15]) ? node24241 : node24238;
															assign node24238 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node24241 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node24244 = (inp[0]) ? node24248 : node24245;
														assign node24245 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node24248 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node24251 = (inp[14]) ? node24279 : node24252;
												assign node24252 = (inp[2]) ? node24266 : node24253;
													assign node24253 = (inp[15]) ? node24261 : node24254;
														assign node24254 = (inp[0]) ? node24258 : node24255;
															assign node24255 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node24258 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node24261 = (inp[0]) ? node24263 : 4'b1110;
															assign node24263 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node24266 = (inp[0]) ? node24274 : node24267;
														assign node24267 = (inp[15]) ? node24271 : node24268;
															assign node24268 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node24271 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node24274 = (inp[5]) ? 4'b1101 : node24275;
															assign node24275 = (inp[3]) ? 4'b1101 : 4'b1101;
												assign node24279 = (inp[15]) ? node24291 : node24280;
													assign node24280 = (inp[0]) ? node24286 : node24281;
														assign node24281 = (inp[3]) ? 4'b1101 : node24282;
															assign node24282 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node24286 = (inp[5]) ? 4'b1111 : node24287;
															assign node24287 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node24291 = (inp[0]) ? node24297 : node24292;
														assign node24292 = (inp[3]) ? 4'b1111 : node24293;
															assign node24293 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node24297 = (inp[3]) ? 4'b1101 : node24298;
															assign node24298 = (inp[5]) ? 4'b1101 : 4'b1111;
										assign node24302 = (inp[8]) ? node24366 : node24303;
											assign node24303 = (inp[2]) ? node24335 : node24304;
												assign node24304 = (inp[14]) ? node24320 : node24305;
													assign node24305 = (inp[5]) ? node24313 : node24306;
														assign node24306 = (inp[15]) ? node24310 : node24307;
															assign node24307 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node24310 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node24313 = (inp[15]) ? node24317 : node24314;
															assign node24314 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node24317 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node24320 = (inp[15]) ? node24328 : node24321;
														assign node24321 = (inp[0]) ? node24325 : node24322;
															assign node24322 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node24325 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node24328 = (inp[0]) ? node24332 : node24329;
															assign node24329 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node24332 = (inp[3]) ? 4'b1101 : 4'b1101;
												assign node24335 = (inp[5]) ? node24351 : node24336;
													assign node24336 = (inp[0]) ? node24344 : node24337;
														assign node24337 = (inp[14]) ? node24341 : node24338;
															assign node24338 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node24341 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node24344 = (inp[15]) ? node24348 : node24345;
															assign node24345 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node24348 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node24351 = (inp[14]) ? node24359 : node24352;
														assign node24352 = (inp[15]) ? node24356 : node24353;
															assign node24353 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node24356 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node24359 = (inp[3]) ? node24363 : node24360;
															assign node24360 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node24363 = (inp[15]) ? 4'b1101 : 4'b1101;
											assign node24366 = (inp[14]) ? node24398 : node24367;
												assign node24367 = (inp[2]) ? node24383 : node24368;
													assign node24368 = (inp[5]) ? node24376 : node24369;
														assign node24369 = (inp[0]) ? node24373 : node24370;
															assign node24370 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node24373 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node24376 = (inp[0]) ? node24380 : node24377;
															assign node24377 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node24380 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node24383 = (inp[5]) ? node24391 : node24384;
														assign node24384 = (inp[0]) ? node24388 : node24385;
															assign node24385 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node24388 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node24391 = (inp[15]) ? node24395 : node24392;
															assign node24392 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node24395 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node24398 = (inp[5]) ? node24412 : node24399;
													assign node24399 = (inp[0]) ? node24405 : node24400;
														assign node24400 = (inp[3]) ? 4'b1110 : node24401;
															assign node24401 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node24405 = (inp[2]) ? node24409 : node24406;
															assign node24406 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node24409 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node24412 = (inp[2]) ? node24420 : node24413;
														assign node24413 = (inp[15]) ? node24417 : node24414;
															assign node24414 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node24417 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node24420 = (inp[15]) ? node24424 : node24421;
															assign node24421 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node24424 = (inp[0]) ? 4'b1100 : 4'b1110;
									assign node24427 = (inp[7]) ? node24533 : node24428;
										assign node24428 = (inp[8]) ? node24480 : node24429;
											assign node24429 = (inp[14]) ? node24457 : node24430;
												assign node24430 = (inp[2]) ? node24444 : node24431;
													assign node24431 = (inp[3]) ? node24437 : node24432;
														assign node24432 = (inp[0]) ? node24434 : 4'b1101;
															assign node24434 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node24437 = (inp[15]) ? node24441 : node24438;
															assign node24438 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node24441 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node24444 = (inp[15]) ? node24452 : node24445;
														assign node24445 = (inp[0]) ? node24449 : node24446;
															assign node24446 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node24449 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node24452 = (inp[5]) ? 4'b1100 : node24453;
															assign node24453 = (inp[0]) ? 4'b1100 : 4'b1100;
												assign node24457 = (inp[0]) ? node24469 : node24458;
													assign node24458 = (inp[15]) ? node24464 : node24459;
														assign node24459 = (inp[3]) ? 4'b1100 : node24460;
															assign node24460 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node24464 = (inp[3]) ? 4'b1110 : node24465;
															assign node24465 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node24469 = (inp[15]) ? node24475 : node24470;
														assign node24470 = (inp[5]) ? 4'b1110 : node24471;
															assign node24471 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node24475 = (inp[2]) ? node24477 : 4'b1100;
															assign node24477 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node24480 = (inp[14]) ? node24510 : node24481;
												assign node24481 = (inp[2]) ? node24497 : node24482;
													assign node24482 = (inp[15]) ? node24490 : node24483;
														assign node24483 = (inp[0]) ? node24487 : node24484;
															assign node24484 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node24487 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node24490 = (inp[0]) ? node24494 : node24491;
															assign node24491 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node24494 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node24497 = (inp[15]) ? node24503 : node24498;
														assign node24498 = (inp[0]) ? node24500 : 4'b0101;
															assign node24500 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node24503 = (inp[0]) ? node24507 : node24504;
															assign node24504 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node24507 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node24510 = (inp[0]) ? node24522 : node24511;
													assign node24511 = (inp[15]) ? node24517 : node24512;
														assign node24512 = (inp[3]) ? 4'b0101 : node24513;
															assign node24513 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node24517 = (inp[5]) ? 4'b0111 : node24518;
															assign node24518 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node24522 = (inp[15]) ? node24528 : node24523;
														assign node24523 = (inp[3]) ? 4'b0111 : node24524;
															assign node24524 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node24528 = (inp[5]) ? 4'b0101 : node24529;
															assign node24529 = (inp[3]) ? 4'b0101 : 4'b0111;
										assign node24533 = (inp[8]) ? node24595 : node24534;
											assign node24534 = (inp[14]) ? node24564 : node24535;
												assign node24535 = (inp[2]) ? node24549 : node24536;
													assign node24536 = (inp[15]) ? node24542 : node24537;
														assign node24537 = (inp[0]) ? node24539 : 4'b1100;
															assign node24539 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node24542 = (inp[0]) ? node24546 : node24543;
															assign node24543 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node24546 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node24549 = (inp[0]) ? node24557 : node24550;
														assign node24550 = (inp[15]) ? node24554 : node24551;
															assign node24551 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node24554 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node24557 = (inp[15]) ? node24561 : node24558;
															assign node24558 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node24561 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node24564 = (inp[3]) ? node24580 : node24565;
													assign node24565 = (inp[5]) ? node24573 : node24566;
														assign node24566 = (inp[0]) ? node24570 : node24567;
															assign node24567 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node24570 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node24573 = (inp[0]) ? node24577 : node24574;
															assign node24574 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node24577 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node24580 = (inp[2]) ? node24588 : node24581;
														assign node24581 = (inp[5]) ? node24585 : node24582;
															assign node24582 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node24585 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node24588 = (inp[15]) ? node24592 : node24589;
															assign node24589 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node24592 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node24595 = (inp[2]) ? node24623 : node24596;
												assign node24596 = (inp[14]) ? node24610 : node24597;
													assign node24597 = (inp[5]) ? node24605 : node24598;
														assign node24598 = (inp[0]) ? node24602 : node24599;
															assign node24599 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node24602 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node24605 = (inp[15]) ? node24607 : 4'b0111;
															assign node24607 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node24610 = (inp[15]) ? node24616 : node24611;
														assign node24611 = (inp[0]) ? node24613 : 4'b0100;
															assign node24613 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node24616 = (inp[0]) ? node24620 : node24617;
															assign node24617 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node24620 = (inp[5]) ? 4'b0100 : 4'b0100;
												assign node24623 = (inp[3]) ? node24637 : node24624;
													assign node24624 = (inp[15]) ? node24630 : node24625;
														assign node24625 = (inp[0]) ? node24627 : 4'b0110;
															assign node24627 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node24630 = (inp[5]) ? node24634 : node24631;
															assign node24631 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node24634 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node24637 = (inp[0]) ? node24641 : node24638;
														assign node24638 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node24641 = (inp[15]) ? 4'b0100 : 4'b0110;
								assign node24644 = (inp[13]) ? node24864 : node24645;
									assign node24645 = (inp[7]) ? node24757 : node24646;
										assign node24646 = (inp[8]) ? node24698 : node24647;
											assign node24647 = (inp[14]) ? node24677 : node24648;
												assign node24648 = (inp[2]) ? node24662 : node24649;
													assign node24649 = (inp[3]) ? node24655 : node24650;
														assign node24650 = (inp[0]) ? 4'b1111 : node24651;
															assign node24651 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node24655 = (inp[0]) ? node24659 : node24656;
															assign node24656 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node24659 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node24662 = (inp[15]) ? node24670 : node24663;
														assign node24663 = (inp[0]) ? node24667 : node24664;
															assign node24664 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node24667 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node24670 = (inp[0]) ? node24674 : node24671;
															assign node24671 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node24674 = (inp[3]) ? 4'b1100 : 4'b1100;
												assign node24677 = (inp[15]) ? node24687 : node24678;
													assign node24678 = (inp[0]) ? node24682 : node24679;
														assign node24679 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node24682 = (inp[3]) ? 4'b1110 : node24683;
															assign node24683 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node24687 = (inp[0]) ? node24693 : node24688;
														assign node24688 = (inp[3]) ? 4'b1110 : node24689;
															assign node24689 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node24693 = (inp[3]) ? 4'b1100 : node24694;
															assign node24694 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node24698 = (inp[14]) ? node24728 : node24699;
												assign node24699 = (inp[2]) ? node24715 : node24700;
													assign node24700 = (inp[3]) ? node24708 : node24701;
														assign node24701 = (inp[15]) ? node24705 : node24702;
															assign node24702 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node24705 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node24708 = (inp[0]) ? node24712 : node24709;
															assign node24709 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node24712 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node24715 = (inp[3]) ? node24721 : node24716;
														assign node24716 = (inp[5]) ? 4'b0101 : node24717;
															assign node24717 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node24721 = (inp[0]) ? node24725 : node24722;
															assign node24722 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node24725 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node24728 = (inp[2]) ? node24744 : node24729;
													assign node24729 = (inp[5]) ? node24737 : node24730;
														assign node24730 = (inp[3]) ? node24734 : node24731;
															assign node24731 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node24734 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node24737 = (inp[3]) ? node24741 : node24738;
															assign node24738 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node24741 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node24744 = (inp[3]) ? node24750 : node24745;
														assign node24745 = (inp[0]) ? 4'b0101 : node24746;
															assign node24746 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node24750 = (inp[15]) ? node24754 : node24751;
															assign node24751 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node24754 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node24757 = (inp[8]) ? node24813 : node24758;
											assign node24758 = (inp[2]) ? node24790 : node24759;
												assign node24759 = (inp[14]) ? node24775 : node24760;
													assign node24760 = (inp[5]) ? node24768 : node24761;
														assign node24761 = (inp[15]) ? node24765 : node24762;
															assign node24762 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node24765 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node24768 = (inp[3]) ? node24772 : node24769;
															assign node24769 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node24772 = (inp[0]) ? 4'b1100 : 4'b1100;
													assign node24775 = (inp[3]) ? node24783 : node24776;
														assign node24776 = (inp[0]) ? node24780 : node24777;
															assign node24777 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node24780 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node24783 = (inp[15]) ? node24787 : node24784;
															assign node24784 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node24787 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node24790 = (inp[5]) ? node24806 : node24791;
													assign node24791 = (inp[0]) ? node24799 : node24792;
														assign node24792 = (inp[15]) ? node24796 : node24793;
															assign node24793 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node24796 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node24799 = (inp[14]) ? node24803 : node24800;
															assign node24800 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node24803 = (inp[3]) ? 4'b0101 : 4'b0101;
													assign node24806 = (inp[0]) ? node24810 : node24807;
														assign node24807 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node24810 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node24813 = (inp[2]) ? node24841 : node24814;
												assign node24814 = (inp[14]) ? node24828 : node24815;
													assign node24815 = (inp[15]) ? node24823 : node24816;
														assign node24816 = (inp[0]) ? node24820 : node24817;
															assign node24817 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node24820 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node24823 = (inp[5]) ? 4'b0101 : node24824;
															assign node24824 = (inp[0]) ? 4'b0101 : 4'b0101;
													assign node24828 = (inp[0]) ? node24836 : node24829;
														assign node24829 = (inp[15]) ? node24833 : node24830;
															assign node24830 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node24833 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node24836 = (inp[15]) ? node24838 : 4'b0110;
															assign node24838 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node24841 = (inp[3]) ? node24857 : node24842;
													assign node24842 = (inp[5]) ? node24850 : node24843;
														assign node24843 = (inp[15]) ? node24847 : node24844;
															assign node24844 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node24847 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node24850 = (inp[15]) ? node24854 : node24851;
															assign node24851 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node24854 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node24857 = (inp[0]) ? node24861 : node24858;
														assign node24858 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node24861 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node24864 = (inp[15]) ? node24974 : node24865;
										assign node24865 = (inp[0]) ? node24919 : node24866;
											assign node24866 = (inp[3]) ? node24896 : node24867;
												assign node24867 = (inp[5]) ? node24883 : node24868;
													assign node24868 = (inp[2]) ? node24876 : node24869;
														assign node24869 = (inp[8]) ? node24873 : node24870;
															assign node24870 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node24873 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node24876 = (inp[14]) ? node24880 : node24877;
															assign node24877 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node24880 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node24883 = (inp[7]) ? node24891 : node24884;
														assign node24884 = (inp[8]) ? node24888 : node24885;
															assign node24885 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node24888 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node24891 = (inp[8]) ? 4'b0100 : node24892;
															assign node24892 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node24896 = (inp[8]) ? node24908 : node24897;
													assign node24897 = (inp[7]) ? node24903 : node24898;
														assign node24898 = (inp[2]) ? 4'b0100 : node24899;
															assign node24899 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node24903 = (inp[2]) ? 4'b0101 : node24904;
															assign node24904 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node24908 = (inp[7]) ? node24914 : node24909;
														assign node24909 = (inp[14]) ? 4'b0101 : node24910;
															assign node24910 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node24914 = (inp[14]) ? 4'b0100 : node24915;
															assign node24915 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node24919 = (inp[5]) ? node24951 : node24920;
												assign node24920 = (inp[3]) ? node24936 : node24921;
													assign node24921 = (inp[14]) ? node24929 : node24922;
														assign node24922 = (inp[2]) ? node24926 : node24923;
															assign node24923 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node24926 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node24929 = (inp[2]) ? node24933 : node24930;
															assign node24930 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node24933 = (inp[7]) ? 4'b0100 : 4'b0100;
													assign node24936 = (inp[2]) ? node24944 : node24937;
														assign node24937 = (inp[8]) ? node24941 : node24938;
															assign node24938 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node24941 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node24944 = (inp[8]) ? node24948 : node24945;
															assign node24945 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node24948 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node24951 = (inp[14]) ? node24967 : node24952;
													assign node24952 = (inp[7]) ? node24960 : node24953;
														assign node24953 = (inp[3]) ? node24957 : node24954;
															assign node24954 = (inp[2]) ? 4'b0110 : 4'b0110;
															assign node24957 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node24960 = (inp[3]) ? node24964 : node24961;
															assign node24961 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node24964 = (inp[2]) ? 4'b0110 : 4'b0110;
													assign node24967 = (inp[8]) ? node24971 : node24968;
														assign node24968 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node24971 = (inp[7]) ? 4'b0110 : 4'b0111;
										assign node24974 = (inp[0]) ? node25030 : node24975;
											assign node24975 = (inp[5]) ? node25007 : node24976;
												assign node24976 = (inp[3]) ? node24992 : node24977;
													assign node24977 = (inp[7]) ? node24985 : node24978;
														assign node24978 = (inp[8]) ? node24982 : node24979;
															assign node24979 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node24982 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node24985 = (inp[8]) ? node24989 : node24986;
															assign node24986 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node24989 = (inp[2]) ? 4'b0100 : 4'b0100;
													assign node24992 = (inp[8]) ? node25000 : node24993;
														assign node24993 = (inp[7]) ? node24997 : node24994;
															assign node24994 = (inp[2]) ? 4'b0110 : 4'b0110;
															assign node24997 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node25000 = (inp[7]) ? node25004 : node25001;
															assign node25001 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node25004 = (inp[2]) ? 4'b0110 : 4'b0110;
												assign node25007 = (inp[7]) ? node25019 : node25008;
													assign node25008 = (inp[8]) ? node25014 : node25009;
														assign node25009 = (inp[2]) ? 4'b0110 : node25010;
															assign node25010 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node25014 = (inp[2]) ? 4'b0111 : node25015;
															assign node25015 = (inp[3]) ? 4'b0111 : 4'b0110;
													assign node25019 = (inp[8]) ? node25025 : node25020;
														assign node25020 = (inp[14]) ? 4'b0111 : node25021;
															assign node25021 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node25025 = (inp[14]) ? 4'b0110 : node25026;
															assign node25026 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node25030 = (inp[3]) ? node25060 : node25031;
												assign node25031 = (inp[5]) ? node25045 : node25032;
													assign node25032 = (inp[2]) ? node25038 : node25033;
														assign node25033 = (inp[7]) ? 4'b0110 : node25034;
															assign node25034 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node25038 = (inp[14]) ? node25042 : node25039;
															assign node25039 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node25042 = (inp[8]) ? 4'b0110 : 4'b0110;
													assign node25045 = (inp[14]) ? node25053 : node25046;
														assign node25046 = (inp[8]) ? node25050 : node25047;
															assign node25047 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node25050 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node25053 = (inp[7]) ? node25057 : node25054;
															assign node25054 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node25057 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node25060 = (inp[8]) ? node25072 : node25061;
													assign node25061 = (inp[7]) ? node25067 : node25062;
														assign node25062 = (inp[14]) ? 4'b0100 : node25063;
															assign node25063 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node25067 = (inp[14]) ? 4'b0101 : node25068;
															assign node25068 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node25072 = (inp[7]) ? node25078 : node25073;
														assign node25073 = (inp[14]) ? 4'b0101 : node25074;
															assign node25074 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node25078 = (inp[14]) ? 4'b0100 : node25079;
															assign node25079 = (inp[2]) ? 4'b0100 : 4'b0101;
					assign node25083 = (inp[15]) ? node26775 : node25084;
						assign node25084 = (inp[0]) ? node25916 : node25085;
							assign node25085 = (inp[3]) ? node25561 : node25086;
								assign node25086 = (inp[5]) ? node25326 : node25087;
									assign node25087 = (inp[8]) ? node25211 : node25088;
										assign node25088 = (inp[7]) ? node25150 : node25089;
											assign node25089 = (inp[14]) ? node25119 : node25090;
												assign node25090 = (inp[2]) ? node25104 : node25091;
													assign node25091 = (inp[13]) ? node25099 : node25092;
														assign node25092 = (inp[1]) ? node25096 : node25093;
															assign node25093 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node25096 = (inp[11]) ? 4'b0111 : 4'b0111;
														assign node25099 = (inp[6]) ? 4'b1111 : node25100;
															assign node25100 = (inp[1]) ? 4'b0111 : 4'b0111;
													assign node25104 = (inp[6]) ? node25112 : node25105;
														assign node25105 = (inp[11]) ? node25109 : node25106;
															assign node25106 = (inp[13]) ? 4'b0110 : 4'b1110;
															assign node25109 = (inp[1]) ? 4'b1110 : 4'b0110;
														assign node25112 = (inp[11]) ? node25116 : node25113;
															assign node25113 = (inp[1]) ? 4'b0110 : 4'b0110;
															assign node25116 = (inp[1]) ? 4'b0110 : 4'b1110;
												assign node25119 = (inp[1]) ? node25135 : node25120;
													assign node25120 = (inp[13]) ? node25128 : node25121;
														assign node25121 = (inp[2]) ? node25125 : node25122;
															assign node25122 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node25125 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node25128 = (inp[2]) ? node25132 : node25129;
															assign node25129 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node25132 = (inp[11]) ? 4'b0110 : 4'b0110;
													assign node25135 = (inp[13]) ? node25143 : node25136;
														assign node25136 = (inp[6]) ? node25140 : node25137;
															assign node25137 = (inp[11]) ? 4'b0110 : 4'b1110;
															assign node25140 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node25143 = (inp[11]) ? node25147 : node25144;
															assign node25144 = (inp[6]) ? 4'b1110 : 4'b0110;
															assign node25147 = (inp[6]) ? 4'b0110 : 4'b1110;
											assign node25150 = (inp[14]) ? node25180 : node25151;
												assign node25151 = (inp[2]) ? node25167 : node25152;
													assign node25152 = (inp[13]) ? node25160 : node25153;
														assign node25153 = (inp[6]) ? node25157 : node25154;
															assign node25154 = (inp[11]) ? 4'b0110 : 4'b1110;
															assign node25157 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node25160 = (inp[11]) ? node25164 : node25161;
															assign node25161 = (inp[1]) ? 4'b0110 : 4'b0110;
															assign node25164 = (inp[6]) ? 4'b0110 : 4'b0110;
													assign node25167 = (inp[6]) ? node25173 : node25168;
														assign node25168 = (inp[11]) ? 4'b1111 : node25169;
															assign node25169 = (inp[13]) ? 4'b0111 : 4'b1111;
														assign node25173 = (inp[11]) ? node25177 : node25174;
															assign node25174 = (inp[13]) ? 4'b1111 : 4'b0111;
															assign node25177 = (inp[13]) ? 4'b0111 : 4'b0111;
												assign node25180 = (inp[1]) ? node25196 : node25181;
													assign node25181 = (inp[6]) ? node25189 : node25182;
														assign node25182 = (inp[11]) ? node25186 : node25183;
															assign node25183 = (inp[13]) ? 4'b0111 : 4'b1111;
															assign node25186 = (inp[13]) ? 4'b1111 : 4'b0111;
														assign node25189 = (inp[2]) ? node25193 : node25190;
															assign node25190 = (inp[13]) ? 4'b0111 : 4'b0111;
															assign node25193 = (inp[13]) ? 4'b0111 : 4'b1111;
													assign node25196 = (inp[13]) ? node25204 : node25197;
														assign node25197 = (inp[2]) ? node25201 : node25198;
															assign node25198 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node25201 = (inp[11]) ? 4'b0111 : 4'b0111;
														assign node25204 = (inp[2]) ? node25208 : node25205;
															assign node25205 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node25208 = (inp[6]) ? 4'b0111 : 4'b0111;
										assign node25211 = (inp[7]) ? node25273 : node25212;
											assign node25212 = (inp[14]) ? node25242 : node25213;
												assign node25213 = (inp[2]) ? node25227 : node25214;
													assign node25214 = (inp[13]) ? node25222 : node25215;
														assign node25215 = (inp[6]) ? node25219 : node25216;
															assign node25216 = (inp[11]) ? 4'b0110 : 4'b1110;
															assign node25219 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node25222 = (inp[6]) ? node25224 : 4'b0110;
															assign node25224 = (inp[11]) ? 4'b0110 : 4'b0110;
													assign node25227 = (inp[6]) ? node25235 : node25228;
														assign node25228 = (inp[11]) ? node25232 : node25229;
															assign node25229 = (inp[1]) ? 4'b0111 : 4'b0111;
															assign node25232 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node25235 = (inp[11]) ? node25239 : node25236;
															assign node25236 = (inp[1]) ? 4'b1111 : 4'b0111;
															assign node25239 = (inp[13]) ? 4'b0111 : 4'b0111;
												assign node25242 = (inp[13]) ? node25258 : node25243;
													assign node25243 = (inp[11]) ? node25251 : node25244;
														assign node25244 = (inp[1]) ? node25248 : node25245;
															assign node25245 = (inp[6]) ? 4'b0111 : 4'b1111;
															assign node25248 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node25251 = (inp[1]) ? node25255 : node25252;
															assign node25252 = (inp[6]) ? 4'b1111 : 4'b0111;
															assign node25255 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node25258 = (inp[2]) ? node25266 : node25259;
														assign node25259 = (inp[1]) ? node25263 : node25260;
															assign node25260 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node25263 = (inp[6]) ? 4'b0111 : 4'b0111;
														assign node25266 = (inp[1]) ? node25270 : node25267;
															assign node25267 = (inp[11]) ? 4'b0111 : 4'b1111;
															assign node25270 = (inp[6]) ? 4'b0111 : 4'b0111;
											assign node25273 = (inp[14]) ? node25303 : node25274;
												assign node25274 = (inp[2]) ? node25288 : node25275;
													assign node25275 = (inp[13]) ? node25283 : node25276;
														assign node25276 = (inp[6]) ? node25280 : node25277;
															assign node25277 = (inp[1]) ? 4'b1111 : 4'b0111;
															assign node25280 = (inp[1]) ? 4'b0111 : 4'b0111;
														assign node25283 = (inp[11]) ? 4'b0111 : node25284;
															assign node25284 = (inp[6]) ? 4'b1111 : 4'b0111;
													assign node25288 = (inp[13]) ? node25296 : node25289;
														assign node25289 = (inp[1]) ? node25293 : node25290;
															assign node25290 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node25293 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node25296 = (inp[6]) ? node25300 : node25297;
															assign node25297 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node25300 = (inp[11]) ? 4'b0110 : 4'b1110;
												assign node25303 = (inp[13]) ? node25319 : node25304;
													assign node25304 = (inp[1]) ? node25312 : node25305;
														assign node25305 = (inp[6]) ? node25309 : node25306;
															assign node25306 = (inp[11]) ? 4'b0110 : 4'b1110;
															assign node25309 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node25312 = (inp[2]) ? node25316 : node25313;
															assign node25313 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node25316 = (inp[11]) ? 4'b0110 : 4'b0110;
													assign node25319 = (inp[6]) ? node25323 : node25320;
														assign node25320 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node25323 = (inp[11]) ? 4'b0110 : 4'b1110;
									assign node25326 = (inp[6]) ? node25438 : node25327;
										assign node25327 = (inp[11]) ? node25389 : node25328;
											assign node25328 = (inp[13]) ? node25358 : node25329;
												assign node25329 = (inp[1]) ? node25345 : node25330;
													assign node25330 = (inp[7]) ? node25338 : node25331;
														assign node25331 = (inp[8]) ? node25335 : node25332;
															assign node25332 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node25335 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node25338 = (inp[8]) ? node25342 : node25339;
															assign node25339 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node25342 = (inp[2]) ? 4'b1100 : 4'b1100;
													assign node25345 = (inp[8]) ? node25351 : node25346;
														assign node25346 = (inp[7]) ? node25348 : 4'b1100;
															assign node25348 = (inp[2]) ? 4'b0101 : 4'b1100;
														assign node25351 = (inp[7]) ? node25355 : node25352;
															assign node25352 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node25355 = (inp[14]) ? 4'b0100 : 4'b0100;
												assign node25358 = (inp[1]) ? node25374 : node25359;
													assign node25359 = (inp[8]) ? node25367 : node25360;
														assign node25360 = (inp[7]) ? node25364 : node25361;
															assign node25361 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node25364 = (inp[2]) ? 4'b0101 : 4'b1100;
														assign node25367 = (inp[7]) ? node25371 : node25368;
															assign node25368 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node25371 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node25374 = (inp[8]) ? node25382 : node25375;
														assign node25375 = (inp[7]) ? node25379 : node25376;
															assign node25376 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node25379 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node25382 = (inp[7]) ? node25386 : node25383;
															assign node25383 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node25386 = (inp[14]) ? 4'b0100 : 4'b0100;
											assign node25389 = (inp[1]) ? node25419 : node25390;
												assign node25390 = (inp[13]) ? node25404 : node25391;
													assign node25391 = (inp[2]) ? node25397 : node25392;
														assign node25392 = (inp[14]) ? node25394 : 4'b0100;
															assign node25394 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node25397 = (inp[7]) ? node25401 : node25398;
															assign node25398 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node25401 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node25404 = (inp[8]) ? node25412 : node25405;
														assign node25405 = (inp[7]) ? node25409 : node25406;
															assign node25406 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node25409 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node25412 = (inp[7]) ? node25416 : node25413;
															assign node25413 = (inp[14]) ? 4'b1101 : 4'b0100;
															assign node25416 = (inp[14]) ? 4'b1100 : 4'b1100;
												assign node25419 = (inp[7]) ? node25431 : node25420;
													assign node25420 = (inp[8]) ? node25426 : node25421;
														assign node25421 = (inp[13]) ? 4'b1100 : node25422;
															assign node25422 = (inp[2]) ? 4'b0100 : 4'b0100;
														assign node25426 = (inp[14]) ? 4'b1101 : node25427;
															assign node25427 = (inp[2]) ? 4'b1101 : 4'b0100;
													assign node25431 = (inp[8]) ? node25433 : 4'b1101;
														assign node25433 = (inp[14]) ? 4'b1100 : node25434;
															assign node25434 = (inp[2]) ? 4'b1100 : 4'b1101;
										assign node25438 = (inp[11]) ? node25502 : node25439;
											assign node25439 = (inp[1]) ? node25471 : node25440;
												assign node25440 = (inp[13]) ? node25456 : node25441;
													assign node25441 = (inp[14]) ? node25449 : node25442;
														assign node25442 = (inp[2]) ? node25446 : node25443;
															assign node25443 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node25446 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node25449 = (inp[2]) ? node25453 : node25450;
															assign node25450 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node25453 = (inp[7]) ? 4'b0100 : 4'b0100;
													assign node25456 = (inp[7]) ? node25464 : node25457;
														assign node25457 = (inp[8]) ? node25461 : node25458;
															assign node25458 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node25461 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node25464 = (inp[8]) ? node25468 : node25465;
															assign node25465 = (inp[2]) ? 4'b1101 : 4'b0100;
															assign node25468 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node25471 = (inp[13]) ? node25487 : node25472;
													assign node25472 = (inp[8]) ? node25480 : node25473;
														assign node25473 = (inp[7]) ? node25477 : node25474;
															assign node25474 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node25477 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node25480 = (inp[7]) ? node25484 : node25481;
															assign node25481 = (inp[2]) ? 4'b1101 : 4'b0100;
															assign node25484 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node25487 = (inp[14]) ? node25495 : node25488;
														assign node25488 = (inp[2]) ? node25492 : node25489;
															assign node25489 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node25492 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node25495 = (inp[2]) ? node25499 : node25496;
															assign node25496 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node25499 = (inp[7]) ? 4'b1100 : 4'b1100;
											assign node25502 = (inp[1]) ? node25532 : node25503;
												assign node25503 = (inp[13]) ? node25517 : node25504;
													assign node25504 = (inp[2]) ? node25510 : node25505;
														assign node25505 = (inp[7]) ? 4'b1101 : node25506;
															assign node25506 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node25510 = (inp[7]) ? node25514 : node25511;
															assign node25511 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node25514 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node25517 = (inp[8]) ? node25525 : node25518;
														assign node25518 = (inp[7]) ? node25522 : node25519;
															assign node25519 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node25522 = (inp[14]) ? 4'b0101 : 4'b1100;
														assign node25525 = (inp[7]) ? node25529 : node25526;
															assign node25526 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node25529 = (inp[14]) ? 4'b0100 : 4'b0100;
												assign node25532 = (inp[13]) ? node25546 : node25533;
													assign node25533 = (inp[8]) ? node25539 : node25534;
														assign node25534 = (inp[7]) ? 4'b0101 : node25535;
															assign node25535 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node25539 = (inp[7]) ? node25543 : node25540;
															assign node25540 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node25543 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node25546 = (inp[8]) ? node25554 : node25547;
														assign node25547 = (inp[7]) ? node25551 : node25548;
															assign node25548 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node25551 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node25554 = (inp[7]) ? node25558 : node25555;
															assign node25555 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node25558 = (inp[2]) ? 4'b0100 : 4'b0100;
								assign node25561 = (inp[1]) ? node25761 : node25562;
									assign node25562 = (inp[11]) ? node25652 : node25563;
										assign node25563 = (inp[6]) ? node25605 : node25564;
											assign node25564 = (inp[13]) ? node25582 : node25565;
												assign node25565 = (inp[8]) ? node25571 : node25566;
													assign node25566 = (inp[7]) ? 4'b1101 : node25567;
														assign node25567 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node25571 = (inp[7]) ? node25577 : node25572;
														assign node25572 = (inp[14]) ? 4'b1101 : node25573;
															assign node25573 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node25577 = (inp[2]) ? 4'b1100 : node25578;
															assign node25578 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node25582 = (inp[7]) ? node25594 : node25583;
													assign node25583 = (inp[8]) ? node25589 : node25584;
														assign node25584 = (inp[2]) ? 4'b1100 : node25585;
															assign node25585 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node25589 = (inp[14]) ? 4'b0101 : node25590;
															assign node25590 = (inp[2]) ? 4'b0101 : 4'b1100;
													assign node25594 = (inp[8]) ? node25600 : node25595;
														assign node25595 = (inp[2]) ? 4'b0101 : node25596;
															assign node25596 = (inp[14]) ? 4'b0101 : 4'b1100;
														assign node25600 = (inp[14]) ? 4'b0100 : node25601;
															assign node25601 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node25605 = (inp[13]) ? node25629 : node25606;
												assign node25606 = (inp[14]) ? node25622 : node25607;
													assign node25607 = (inp[8]) ? node25615 : node25608;
														assign node25608 = (inp[7]) ? node25612 : node25609;
															assign node25609 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node25612 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node25615 = (inp[2]) ? node25619 : node25616;
															assign node25616 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node25619 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node25622 = (inp[7]) ? node25626 : node25623;
														assign node25623 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node25626 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node25629 = (inp[7]) ? node25641 : node25630;
													assign node25630 = (inp[8]) ? node25636 : node25631;
														assign node25631 = (inp[2]) ? 4'b0100 : node25632;
															assign node25632 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node25636 = (inp[2]) ? 4'b1101 : node25637;
															assign node25637 = (inp[14]) ? 4'b1101 : 4'b0100;
													assign node25641 = (inp[8]) ? node25647 : node25642;
														assign node25642 = (inp[14]) ? 4'b1101 : node25643;
															assign node25643 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node25647 = (inp[14]) ? 4'b1100 : node25648;
															assign node25648 = (inp[2]) ? 4'b1100 : 4'b1101;
										assign node25652 = (inp[6]) ? node25706 : node25653;
											assign node25653 = (inp[13]) ? node25683 : node25654;
												assign node25654 = (inp[5]) ? node25670 : node25655;
													assign node25655 = (inp[2]) ? node25663 : node25656;
														assign node25656 = (inp[14]) ? node25660 : node25657;
															assign node25657 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node25660 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node25663 = (inp[14]) ? node25667 : node25664;
															assign node25664 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node25667 = (inp[8]) ? 4'b0100 : 4'b0100;
													assign node25670 = (inp[14]) ? node25676 : node25671;
														assign node25671 = (inp[2]) ? node25673 : 4'b0101;
															assign node25673 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node25676 = (inp[2]) ? node25680 : node25677;
															assign node25677 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node25680 = (inp[7]) ? 4'b0100 : 4'b0100;
												assign node25683 = (inp[8]) ? node25695 : node25684;
													assign node25684 = (inp[7]) ? node25690 : node25685;
														assign node25685 = (inp[14]) ? 4'b0100 : node25686;
															assign node25686 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node25690 = (inp[2]) ? 4'b1101 : node25691;
															assign node25691 = (inp[14]) ? 4'b1101 : 4'b0100;
													assign node25695 = (inp[7]) ? node25701 : node25696;
														assign node25696 = (inp[2]) ? 4'b1101 : node25697;
															assign node25697 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node25701 = (inp[14]) ? 4'b1100 : node25702;
															assign node25702 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node25706 = (inp[13]) ? node25738 : node25707;
												assign node25707 = (inp[2]) ? node25723 : node25708;
													assign node25708 = (inp[14]) ? node25716 : node25709;
														assign node25709 = (inp[8]) ? node25713 : node25710;
															assign node25710 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node25713 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node25716 = (inp[7]) ? node25720 : node25717;
															assign node25717 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node25720 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node25723 = (inp[5]) ? node25731 : node25724;
														assign node25724 = (inp[14]) ? node25728 : node25725;
															assign node25725 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node25728 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node25731 = (inp[7]) ? node25735 : node25732;
															assign node25732 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node25735 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node25738 = (inp[8]) ? node25750 : node25739;
													assign node25739 = (inp[7]) ? node25745 : node25740;
														assign node25740 = (inp[14]) ? 4'b1100 : node25741;
															assign node25741 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node25745 = (inp[14]) ? 4'b0101 : node25746;
															assign node25746 = (inp[2]) ? 4'b0101 : 4'b1100;
													assign node25750 = (inp[7]) ? node25756 : node25751;
														assign node25751 = (inp[14]) ? 4'b0101 : node25752;
															assign node25752 = (inp[2]) ? 4'b0101 : 4'b1100;
														assign node25756 = (inp[14]) ? 4'b0100 : node25757;
															assign node25757 = (inp[2]) ? 4'b0100 : 4'b0101;
									assign node25761 = (inp[8]) ? node25855 : node25762;
										assign node25762 = (inp[7]) ? node25824 : node25763;
											assign node25763 = (inp[14]) ? node25793 : node25764;
												assign node25764 = (inp[2]) ? node25778 : node25765;
													assign node25765 = (inp[11]) ? node25773 : node25766;
														assign node25766 = (inp[5]) ? node25770 : node25767;
															assign node25767 = (inp[6]) ? 4'b1101 : 4'b0101;
															assign node25770 = (inp[6]) ? 4'b0101 : 4'b0101;
														assign node25773 = (inp[13]) ? node25775 : 4'b0101;
															assign node25775 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node25778 = (inp[6]) ? node25786 : node25779;
														assign node25779 = (inp[5]) ? node25783 : node25780;
															assign node25780 = (inp[11]) ? 4'b0100 : 4'b0100;
															assign node25783 = (inp[13]) ? 4'b0100 : 4'b0100;
														assign node25786 = (inp[13]) ? node25790 : node25787;
															assign node25787 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node25790 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node25793 = (inp[13]) ? node25809 : node25794;
													assign node25794 = (inp[2]) ? node25802 : node25795;
														assign node25795 = (inp[6]) ? node25799 : node25796;
															assign node25796 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node25799 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node25802 = (inp[11]) ? node25806 : node25803;
															assign node25803 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node25806 = (inp[6]) ? 4'b1100 : 4'b0100;
													assign node25809 = (inp[5]) ? node25817 : node25810;
														assign node25810 = (inp[2]) ? node25814 : node25811;
															assign node25811 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node25814 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node25817 = (inp[11]) ? node25821 : node25818;
															assign node25818 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node25821 = (inp[6]) ? 4'b0100 : 4'b1100;
											assign node25824 = (inp[2]) ? node25848 : node25825;
												assign node25825 = (inp[14]) ? node25841 : node25826;
													assign node25826 = (inp[5]) ? node25834 : node25827;
														assign node25827 = (inp[6]) ? node25831 : node25828;
															assign node25828 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node25831 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node25834 = (inp[11]) ? node25838 : node25835;
															assign node25835 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node25838 = (inp[13]) ? 4'b0100 : 4'b0100;
													assign node25841 = (inp[6]) ? node25845 : node25842;
														assign node25842 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node25845 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node25848 = (inp[6]) ? node25852 : node25849;
													assign node25849 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node25852 = (inp[11]) ? 4'b0101 : 4'b1101;
										assign node25855 = (inp[7]) ? node25885 : node25856;
											assign node25856 = (inp[14]) ? node25878 : node25857;
												assign node25857 = (inp[2]) ? node25871 : node25858;
													assign node25858 = (inp[5]) ? node25866 : node25859;
														assign node25859 = (inp[13]) ? node25863 : node25860;
															assign node25860 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node25863 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node25866 = (inp[13]) ? 4'b0100 : node25867;
															assign node25867 = (inp[11]) ? 4'b0100 : 4'b0100;
													assign node25871 = (inp[11]) ? node25875 : node25872;
														assign node25872 = (inp[6]) ? 4'b1101 : 4'b0101;
														assign node25875 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node25878 = (inp[6]) ? node25882 : node25879;
													assign node25879 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node25882 = (inp[11]) ? 4'b0101 : 4'b1101;
											assign node25885 = (inp[14]) ? node25909 : node25886;
												assign node25886 = (inp[2]) ? node25894 : node25887;
													assign node25887 = (inp[11]) ? node25891 : node25888;
														assign node25888 = (inp[6]) ? 4'b1101 : 4'b0101;
														assign node25891 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node25894 = (inp[13]) ? node25902 : node25895;
														assign node25895 = (inp[5]) ? node25899 : node25896;
															assign node25896 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node25899 = (inp[11]) ? 4'b0100 : 4'b1100;
														assign node25902 = (inp[6]) ? node25906 : node25903;
															assign node25903 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node25906 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node25909 = (inp[11]) ? node25913 : node25910;
													assign node25910 = (inp[6]) ? 4'b1100 : 4'b0100;
													assign node25913 = (inp[6]) ? 4'b0100 : 4'b1100;
							assign node25916 = (inp[5]) ? node26394 : node25917;
								assign node25917 = (inp[3]) ? node26159 : node25918;
									assign node25918 = (inp[13]) ? node26040 : node25919;
										assign node25919 = (inp[7]) ? node25979 : node25920;
											assign node25920 = (inp[8]) ? node25948 : node25921;
												assign node25921 = (inp[2]) ? node25935 : node25922;
													assign node25922 = (inp[14]) ? node25930 : node25923;
														assign node25923 = (inp[1]) ? node25927 : node25924;
															assign node25924 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node25927 = (inp[6]) ? 4'b0101 : 4'b0101;
														assign node25930 = (inp[11]) ? 4'b1100 : node25931;
															assign node25931 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node25935 = (inp[14]) ? node25943 : node25936;
														assign node25936 = (inp[6]) ? node25940 : node25937;
															assign node25937 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node25940 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node25943 = (inp[6]) ? 4'b0100 : node25944;
															assign node25944 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node25948 = (inp[2]) ? node25964 : node25949;
													assign node25949 = (inp[14]) ? node25957 : node25950;
														assign node25950 = (inp[6]) ? node25954 : node25951;
															assign node25951 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node25954 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node25957 = (inp[6]) ? node25961 : node25958;
															assign node25958 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node25961 = (inp[1]) ? 4'b0101 : 4'b0101;
													assign node25964 = (inp[11]) ? node25972 : node25965;
														assign node25965 = (inp[14]) ? node25969 : node25966;
															assign node25966 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node25969 = (inp[1]) ? 4'b0101 : 4'b0101;
														assign node25972 = (inp[6]) ? node25976 : node25973;
															assign node25973 = (inp[1]) ? 4'b1101 : 4'b0101;
															assign node25976 = (inp[1]) ? 4'b0101 : 4'b1101;
											assign node25979 = (inp[8]) ? node26011 : node25980;
												assign node25980 = (inp[2]) ? node25996 : node25981;
													assign node25981 = (inp[14]) ? node25989 : node25982;
														assign node25982 = (inp[1]) ? node25986 : node25983;
															assign node25983 = (inp[11]) ? 4'b0100 : 4'b0100;
															assign node25986 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node25989 = (inp[11]) ? node25993 : node25990;
															assign node25990 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node25993 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node25996 = (inp[1]) ? node26004 : node25997;
														assign node25997 = (inp[14]) ? node26001 : node25998;
															assign node25998 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node26001 = (inp[11]) ? 4'b0101 : 4'b0101;
														assign node26004 = (inp[14]) ? node26008 : node26005;
															assign node26005 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node26008 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node26011 = (inp[2]) ? node26025 : node26012;
													assign node26012 = (inp[14]) ? node26018 : node26013;
														assign node26013 = (inp[11]) ? 4'b0101 : node26014;
															assign node26014 = (inp[1]) ? 4'b0101 : 4'b0101;
														assign node26018 = (inp[1]) ? node26022 : node26019;
															assign node26019 = (inp[11]) ? 4'b0100 : 4'b0100;
															assign node26022 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node26025 = (inp[11]) ? node26033 : node26026;
														assign node26026 = (inp[1]) ? node26030 : node26027;
															assign node26027 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node26030 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node26033 = (inp[14]) ? node26037 : node26034;
															assign node26034 = (inp[1]) ? 4'b0100 : 4'b0100;
															assign node26037 = (inp[6]) ? 4'b0100 : 4'b0100;
										assign node26040 = (inp[6]) ? node26100 : node26041;
											assign node26041 = (inp[11]) ? node26073 : node26042;
												assign node26042 = (inp[1]) ? node26058 : node26043;
													assign node26043 = (inp[8]) ? node26051 : node26044;
														assign node26044 = (inp[7]) ? node26048 : node26045;
															assign node26045 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node26048 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node26051 = (inp[7]) ? node26055 : node26052;
															assign node26052 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node26055 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node26058 = (inp[2]) ? node26066 : node26059;
														assign node26059 = (inp[7]) ? node26063 : node26060;
															assign node26060 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node26063 = (inp[14]) ? 4'b0100 : 4'b0100;
														assign node26066 = (inp[8]) ? node26070 : node26067;
															assign node26067 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node26070 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node26073 = (inp[1]) ? node26087 : node26074;
													assign node26074 = (inp[7]) ? node26082 : node26075;
														assign node26075 = (inp[8]) ? node26079 : node26076;
															assign node26076 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node26079 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node26082 = (inp[8]) ? node26084 : 4'b1101;
															assign node26084 = (inp[2]) ? 4'b1100 : 4'b1100;
													assign node26087 = (inp[14]) ? node26095 : node26088;
														assign node26088 = (inp[2]) ? node26092 : node26089;
															assign node26089 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node26092 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node26095 = (inp[7]) ? 4'b1100 : node26096;
															assign node26096 = (inp[8]) ? 4'b1101 : 4'b1100;
											assign node26100 = (inp[11]) ? node26128 : node26101;
												assign node26101 = (inp[1]) ? node26117 : node26102;
													assign node26102 = (inp[8]) ? node26110 : node26103;
														assign node26103 = (inp[7]) ? node26107 : node26104;
															assign node26104 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node26107 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node26110 = (inp[7]) ? node26114 : node26111;
															assign node26111 = (inp[2]) ? 4'b1101 : 4'b0100;
															assign node26114 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node26117 = (inp[8]) ? node26123 : node26118;
														assign node26118 = (inp[7]) ? node26120 : 4'b1100;
															assign node26120 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node26123 = (inp[7]) ? node26125 : 4'b1101;
															assign node26125 = (inp[2]) ? 4'b1100 : 4'b1100;
												assign node26128 = (inp[1]) ? node26144 : node26129;
													assign node26129 = (inp[8]) ? node26137 : node26130;
														assign node26130 = (inp[7]) ? node26134 : node26131;
															assign node26131 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node26134 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node26137 = (inp[7]) ? node26141 : node26138;
															assign node26138 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node26141 = (inp[2]) ? 4'b0100 : 4'b0100;
													assign node26144 = (inp[14]) ? node26152 : node26145;
														assign node26145 = (inp[8]) ? node26149 : node26146;
															assign node26146 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node26149 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node26152 = (inp[8]) ? node26156 : node26153;
															assign node26153 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node26156 = (inp[7]) ? 4'b0100 : 4'b0101;
									assign node26159 = (inp[1]) ? node26277 : node26160;
										assign node26160 = (inp[8]) ? node26216 : node26161;
											assign node26161 = (inp[7]) ? node26185 : node26162;
												assign node26162 = (inp[14]) ? node26178 : node26163;
													assign node26163 = (inp[2]) ? node26171 : node26164;
														assign node26164 = (inp[6]) ? node26168 : node26165;
															assign node26165 = (inp[11]) ? 4'b0111 : 4'b1111;
															assign node26168 = (inp[11]) ? 4'b1111 : 4'b0111;
														assign node26171 = (inp[13]) ? node26175 : node26172;
															assign node26172 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node26175 = (inp[11]) ? 4'b0110 : 4'b0110;
													assign node26178 = (inp[6]) ? node26182 : node26179;
														assign node26179 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node26182 = (inp[11]) ? 4'b1110 : 4'b0110;
												assign node26185 = (inp[14]) ? node26201 : node26186;
													assign node26186 = (inp[2]) ? node26194 : node26187;
														assign node26187 = (inp[13]) ? node26191 : node26188;
															assign node26188 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node26191 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node26194 = (inp[11]) ? node26198 : node26195;
															assign node26195 = (inp[13]) ? 4'b0111 : 4'b0111;
															assign node26198 = (inp[13]) ? 4'b1111 : 4'b0111;
													assign node26201 = (inp[11]) ? node26209 : node26202;
														assign node26202 = (inp[2]) ? node26206 : node26203;
															assign node26203 = (inp[13]) ? 4'b0111 : 4'b0111;
															assign node26206 = (inp[13]) ? 4'b0111 : 4'b0111;
														assign node26209 = (inp[2]) ? node26213 : node26210;
															assign node26210 = (inp[13]) ? 4'b0111 : 4'b0111;
															assign node26213 = (inp[13]) ? 4'b0111 : 4'b0111;
											assign node26216 = (inp[7]) ? node26246 : node26217;
												assign node26217 = (inp[2]) ? node26233 : node26218;
													assign node26218 = (inp[14]) ? node26226 : node26219;
														assign node26219 = (inp[13]) ? node26223 : node26220;
															assign node26220 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node26223 = (inp[6]) ? 4'b0110 : 4'b0110;
														assign node26226 = (inp[13]) ? node26230 : node26227;
															assign node26227 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node26230 = (inp[6]) ? 4'b0111 : 4'b0111;
													assign node26233 = (inp[13]) ? node26239 : node26234;
														assign node26234 = (inp[14]) ? 4'b0111 : node26235;
															assign node26235 = (inp[11]) ? 4'b0111 : 4'b0111;
														assign node26239 = (inp[11]) ? node26243 : node26240;
															assign node26240 = (inp[6]) ? 4'b1111 : 4'b0111;
															assign node26243 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node26246 = (inp[14]) ? node26262 : node26247;
													assign node26247 = (inp[2]) ? node26255 : node26248;
														assign node26248 = (inp[6]) ? node26252 : node26249;
															assign node26249 = (inp[13]) ? 4'b0111 : 4'b0111;
															assign node26252 = (inp[11]) ? 4'b0111 : 4'b0111;
														assign node26255 = (inp[13]) ? node26259 : node26256;
															assign node26256 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node26259 = (inp[11]) ? 4'b0110 : 4'b0110;
													assign node26262 = (inp[2]) ? node26270 : node26263;
														assign node26263 = (inp[11]) ? node26267 : node26264;
															assign node26264 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node26267 = (inp[6]) ? 4'b0110 : 4'b0110;
														assign node26270 = (inp[11]) ? node26274 : node26271;
															assign node26271 = (inp[13]) ? 4'b0110 : 4'b0110;
															assign node26274 = (inp[13]) ? 4'b0110 : 4'b0110;
										assign node26277 = (inp[13]) ? node26333 : node26278;
											assign node26278 = (inp[6]) ? node26306 : node26279;
												assign node26279 = (inp[11]) ? node26293 : node26280;
													assign node26280 = (inp[7]) ? node26288 : node26281;
														assign node26281 = (inp[8]) ? node26285 : node26282;
															assign node26282 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node26285 = (inp[14]) ? 4'b0111 : 4'b1110;
														assign node26288 = (inp[8]) ? 4'b0110 : node26289;
															assign node26289 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node26293 = (inp[7]) ? node26299 : node26294;
														assign node26294 = (inp[8]) ? node26296 : 4'b0110;
															assign node26296 = (inp[14]) ? 4'b1111 : 4'b0110;
														assign node26299 = (inp[8]) ? node26303 : node26300;
															assign node26300 = (inp[14]) ? 4'b1111 : 4'b0110;
															assign node26303 = (inp[14]) ? 4'b1110 : 4'b1110;
												assign node26306 = (inp[11]) ? node26320 : node26307;
													assign node26307 = (inp[8]) ? node26315 : node26308;
														assign node26308 = (inp[7]) ? node26312 : node26309;
															assign node26309 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node26312 = (inp[14]) ? 4'b1111 : 4'b0110;
														assign node26315 = (inp[7]) ? node26317 : 4'b1111;
															assign node26317 = (inp[14]) ? 4'b1110 : 4'b1110;
													assign node26320 = (inp[7]) ? node26326 : node26321;
														assign node26321 = (inp[8]) ? node26323 : 4'b1110;
															assign node26323 = (inp[2]) ? 4'b0111 : 4'b1110;
														assign node26326 = (inp[8]) ? node26330 : node26327;
															assign node26327 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node26330 = (inp[2]) ? 4'b0110 : 4'b0110;
											assign node26333 = (inp[6]) ? node26363 : node26334;
												assign node26334 = (inp[11]) ? node26350 : node26335;
													assign node26335 = (inp[14]) ? node26343 : node26336;
														assign node26336 = (inp[7]) ? node26340 : node26337;
															assign node26337 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node26340 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node26343 = (inp[2]) ? node26347 : node26344;
															assign node26344 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node26347 = (inp[8]) ? 4'b0110 : 4'b0110;
													assign node26350 = (inp[14]) ? node26356 : node26351;
														assign node26351 = (inp[2]) ? node26353 : 4'b1111;
															assign node26353 = (inp[7]) ? 4'b1110 : 4'b1110;
														assign node26356 = (inp[2]) ? node26360 : node26357;
															assign node26357 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node26360 = (inp[8]) ? 4'b1110 : 4'b1110;
												assign node26363 = (inp[11]) ? node26379 : node26364;
													assign node26364 = (inp[14]) ? node26372 : node26365;
														assign node26365 = (inp[2]) ? node26369 : node26366;
															assign node26366 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node26369 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node26372 = (inp[8]) ? node26376 : node26373;
															assign node26373 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node26376 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node26379 = (inp[14]) ? node26387 : node26380;
														assign node26380 = (inp[2]) ? node26384 : node26381;
															assign node26381 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node26384 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node26387 = (inp[7]) ? node26391 : node26388;
															assign node26388 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node26391 = (inp[8]) ? 4'b0110 : 4'b0111;
								assign node26394 = (inp[7]) ? node26566 : node26395;
									assign node26395 = (inp[8]) ? node26471 : node26396;
										assign node26396 = (inp[14]) ? node26448 : node26397;
											assign node26397 = (inp[2]) ? node26421 : node26398;
												assign node26398 = (inp[6]) ? node26410 : node26399;
													assign node26399 = (inp[11]) ? node26405 : node26400;
														assign node26400 = (inp[1]) ? node26402 : 4'b1111;
															assign node26402 = (inp[13]) ? 4'b0111 : 4'b1111;
														assign node26405 = (inp[1]) ? node26407 : 4'b0111;
															assign node26407 = (inp[13]) ? 4'b1111 : 4'b0111;
													assign node26410 = (inp[11]) ? node26416 : node26411;
														assign node26411 = (inp[1]) ? node26413 : 4'b0111;
															assign node26413 = (inp[13]) ? 4'b1111 : 4'b0111;
														assign node26416 = (inp[1]) ? node26418 : 4'b1111;
															assign node26418 = (inp[13]) ? 4'b0111 : 4'b1111;
												assign node26421 = (inp[3]) ? node26435 : node26422;
													assign node26422 = (inp[11]) ? node26428 : node26423;
														assign node26423 = (inp[13]) ? 4'b0110 : node26424;
															assign node26424 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node26428 = (inp[6]) ? node26432 : node26429;
															assign node26429 = (inp[13]) ? 4'b0110 : 4'b0110;
															assign node26432 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node26435 = (inp[11]) ? node26441 : node26436;
														assign node26436 = (inp[6]) ? node26438 : 4'b1110;
															assign node26438 = (inp[1]) ? 4'b1110 : 4'b0110;
														assign node26441 = (inp[6]) ? node26445 : node26442;
															assign node26442 = (inp[13]) ? 4'b0110 : 4'b0110;
															assign node26445 = (inp[13]) ? 4'b0110 : 4'b1110;
											assign node26448 = (inp[6]) ? node26460 : node26449;
												assign node26449 = (inp[11]) ? node26455 : node26450;
													assign node26450 = (inp[1]) ? node26452 : 4'b1110;
														assign node26452 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node26455 = (inp[1]) ? node26457 : 4'b0110;
														assign node26457 = (inp[13]) ? 4'b1110 : 4'b0110;
												assign node26460 = (inp[11]) ? node26466 : node26461;
													assign node26461 = (inp[1]) ? node26463 : 4'b0110;
														assign node26463 = (inp[13]) ? 4'b1110 : 4'b0110;
													assign node26466 = (inp[1]) ? node26468 : 4'b1110;
														assign node26468 = (inp[13]) ? 4'b0110 : 4'b1110;
										assign node26471 = (inp[14]) ? node26535 : node26472;
											assign node26472 = (inp[2]) ? node26504 : node26473;
												assign node26473 = (inp[1]) ? node26489 : node26474;
													assign node26474 = (inp[13]) ? node26482 : node26475;
														assign node26475 = (inp[3]) ? node26479 : node26476;
															assign node26476 = (inp[6]) ? 4'b1110 : 4'b0110;
															assign node26479 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node26482 = (inp[3]) ? node26486 : node26483;
															assign node26483 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node26486 = (inp[6]) ? 4'b0110 : 4'b0110;
													assign node26489 = (inp[13]) ? node26497 : node26490;
														assign node26490 = (inp[3]) ? node26494 : node26491;
															assign node26491 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node26494 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node26497 = (inp[11]) ? node26501 : node26498;
															assign node26498 = (inp[6]) ? 4'b1110 : 4'b0110;
															assign node26501 = (inp[6]) ? 4'b0110 : 4'b1110;
												assign node26504 = (inp[3]) ? node26520 : node26505;
													assign node26505 = (inp[6]) ? node26513 : node26506;
														assign node26506 = (inp[11]) ? node26510 : node26507;
															assign node26507 = (inp[1]) ? 4'b0111 : 4'b0111;
															assign node26510 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node26513 = (inp[11]) ? node26517 : node26514;
															assign node26514 = (inp[1]) ? 4'b1111 : 4'b0111;
															assign node26517 = (inp[1]) ? 4'b0111 : 4'b0111;
													assign node26520 = (inp[1]) ? node26528 : node26521;
														assign node26521 = (inp[11]) ? node26525 : node26522;
															assign node26522 = (inp[13]) ? 4'b0111 : 4'b0111;
															assign node26525 = (inp[13]) ? 4'b0111 : 4'b0111;
														assign node26528 = (inp[6]) ? node26532 : node26529;
															assign node26529 = (inp[11]) ? 4'b1111 : 4'b0111;
															assign node26532 = (inp[11]) ? 4'b0111 : 4'b1111;
											assign node26535 = (inp[1]) ? node26551 : node26536;
												assign node26536 = (inp[11]) ? node26544 : node26537;
													assign node26537 = (inp[6]) ? node26541 : node26538;
														assign node26538 = (inp[13]) ? 4'b0111 : 4'b1111;
														assign node26541 = (inp[13]) ? 4'b1111 : 4'b0111;
													assign node26544 = (inp[13]) ? node26548 : node26545;
														assign node26545 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node26548 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node26551 = (inp[3]) ? node26559 : node26552;
													assign node26552 = (inp[6]) ? node26556 : node26553;
														assign node26553 = (inp[11]) ? 4'b1111 : 4'b0111;
														assign node26556 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node26559 = (inp[6]) ? node26563 : node26560;
														assign node26560 = (inp[11]) ? 4'b1111 : 4'b0111;
														assign node26563 = (inp[11]) ? 4'b0111 : 4'b1111;
									assign node26566 = (inp[8]) ? node26666 : node26567;
										assign node26567 = (inp[2]) ? node26623 : node26568;
											assign node26568 = (inp[14]) ? node26600 : node26569;
												assign node26569 = (inp[1]) ? node26585 : node26570;
													assign node26570 = (inp[3]) ? node26578 : node26571;
														assign node26571 = (inp[11]) ? node26575 : node26572;
															assign node26572 = (inp[6]) ? 4'b0110 : 4'b1110;
															assign node26575 = (inp[6]) ? 4'b1110 : 4'b0110;
														assign node26578 = (inp[13]) ? node26582 : node26579;
															assign node26579 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node26582 = (inp[6]) ? 4'b0110 : 4'b0110;
													assign node26585 = (inp[3]) ? node26593 : node26586;
														assign node26586 = (inp[11]) ? node26590 : node26587;
															assign node26587 = (inp[13]) ? 4'b0110 : 4'b0110;
															assign node26590 = (inp[6]) ? 4'b0110 : 4'b0110;
														assign node26593 = (inp[6]) ? node26597 : node26594;
															assign node26594 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node26597 = (inp[11]) ? 4'b0110 : 4'b0110;
												assign node26600 = (inp[6]) ? node26612 : node26601;
													assign node26601 = (inp[11]) ? node26607 : node26602;
														assign node26602 = (inp[13]) ? 4'b0111 : node26603;
															assign node26603 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node26607 = (inp[1]) ? 4'b1111 : node26608;
															assign node26608 = (inp[13]) ? 4'b1111 : 4'b0111;
													assign node26612 = (inp[11]) ? node26618 : node26613;
														assign node26613 = (inp[13]) ? 4'b1111 : node26614;
															assign node26614 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node26618 = (inp[13]) ? 4'b0111 : node26619;
															assign node26619 = (inp[1]) ? 4'b0111 : 4'b1111;
											assign node26623 = (inp[14]) ? node26647 : node26624;
												assign node26624 = (inp[6]) ? node26636 : node26625;
													assign node26625 = (inp[11]) ? node26631 : node26626;
														assign node26626 = (inp[1]) ? 4'b0111 : node26627;
															assign node26627 = (inp[13]) ? 4'b0111 : 4'b1111;
														assign node26631 = (inp[13]) ? 4'b1111 : node26632;
															assign node26632 = (inp[1]) ? 4'b1111 : 4'b0111;
													assign node26636 = (inp[11]) ? node26642 : node26637;
														assign node26637 = (inp[1]) ? 4'b1111 : node26638;
															assign node26638 = (inp[13]) ? 4'b1111 : 4'b0111;
														assign node26642 = (inp[13]) ? 4'b0111 : node26643;
															assign node26643 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node26647 = (inp[6]) ? node26655 : node26648;
													assign node26648 = (inp[11]) ? 4'b1111 : node26649;
														assign node26649 = (inp[3]) ? node26651 : 4'b0111;
															assign node26651 = (inp[1]) ? 4'b0111 : 4'b0111;
													assign node26655 = (inp[11]) ? node26661 : node26656;
														assign node26656 = (inp[13]) ? 4'b1111 : node26657;
															assign node26657 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node26661 = (inp[13]) ? 4'b0111 : node26662;
															assign node26662 = (inp[1]) ? 4'b0111 : 4'b1111;
										assign node26666 = (inp[14]) ? node26722 : node26667;
											assign node26667 = (inp[2]) ? node26699 : node26668;
												assign node26668 = (inp[13]) ? node26684 : node26669;
													assign node26669 = (inp[11]) ? node26677 : node26670;
														assign node26670 = (inp[3]) ? node26674 : node26671;
															assign node26671 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node26674 = (inp[1]) ? 4'b0111 : 4'b0111;
														assign node26677 = (inp[1]) ? node26681 : node26678;
															assign node26678 = (inp[6]) ? 4'b1111 : 4'b0111;
															assign node26681 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node26684 = (inp[3]) ? node26692 : node26685;
														assign node26685 = (inp[6]) ? node26689 : node26686;
															assign node26686 = (inp[11]) ? 4'b1111 : 4'b0111;
															assign node26689 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node26692 = (inp[6]) ? node26696 : node26693;
															assign node26693 = (inp[11]) ? 4'b1111 : 4'b0111;
															assign node26696 = (inp[11]) ? 4'b0111 : 4'b1111;
												assign node26699 = (inp[11]) ? node26711 : node26700;
													assign node26700 = (inp[6]) ? node26706 : node26701;
														assign node26701 = (inp[1]) ? 4'b0110 : node26702;
															assign node26702 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node26706 = (inp[13]) ? 4'b1110 : node26707;
															assign node26707 = (inp[1]) ? 4'b1110 : 4'b0110;
													assign node26711 = (inp[6]) ? node26717 : node26712;
														assign node26712 = (inp[13]) ? 4'b1110 : node26713;
															assign node26713 = (inp[1]) ? 4'b1110 : 4'b0110;
														assign node26717 = (inp[13]) ? 4'b0110 : node26718;
															assign node26718 = (inp[1]) ? 4'b0110 : 4'b1110;
											assign node26722 = (inp[3]) ? node26746 : node26723;
												assign node26723 = (inp[1]) ? node26739 : node26724;
													assign node26724 = (inp[6]) ? node26732 : node26725;
														assign node26725 = (inp[13]) ? node26729 : node26726;
															assign node26726 = (inp[11]) ? 4'b0110 : 4'b1110;
															assign node26729 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node26732 = (inp[11]) ? node26736 : node26733;
															assign node26733 = (inp[13]) ? 4'b1110 : 4'b0110;
															assign node26736 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node26739 = (inp[6]) ? node26743 : node26740;
														assign node26740 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node26743 = (inp[11]) ? 4'b0110 : 4'b1110;
												assign node26746 = (inp[13]) ? node26760 : node26747;
													assign node26747 = (inp[2]) ? node26755 : node26748;
														assign node26748 = (inp[1]) ? node26752 : node26749;
															assign node26749 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node26752 = (inp[6]) ? 4'b0110 : 4'b0110;
														assign node26755 = (inp[11]) ? node26757 : 4'b1110;
															assign node26757 = (inp[1]) ? 4'b0110 : 4'b0110;
													assign node26760 = (inp[1]) ? node26768 : node26761;
														assign node26761 = (inp[6]) ? node26765 : node26762;
															assign node26762 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node26765 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node26768 = (inp[11]) ? node26772 : node26769;
															assign node26769 = (inp[6]) ? 4'b1110 : 4'b0110;
															assign node26772 = (inp[6]) ? 4'b0110 : 4'b1110;
						assign node26775 = (inp[0]) ? node27669 : node26776;
							assign node26776 = (inp[5]) ? node27244 : node26777;
								assign node26777 = (inp[3]) ? node27009 : node26778;
									assign node26778 = (inp[1]) ? node26902 : node26779;
										assign node26779 = (inp[7]) ? node26841 : node26780;
											assign node26780 = (inp[8]) ? node26810 : node26781;
												assign node26781 = (inp[2]) ? node26797 : node26782;
													assign node26782 = (inp[14]) ? node26790 : node26783;
														assign node26783 = (inp[11]) ? node26787 : node26784;
															assign node26784 = (inp[6]) ? 4'b0101 : 4'b1101;
															assign node26787 = (inp[6]) ? 4'b1101 : 4'b0101;
														assign node26790 = (inp[13]) ? node26794 : node26791;
															assign node26791 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node26794 = (inp[11]) ? 4'b0100 : 4'b0100;
													assign node26797 = (inp[14]) ? node26805 : node26798;
														assign node26798 = (inp[11]) ? node26802 : node26799;
															assign node26799 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node26802 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node26805 = (inp[13]) ? node26807 : 4'b1100;
															assign node26807 = (inp[11]) ? 4'b0100 : 4'b0100;
												assign node26810 = (inp[2]) ? node26826 : node26811;
													assign node26811 = (inp[14]) ? node26819 : node26812;
														assign node26812 = (inp[6]) ? node26816 : node26813;
															assign node26813 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node26816 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node26819 = (inp[11]) ? node26823 : node26820;
															assign node26820 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node26823 = (inp[13]) ? 4'b1101 : 4'b0101;
													assign node26826 = (inp[11]) ? node26834 : node26827;
														assign node26827 = (inp[14]) ? node26831 : node26828;
															assign node26828 = (inp[13]) ? 4'b0101 : 4'b0101;
															assign node26831 = (inp[6]) ? 4'b0101 : 4'b0101;
														assign node26834 = (inp[6]) ? node26838 : node26835;
															assign node26835 = (inp[13]) ? 4'b1101 : 4'b0101;
															assign node26838 = (inp[13]) ? 4'b0101 : 4'b1101;
											assign node26841 = (inp[8]) ? node26873 : node26842;
												assign node26842 = (inp[2]) ? node26858 : node26843;
													assign node26843 = (inp[14]) ? node26851 : node26844;
														assign node26844 = (inp[13]) ? node26848 : node26845;
															assign node26845 = (inp[11]) ? 4'b0100 : 4'b0100;
															assign node26848 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node26851 = (inp[13]) ? node26855 : node26852;
															assign node26852 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node26855 = (inp[6]) ? 4'b0101 : 4'b0101;
													assign node26858 = (inp[6]) ? node26866 : node26859;
														assign node26859 = (inp[13]) ? node26863 : node26860;
															assign node26860 = (inp[11]) ? 4'b0101 : 4'b1101;
															assign node26863 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node26866 = (inp[14]) ? node26870 : node26867;
															assign node26867 = (inp[13]) ? 4'b0101 : 4'b0101;
															assign node26870 = (inp[11]) ? 4'b0101 : 4'b0101;
												assign node26873 = (inp[2]) ? node26887 : node26874;
													assign node26874 = (inp[14]) ? node26882 : node26875;
														assign node26875 = (inp[6]) ? node26879 : node26876;
															assign node26876 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node26879 = (inp[13]) ? 4'b0101 : 4'b0101;
														assign node26882 = (inp[13]) ? 4'b1100 : node26883;
															assign node26883 = (inp[6]) ? 4'b0100 : 4'b0100;
													assign node26887 = (inp[11]) ? node26895 : node26888;
														assign node26888 = (inp[6]) ? node26892 : node26889;
															assign node26889 = (inp[13]) ? 4'b0100 : 4'b1100;
															assign node26892 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node26895 = (inp[13]) ? node26899 : node26896;
															assign node26896 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node26899 = (inp[6]) ? 4'b0100 : 4'b1100;
										assign node26902 = (inp[7]) ? node26958 : node26903;
											assign node26903 = (inp[8]) ? node26935 : node26904;
												assign node26904 = (inp[2]) ? node26920 : node26905;
													assign node26905 = (inp[14]) ? node26913 : node26906;
														assign node26906 = (inp[6]) ? node26910 : node26907;
															assign node26907 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node26910 = (inp[13]) ? 4'b0101 : 4'b0101;
														assign node26913 = (inp[13]) ? node26917 : node26914;
															assign node26914 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node26917 = (inp[11]) ? 4'b0100 : 4'b0100;
													assign node26920 = (inp[11]) ? node26928 : node26921;
														assign node26921 = (inp[6]) ? node26925 : node26922;
															assign node26922 = (inp[13]) ? 4'b0100 : 4'b1100;
															assign node26925 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node26928 = (inp[6]) ? node26932 : node26929;
															assign node26929 = (inp[13]) ? 4'b1100 : 4'b0100;
															assign node26932 = (inp[13]) ? 4'b0100 : 4'b1100;
												assign node26935 = (inp[14]) ? node26951 : node26936;
													assign node26936 = (inp[2]) ? node26944 : node26937;
														assign node26937 = (inp[13]) ? node26941 : node26938;
															assign node26938 = (inp[11]) ? 4'b0100 : 4'b0100;
															assign node26941 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node26944 = (inp[6]) ? node26948 : node26945;
															assign node26945 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node26948 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node26951 = (inp[6]) ? node26955 : node26952;
														assign node26952 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node26955 = (inp[11]) ? 4'b0101 : 4'b1101;
											assign node26958 = (inp[8]) ? node26980 : node26959;
												assign node26959 = (inp[14]) ? node26973 : node26960;
													assign node26960 = (inp[2]) ? node26966 : node26961;
														assign node26961 = (inp[11]) ? node26963 : 4'b0100;
															assign node26963 = (inp[6]) ? 4'b0100 : 4'b0100;
														assign node26966 = (inp[11]) ? node26970 : node26967;
															assign node26967 = (inp[6]) ? 4'b1101 : 4'b0101;
															assign node26970 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node26973 = (inp[6]) ? node26977 : node26974;
														assign node26974 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node26977 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node26980 = (inp[2]) ? node26994 : node26981;
													assign node26981 = (inp[14]) ? node26989 : node26982;
														assign node26982 = (inp[6]) ? node26986 : node26983;
															assign node26983 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node26986 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node26989 = (inp[6]) ? 4'b0100 : node26990;
															assign node26990 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node26994 = (inp[14]) ? node27002 : node26995;
														assign node26995 = (inp[13]) ? node26999 : node26996;
															assign node26996 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node26999 = (inp[6]) ? 4'b0100 : 4'b0100;
														assign node27002 = (inp[13]) ? node27006 : node27003;
															assign node27003 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node27006 = (inp[6]) ? 4'b0100 : 4'b0100;
									assign node27009 = (inp[1]) ? node27129 : node27010;
										assign node27010 = (inp[6]) ? node27070 : node27011;
											assign node27011 = (inp[11]) ? node27041 : node27012;
												assign node27012 = (inp[13]) ? node27026 : node27013;
													assign node27013 = (inp[2]) ? node27021 : node27014;
														assign node27014 = (inp[8]) ? node27018 : node27015;
															assign node27015 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node27018 = (inp[14]) ? 4'b1110 : 4'b1110;
														assign node27021 = (inp[14]) ? 4'b1111 : node27022;
															assign node27022 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node27026 = (inp[7]) ? node27034 : node27027;
														assign node27027 = (inp[8]) ? node27031 : node27028;
															assign node27028 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node27031 = (inp[2]) ? 4'b0111 : 4'b1110;
														assign node27034 = (inp[8]) ? node27038 : node27035;
															assign node27035 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node27038 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node27041 = (inp[13]) ? node27057 : node27042;
													assign node27042 = (inp[14]) ? node27050 : node27043;
														assign node27043 = (inp[7]) ? node27047 : node27044;
															assign node27044 = (inp[2]) ? 4'b0110 : 4'b0110;
															assign node27047 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node27050 = (inp[7]) ? node27054 : node27051;
															assign node27051 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node27054 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node27057 = (inp[7]) ? node27063 : node27058;
														assign node27058 = (inp[8]) ? node27060 : 4'b0110;
															assign node27060 = (inp[2]) ? 4'b1111 : 4'b0110;
														assign node27063 = (inp[8]) ? node27067 : node27064;
															assign node27064 = (inp[2]) ? 4'b1111 : 4'b0110;
															assign node27067 = (inp[2]) ? 4'b1110 : 4'b1110;
											assign node27070 = (inp[11]) ? node27098 : node27071;
												assign node27071 = (inp[13]) ? node27085 : node27072;
													assign node27072 = (inp[7]) ? node27080 : node27073;
														assign node27073 = (inp[8]) ? node27077 : node27074;
															assign node27074 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node27077 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node27080 = (inp[2]) ? 4'b0110 : node27081;
															assign node27081 = (inp[8]) ? 4'b0110 : 4'b0110;
													assign node27085 = (inp[8]) ? node27093 : node27086;
														assign node27086 = (inp[2]) ? node27090 : node27087;
															assign node27087 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node27090 = (inp[7]) ? 4'b1111 : 4'b0110;
														assign node27093 = (inp[7]) ? 4'b1110 : node27094;
															assign node27094 = (inp[2]) ? 4'b1111 : 4'b0110;
												assign node27098 = (inp[13]) ? node27114 : node27099;
													assign node27099 = (inp[7]) ? node27107 : node27100;
														assign node27100 = (inp[8]) ? node27104 : node27101;
															assign node27101 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node27104 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node27107 = (inp[8]) ? node27111 : node27108;
															assign node27108 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node27111 = (inp[14]) ? 4'b1110 : 4'b1110;
													assign node27114 = (inp[8]) ? node27122 : node27115;
														assign node27115 = (inp[7]) ? node27119 : node27116;
															assign node27116 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node27119 = (inp[14]) ? 4'b0111 : 4'b1110;
														assign node27122 = (inp[2]) ? node27126 : node27123;
															assign node27123 = (inp[14]) ? 4'b0110 : 4'b1110;
															assign node27126 = (inp[7]) ? 4'b0110 : 4'b0111;
										assign node27129 = (inp[7]) ? node27183 : node27130;
											assign node27130 = (inp[8]) ? node27162 : node27131;
												assign node27131 = (inp[2]) ? node27147 : node27132;
													assign node27132 = (inp[14]) ? node27140 : node27133;
														assign node27133 = (inp[6]) ? node27137 : node27134;
															assign node27134 = (inp[13]) ? 4'b0111 : 4'b1111;
															assign node27137 = (inp[13]) ? 4'b0111 : 4'b0111;
														assign node27140 = (inp[11]) ? node27144 : node27141;
															assign node27141 = (inp[13]) ? 4'b0110 : 4'b0110;
															assign node27144 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node27147 = (inp[13]) ? node27155 : node27148;
														assign node27148 = (inp[6]) ? node27152 : node27149;
															assign node27149 = (inp[11]) ? 4'b0110 : 4'b1110;
															assign node27152 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node27155 = (inp[6]) ? node27159 : node27156;
															assign node27156 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node27159 = (inp[11]) ? 4'b0110 : 4'b1110;
												assign node27162 = (inp[2]) ? node27176 : node27163;
													assign node27163 = (inp[14]) ? node27171 : node27164;
														assign node27164 = (inp[6]) ? node27168 : node27165;
															assign node27165 = (inp[13]) ? 4'b0110 : 4'b0110;
															assign node27168 = (inp[13]) ? 4'b0110 : 4'b0110;
														assign node27171 = (inp[13]) ? node27173 : 4'b1111;
															assign node27173 = (inp[6]) ? 4'b0111 : 4'b0111;
													assign node27176 = (inp[11]) ? node27180 : node27177;
														assign node27177 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node27180 = (inp[6]) ? 4'b0111 : 4'b1111;
											assign node27183 = (inp[8]) ? node27215 : node27184;
												assign node27184 = (inp[14]) ? node27200 : node27185;
													assign node27185 = (inp[2]) ? node27193 : node27186;
														assign node27186 = (inp[11]) ? node27190 : node27187;
															assign node27187 = (inp[13]) ? 4'b1110 : 4'b0110;
															assign node27190 = (inp[6]) ? 4'b0110 : 4'b0110;
														assign node27193 = (inp[6]) ? node27197 : node27194;
															assign node27194 = (inp[11]) ? 4'b1111 : 4'b0111;
															assign node27197 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node27200 = (inp[2]) ? node27208 : node27201;
														assign node27201 = (inp[6]) ? node27205 : node27202;
															assign node27202 = (inp[11]) ? 4'b1111 : 4'b0111;
															assign node27205 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node27208 = (inp[11]) ? node27212 : node27209;
															assign node27209 = (inp[6]) ? 4'b1111 : 4'b0111;
															assign node27212 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node27215 = (inp[2]) ? node27231 : node27216;
													assign node27216 = (inp[14]) ? node27224 : node27217;
														assign node27217 = (inp[13]) ? node27221 : node27218;
															assign node27218 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node27221 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node27224 = (inp[11]) ? node27228 : node27225;
															assign node27225 = (inp[6]) ? 4'b1110 : 4'b0110;
															assign node27228 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node27231 = (inp[14]) ? node27239 : node27232;
														assign node27232 = (inp[13]) ? node27236 : node27233;
															assign node27233 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node27236 = (inp[6]) ? 4'b0110 : 4'b0110;
														assign node27239 = (inp[11]) ? 4'b0110 : node27240;
															assign node27240 = (inp[6]) ? 4'b1110 : 4'b0110;
								assign node27244 = (inp[1]) ? node27442 : node27245;
									assign node27245 = (inp[11]) ? node27345 : node27246;
										assign node27246 = (inp[6]) ? node27298 : node27247;
											assign node27247 = (inp[13]) ? node27277 : node27248;
												assign node27248 = (inp[3]) ? node27264 : node27249;
													assign node27249 = (inp[7]) ? node27257 : node27250;
														assign node27250 = (inp[8]) ? node27254 : node27251;
															assign node27251 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node27254 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node27257 = (inp[8]) ? node27261 : node27258;
															assign node27258 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node27261 = (inp[2]) ? 4'b1110 : 4'b1110;
													assign node27264 = (inp[8]) ? node27272 : node27265;
														assign node27265 = (inp[7]) ? node27269 : node27266;
															assign node27266 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node27269 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node27272 = (inp[7]) ? 4'b1110 : node27273;
															assign node27273 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node27277 = (inp[7]) ? node27287 : node27278;
													assign node27278 = (inp[8]) ? node27284 : node27279;
														assign node27279 = (inp[2]) ? 4'b1110 : node27280;
															assign node27280 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node27284 = (inp[2]) ? 4'b0111 : 4'b1110;
													assign node27287 = (inp[8]) ? node27293 : node27288;
														assign node27288 = (inp[2]) ? 4'b0111 : node27289;
															assign node27289 = (inp[14]) ? 4'b0111 : 4'b1110;
														assign node27293 = (inp[14]) ? 4'b0110 : node27294;
															assign node27294 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node27298 = (inp[13]) ? node27322 : node27299;
												assign node27299 = (inp[8]) ? node27311 : node27300;
													assign node27300 = (inp[7]) ? node27306 : node27301;
														assign node27301 = (inp[14]) ? 4'b0110 : node27302;
															assign node27302 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node27306 = (inp[14]) ? 4'b0111 : node27307;
															assign node27307 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node27311 = (inp[7]) ? node27317 : node27312;
														assign node27312 = (inp[2]) ? 4'b0111 : node27313;
															assign node27313 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node27317 = (inp[14]) ? 4'b0110 : node27318;
															assign node27318 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node27322 = (inp[8]) ? node27334 : node27323;
													assign node27323 = (inp[7]) ? node27329 : node27324;
														assign node27324 = (inp[2]) ? 4'b0110 : node27325;
															assign node27325 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node27329 = (inp[2]) ? 4'b1111 : node27330;
															assign node27330 = (inp[14]) ? 4'b1111 : 4'b0110;
													assign node27334 = (inp[7]) ? node27340 : node27335;
														assign node27335 = (inp[2]) ? 4'b1111 : node27336;
															assign node27336 = (inp[14]) ? 4'b1111 : 4'b0110;
														assign node27340 = (inp[2]) ? 4'b1110 : node27341;
															assign node27341 = (inp[14]) ? 4'b1110 : 4'b1111;
										assign node27345 = (inp[6]) ? node27399 : node27346;
											assign node27346 = (inp[13]) ? node27376 : node27347;
												assign node27347 = (inp[3]) ? node27363 : node27348;
													assign node27348 = (inp[14]) ? node27356 : node27349;
														assign node27349 = (inp[8]) ? node27353 : node27350;
															assign node27350 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node27353 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node27356 = (inp[8]) ? node27360 : node27357;
															assign node27357 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node27360 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node27363 = (inp[2]) ? node27371 : node27364;
														assign node27364 = (inp[7]) ? node27368 : node27365;
															assign node27365 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node27368 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node27371 = (inp[7]) ? 4'b0111 : node27372;
															assign node27372 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node27376 = (inp[8]) ? node27388 : node27377;
													assign node27377 = (inp[7]) ? node27383 : node27378;
														assign node27378 = (inp[14]) ? 4'b0110 : node27379;
															assign node27379 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node27383 = (inp[2]) ? 4'b1111 : node27384;
															assign node27384 = (inp[14]) ? 4'b1111 : 4'b0110;
													assign node27388 = (inp[7]) ? node27394 : node27389;
														assign node27389 = (inp[2]) ? 4'b1111 : node27390;
															assign node27390 = (inp[3]) ? 4'b0110 : 4'b1111;
														assign node27394 = (inp[2]) ? 4'b1110 : node27395;
															assign node27395 = (inp[14]) ? 4'b1110 : 4'b1111;
											assign node27399 = (inp[13]) ? node27419 : node27400;
												assign node27400 = (inp[7]) ? node27412 : node27401;
													assign node27401 = (inp[8]) ? node27407 : node27402;
														assign node27402 = (inp[2]) ? 4'b1110 : node27403;
															assign node27403 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node27407 = (inp[2]) ? 4'b1111 : node27408;
															assign node27408 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node27412 = (inp[8]) ? node27414 : 4'b1111;
														assign node27414 = (inp[14]) ? 4'b1110 : node27415;
															assign node27415 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node27419 = (inp[8]) ? node27431 : node27420;
													assign node27420 = (inp[7]) ? node27426 : node27421;
														assign node27421 = (inp[14]) ? 4'b1110 : node27422;
															assign node27422 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node27426 = (inp[2]) ? 4'b0111 : node27427;
															assign node27427 = (inp[14]) ? 4'b0111 : 4'b1110;
													assign node27431 = (inp[7]) ? node27437 : node27432;
														assign node27432 = (inp[2]) ? 4'b0111 : node27433;
															assign node27433 = (inp[14]) ? 4'b0111 : 4'b1110;
														assign node27437 = (inp[14]) ? 4'b0110 : node27438;
															assign node27438 = (inp[2]) ? 4'b0110 : 4'b0111;
									assign node27442 = (inp[13]) ? node27566 : node27443;
										assign node27443 = (inp[3]) ? node27503 : node27444;
											assign node27444 = (inp[14]) ? node27476 : node27445;
												assign node27445 = (inp[8]) ? node27461 : node27446;
													assign node27446 = (inp[2]) ? node27454 : node27447;
														assign node27447 = (inp[7]) ? node27451 : node27448;
															assign node27448 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node27451 = (inp[6]) ? 4'b0110 : 4'b0110;
														assign node27454 = (inp[7]) ? node27458 : node27455;
															assign node27455 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node27458 = (inp[11]) ? 4'b0111 : 4'b0111;
													assign node27461 = (inp[11]) ? node27469 : node27462;
														assign node27462 = (inp[6]) ? node27466 : node27463;
															assign node27463 = (inp[2]) ? 4'b0110 : 4'b1110;
															assign node27466 = (inp[7]) ? 4'b1110 : 4'b0110;
														assign node27469 = (inp[6]) ? node27473 : node27470;
															assign node27470 = (inp[7]) ? 4'b1110 : 4'b0110;
															assign node27473 = (inp[7]) ? 4'b0110 : 4'b1110;
												assign node27476 = (inp[11]) ? node27492 : node27477;
													assign node27477 = (inp[6]) ? node27485 : node27478;
														assign node27478 = (inp[8]) ? node27482 : node27479;
															assign node27479 = (inp[7]) ? 4'b0111 : 4'b1110;
															assign node27482 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node27485 = (inp[8]) ? node27489 : node27486;
															assign node27486 = (inp[7]) ? 4'b1111 : 4'b0110;
															assign node27489 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node27492 = (inp[6]) ? node27498 : node27493;
														assign node27493 = (inp[7]) ? node27495 : 4'b1111;
															assign node27495 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node27498 = (inp[8]) ? node27500 : 4'b1110;
															assign node27500 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node27503 = (inp[7]) ? node27535 : node27504;
												assign node27504 = (inp[8]) ? node27520 : node27505;
													assign node27505 = (inp[2]) ? node27513 : node27506;
														assign node27506 = (inp[14]) ? node27510 : node27507;
															assign node27507 = (inp[6]) ? 4'b1111 : 4'b0111;
															assign node27510 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node27513 = (inp[11]) ? node27517 : node27514;
															assign node27514 = (inp[6]) ? 4'b0110 : 4'b1110;
															assign node27517 = (inp[6]) ? 4'b1110 : 4'b0110;
													assign node27520 = (inp[14]) ? node27528 : node27521;
														assign node27521 = (inp[2]) ? node27525 : node27522;
															assign node27522 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node27525 = (inp[11]) ? 4'b1111 : 4'b0111;
														assign node27528 = (inp[2]) ? node27532 : node27529;
															assign node27529 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node27532 = (inp[11]) ? 4'b1111 : 4'b0111;
												assign node27535 = (inp[8]) ? node27551 : node27536;
													assign node27536 = (inp[14]) ? node27544 : node27537;
														assign node27537 = (inp[2]) ? node27541 : node27538;
															assign node27538 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node27541 = (inp[6]) ? 4'b0111 : 4'b1111;
														assign node27544 = (inp[2]) ? node27548 : node27545;
															assign node27545 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node27548 = (inp[11]) ? 4'b0111 : 4'b0111;
													assign node27551 = (inp[14]) ? node27559 : node27552;
														assign node27552 = (inp[2]) ? node27556 : node27553;
															assign node27553 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node27556 = (inp[6]) ? 4'b0110 : 4'b0110;
														assign node27559 = (inp[2]) ? node27563 : node27560;
															assign node27560 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node27563 = (inp[11]) ? 4'b0110 : 4'b0110;
										assign node27566 = (inp[6]) ? node27622 : node27567;
											assign node27567 = (inp[11]) ? node27595 : node27568;
												assign node27568 = (inp[3]) ? node27582 : node27569;
													assign node27569 = (inp[2]) ? node27575 : node27570;
														assign node27570 = (inp[7]) ? 4'b0111 : node27571;
															assign node27571 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node27575 = (inp[14]) ? node27579 : node27576;
															assign node27576 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node27579 = (inp[8]) ? 4'b0110 : 4'b0110;
													assign node27582 = (inp[8]) ? node27590 : node27583;
														assign node27583 = (inp[14]) ? node27587 : node27584;
															assign node27584 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node27587 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node27590 = (inp[7]) ? 4'b0110 : node27591;
															assign node27591 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node27595 = (inp[3]) ? node27607 : node27596;
													assign node27596 = (inp[14]) ? node27602 : node27597;
														assign node27597 = (inp[8]) ? 4'b1110 : node27598;
															assign node27598 = (inp[7]) ? 4'b1110 : 4'b1110;
														assign node27602 = (inp[8]) ? node27604 : 4'b1110;
															assign node27604 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node27607 = (inp[8]) ? node27615 : node27608;
														assign node27608 = (inp[7]) ? node27612 : node27609;
															assign node27609 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node27612 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node27615 = (inp[7]) ? node27619 : node27616;
															assign node27616 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node27619 = (inp[14]) ? 4'b1110 : 4'b1110;
											assign node27622 = (inp[11]) ? node27646 : node27623;
												assign node27623 = (inp[7]) ? node27635 : node27624;
													assign node27624 = (inp[8]) ? node27630 : node27625;
														assign node27625 = (inp[2]) ? 4'b1110 : node27626;
															assign node27626 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node27630 = (inp[2]) ? 4'b1111 : node27631;
															assign node27631 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node27635 = (inp[8]) ? node27641 : node27636;
														assign node27636 = (inp[2]) ? 4'b1111 : node27637;
															assign node27637 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node27641 = (inp[14]) ? 4'b1110 : node27642;
															assign node27642 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node27646 = (inp[7]) ? node27658 : node27647;
													assign node27647 = (inp[8]) ? node27653 : node27648;
														assign node27648 = (inp[14]) ? 4'b0110 : node27649;
															assign node27649 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node27653 = (inp[2]) ? 4'b0111 : node27654;
															assign node27654 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node27658 = (inp[8]) ? node27664 : node27659;
														assign node27659 = (inp[14]) ? 4'b0111 : node27660;
															assign node27660 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node27664 = (inp[2]) ? 4'b0110 : node27665;
															assign node27665 = (inp[14]) ? 4'b0110 : 4'b0111;
							assign node27669 = (inp[3]) ? node28145 : node27670;
								assign node27670 = (inp[5]) ? node27908 : node27671;
									assign node27671 = (inp[11]) ? node27789 : node27672;
										assign node27672 = (inp[6]) ? node27732 : node27673;
											assign node27673 = (inp[1]) ? node27703 : node27674;
												assign node27674 = (inp[13]) ? node27690 : node27675;
													assign node27675 = (inp[14]) ? node27683 : node27676;
														assign node27676 = (inp[7]) ? node27680 : node27677;
															assign node27677 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node27680 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node27683 = (inp[8]) ? node27687 : node27684;
															assign node27684 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node27687 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node27690 = (inp[8]) ? node27698 : node27691;
														assign node27691 = (inp[7]) ? node27695 : node27692;
															assign node27692 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node27695 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node27698 = (inp[7]) ? node27700 : 4'b0111;
															assign node27700 = (inp[14]) ? 4'b0110 : 4'b0110;
												assign node27703 = (inp[13]) ? node27717 : node27704;
													assign node27704 = (inp[7]) ? node27712 : node27705;
														assign node27705 = (inp[8]) ? node27709 : node27706;
															assign node27706 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node27709 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node27712 = (inp[8]) ? node27714 : 4'b0111;
															assign node27714 = (inp[14]) ? 4'b0110 : 4'b0110;
													assign node27717 = (inp[14]) ? node27725 : node27718;
														assign node27718 = (inp[8]) ? node27722 : node27719;
															assign node27719 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node27722 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node27725 = (inp[8]) ? node27729 : node27726;
															assign node27726 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node27729 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node27732 = (inp[1]) ? node27762 : node27733;
												assign node27733 = (inp[13]) ? node27749 : node27734;
													assign node27734 = (inp[7]) ? node27742 : node27735;
														assign node27735 = (inp[8]) ? node27739 : node27736;
															assign node27736 = (inp[2]) ? 4'b0110 : 4'b0110;
															assign node27739 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node27742 = (inp[8]) ? node27746 : node27743;
															assign node27743 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node27746 = (inp[14]) ? 4'b0110 : 4'b0110;
													assign node27749 = (inp[8]) ? node27755 : node27750;
														assign node27750 = (inp[14]) ? 4'b0110 : node27751;
															assign node27751 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node27755 = (inp[7]) ? node27759 : node27756;
															assign node27756 = (inp[14]) ? 4'b1111 : 4'b0110;
															assign node27759 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node27762 = (inp[13]) ? node27778 : node27763;
													assign node27763 = (inp[8]) ? node27771 : node27764;
														assign node27764 = (inp[7]) ? node27768 : node27765;
															assign node27765 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node27768 = (inp[14]) ? 4'b1111 : 4'b0110;
														assign node27771 = (inp[7]) ? node27775 : node27772;
															assign node27772 = (inp[2]) ? 4'b1111 : 4'b0110;
															assign node27775 = (inp[14]) ? 4'b1110 : 4'b1110;
													assign node27778 = (inp[8]) ? node27784 : node27779;
														assign node27779 = (inp[7]) ? 4'b1111 : node27780;
															assign node27780 = (inp[2]) ? 4'b1110 : 4'b1110;
														assign node27784 = (inp[14]) ? 4'b1110 : node27785;
															assign node27785 = (inp[7]) ? 4'b1110 : 4'b1110;
										assign node27789 = (inp[6]) ? node27847 : node27790;
											assign node27790 = (inp[13]) ? node27820 : node27791;
												assign node27791 = (inp[1]) ? node27805 : node27792;
													assign node27792 = (inp[7]) ? node27800 : node27793;
														assign node27793 = (inp[8]) ? node27797 : node27794;
															assign node27794 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node27797 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node27800 = (inp[8]) ? node27802 : 4'b0111;
															assign node27802 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node27805 = (inp[8]) ? node27813 : node27806;
														assign node27806 = (inp[7]) ? node27810 : node27807;
															assign node27807 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node27810 = (inp[2]) ? 4'b1111 : 4'b0110;
														assign node27813 = (inp[7]) ? node27817 : node27814;
															assign node27814 = (inp[14]) ? 4'b1111 : 4'b0110;
															assign node27817 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node27820 = (inp[1]) ? node27832 : node27821;
													assign node27821 = (inp[8]) ? node27827 : node27822;
														assign node27822 = (inp[7]) ? node27824 : 4'b0110;
															assign node27824 = (inp[14]) ? 4'b1111 : 4'b0110;
														assign node27827 = (inp[7]) ? node27829 : 4'b1111;
															assign node27829 = (inp[2]) ? 4'b1110 : 4'b1110;
													assign node27832 = (inp[2]) ? node27840 : node27833;
														assign node27833 = (inp[14]) ? node27837 : node27834;
															assign node27834 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node27837 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node27840 = (inp[14]) ? node27844 : node27841;
															assign node27841 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node27844 = (inp[7]) ? 4'b1111 : 4'b1110;
											assign node27847 = (inp[13]) ? node27879 : node27848;
												assign node27848 = (inp[1]) ? node27864 : node27849;
													assign node27849 = (inp[14]) ? node27857 : node27850;
														assign node27850 = (inp[8]) ? node27854 : node27851;
															assign node27851 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node27854 = (inp[2]) ? 4'b1110 : 4'b1110;
														assign node27857 = (inp[7]) ? node27861 : node27858;
															assign node27858 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node27861 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node27864 = (inp[7]) ? node27872 : node27865;
														assign node27865 = (inp[8]) ? node27869 : node27866;
															assign node27866 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node27869 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node27872 = (inp[8]) ? node27876 : node27873;
															assign node27873 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node27876 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node27879 = (inp[1]) ? node27895 : node27880;
													assign node27880 = (inp[7]) ? node27888 : node27881;
														assign node27881 = (inp[8]) ? node27885 : node27882;
															assign node27882 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node27885 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node27888 = (inp[8]) ? node27892 : node27889;
															assign node27889 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node27892 = (inp[14]) ? 4'b0110 : 4'b0110;
													assign node27895 = (inp[7]) ? node27903 : node27896;
														assign node27896 = (inp[8]) ? node27900 : node27897;
															assign node27897 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node27900 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node27903 = (inp[14]) ? 4'b0111 : node27904;
															assign node27904 = (inp[2]) ? 4'b0110 : 4'b0110;
									assign node27908 = (inp[13]) ? node28024 : node27909;
										assign node27909 = (inp[14]) ? node27971 : node27910;
											assign node27910 = (inp[6]) ? node27940 : node27911;
												assign node27911 = (inp[11]) ? node27927 : node27912;
													assign node27912 = (inp[1]) ? node27920 : node27913;
														assign node27913 = (inp[2]) ? node27917 : node27914;
															assign node27914 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node27917 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node27920 = (inp[2]) ? node27924 : node27921;
															assign node27921 = (inp[8]) ? 4'b0100 : 4'b1100;
															assign node27924 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node27927 = (inp[2]) ? node27935 : node27928;
														assign node27928 = (inp[8]) ? node27932 : node27929;
															assign node27929 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node27932 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node27935 = (inp[1]) ? 4'b1101 : node27936;
															assign node27936 = (inp[8]) ? 4'b0100 : 4'b0100;
												assign node27940 = (inp[11]) ? node27956 : node27941;
													assign node27941 = (inp[1]) ? node27949 : node27942;
														assign node27942 = (inp[8]) ? node27946 : node27943;
															assign node27943 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node27946 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node27949 = (inp[7]) ? node27953 : node27950;
															assign node27950 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node27953 = (inp[8]) ? 4'b1100 : 4'b0100;
													assign node27956 = (inp[1]) ? node27964 : node27957;
														assign node27957 = (inp[2]) ? node27961 : node27958;
															assign node27958 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node27961 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node27964 = (inp[7]) ? node27968 : node27965;
															assign node27965 = (inp[2]) ? 4'b0100 : 4'b1100;
															assign node27968 = (inp[2]) ? 4'b0100 : 4'b0100;
											assign node27971 = (inp[8]) ? node27995 : node27972;
												assign node27972 = (inp[7]) ? node27980 : node27973;
													assign node27973 = (inp[6]) ? node27977 : node27974;
														assign node27974 = (inp[11]) ? 4'b0100 : 4'b1100;
														assign node27977 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node27980 = (inp[6]) ? node27988 : node27981;
														assign node27981 = (inp[2]) ? node27985 : node27982;
															assign node27982 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node27985 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node27988 = (inp[2]) ? node27992 : node27989;
															assign node27989 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node27992 = (inp[11]) ? 4'b0101 : 4'b0101;
												assign node27995 = (inp[7]) ? node28009 : node27996;
													assign node27996 = (inp[6]) ? node28004 : node27997;
														assign node27997 = (inp[11]) ? node28001 : node27998;
															assign node27998 = (inp[1]) ? 4'b0101 : 4'b1101;
															assign node28001 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node28004 = (inp[1]) ? 4'b0101 : node28005;
															assign node28005 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node28009 = (inp[6]) ? node28017 : node28010;
														assign node28010 = (inp[1]) ? node28014 : node28011;
															assign node28011 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node28014 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node28017 = (inp[1]) ? node28021 : node28018;
															assign node28018 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node28021 = (inp[11]) ? 4'b0100 : 4'b1100;
										assign node28024 = (inp[6]) ? node28086 : node28025;
											assign node28025 = (inp[11]) ? node28055 : node28026;
												assign node28026 = (inp[1]) ? node28040 : node28027;
													assign node28027 = (inp[7]) ? node28035 : node28028;
														assign node28028 = (inp[8]) ? node28032 : node28029;
															assign node28029 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node28032 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node28035 = (inp[8]) ? node28037 : 4'b0101;
															assign node28037 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node28040 = (inp[8]) ? node28048 : node28041;
														assign node28041 = (inp[7]) ? node28045 : node28042;
															assign node28042 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node28045 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node28048 = (inp[7]) ? node28052 : node28049;
															assign node28049 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node28052 = (inp[14]) ? 4'b0100 : 4'b0100;
												assign node28055 = (inp[1]) ? node28071 : node28056;
													assign node28056 = (inp[7]) ? node28064 : node28057;
														assign node28057 = (inp[8]) ? node28061 : node28058;
															assign node28058 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node28061 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node28064 = (inp[8]) ? node28068 : node28065;
															assign node28065 = (inp[2]) ? 4'b1101 : 4'b0100;
															assign node28068 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node28071 = (inp[14]) ? node28079 : node28072;
														assign node28072 = (inp[8]) ? node28076 : node28073;
															assign node28073 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node28076 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node28079 = (inp[8]) ? node28083 : node28080;
															assign node28080 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node28083 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node28086 = (inp[11]) ? node28116 : node28087;
												assign node28087 = (inp[1]) ? node28103 : node28088;
													assign node28088 = (inp[8]) ? node28096 : node28089;
														assign node28089 = (inp[7]) ? node28093 : node28090;
															assign node28090 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node28093 = (inp[2]) ? 4'b1101 : 4'b0100;
														assign node28096 = (inp[7]) ? node28100 : node28097;
															assign node28097 = (inp[2]) ? 4'b1101 : 4'b0100;
															assign node28100 = (inp[2]) ? 4'b1100 : 4'b1100;
													assign node28103 = (inp[8]) ? node28111 : node28104;
														assign node28104 = (inp[7]) ? node28108 : node28105;
															assign node28105 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node28108 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node28111 = (inp[7]) ? node28113 : 4'b1101;
															assign node28113 = (inp[2]) ? 4'b1100 : 4'b1100;
												assign node28116 = (inp[1]) ? node28132 : node28117;
													assign node28117 = (inp[8]) ? node28125 : node28118;
														assign node28118 = (inp[7]) ? node28122 : node28119;
															assign node28119 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node28122 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node28125 = (inp[7]) ? node28129 : node28126;
															assign node28126 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node28129 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node28132 = (inp[7]) ? node28140 : node28133;
														assign node28133 = (inp[8]) ? node28137 : node28134;
															assign node28134 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node28137 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node28140 = (inp[8]) ? node28142 : 4'b0101;
															assign node28142 = (inp[14]) ? 4'b0100 : 4'b0101;
								assign node28145 = (inp[8]) ? node28327 : node28146;
									assign node28146 = (inp[7]) ? node28252 : node28147;
										assign node28147 = (inp[14]) ? node28199 : node28148;
											assign node28148 = (inp[2]) ? node28172 : node28149;
												assign node28149 = (inp[13]) ? node28157 : node28150;
													assign node28150 = (inp[6]) ? node28154 : node28151;
														assign node28151 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node28154 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node28157 = (inp[6]) ? node28165 : node28158;
														assign node28158 = (inp[11]) ? node28162 : node28159;
															assign node28159 = (inp[1]) ? 4'b0101 : 4'b1101;
															assign node28162 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node28165 = (inp[5]) ? node28169 : node28166;
															assign node28166 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node28169 = (inp[11]) ? 4'b0101 : 4'b0101;
												assign node28172 = (inp[5]) ? node28186 : node28173;
													assign node28173 = (inp[6]) ? node28179 : node28174;
														assign node28174 = (inp[1]) ? node28176 : 4'b1100;
															assign node28176 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node28179 = (inp[11]) ? node28183 : node28180;
															assign node28180 = (inp[13]) ? 4'b1100 : 4'b0100;
															assign node28183 = (inp[1]) ? 4'b0100 : 4'b1100;
													assign node28186 = (inp[11]) ? node28194 : node28187;
														assign node28187 = (inp[6]) ? node28191 : node28188;
															assign node28188 = (inp[1]) ? 4'b0100 : 4'b1100;
															assign node28191 = (inp[13]) ? 4'b0100 : 4'b0100;
														assign node28194 = (inp[1]) ? node28196 : 4'b0100;
															assign node28196 = (inp[6]) ? 4'b0100 : 4'b0100;
											assign node28199 = (inp[2]) ? node28229 : node28200;
												assign node28200 = (inp[1]) ? node28214 : node28201;
													assign node28201 = (inp[13]) ? node28209 : node28202;
														assign node28202 = (inp[11]) ? node28206 : node28203;
															assign node28203 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node28206 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node28209 = (inp[5]) ? 4'b0100 : node28210;
															assign node28210 = (inp[6]) ? 4'b0100 : 4'b0100;
													assign node28214 = (inp[5]) ? node28222 : node28215;
														assign node28215 = (inp[13]) ? node28219 : node28216;
															assign node28216 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node28219 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node28222 = (inp[11]) ? node28226 : node28223;
															assign node28223 = (inp[13]) ? 4'b1100 : 4'b0100;
															assign node28226 = (inp[6]) ? 4'b0100 : 4'b0100;
												assign node28229 = (inp[11]) ? node28241 : node28230;
													assign node28230 = (inp[6]) ? node28236 : node28231;
														assign node28231 = (inp[1]) ? node28233 : 4'b1100;
															assign node28233 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node28236 = (inp[1]) ? node28238 : 4'b0100;
															assign node28238 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node28241 = (inp[6]) ? node28247 : node28242;
														assign node28242 = (inp[13]) ? node28244 : 4'b0100;
															assign node28244 = (inp[1]) ? 4'b1100 : 4'b0100;
														assign node28247 = (inp[1]) ? node28249 : 4'b1100;
															assign node28249 = (inp[13]) ? 4'b0100 : 4'b1100;
										assign node28252 = (inp[14]) ? node28304 : node28253;
											assign node28253 = (inp[2]) ? node28285 : node28254;
												assign node28254 = (inp[13]) ? node28270 : node28255;
													assign node28255 = (inp[5]) ? node28263 : node28256;
														assign node28256 = (inp[1]) ? node28260 : node28257;
															assign node28257 = (inp[11]) ? 4'b0100 : 4'b0100;
															assign node28260 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node28263 = (inp[1]) ? node28267 : node28264;
															assign node28264 = (inp[11]) ? 4'b0100 : 4'b0100;
															assign node28267 = (inp[11]) ? 4'b0100 : 4'b0100;
													assign node28270 = (inp[6]) ? node28278 : node28271;
														assign node28271 = (inp[5]) ? node28275 : node28272;
															assign node28272 = (inp[1]) ? 4'b0100 : 4'b0100;
															assign node28275 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node28278 = (inp[11]) ? node28282 : node28279;
															assign node28279 = (inp[1]) ? 4'b1100 : 4'b0100;
															assign node28282 = (inp[1]) ? 4'b0100 : 4'b1100;
												assign node28285 = (inp[11]) ? node28293 : node28286;
													assign node28286 = (inp[6]) ? node28288 : 4'b0101;
														assign node28288 = (inp[13]) ? 4'b1101 : node28289;
															assign node28289 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node28293 = (inp[6]) ? node28299 : node28294;
														assign node28294 = (inp[13]) ? 4'b1101 : node28295;
															assign node28295 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node28299 = (inp[1]) ? 4'b0101 : node28300;
															assign node28300 = (inp[13]) ? 4'b0101 : 4'b1101;
											assign node28304 = (inp[11]) ? node28316 : node28305;
												assign node28305 = (inp[6]) ? node28311 : node28306;
													assign node28306 = (inp[1]) ? 4'b0101 : node28307;
														assign node28307 = (inp[13]) ? 4'b0101 : 4'b1101;
													assign node28311 = (inp[1]) ? 4'b1101 : node28312;
														assign node28312 = (inp[13]) ? 4'b1101 : 4'b0101;
												assign node28316 = (inp[6]) ? node28322 : node28317;
													assign node28317 = (inp[13]) ? 4'b1101 : node28318;
														assign node28318 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node28322 = (inp[1]) ? 4'b0101 : node28323;
														assign node28323 = (inp[13]) ? 4'b0101 : 4'b1101;
									assign node28327 = (inp[7]) ? node28435 : node28328;
										assign node28328 = (inp[2]) ? node28388 : node28329;
											assign node28329 = (inp[14]) ? node28361 : node28330;
												assign node28330 = (inp[5]) ? node28346 : node28331;
													assign node28331 = (inp[11]) ? node28339 : node28332;
														assign node28332 = (inp[6]) ? node28336 : node28333;
															assign node28333 = (inp[13]) ? 4'b0100 : 4'b1100;
															assign node28336 = (inp[1]) ? 4'b0100 : 4'b0100;
														assign node28339 = (inp[6]) ? node28343 : node28340;
															assign node28340 = (inp[13]) ? 4'b0100 : 4'b0100;
															assign node28343 = (inp[13]) ? 4'b0100 : 4'b1100;
													assign node28346 = (inp[6]) ? node28354 : node28347;
														assign node28347 = (inp[11]) ? node28351 : node28348;
															assign node28348 = (inp[13]) ? 4'b0100 : 4'b1100;
															assign node28351 = (inp[13]) ? 4'b0100 : 4'b0100;
														assign node28354 = (inp[11]) ? node28358 : node28355;
															assign node28355 = (inp[1]) ? 4'b0100 : 4'b0100;
															assign node28358 = (inp[13]) ? 4'b0100 : 4'b1100;
												assign node28361 = (inp[5]) ? node28375 : node28362;
													assign node28362 = (inp[1]) ? node28368 : node28363;
														assign node28363 = (inp[11]) ? node28365 : 4'b0101;
															assign node28365 = (inp[6]) ? 4'b0101 : 4'b0101;
														assign node28368 = (inp[11]) ? node28372 : node28369;
															assign node28369 = (inp[6]) ? 4'b1101 : 4'b0101;
															assign node28372 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node28375 = (inp[6]) ? node28383 : node28376;
														assign node28376 = (inp[11]) ? node28380 : node28377;
															assign node28377 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node28380 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node28383 = (inp[11]) ? 4'b0101 : node28384;
															assign node28384 = (inp[1]) ? 4'b1101 : 4'b0101;
											assign node28388 = (inp[5]) ? node28412 : node28389;
												assign node28389 = (inp[6]) ? node28401 : node28390;
													assign node28390 = (inp[11]) ? node28396 : node28391;
														assign node28391 = (inp[1]) ? 4'b0101 : node28392;
															assign node28392 = (inp[13]) ? 4'b0101 : 4'b1101;
														assign node28396 = (inp[13]) ? 4'b1101 : node28397;
															assign node28397 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node28401 = (inp[11]) ? node28407 : node28402;
														assign node28402 = (inp[1]) ? 4'b1101 : node28403;
															assign node28403 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node28407 = (inp[1]) ? 4'b0101 : node28408;
															assign node28408 = (inp[13]) ? 4'b0101 : 4'b1101;
												assign node28412 = (inp[13]) ? node28428 : node28413;
													assign node28413 = (inp[14]) ? node28421 : node28414;
														assign node28414 = (inp[11]) ? node28418 : node28415;
															assign node28415 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node28418 = (inp[1]) ? 4'b0101 : 4'b0101;
														assign node28421 = (inp[11]) ? node28425 : node28422;
															assign node28422 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node28425 = (inp[6]) ? 4'b0101 : 4'b0101;
													assign node28428 = (inp[6]) ? node28432 : node28429;
														assign node28429 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node28432 = (inp[11]) ? 4'b0101 : 4'b1101;
										assign node28435 = (inp[2]) ? node28489 : node28436;
											assign node28436 = (inp[14]) ? node28466 : node28437;
												assign node28437 = (inp[5]) ? node28453 : node28438;
													assign node28438 = (inp[1]) ? node28446 : node28439;
														assign node28439 = (inp[6]) ? node28443 : node28440;
															assign node28440 = (inp[13]) ? 4'b0101 : 4'b0101;
															assign node28443 = (inp[13]) ? 4'b0101 : 4'b0101;
														assign node28446 = (inp[13]) ? node28450 : node28447;
															assign node28447 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node28450 = (inp[11]) ? 4'b0101 : 4'b0101;
													assign node28453 = (inp[6]) ? node28459 : node28454;
														assign node28454 = (inp[13]) ? 4'b1101 : node28455;
															assign node28455 = (inp[11]) ? 4'b0101 : 4'b0101;
														assign node28459 = (inp[11]) ? node28463 : node28460;
															assign node28460 = (inp[13]) ? 4'b1101 : 4'b0101;
															assign node28463 = (inp[1]) ? 4'b0101 : 4'b0101;
												assign node28466 = (inp[11]) ? node28478 : node28467;
													assign node28467 = (inp[6]) ? node28473 : node28468;
														assign node28468 = (inp[1]) ? 4'b0100 : node28469;
															assign node28469 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node28473 = (inp[13]) ? 4'b1100 : node28474;
															assign node28474 = (inp[1]) ? 4'b1100 : 4'b0100;
													assign node28478 = (inp[6]) ? node28484 : node28479;
														assign node28479 = (inp[1]) ? 4'b1100 : node28480;
															assign node28480 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node28484 = (inp[1]) ? 4'b0100 : node28485;
															assign node28485 = (inp[13]) ? 4'b0100 : 4'b1100;
											assign node28489 = (inp[1]) ? node28521 : node28490;
												assign node28490 = (inp[5]) ? node28506 : node28491;
													assign node28491 = (inp[13]) ? node28499 : node28492;
														assign node28492 = (inp[6]) ? node28496 : node28493;
															assign node28493 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node28496 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node28499 = (inp[11]) ? node28503 : node28500;
															assign node28500 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node28503 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node28506 = (inp[13]) ? node28514 : node28507;
														assign node28507 = (inp[6]) ? node28511 : node28508;
															assign node28508 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node28511 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node28514 = (inp[6]) ? node28518 : node28515;
															assign node28515 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node28518 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node28521 = (inp[14]) ? node28529 : node28522;
													assign node28522 = (inp[6]) ? node28526 : node28523;
														assign node28523 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node28526 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node28529 = (inp[11]) ? node28533 : node28530;
														assign node28530 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node28533 = (inp[6]) ? 4'b0100 : 4'b1100;
		assign node28536 = (inp[4]) ? node43066 : node28537;
			assign node28537 = (inp[10]) ? node35657 : node28538;
				assign node28538 = (inp[12]) ? node31996 : node28539;
					assign node28539 = (inp[8]) ? node30227 : node28540;
						assign node28540 = (inp[7]) ? node29308 : node28541;
							assign node28541 = (inp[2]) ? node29009 : node28542;
								assign node28542 = (inp[14]) ? node28778 : node28543;
									assign node28543 = (inp[3]) ? node28653 : node28544;
										assign node28544 = (inp[15]) ? node28600 : node28545;
											assign node28545 = (inp[0]) ? node28577 : node28546;
												assign node28546 = (inp[13]) ? node28562 : node28547;
													assign node28547 = (inp[1]) ? node28555 : node28548;
														assign node28548 = (inp[6]) ? node28552 : node28549;
															assign node28549 = (inp[11]) ? 4'b0011 : 4'b1011;
															assign node28552 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node28555 = (inp[11]) ? node28559 : node28556;
															assign node28556 = (inp[6]) ? 4'b0011 : 4'b1011;
															assign node28559 = (inp[6]) ? 4'b1011 : 4'b0011;
													assign node28562 = (inp[11]) ? node28570 : node28563;
														assign node28563 = (inp[1]) ? node28567 : node28564;
															assign node28564 = (inp[6]) ? 4'b0011 : 4'b1011;
															assign node28567 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node28570 = (inp[6]) ? node28574 : node28571;
															assign node28571 = (inp[1]) ? 4'b1011 : 4'b0011;
															assign node28574 = (inp[1]) ? 4'b0011 : 4'b1011;
												assign node28577 = (inp[6]) ? node28589 : node28578;
													assign node28578 = (inp[11]) ? node28584 : node28579;
														assign node28579 = (inp[13]) ? node28581 : 4'b1001;
															assign node28581 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node28584 = (inp[13]) ? node28586 : 4'b0001;
															assign node28586 = (inp[5]) ? 4'b1001 : 4'b0001;
													assign node28589 = (inp[11]) ? node28595 : node28590;
														assign node28590 = (inp[13]) ? node28592 : 4'b0001;
															assign node28592 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node28595 = (inp[13]) ? node28597 : 4'b1001;
															assign node28597 = (inp[1]) ? 4'b0001 : 4'b1001;
											assign node28600 = (inp[0]) ? node28630 : node28601;
												assign node28601 = (inp[5]) ? node28615 : node28602;
													assign node28602 = (inp[1]) ? node28610 : node28603;
														assign node28603 = (inp[11]) ? node28607 : node28604;
															assign node28604 = (inp[6]) ? 4'b0001 : 4'b1001;
															assign node28607 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node28610 = (inp[13]) ? node28612 : 4'b1001;
															assign node28612 = (inp[11]) ? 4'b0001 : 4'b0001;
													assign node28615 = (inp[1]) ? node28623 : node28616;
														assign node28616 = (inp[13]) ? node28620 : node28617;
															assign node28617 = (inp[11]) ? 4'b0001 : 4'b0001;
															assign node28620 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node28623 = (inp[11]) ? node28627 : node28624;
															assign node28624 = (inp[13]) ? 4'b0001 : 4'b0001;
															assign node28627 = (inp[6]) ? 4'b0001 : 4'b0001;
												assign node28630 = (inp[11]) ? node28642 : node28631;
													assign node28631 = (inp[6]) ? node28637 : node28632;
														assign node28632 = (inp[1]) ? node28634 : 4'b1011;
															assign node28634 = (inp[13]) ? 4'b0011 : 4'b1011;
														assign node28637 = (inp[1]) ? node28639 : 4'b0011;
															assign node28639 = (inp[13]) ? 4'b1011 : 4'b0011;
													assign node28642 = (inp[6]) ? node28648 : node28643;
														assign node28643 = (inp[1]) ? node28645 : 4'b0011;
															assign node28645 = (inp[13]) ? 4'b1011 : 4'b0011;
														assign node28648 = (inp[1]) ? node28650 : 4'b1011;
															assign node28650 = (inp[13]) ? 4'b0011 : 4'b1011;
										assign node28653 = (inp[11]) ? node28715 : node28654;
											assign node28654 = (inp[6]) ? node28686 : node28655;
												assign node28655 = (inp[13]) ? node28671 : node28656;
													assign node28656 = (inp[0]) ? node28664 : node28657;
														assign node28657 = (inp[5]) ? node28661 : node28658;
															assign node28658 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node28661 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node28664 = (inp[15]) ? node28668 : node28665;
															assign node28665 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node28668 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node28671 = (inp[1]) ? node28679 : node28672;
														assign node28672 = (inp[15]) ? node28676 : node28673;
															assign node28673 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node28676 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node28679 = (inp[0]) ? node28683 : node28680;
															assign node28680 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node28683 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node28686 = (inp[13]) ? node28700 : node28687;
													assign node28687 = (inp[1]) ? node28693 : node28688;
														assign node28688 = (inp[5]) ? node28690 : 4'b0011;
															assign node28690 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node28693 = (inp[15]) ? node28697 : node28694;
															assign node28694 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node28697 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node28700 = (inp[1]) ? node28708 : node28701;
														assign node28701 = (inp[0]) ? node28705 : node28702;
															assign node28702 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node28705 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node28708 = (inp[0]) ? node28712 : node28709;
															assign node28709 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node28712 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node28715 = (inp[6]) ? node28747 : node28716;
												assign node28716 = (inp[13]) ? node28732 : node28717;
													assign node28717 = (inp[15]) ? node28725 : node28718;
														assign node28718 = (inp[0]) ? node28722 : node28719;
															assign node28719 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node28722 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node28725 = (inp[5]) ? node28729 : node28726;
															assign node28726 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node28729 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node28732 = (inp[1]) ? node28740 : node28733;
														assign node28733 = (inp[15]) ? node28737 : node28734;
															assign node28734 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node28737 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node28740 = (inp[0]) ? node28744 : node28741;
															assign node28741 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node28744 = (inp[15]) ? 4'b1001 : 4'b1001;
												assign node28747 = (inp[1]) ? node28763 : node28748;
													assign node28748 = (inp[5]) ? node28756 : node28749;
														assign node28749 = (inp[13]) ? node28753 : node28750;
															assign node28750 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node28753 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node28756 = (inp[0]) ? node28760 : node28757;
															assign node28757 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node28760 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node28763 = (inp[13]) ? node28771 : node28764;
														assign node28764 = (inp[15]) ? node28768 : node28765;
															assign node28765 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node28768 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node28771 = (inp[5]) ? node28775 : node28772;
															assign node28772 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node28775 = (inp[15]) ? 4'b0001 : 4'b0001;
									assign node28778 = (inp[0]) ? node28892 : node28779;
										assign node28779 = (inp[15]) ? node28839 : node28780;
											assign node28780 = (inp[5]) ? node28810 : node28781;
												assign node28781 = (inp[3]) ? node28795 : node28782;
													assign node28782 = (inp[6]) ? node28790 : node28783;
														assign node28783 = (inp[11]) ? node28787 : node28784;
															assign node28784 = (inp[13]) ? 4'b0010 : 4'b1010;
															assign node28787 = (inp[13]) ? 4'b0010 : 4'b0010;
														assign node28790 = (inp[11]) ? node28792 : 4'b0010;
															assign node28792 = (inp[13]) ? 4'b0010 : 4'b1010;
													assign node28795 = (inp[1]) ? node28803 : node28796;
														assign node28796 = (inp[13]) ? node28800 : node28797;
															assign node28797 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node28800 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node28803 = (inp[11]) ? node28807 : node28804;
															assign node28804 = (inp[13]) ? 4'b0010 : 4'b0010;
															assign node28807 = (inp[13]) ? 4'b0010 : 4'b0010;
												assign node28810 = (inp[3]) ? node28826 : node28811;
													assign node28811 = (inp[13]) ? node28819 : node28812;
														assign node28812 = (inp[1]) ? node28816 : node28813;
															assign node28813 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node28816 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node28819 = (inp[11]) ? node28823 : node28820;
															assign node28820 = (inp[1]) ? 4'b0010 : 4'b1010;
															assign node28823 = (inp[6]) ? 4'b0010 : 4'b0010;
													assign node28826 = (inp[1]) ? node28834 : node28827;
														assign node28827 = (inp[11]) ? node28831 : node28828;
															assign node28828 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node28831 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node28834 = (inp[11]) ? 4'b0000 : node28835;
															assign node28835 = (inp[6]) ? 4'b0000 : 4'b0000;
											assign node28839 = (inp[3]) ? node28861 : node28840;
												assign node28840 = (inp[11]) ? node28852 : node28841;
													assign node28841 = (inp[6]) ? node28847 : node28842;
														assign node28842 = (inp[13]) ? node28844 : 4'b1000;
															assign node28844 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node28847 = (inp[13]) ? node28849 : 4'b0000;
															assign node28849 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node28852 = (inp[6]) ? node28858 : node28853;
														assign node28853 = (inp[13]) ? node28855 : 4'b0000;
															assign node28855 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node28858 = (inp[1]) ? 4'b0000 : 4'b1000;
												assign node28861 = (inp[5]) ? node28877 : node28862;
													assign node28862 = (inp[13]) ? node28870 : node28863;
														assign node28863 = (inp[1]) ? node28867 : node28864;
															assign node28864 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node28867 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node28870 = (inp[11]) ? node28874 : node28871;
															assign node28871 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node28874 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node28877 = (inp[6]) ? node28885 : node28878;
														assign node28878 = (inp[11]) ? node28882 : node28879;
															assign node28879 = (inp[13]) ? 4'b0010 : 4'b1010;
															assign node28882 = (inp[13]) ? 4'b0010 : 4'b0010;
														assign node28885 = (inp[11]) ? node28889 : node28886;
															assign node28886 = (inp[13]) ? 4'b0010 : 4'b0010;
															assign node28889 = (inp[13]) ? 4'b0010 : 4'b1010;
										assign node28892 = (inp[15]) ? node28950 : node28893;
											assign node28893 = (inp[5]) ? node28925 : node28894;
												assign node28894 = (inp[13]) ? node28910 : node28895;
													assign node28895 = (inp[3]) ? node28903 : node28896;
														assign node28896 = (inp[6]) ? node28900 : node28897;
															assign node28897 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node28900 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node28903 = (inp[6]) ? node28907 : node28904;
															assign node28904 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node28907 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node28910 = (inp[6]) ? node28918 : node28911;
														assign node28911 = (inp[1]) ? node28915 : node28912;
															assign node28912 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node28915 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node28918 = (inp[3]) ? node28922 : node28919;
															assign node28919 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node28922 = (inp[11]) ? 4'b0000 : 4'b0000;
												assign node28925 = (inp[3]) ? node28939 : node28926;
													assign node28926 = (inp[13]) ? node28934 : node28927;
														assign node28927 = (inp[11]) ? node28931 : node28928;
															assign node28928 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node28931 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node28934 = (inp[11]) ? 4'b0000 : node28935;
															assign node28935 = (inp[6]) ? 4'b0000 : 4'b0000;
													assign node28939 = (inp[11]) ? node28945 : node28940;
														assign node28940 = (inp[6]) ? 4'b0010 : node28941;
															assign node28941 = (inp[1]) ? 4'b0010 : 4'b1010;
														assign node28945 = (inp[6]) ? 4'b1010 : node28946;
															assign node28946 = (inp[13]) ? 4'b0010 : 4'b0010;
											assign node28950 = (inp[5]) ? node28982 : node28951;
												assign node28951 = (inp[3]) ? node28967 : node28952;
													assign node28952 = (inp[1]) ? node28960 : node28953;
														assign node28953 = (inp[11]) ? node28957 : node28954;
															assign node28954 = (inp[6]) ? 4'b0010 : 4'b1010;
															assign node28957 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node28960 = (inp[6]) ? node28964 : node28961;
															assign node28961 = (inp[13]) ? 4'b0010 : 4'b0010;
															assign node28964 = (inp[11]) ? 4'b0010 : 4'b1010;
													assign node28967 = (inp[13]) ? node28975 : node28968;
														assign node28968 = (inp[6]) ? node28972 : node28969;
															assign node28969 = (inp[11]) ? 4'b0010 : 4'b1010;
															assign node28972 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node28975 = (inp[6]) ? node28979 : node28976;
															assign node28976 = (inp[1]) ? 4'b0010 : 4'b0010;
															assign node28979 = (inp[1]) ? 4'b0010 : 4'b0010;
												assign node28982 = (inp[3]) ? node28996 : node28983;
													assign node28983 = (inp[1]) ? node28991 : node28984;
														assign node28984 = (inp[11]) ? node28988 : node28985;
															assign node28985 = (inp[6]) ? 4'b0010 : 4'b1010;
															assign node28988 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node28991 = (inp[6]) ? 4'b1010 : node28992;
															assign node28992 = (inp[11]) ? 4'b0010 : 4'b0010;
													assign node28996 = (inp[11]) ? node29004 : node28997;
														assign node28997 = (inp[6]) ? node29001 : node28998;
															assign node28998 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node29001 = (inp[13]) ? 4'b0000 : 4'b0000;
														assign node29004 = (inp[6]) ? 4'b1000 : node29005;
															assign node29005 = (inp[1]) ? 4'b1000 : 4'b0000;
								assign node29009 = (inp[11]) ? node29163 : node29010;
									assign node29010 = (inp[6]) ? node29086 : node29011;
										assign node29011 = (inp[13]) ? node29035 : node29012;
											assign node29012 = (inp[15]) ? node29024 : node29013;
												assign node29013 = (inp[0]) ? node29019 : node29014;
													assign node29014 = (inp[5]) ? node29016 : 4'b1010;
														assign node29016 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node29019 = (inp[3]) ? node29021 : 4'b1000;
														assign node29021 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node29024 = (inp[0]) ? node29030 : node29025;
													assign node29025 = (inp[5]) ? node29027 : 4'b1000;
														assign node29027 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node29030 = (inp[5]) ? node29032 : 4'b1010;
														assign node29032 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node29035 = (inp[1]) ? node29063 : node29036;
												assign node29036 = (inp[14]) ? node29050 : node29037;
													assign node29037 = (inp[5]) ? node29045 : node29038;
														assign node29038 = (inp[0]) ? node29042 : node29039;
															assign node29039 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node29042 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node29045 = (inp[15]) ? 4'b1010 : node29046;
															assign node29046 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node29050 = (inp[3]) ? node29058 : node29051;
														assign node29051 = (inp[15]) ? node29055 : node29052;
															assign node29052 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node29055 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node29058 = (inp[5]) ? node29060 : 4'b1000;
															assign node29060 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node29063 = (inp[0]) ? node29075 : node29064;
													assign node29064 = (inp[15]) ? node29070 : node29065;
														assign node29065 = (inp[3]) ? node29067 : 4'b0010;
															assign node29067 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node29070 = (inp[5]) ? node29072 : 4'b0000;
															assign node29072 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node29075 = (inp[15]) ? node29081 : node29076;
														assign node29076 = (inp[3]) ? node29078 : 4'b0000;
															assign node29078 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node29081 = (inp[3]) ? node29083 : 4'b0010;
															assign node29083 = (inp[5]) ? 4'b0000 : 4'b0010;
										assign node29086 = (inp[1]) ? node29110 : node29087;
											assign node29087 = (inp[0]) ? node29099 : node29088;
												assign node29088 = (inp[15]) ? node29094 : node29089;
													assign node29089 = (inp[5]) ? node29091 : 4'b0010;
														assign node29091 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node29094 = (inp[3]) ? node29096 : 4'b0000;
														assign node29096 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node29099 = (inp[15]) ? node29105 : node29100;
													assign node29100 = (inp[5]) ? node29102 : 4'b0000;
														assign node29102 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node29105 = (inp[5]) ? node29107 : 4'b0010;
														assign node29107 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node29110 = (inp[13]) ? node29134 : node29111;
												assign node29111 = (inp[15]) ? node29123 : node29112;
													assign node29112 = (inp[0]) ? node29118 : node29113;
														assign node29113 = (inp[3]) ? node29115 : 4'b0010;
															assign node29115 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node29118 = (inp[5]) ? node29120 : 4'b0000;
															assign node29120 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node29123 = (inp[0]) ? node29129 : node29124;
														assign node29124 = (inp[3]) ? node29126 : 4'b0000;
															assign node29126 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node29129 = (inp[3]) ? node29131 : 4'b0010;
															assign node29131 = (inp[14]) ? 4'b0010 : 4'b0000;
												assign node29134 = (inp[3]) ? node29150 : node29135;
													assign node29135 = (inp[5]) ? node29143 : node29136;
														assign node29136 = (inp[15]) ? node29140 : node29137;
															assign node29137 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node29140 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node29143 = (inp[14]) ? node29147 : node29144;
															assign node29144 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node29147 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node29150 = (inp[15]) ? node29156 : node29151;
														assign node29151 = (inp[0]) ? 4'b1010 : node29152;
															assign node29152 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node29156 = (inp[0]) ? node29160 : node29157;
															assign node29157 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node29160 = (inp[5]) ? 4'b1000 : 4'b1010;
									assign node29163 = (inp[6]) ? node29239 : node29164;
										assign node29164 = (inp[1]) ? node29188 : node29165;
											assign node29165 = (inp[0]) ? node29177 : node29166;
												assign node29166 = (inp[15]) ? node29172 : node29167;
													assign node29167 = (inp[5]) ? node29169 : 4'b0010;
														assign node29169 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node29172 = (inp[3]) ? node29174 : 4'b0000;
														assign node29174 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node29177 = (inp[15]) ? node29183 : node29178;
													assign node29178 = (inp[3]) ? node29180 : 4'b0000;
														assign node29180 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node29183 = (inp[3]) ? node29185 : 4'b0010;
														assign node29185 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node29188 = (inp[13]) ? node29216 : node29189;
												assign node29189 = (inp[14]) ? node29203 : node29190;
													assign node29190 = (inp[15]) ? node29198 : node29191;
														assign node29191 = (inp[0]) ? node29195 : node29192;
															assign node29192 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node29195 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node29198 = (inp[0]) ? node29200 : 4'b0000;
															assign node29200 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node29203 = (inp[0]) ? node29211 : node29204;
														assign node29204 = (inp[15]) ? node29208 : node29205;
															assign node29205 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node29208 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node29211 = (inp[5]) ? node29213 : 4'b0010;
															assign node29213 = (inp[3]) ? 4'b0000 : 4'b0000;
												assign node29216 = (inp[0]) ? node29228 : node29217;
													assign node29217 = (inp[15]) ? node29223 : node29218;
														assign node29218 = (inp[5]) ? node29220 : 4'b1010;
															assign node29220 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node29223 = (inp[3]) ? node29225 : 4'b1000;
															assign node29225 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node29228 = (inp[15]) ? node29234 : node29229;
														assign node29229 = (inp[3]) ? node29231 : 4'b1000;
															assign node29231 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node29234 = (inp[5]) ? node29236 : 4'b1010;
															assign node29236 = (inp[3]) ? 4'b1000 : 4'b1010;
										assign node29239 = (inp[1]) ? node29263 : node29240;
											assign node29240 = (inp[0]) ? node29252 : node29241;
												assign node29241 = (inp[15]) ? node29247 : node29242;
													assign node29242 = (inp[3]) ? node29244 : 4'b1010;
														assign node29244 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node29247 = (inp[5]) ? node29249 : 4'b1000;
														assign node29249 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node29252 = (inp[15]) ? node29258 : node29253;
													assign node29253 = (inp[3]) ? node29255 : 4'b1000;
														assign node29255 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node29258 = (inp[5]) ? node29260 : 4'b1010;
														assign node29260 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node29263 = (inp[13]) ? node29285 : node29264;
												assign node29264 = (inp[5]) ? node29272 : node29265;
													assign node29265 = (inp[0]) ? node29269 : node29266;
														assign node29266 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node29269 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node29272 = (inp[3]) ? node29278 : node29273;
														assign node29273 = (inp[14]) ? 4'b1000 : node29274;
															assign node29274 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node29278 = (inp[14]) ? node29282 : node29279;
															assign node29279 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node29282 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node29285 = (inp[0]) ? node29297 : node29286;
													assign node29286 = (inp[15]) ? node29292 : node29287;
														assign node29287 = (inp[5]) ? node29289 : 4'b0010;
															assign node29289 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node29292 = (inp[5]) ? node29294 : 4'b0000;
															assign node29294 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node29297 = (inp[15]) ? node29303 : node29298;
														assign node29298 = (inp[5]) ? node29300 : 4'b0000;
															assign node29300 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node29303 = (inp[5]) ? node29305 : 4'b0010;
															assign node29305 = (inp[3]) ? 4'b0000 : 4'b0010;
							assign node29308 = (inp[2]) ? node29760 : node29309;
								assign node29309 = (inp[14]) ? node29549 : node29310;
									assign node29310 = (inp[1]) ? node29428 : node29311;
										assign node29311 = (inp[3]) ? node29365 : node29312;
											assign node29312 = (inp[11]) ? node29342 : node29313;
												assign node29313 = (inp[6]) ? node29327 : node29314;
													assign node29314 = (inp[13]) ? node29320 : node29315;
														assign node29315 = (inp[0]) ? node29317 : 4'b1010;
															assign node29317 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node29320 = (inp[0]) ? node29324 : node29321;
															assign node29321 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node29324 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node29327 = (inp[5]) ? node29335 : node29328;
														assign node29328 = (inp[15]) ? node29332 : node29329;
															assign node29329 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node29332 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node29335 = (inp[13]) ? node29339 : node29336;
															assign node29336 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node29339 = (inp[0]) ? 4'b0000 : 4'b0000;
												assign node29342 = (inp[6]) ? node29350 : node29343;
													assign node29343 = (inp[15]) ? node29347 : node29344;
														assign node29344 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node29347 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node29350 = (inp[13]) ? node29358 : node29351;
														assign node29351 = (inp[5]) ? node29355 : node29352;
															assign node29352 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node29355 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node29358 = (inp[5]) ? node29362 : node29359;
															assign node29359 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node29362 = (inp[15]) ? 4'b1000 : 4'b1000;
											assign node29365 = (inp[5]) ? node29397 : node29366;
												assign node29366 = (inp[15]) ? node29382 : node29367;
													assign node29367 = (inp[0]) ? node29375 : node29368;
														assign node29368 = (inp[13]) ? node29372 : node29369;
															assign node29369 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node29372 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node29375 = (inp[13]) ? node29379 : node29376;
															assign node29376 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node29379 = (inp[11]) ? 4'b0000 : 4'b0000;
													assign node29382 = (inp[0]) ? node29390 : node29383;
														assign node29383 = (inp[13]) ? node29387 : node29384;
															assign node29384 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node29387 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node29390 = (inp[13]) ? node29394 : node29391;
															assign node29391 = (inp[6]) ? 4'b0010 : 4'b1010;
															assign node29394 = (inp[6]) ? 4'b1010 : 4'b0010;
												assign node29397 = (inp[13]) ? node29413 : node29398;
													assign node29398 = (inp[6]) ? node29406 : node29399;
														assign node29399 = (inp[11]) ? node29403 : node29400;
															assign node29400 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node29403 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node29406 = (inp[11]) ? node29410 : node29407;
															assign node29407 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node29410 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node29413 = (inp[6]) ? node29421 : node29414;
														assign node29414 = (inp[11]) ? node29418 : node29415;
															assign node29415 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node29418 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node29421 = (inp[11]) ? node29425 : node29422;
															assign node29422 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node29425 = (inp[0]) ? 4'b1000 : 4'b1000;
										assign node29428 = (inp[15]) ? node29492 : node29429;
											assign node29429 = (inp[0]) ? node29461 : node29430;
												assign node29430 = (inp[5]) ? node29446 : node29431;
													assign node29431 = (inp[13]) ? node29439 : node29432;
														assign node29432 = (inp[3]) ? node29436 : node29433;
															assign node29433 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node29436 = (inp[11]) ? 4'b0010 : 4'b0010;
														assign node29439 = (inp[6]) ? node29443 : node29440;
															assign node29440 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node29443 = (inp[11]) ? 4'b0010 : 4'b1010;
													assign node29446 = (inp[3]) ? node29454 : node29447;
														assign node29447 = (inp[13]) ? node29451 : node29448;
															assign node29448 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node29451 = (inp[6]) ? 4'b0010 : 4'b1010;
														assign node29454 = (inp[11]) ? node29458 : node29455;
															assign node29455 = (inp[13]) ? 4'b0000 : 4'b0000;
															assign node29458 = (inp[13]) ? 4'b0000 : 4'b0000;
												assign node29461 = (inp[3]) ? node29477 : node29462;
													assign node29462 = (inp[5]) ? node29470 : node29463;
														assign node29463 = (inp[6]) ? node29467 : node29464;
															assign node29464 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node29467 = (inp[11]) ? 4'b0000 : 4'b0000;
														assign node29470 = (inp[6]) ? node29474 : node29471;
															assign node29471 = (inp[13]) ? 4'b0000 : 4'b0000;
															assign node29474 = (inp[13]) ? 4'b0000 : 4'b0000;
													assign node29477 = (inp[5]) ? node29485 : node29478;
														assign node29478 = (inp[11]) ? node29482 : node29479;
															assign node29479 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node29482 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node29485 = (inp[13]) ? node29489 : node29486;
															assign node29486 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node29489 = (inp[11]) ? 4'b0010 : 4'b0010;
											assign node29492 = (inp[0]) ? node29520 : node29493;
												assign node29493 = (inp[5]) ? node29507 : node29494;
													assign node29494 = (inp[13]) ? node29502 : node29495;
														assign node29495 = (inp[11]) ? node29499 : node29496;
															assign node29496 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node29499 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node29502 = (inp[3]) ? node29504 : 4'b0000;
															assign node29504 = (inp[6]) ? 4'b0000 : 4'b0000;
													assign node29507 = (inp[3]) ? node29513 : node29508;
														assign node29508 = (inp[11]) ? node29510 : 4'b1000;
															assign node29510 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node29513 = (inp[13]) ? node29517 : node29514;
															assign node29514 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node29517 = (inp[11]) ? 4'b0010 : 4'b0010;
												assign node29520 = (inp[5]) ? node29536 : node29521;
													assign node29521 = (inp[3]) ? node29529 : node29522;
														assign node29522 = (inp[11]) ? node29526 : node29523;
															assign node29523 = (inp[13]) ? 4'b0010 : 4'b0010;
															assign node29526 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node29529 = (inp[13]) ? node29533 : node29530;
															assign node29530 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node29533 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node29536 = (inp[3]) ? node29544 : node29537;
														assign node29537 = (inp[13]) ? node29541 : node29538;
															assign node29538 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node29541 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node29544 = (inp[6]) ? node29546 : 4'b0000;
															assign node29546 = (inp[11]) ? 4'b0000 : 4'b1000;
									assign node29549 = (inp[1]) ? node29659 : node29550;
										assign node29550 = (inp[0]) ? node29602 : node29551;
											assign node29551 = (inp[15]) ? node29579 : node29552;
												assign node29552 = (inp[3]) ? node29568 : node29553;
													assign node29553 = (inp[5]) ? node29561 : node29554;
														assign node29554 = (inp[13]) ? node29558 : node29555;
															assign node29555 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node29558 = (inp[6]) ? 4'b0011 : 4'b0011;
														assign node29561 = (inp[13]) ? node29565 : node29562;
															assign node29562 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node29565 = (inp[11]) ? 4'b0011 : 4'b0011;
													assign node29568 = (inp[5]) ? node29574 : node29569;
														assign node29569 = (inp[11]) ? node29571 : 4'b1011;
															assign node29571 = (inp[6]) ? 4'b0011 : 4'b0011;
														assign node29574 = (inp[11]) ? node29576 : 4'b1001;
															assign node29576 = (inp[13]) ? 4'b0001 : 4'b0001;
												assign node29579 = (inp[5]) ? node29589 : node29580;
													assign node29580 = (inp[11]) ? node29582 : 4'b1001;
														assign node29582 = (inp[3]) ? node29586 : node29583;
															assign node29583 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node29586 = (inp[13]) ? 4'b0001 : 4'b0001;
													assign node29589 = (inp[3]) ? node29595 : node29590;
														assign node29590 = (inp[6]) ? 4'b0001 : node29591;
															assign node29591 = (inp[11]) ? 4'b0001 : 4'b0001;
														assign node29595 = (inp[11]) ? node29599 : node29596;
															assign node29596 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node29599 = (inp[6]) ? 4'b0011 : 4'b0011;
											assign node29602 = (inp[15]) ? node29632 : node29603;
												assign node29603 = (inp[3]) ? node29617 : node29604;
													assign node29604 = (inp[5]) ? node29610 : node29605;
														assign node29605 = (inp[6]) ? 4'b0001 : node29606;
															assign node29606 = (inp[11]) ? 4'b0001 : 4'b0001;
														assign node29610 = (inp[11]) ? node29614 : node29611;
															assign node29611 = (inp[13]) ? 4'b0001 : 4'b0001;
															assign node29614 = (inp[6]) ? 4'b0001 : 4'b0001;
													assign node29617 = (inp[5]) ? node29625 : node29618;
														assign node29618 = (inp[11]) ? node29622 : node29619;
															assign node29619 = (inp[13]) ? 4'b0001 : 4'b0001;
															assign node29622 = (inp[6]) ? 4'b0001 : 4'b0001;
														assign node29625 = (inp[6]) ? node29629 : node29626;
															assign node29626 = (inp[13]) ? 4'b0011 : 4'b0011;
															assign node29629 = (inp[13]) ? 4'b0011 : 4'b0011;
												assign node29632 = (inp[3]) ? node29646 : node29633;
													assign node29633 = (inp[5]) ? node29639 : node29634;
														assign node29634 = (inp[13]) ? node29636 : 4'b0011;
															assign node29636 = (inp[11]) ? 4'b0011 : 4'b0011;
														assign node29639 = (inp[11]) ? node29643 : node29640;
															assign node29640 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node29643 = (inp[6]) ? 4'b0011 : 4'b0011;
													assign node29646 = (inp[5]) ? node29654 : node29647;
														assign node29647 = (inp[13]) ? node29651 : node29648;
															assign node29648 = (inp[11]) ? 4'b0011 : 4'b0011;
															assign node29651 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node29654 = (inp[13]) ? node29656 : 4'b1001;
															assign node29656 = (inp[6]) ? 4'b0001 : 4'b0001;
										assign node29659 = (inp[11]) ? node29707 : node29660;
											assign node29660 = (inp[6]) ? node29684 : node29661;
												assign node29661 = (inp[15]) ? node29673 : node29662;
													assign node29662 = (inp[0]) ? node29668 : node29663;
														assign node29663 = (inp[3]) ? node29665 : 4'b0011;
															assign node29665 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node29668 = (inp[3]) ? node29670 : 4'b0001;
															assign node29670 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node29673 = (inp[0]) ? node29679 : node29674;
														assign node29674 = (inp[3]) ? node29676 : 4'b0001;
															assign node29676 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node29679 = (inp[3]) ? node29681 : 4'b0011;
															assign node29681 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node29684 = (inp[15]) ? node29696 : node29685;
													assign node29685 = (inp[0]) ? node29691 : node29686;
														assign node29686 = (inp[5]) ? node29688 : 4'b1011;
															assign node29688 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node29691 = (inp[3]) ? node29693 : 4'b1001;
															assign node29693 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node29696 = (inp[0]) ? node29702 : node29697;
														assign node29697 = (inp[5]) ? node29699 : 4'b1001;
															assign node29699 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node29702 = (inp[5]) ? node29704 : 4'b1011;
															assign node29704 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node29707 = (inp[6]) ? node29731 : node29708;
												assign node29708 = (inp[13]) ? node29722 : node29709;
													assign node29709 = (inp[3]) ? node29717 : node29710;
														assign node29710 = (inp[5]) ? node29714 : node29711;
															assign node29711 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node29714 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node29717 = (inp[15]) ? node29719 : 4'b1001;
															assign node29719 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node29722 = (inp[3]) ? node29724 : 4'b1001;
														assign node29724 = (inp[0]) ? node29728 : node29725;
															assign node29725 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node29728 = (inp[5]) ? 4'b1001 : 4'b1001;
												assign node29731 = (inp[13]) ? node29745 : node29732;
													assign node29732 = (inp[15]) ? node29740 : node29733;
														assign node29733 = (inp[0]) ? node29737 : node29734;
															assign node29734 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node29737 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node29740 = (inp[0]) ? node29742 : 4'b0001;
															assign node29742 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node29745 = (inp[15]) ? node29753 : node29746;
														assign node29746 = (inp[0]) ? node29750 : node29747;
															assign node29747 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node29750 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node29753 = (inp[0]) ? node29757 : node29754;
															assign node29754 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node29757 = (inp[3]) ? 4'b0001 : 4'b0011;
								assign node29760 = (inp[14]) ? node29996 : node29761;
									assign node29761 = (inp[15]) ? node29873 : node29762;
										assign node29762 = (inp[0]) ? node29814 : node29763;
											assign node29763 = (inp[5]) ? node29785 : node29764;
												assign node29764 = (inp[1]) ? node29778 : node29765;
													assign node29765 = (inp[13]) ? node29771 : node29766;
														assign node29766 = (inp[6]) ? 4'b1011 : node29767;
															assign node29767 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node29771 = (inp[11]) ? node29775 : node29772;
															assign node29772 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node29775 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node29778 = (inp[6]) ? node29782 : node29779;
														assign node29779 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node29782 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node29785 = (inp[3]) ? node29801 : node29786;
													assign node29786 = (inp[11]) ? node29794 : node29787;
														assign node29787 = (inp[6]) ? node29791 : node29788;
															assign node29788 = (inp[1]) ? 4'b0011 : 4'b1011;
															assign node29791 = (inp[13]) ? 4'b1011 : 4'b0011;
														assign node29794 = (inp[6]) ? node29798 : node29795;
															assign node29795 = (inp[1]) ? 4'b1011 : 4'b0011;
															assign node29798 = (inp[1]) ? 4'b0011 : 4'b0011;
													assign node29801 = (inp[11]) ? node29809 : node29802;
														assign node29802 = (inp[6]) ? node29806 : node29803;
															assign node29803 = (inp[1]) ? 4'b0001 : 4'b0001;
															assign node29806 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node29809 = (inp[6]) ? node29811 : 4'b1001;
															assign node29811 = (inp[13]) ? 4'b0001 : 4'b1001;
											assign node29814 = (inp[3]) ? node29846 : node29815;
												assign node29815 = (inp[5]) ? node29831 : node29816;
													assign node29816 = (inp[11]) ? node29824 : node29817;
														assign node29817 = (inp[6]) ? node29821 : node29818;
															assign node29818 = (inp[13]) ? 4'b0001 : 4'b0001;
															assign node29821 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node29824 = (inp[6]) ? node29828 : node29825;
															assign node29825 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node29828 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node29831 = (inp[1]) ? node29839 : node29832;
														assign node29832 = (inp[13]) ? node29836 : node29833;
															assign node29833 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node29836 = (inp[11]) ? 4'b0001 : 4'b0001;
														assign node29839 = (inp[13]) ? node29843 : node29840;
															assign node29840 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node29843 = (inp[6]) ? 4'b0001 : 4'b0001;
												assign node29846 = (inp[5]) ? node29858 : node29847;
													assign node29847 = (inp[11]) ? node29853 : node29848;
														assign node29848 = (inp[6]) ? 4'b1001 : node29849;
															assign node29849 = (inp[1]) ? 4'b0001 : 4'b0001;
														assign node29853 = (inp[6]) ? 4'b0001 : node29854;
															assign node29854 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node29858 = (inp[6]) ? node29866 : node29859;
														assign node29859 = (inp[11]) ? node29863 : node29860;
															assign node29860 = (inp[13]) ? 4'b0011 : 4'b0011;
															assign node29863 = (inp[13]) ? 4'b1011 : 4'b0011;
														assign node29866 = (inp[11]) ? node29870 : node29867;
															assign node29867 = (inp[1]) ? 4'b1011 : 4'b0011;
															assign node29870 = (inp[13]) ? 4'b0011 : 4'b1011;
										assign node29873 = (inp[0]) ? node29937 : node29874;
											assign node29874 = (inp[3]) ? node29906 : node29875;
												assign node29875 = (inp[13]) ? node29891 : node29876;
													assign node29876 = (inp[1]) ? node29884 : node29877;
														assign node29877 = (inp[11]) ? node29881 : node29878;
															assign node29878 = (inp[6]) ? 4'b0001 : 4'b1001;
															assign node29881 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node29884 = (inp[5]) ? node29888 : node29885;
															assign node29885 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node29888 = (inp[11]) ? 4'b0001 : 4'b0001;
													assign node29891 = (inp[1]) ? node29899 : node29892;
														assign node29892 = (inp[6]) ? node29896 : node29893;
															assign node29893 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node29896 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node29899 = (inp[5]) ? node29903 : node29900;
															assign node29900 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node29903 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node29906 = (inp[5]) ? node29922 : node29907;
													assign node29907 = (inp[13]) ? node29915 : node29908;
														assign node29908 = (inp[11]) ? node29912 : node29909;
															assign node29909 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node29912 = (inp[6]) ? 4'b0001 : 4'b0001;
														assign node29915 = (inp[6]) ? node29919 : node29916;
															assign node29916 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node29919 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node29922 = (inp[13]) ? node29930 : node29923;
														assign node29923 = (inp[11]) ? node29927 : node29924;
															assign node29924 = (inp[1]) ? 4'b0011 : 4'b0011;
															assign node29927 = (inp[1]) ? 4'b0011 : 4'b0011;
														assign node29930 = (inp[11]) ? node29934 : node29931;
															assign node29931 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node29934 = (inp[6]) ? 4'b0011 : 4'b1011;
											assign node29937 = (inp[3]) ? node29967 : node29938;
												assign node29938 = (inp[13]) ? node29952 : node29939;
													assign node29939 = (inp[5]) ? node29945 : node29940;
														assign node29940 = (inp[11]) ? node29942 : 4'b0011;
															assign node29942 = (inp[1]) ? 4'b0011 : 4'b0011;
														assign node29945 = (inp[11]) ? node29949 : node29946;
															assign node29946 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node29949 = (inp[1]) ? 4'b0011 : 4'b0011;
													assign node29952 = (inp[1]) ? node29960 : node29953;
														assign node29953 = (inp[5]) ? node29957 : node29954;
															assign node29954 = (inp[11]) ? 4'b0011 : 4'b0011;
															assign node29957 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node29960 = (inp[11]) ? node29964 : node29961;
															assign node29961 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node29964 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node29967 = (inp[5]) ? node29983 : node29968;
													assign node29968 = (inp[1]) ? node29976 : node29969;
														assign node29969 = (inp[13]) ? node29973 : node29970;
															assign node29970 = (inp[11]) ? 4'b0011 : 4'b1011;
															assign node29973 = (inp[6]) ? 4'b0011 : 4'b0011;
														assign node29976 = (inp[11]) ? node29980 : node29977;
															assign node29977 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node29980 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node29983 = (inp[11]) ? node29989 : node29984;
														assign node29984 = (inp[6]) ? node29986 : 4'b0001;
															assign node29986 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node29989 = (inp[6]) ? node29993 : node29990;
															assign node29990 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node29993 = (inp[1]) ? 4'b0001 : 4'b0001;
									assign node29996 = (inp[13]) ? node30120 : node29997;
										assign node29997 = (inp[11]) ? node30059 : node29998;
											assign node29998 = (inp[3]) ? node30028 : node29999;
												assign node29999 = (inp[1]) ? node30013 : node30000;
													assign node30000 = (inp[6]) ? node30008 : node30001;
														assign node30001 = (inp[5]) ? node30005 : node30002;
															assign node30002 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node30005 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node30008 = (inp[15]) ? 4'b0011 : node30009;
															assign node30009 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node30013 = (inp[6]) ? node30021 : node30014;
														assign node30014 = (inp[15]) ? node30018 : node30015;
															assign node30015 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node30018 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node30021 = (inp[5]) ? node30025 : node30022;
															assign node30022 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node30025 = (inp[15]) ? 4'b1001 : 4'b1001;
												assign node30028 = (inp[5]) ? node30044 : node30029;
													assign node30029 = (inp[15]) ? node30037 : node30030;
														assign node30030 = (inp[0]) ? node30034 : node30031;
															assign node30031 = (inp[1]) ? 4'b0011 : 4'b0011;
															assign node30034 = (inp[6]) ? 4'b0001 : 4'b0001;
														assign node30037 = (inp[0]) ? node30041 : node30038;
															assign node30038 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node30041 = (inp[6]) ? 4'b0011 : 4'b0011;
													assign node30044 = (inp[1]) ? node30052 : node30045;
														assign node30045 = (inp[6]) ? node30049 : node30046;
															assign node30046 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node30049 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node30052 = (inp[6]) ? node30056 : node30053;
															assign node30053 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node30056 = (inp[15]) ? 4'b1001 : 4'b1001;
											assign node30059 = (inp[15]) ? node30091 : node30060;
												assign node30060 = (inp[0]) ? node30076 : node30061;
													assign node30061 = (inp[3]) ? node30069 : node30062;
														assign node30062 = (inp[1]) ? node30066 : node30063;
															assign node30063 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node30066 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node30069 = (inp[5]) ? node30073 : node30070;
															assign node30070 = (inp[6]) ? 4'b0011 : 4'b1011;
															assign node30073 = (inp[6]) ? 4'b0001 : 4'b0001;
													assign node30076 = (inp[5]) ? node30084 : node30077;
														assign node30077 = (inp[1]) ? node30081 : node30078;
															assign node30078 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node30081 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node30084 = (inp[3]) ? node30088 : node30085;
															assign node30085 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node30088 = (inp[6]) ? 4'b0011 : 4'b0011;
												assign node30091 = (inp[0]) ? node30105 : node30092;
													assign node30092 = (inp[3]) ? node30100 : node30093;
														assign node30093 = (inp[5]) ? node30097 : node30094;
															assign node30094 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node30097 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node30100 = (inp[5]) ? 4'b1011 : node30101;
															assign node30101 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node30105 = (inp[3]) ? node30113 : node30106;
														assign node30106 = (inp[1]) ? node30110 : node30107;
															assign node30107 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node30110 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node30113 = (inp[5]) ? node30117 : node30114;
															assign node30114 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node30117 = (inp[1]) ? 4'b0001 : 4'b0001;
										assign node30120 = (inp[15]) ? node30174 : node30121;
											assign node30121 = (inp[0]) ? node30151 : node30122;
												assign node30122 = (inp[3]) ? node30138 : node30123;
													assign node30123 = (inp[1]) ? node30131 : node30124;
														assign node30124 = (inp[6]) ? node30128 : node30125;
															assign node30125 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node30128 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node30131 = (inp[11]) ? node30135 : node30132;
															assign node30132 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node30135 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node30138 = (inp[5]) ? node30146 : node30139;
														assign node30139 = (inp[1]) ? node30143 : node30140;
															assign node30140 = (inp[11]) ? 4'b0011 : 4'b0011;
															assign node30143 = (inp[6]) ? 4'b0011 : 4'b0011;
														assign node30146 = (inp[1]) ? node30148 : 4'b0001;
															assign node30148 = (inp[11]) ? 4'b0001 : 4'b0001;
												assign node30151 = (inp[3]) ? node30161 : node30152;
													assign node30152 = (inp[1]) ? 4'b1001 : node30153;
														assign node30153 = (inp[6]) ? node30157 : node30154;
															assign node30154 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node30157 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node30161 = (inp[5]) ? node30167 : node30162;
														assign node30162 = (inp[6]) ? node30164 : 4'b1001;
															assign node30164 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node30167 = (inp[1]) ? node30171 : node30168;
															assign node30168 = (inp[11]) ? 4'b0011 : 4'b0011;
															assign node30171 = (inp[6]) ? 4'b0011 : 4'b0011;
											assign node30174 = (inp[0]) ? node30204 : node30175;
												assign node30175 = (inp[3]) ? node30191 : node30176;
													assign node30176 = (inp[5]) ? node30184 : node30177;
														assign node30177 = (inp[11]) ? node30181 : node30178;
															assign node30178 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node30181 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node30184 = (inp[11]) ? node30188 : node30185;
															assign node30185 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node30188 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node30191 = (inp[5]) ? node30197 : node30192;
														assign node30192 = (inp[11]) ? 4'b1001 : node30193;
															assign node30193 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node30197 = (inp[11]) ? node30201 : node30198;
															assign node30198 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node30201 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node30204 = (inp[5]) ? node30212 : node30205;
													assign node30205 = (inp[6]) ? node30209 : node30206;
														assign node30206 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node30209 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node30212 = (inp[3]) ? node30220 : node30213;
														assign node30213 = (inp[1]) ? node30217 : node30214;
															assign node30214 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node30217 = (inp[6]) ? 4'b0011 : 4'b0011;
														assign node30220 = (inp[11]) ? node30224 : node30221;
															assign node30221 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node30224 = (inp[6]) ? 4'b0001 : 4'b1001;
						assign node30227 = (inp[7]) ? node31079 : node30228;
							assign node30228 = (inp[14]) ? node30662 : node30229;
								assign node30229 = (inp[2]) ? node30439 : node30230;
									assign node30230 = (inp[13]) ? node30320 : node30231;
										assign node30231 = (inp[0]) ? node30279 : node30232;
											assign node30232 = (inp[15]) ? node30256 : node30233;
												assign node30233 = (inp[3]) ? node30241 : node30234;
													assign node30234 = (inp[11]) ? node30238 : node30235;
														assign node30235 = (inp[6]) ? 4'b0010 : 4'b1010;
														assign node30238 = (inp[6]) ? 4'b1010 : 4'b0010;
													assign node30241 = (inp[5]) ? node30249 : node30242;
														assign node30242 = (inp[1]) ? node30246 : node30243;
															assign node30243 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node30246 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node30249 = (inp[6]) ? node30253 : node30250;
															assign node30250 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node30253 = (inp[11]) ? 4'b1000 : 4'b0000;
												assign node30256 = (inp[5]) ? node30264 : node30257;
													assign node30257 = (inp[11]) ? node30261 : node30258;
														assign node30258 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node30261 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node30264 = (inp[3]) ? node30272 : node30265;
														assign node30265 = (inp[11]) ? node30269 : node30266;
															assign node30266 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node30269 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node30272 = (inp[6]) ? node30276 : node30273;
															assign node30273 = (inp[11]) ? 4'b0010 : 4'b1010;
															assign node30276 = (inp[11]) ? 4'b1010 : 4'b0010;
											assign node30279 = (inp[15]) ? node30299 : node30280;
												assign node30280 = (inp[5]) ? node30288 : node30281;
													assign node30281 = (inp[6]) ? node30285 : node30282;
														assign node30282 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node30285 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node30288 = (inp[3]) ? node30296 : node30289;
														assign node30289 = (inp[6]) ? node30293 : node30290;
															assign node30290 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node30293 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node30296 = (inp[11]) ? 4'b1010 : 4'b0010;
												assign node30299 = (inp[3]) ? node30307 : node30300;
													assign node30300 = (inp[6]) ? node30304 : node30301;
														assign node30301 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node30304 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node30307 = (inp[5]) ? node30315 : node30308;
														assign node30308 = (inp[1]) ? node30312 : node30309;
															assign node30309 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node30312 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node30315 = (inp[1]) ? node30317 : 4'b1000;
															assign node30317 = (inp[11]) ? 4'b0000 : 4'b0000;
										assign node30320 = (inp[11]) ? node30382 : node30321;
											assign node30321 = (inp[6]) ? node30353 : node30322;
												assign node30322 = (inp[1]) ? node30338 : node30323;
													assign node30323 = (inp[0]) ? node30331 : node30324;
														assign node30324 = (inp[15]) ? node30328 : node30325;
															assign node30325 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node30328 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node30331 = (inp[15]) ? node30335 : node30332;
															assign node30332 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node30335 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node30338 = (inp[15]) ? node30346 : node30339;
														assign node30339 = (inp[0]) ? node30343 : node30340;
															assign node30340 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node30343 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node30346 = (inp[0]) ? node30350 : node30347;
															assign node30347 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node30350 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node30353 = (inp[1]) ? node30367 : node30354;
													assign node30354 = (inp[3]) ? node30360 : node30355;
														assign node30355 = (inp[5]) ? node30357 : 4'b0000;
															assign node30357 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node30360 = (inp[0]) ? node30364 : node30361;
															assign node30361 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node30364 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node30367 = (inp[0]) ? node30375 : node30368;
														assign node30368 = (inp[15]) ? node30372 : node30369;
															assign node30369 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node30372 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node30375 = (inp[15]) ? node30379 : node30376;
															assign node30376 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node30379 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node30382 = (inp[6]) ? node30412 : node30383;
												assign node30383 = (inp[1]) ? node30397 : node30384;
													assign node30384 = (inp[3]) ? node30392 : node30385;
														assign node30385 = (inp[0]) ? node30389 : node30386;
															assign node30386 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node30389 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node30392 = (inp[5]) ? node30394 : 4'b0010;
															assign node30394 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node30397 = (inp[3]) ? node30405 : node30398;
														assign node30398 = (inp[15]) ? node30402 : node30399;
															assign node30399 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node30402 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node30405 = (inp[15]) ? node30409 : node30406;
															assign node30406 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node30409 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node30412 = (inp[1]) ? node30424 : node30413;
													assign node30413 = (inp[0]) ? node30419 : node30414;
														assign node30414 = (inp[15]) ? node30416 : 4'b1010;
															assign node30416 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node30419 = (inp[15]) ? 4'b1010 : node30420;
															assign node30420 = (inp[3]) ? 4'b1000 : 4'b1000;
													assign node30424 = (inp[0]) ? node30432 : node30425;
														assign node30425 = (inp[15]) ? node30429 : node30426;
															assign node30426 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node30429 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node30432 = (inp[15]) ? node30436 : node30433;
															assign node30433 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node30436 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node30439 = (inp[5]) ? node30537 : node30440;
										assign node30440 = (inp[0]) ? node30488 : node30441;
											assign node30441 = (inp[15]) ? node30465 : node30442;
												assign node30442 = (inp[1]) ? node30458 : node30443;
													assign node30443 = (inp[11]) ? node30451 : node30444;
														assign node30444 = (inp[6]) ? node30448 : node30445;
															assign node30445 = (inp[13]) ? 4'b0011 : 4'b1011;
															assign node30448 = (inp[13]) ? 4'b1011 : 4'b0011;
														assign node30451 = (inp[13]) ? node30455 : node30452;
															assign node30452 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node30455 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node30458 = (inp[11]) ? node30462 : node30459;
														assign node30459 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node30462 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node30465 = (inp[1]) ? node30481 : node30466;
													assign node30466 = (inp[6]) ? node30474 : node30467;
														assign node30467 = (inp[3]) ? node30471 : node30468;
															assign node30468 = (inp[11]) ? 4'b0001 : 4'b0001;
															assign node30471 = (inp[13]) ? 4'b0001 : 4'b0001;
														assign node30474 = (inp[11]) ? node30478 : node30475;
															assign node30475 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node30478 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node30481 = (inp[6]) ? node30485 : node30482;
														assign node30482 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node30485 = (inp[11]) ? 4'b0001 : 4'b1001;
											assign node30488 = (inp[15]) ? node30512 : node30489;
												assign node30489 = (inp[1]) ? node30505 : node30490;
													assign node30490 = (inp[11]) ? node30498 : node30491;
														assign node30491 = (inp[6]) ? node30495 : node30492;
															assign node30492 = (inp[13]) ? 4'b0001 : 4'b1001;
															assign node30495 = (inp[13]) ? 4'b1001 : 4'b0001;
														assign node30498 = (inp[6]) ? node30502 : node30499;
															assign node30499 = (inp[13]) ? 4'b1001 : 4'b0001;
															assign node30502 = (inp[13]) ? 4'b0001 : 4'b1001;
													assign node30505 = (inp[11]) ? node30509 : node30506;
														assign node30506 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node30509 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node30512 = (inp[3]) ? node30526 : node30513;
													assign node30513 = (inp[6]) ? node30521 : node30514;
														assign node30514 = (inp[11]) ? node30518 : node30515;
															assign node30515 = (inp[13]) ? 4'b0011 : 4'b0011;
															assign node30518 = (inp[1]) ? 4'b1011 : 4'b0011;
														assign node30521 = (inp[11]) ? node30523 : 4'b1011;
															assign node30523 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node30526 = (inp[1]) ? node30532 : node30527;
														assign node30527 = (inp[6]) ? 4'b1011 : node30528;
															assign node30528 = (inp[13]) ? 4'b0011 : 4'b0011;
														assign node30532 = (inp[6]) ? node30534 : 4'b1011;
															assign node30534 = (inp[11]) ? 4'b0011 : 4'b1011;
										assign node30537 = (inp[1]) ? node30601 : node30538;
											assign node30538 = (inp[6]) ? node30570 : node30539;
												assign node30539 = (inp[15]) ? node30555 : node30540;
													assign node30540 = (inp[11]) ? node30548 : node30541;
														assign node30541 = (inp[13]) ? node30545 : node30542;
															assign node30542 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node30545 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node30548 = (inp[13]) ? node30552 : node30549;
															assign node30549 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node30552 = (inp[3]) ? 4'b1001 : 4'b1001;
													assign node30555 = (inp[3]) ? node30563 : node30556;
														assign node30556 = (inp[0]) ? node30560 : node30557;
															assign node30557 = (inp[11]) ? 4'b0001 : 4'b0001;
															assign node30560 = (inp[13]) ? 4'b0011 : 4'b0011;
														assign node30563 = (inp[0]) ? node30567 : node30564;
															assign node30564 = (inp[13]) ? 4'b0011 : 4'b0011;
															assign node30567 = (inp[11]) ? 4'b0001 : 4'b0001;
												assign node30570 = (inp[15]) ? node30586 : node30571;
													assign node30571 = (inp[13]) ? node30579 : node30572;
														assign node30572 = (inp[11]) ? node30576 : node30573;
															assign node30573 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node30576 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node30579 = (inp[11]) ? node30583 : node30580;
															assign node30580 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node30583 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node30586 = (inp[13]) ? node30594 : node30587;
														assign node30587 = (inp[11]) ? node30591 : node30588;
															assign node30588 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node30591 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node30594 = (inp[11]) ? node30598 : node30595;
															assign node30595 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node30598 = (inp[3]) ? 4'b0001 : 4'b0001;
											assign node30601 = (inp[6]) ? node30633 : node30602;
												assign node30602 = (inp[11]) ? node30618 : node30603;
													assign node30603 = (inp[0]) ? node30611 : node30604;
														assign node30604 = (inp[3]) ? node30608 : node30605;
															assign node30605 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node30608 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node30611 = (inp[15]) ? node30615 : node30612;
															assign node30612 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node30615 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node30618 = (inp[15]) ? node30626 : node30619;
														assign node30619 = (inp[0]) ? node30623 : node30620;
															assign node30620 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node30623 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node30626 = (inp[0]) ? node30630 : node30627;
															assign node30627 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node30630 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node30633 = (inp[11]) ? node30649 : node30634;
													assign node30634 = (inp[0]) ? node30642 : node30635;
														assign node30635 = (inp[3]) ? node30639 : node30636;
															assign node30636 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node30639 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node30642 = (inp[15]) ? node30646 : node30643;
															assign node30643 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node30646 = (inp[13]) ? 4'b1011 : 4'b1001;
													assign node30649 = (inp[15]) ? node30655 : node30650;
														assign node30650 = (inp[0]) ? 4'b0001 : node30651;
															assign node30651 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node30655 = (inp[0]) ? node30659 : node30656;
															assign node30656 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node30659 = (inp[3]) ? 4'b0001 : 4'b0011;
								assign node30662 = (inp[13]) ? node30898 : node30663;
									assign node30663 = (inp[11]) ? node30781 : node30664;
										assign node30664 = (inp[5]) ? node30718 : node30665;
											assign node30665 = (inp[6]) ? node30689 : node30666;
												assign node30666 = (inp[1]) ? node30674 : node30667;
													assign node30667 = (inp[15]) ? node30671 : node30668;
														assign node30668 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node30671 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node30674 = (inp[3]) ? node30682 : node30675;
														assign node30675 = (inp[15]) ? node30679 : node30676;
															assign node30676 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node30679 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node30682 = (inp[0]) ? node30686 : node30683;
															assign node30683 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node30686 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node30689 = (inp[1]) ? node30705 : node30690;
													assign node30690 = (inp[3]) ? node30698 : node30691;
														assign node30691 = (inp[2]) ? node30695 : node30692;
															assign node30692 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node30695 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node30698 = (inp[0]) ? node30702 : node30699;
															assign node30699 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node30702 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node30705 = (inp[3]) ? node30711 : node30706;
														assign node30706 = (inp[0]) ? 4'b1011 : node30707;
															assign node30707 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node30711 = (inp[2]) ? node30715 : node30712;
															assign node30712 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node30715 = (inp[15]) ? 4'b1001 : 4'b1001;
											assign node30718 = (inp[6]) ? node30750 : node30719;
												assign node30719 = (inp[1]) ? node30735 : node30720;
													assign node30720 = (inp[3]) ? node30728 : node30721;
														assign node30721 = (inp[0]) ? node30725 : node30722;
															assign node30722 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node30725 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node30728 = (inp[15]) ? node30732 : node30729;
															assign node30729 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node30732 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node30735 = (inp[2]) ? node30743 : node30736;
														assign node30736 = (inp[0]) ? node30740 : node30737;
															assign node30737 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node30740 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node30743 = (inp[15]) ? node30747 : node30744;
															assign node30744 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node30747 = (inp[0]) ? 4'b0001 : 4'b0001;
												assign node30750 = (inp[1]) ? node30766 : node30751;
													assign node30751 = (inp[0]) ? node30759 : node30752;
														assign node30752 = (inp[3]) ? node30756 : node30753;
															assign node30753 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node30756 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node30759 = (inp[3]) ? node30763 : node30760;
															assign node30760 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node30763 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node30766 = (inp[0]) ? node30774 : node30767;
														assign node30767 = (inp[3]) ? node30771 : node30768;
															assign node30768 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node30771 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node30774 = (inp[2]) ? node30778 : node30775;
															assign node30775 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node30778 = (inp[3]) ? 4'b1001 : 4'b1001;
										assign node30781 = (inp[1]) ? node30843 : node30782;
											assign node30782 = (inp[6]) ? node30812 : node30783;
												assign node30783 = (inp[3]) ? node30799 : node30784;
													assign node30784 = (inp[5]) ? node30792 : node30785;
														assign node30785 = (inp[2]) ? node30789 : node30786;
															assign node30786 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node30789 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node30792 = (inp[15]) ? node30796 : node30793;
															assign node30793 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node30796 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node30799 = (inp[2]) ? node30805 : node30800;
														assign node30800 = (inp[15]) ? node30802 : 4'b0001;
															assign node30802 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node30805 = (inp[15]) ? node30809 : node30806;
															assign node30806 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node30809 = (inp[0]) ? 4'b0001 : 4'b0001;
												assign node30812 = (inp[2]) ? node30828 : node30813;
													assign node30813 = (inp[5]) ? node30821 : node30814;
														assign node30814 = (inp[3]) ? node30818 : node30815;
															assign node30815 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node30818 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node30821 = (inp[15]) ? node30825 : node30822;
															assign node30822 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node30825 = (inp[3]) ? 4'b1001 : 4'b1001;
													assign node30828 = (inp[15]) ? node30836 : node30829;
														assign node30829 = (inp[0]) ? node30833 : node30830;
															assign node30830 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node30833 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node30836 = (inp[0]) ? node30840 : node30837;
															assign node30837 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node30840 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node30843 = (inp[6]) ? node30875 : node30844;
												assign node30844 = (inp[2]) ? node30860 : node30845;
													assign node30845 = (inp[15]) ? node30853 : node30846;
														assign node30846 = (inp[0]) ? node30850 : node30847;
															assign node30847 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node30850 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node30853 = (inp[0]) ? node30857 : node30854;
															assign node30854 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node30857 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node30860 = (inp[5]) ? node30868 : node30861;
														assign node30861 = (inp[0]) ? node30865 : node30862;
															assign node30862 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node30865 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node30868 = (inp[0]) ? node30872 : node30869;
															assign node30869 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node30872 = (inp[3]) ? 4'b1001 : 4'b1001;
												assign node30875 = (inp[0]) ? node30887 : node30876;
													assign node30876 = (inp[15]) ? node30882 : node30877;
														assign node30877 = (inp[3]) ? node30879 : 4'b0011;
															assign node30879 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node30882 = (inp[5]) ? node30884 : 4'b0001;
															assign node30884 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node30887 = (inp[15]) ? node30893 : node30888;
														assign node30888 = (inp[3]) ? node30890 : 4'b0001;
															assign node30890 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node30893 = (inp[3]) ? node30895 : 4'b0011;
															assign node30895 = (inp[5]) ? 4'b0001 : 4'b0011;
									assign node30898 = (inp[0]) ? node30992 : node30899;
										assign node30899 = (inp[15]) ? node30939 : node30900;
											assign node30900 = (inp[5]) ? node30916 : node30901;
												assign node30901 = (inp[2]) ? node30909 : node30902;
													assign node30902 = (inp[6]) ? node30906 : node30903;
														assign node30903 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node30906 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node30909 = (inp[11]) ? node30913 : node30910;
														assign node30910 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node30913 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node30916 = (inp[3]) ? node30924 : node30917;
													assign node30917 = (inp[11]) ? node30921 : node30918;
														assign node30918 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node30921 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node30924 = (inp[2]) ? node30932 : node30925;
														assign node30925 = (inp[1]) ? node30929 : node30926;
															assign node30926 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node30929 = (inp[11]) ? 4'b0001 : 4'b0001;
														assign node30932 = (inp[1]) ? node30936 : node30933;
															assign node30933 = (inp[11]) ? 4'b0001 : 4'b0001;
															assign node30936 = (inp[6]) ? 4'b0001 : 4'b0001;
											assign node30939 = (inp[5]) ? node30969 : node30940;
												assign node30940 = (inp[3]) ? node30954 : node30941;
													assign node30941 = (inp[2]) ? node30949 : node30942;
														assign node30942 = (inp[1]) ? node30946 : node30943;
															assign node30943 = (inp[11]) ? 4'b0001 : 4'b0001;
															assign node30946 = (inp[6]) ? 4'b0001 : 4'b0001;
														assign node30949 = (inp[6]) ? 4'b1001 : node30950;
															assign node30950 = (inp[11]) ? 4'b1001 : 4'b0001;
													assign node30954 = (inp[2]) ? node30962 : node30955;
														assign node30955 = (inp[1]) ? node30959 : node30956;
															assign node30956 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node30959 = (inp[11]) ? 4'b0001 : 4'b0001;
														assign node30962 = (inp[11]) ? node30966 : node30963;
															assign node30963 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node30966 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node30969 = (inp[3]) ? node30977 : node30970;
													assign node30970 = (inp[11]) ? node30974 : node30971;
														assign node30971 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node30974 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node30977 = (inp[2]) ? node30985 : node30978;
														assign node30978 = (inp[1]) ? node30982 : node30979;
															assign node30979 = (inp[11]) ? 4'b0011 : 4'b0011;
															assign node30982 = (inp[11]) ? 4'b0011 : 4'b0011;
														assign node30985 = (inp[11]) ? node30989 : node30986;
															assign node30986 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node30989 = (inp[6]) ? 4'b0011 : 4'b1011;
										assign node30992 = (inp[15]) ? node31040 : node30993;
											assign node30993 = (inp[3]) ? node31017 : node30994;
												assign node30994 = (inp[2]) ? node31010 : node30995;
													assign node30995 = (inp[1]) ? node31003 : node30996;
														assign node30996 = (inp[11]) ? node31000 : node30997;
															assign node30997 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node31000 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node31003 = (inp[6]) ? node31007 : node31004;
															assign node31004 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node31007 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node31010 = (inp[11]) ? node31014 : node31011;
														assign node31011 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node31014 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node31017 = (inp[5]) ? node31033 : node31018;
													assign node31018 = (inp[2]) ? node31026 : node31019;
														assign node31019 = (inp[11]) ? node31023 : node31020;
															assign node31020 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node31023 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node31026 = (inp[1]) ? node31030 : node31027;
															assign node31027 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node31030 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node31033 = (inp[6]) ? node31037 : node31034;
														assign node31034 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node31037 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node31040 = (inp[3]) ? node31064 : node31041;
												assign node31041 = (inp[5]) ? node31049 : node31042;
													assign node31042 = (inp[11]) ? node31046 : node31043;
														assign node31043 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node31046 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node31049 = (inp[1]) ? node31057 : node31050;
														assign node31050 = (inp[11]) ? node31054 : node31051;
															assign node31051 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node31054 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node31057 = (inp[11]) ? node31061 : node31058;
															assign node31058 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node31061 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node31064 = (inp[5]) ? node31072 : node31065;
													assign node31065 = (inp[6]) ? node31069 : node31066;
														assign node31066 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node31069 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node31072 = (inp[6]) ? node31076 : node31073;
														assign node31073 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node31076 = (inp[11]) ? 4'b0001 : 4'b1001;
							assign node31079 = (inp[14]) ? node31513 : node31080;
								assign node31080 = (inp[2]) ? node31312 : node31081;
									assign node31081 = (inp[13]) ? node31203 : node31082;
										assign node31082 = (inp[1]) ? node31142 : node31083;
											assign node31083 = (inp[5]) ? node31111 : node31084;
												assign node31084 = (inp[11]) ? node31096 : node31085;
													assign node31085 = (inp[6]) ? node31091 : node31086;
														assign node31086 = (inp[3]) ? 4'b1001 : node31087;
															assign node31087 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node31091 = (inp[0]) ? 4'b0001 : node31092;
															assign node31092 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node31096 = (inp[6]) ? node31104 : node31097;
														assign node31097 = (inp[0]) ? node31101 : node31098;
															assign node31098 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node31101 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node31104 = (inp[15]) ? node31108 : node31105;
															assign node31105 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node31108 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node31111 = (inp[15]) ? node31127 : node31112;
													assign node31112 = (inp[3]) ? node31120 : node31113;
														assign node31113 = (inp[0]) ? node31117 : node31114;
															assign node31114 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node31117 = (inp[11]) ? 4'b0001 : 4'b0001;
														assign node31120 = (inp[0]) ? node31124 : node31121;
															assign node31121 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node31124 = (inp[11]) ? 4'b0011 : 4'b0011;
													assign node31127 = (inp[0]) ? node31135 : node31128;
														assign node31128 = (inp[3]) ? node31132 : node31129;
															assign node31129 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node31132 = (inp[6]) ? 4'b0011 : 4'b0011;
														assign node31135 = (inp[3]) ? node31139 : node31136;
															assign node31136 = (inp[11]) ? 4'b0011 : 4'b0011;
															assign node31139 = (inp[6]) ? 4'b0001 : 4'b0001;
											assign node31142 = (inp[6]) ? node31172 : node31143;
												assign node31143 = (inp[11]) ? node31157 : node31144;
													assign node31144 = (inp[3]) ? node31152 : node31145;
														assign node31145 = (inp[5]) ? node31149 : node31146;
															assign node31146 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node31149 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node31152 = (inp[5]) ? 4'b0011 : node31153;
															assign node31153 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node31157 = (inp[3]) ? node31165 : node31158;
														assign node31158 = (inp[5]) ? node31162 : node31159;
															assign node31159 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node31162 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node31165 = (inp[15]) ? node31169 : node31166;
															assign node31166 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node31169 = (inp[5]) ? 4'b1001 : 4'b1001;
												assign node31172 = (inp[11]) ? node31188 : node31173;
													assign node31173 = (inp[5]) ? node31181 : node31174;
														assign node31174 = (inp[15]) ? node31178 : node31175;
															assign node31175 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node31178 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node31181 = (inp[3]) ? node31185 : node31182;
															assign node31182 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node31185 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node31188 = (inp[0]) ? node31196 : node31189;
														assign node31189 = (inp[15]) ? node31193 : node31190;
															assign node31190 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node31193 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node31196 = (inp[15]) ? node31200 : node31197;
															assign node31197 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node31200 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node31203 = (inp[0]) ? node31257 : node31204;
											assign node31204 = (inp[15]) ? node31236 : node31205;
												assign node31205 = (inp[5]) ? node31221 : node31206;
													assign node31206 = (inp[1]) ? node31214 : node31207;
														assign node31207 = (inp[6]) ? node31211 : node31208;
															assign node31208 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node31211 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node31214 = (inp[6]) ? node31218 : node31215;
															assign node31215 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node31218 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node31221 = (inp[3]) ? node31229 : node31222;
														assign node31222 = (inp[6]) ? node31226 : node31223;
															assign node31223 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node31226 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node31229 = (inp[1]) ? node31233 : node31230;
															assign node31230 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node31233 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node31236 = (inp[3]) ? node31244 : node31237;
													assign node31237 = (inp[11]) ? node31241 : node31238;
														assign node31238 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node31241 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node31244 = (inp[5]) ? node31250 : node31245;
														assign node31245 = (inp[1]) ? node31247 : 4'b1001;
															assign node31247 = (inp[6]) ? 4'b0001 : 4'b0001;
														assign node31250 = (inp[1]) ? node31254 : node31251;
															assign node31251 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node31254 = (inp[11]) ? 4'b0011 : 4'b0011;
											assign node31257 = (inp[15]) ? node31289 : node31258;
												assign node31258 = (inp[5]) ? node31274 : node31259;
													assign node31259 = (inp[3]) ? node31267 : node31260;
														assign node31260 = (inp[1]) ? node31264 : node31261;
															assign node31261 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node31264 = (inp[6]) ? 4'b0001 : 4'b0001;
														assign node31267 = (inp[1]) ? node31271 : node31268;
															assign node31268 = (inp[11]) ? 4'b0001 : 4'b0001;
															assign node31271 = (inp[11]) ? 4'b0001 : 4'b0001;
													assign node31274 = (inp[3]) ? node31282 : node31275;
														assign node31275 = (inp[1]) ? node31279 : node31276;
															assign node31276 = (inp[11]) ? 4'b0001 : 4'b0001;
															assign node31279 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node31282 = (inp[6]) ? node31286 : node31283;
															assign node31283 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node31286 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node31289 = (inp[5]) ? node31297 : node31290;
													assign node31290 = (inp[6]) ? node31294 : node31291;
														assign node31291 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node31294 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node31297 = (inp[3]) ? node31305 : node31298;
														assign node31298 = (inp[1]) ? node31302 : node31299;
															assign node31299 = (inp[6]) ? 4'b0011 : 4'b1011;
															assign node31302 = (inp[11]) ? 4'b0011 : 4'b0011;
														assign node31305 = (inp[1]) ? node31309 : node31306;
															assign node31306 = (inp[11]) ? 4'b0001 : 4'b0001;
															assign node31309 = (inp[6]) ? 4'b1001 : 4'b0001;
									assign node31312 = (inp[0]) ? node31410 : node31313;
										assign node31313 = (inp[15]) ? node31365 : node31314;
											assign node31314 = (inp[5]) ? node31338 : node31315;
												assign node31315 = (inp[1]) ? node31331 : node31316;
													assign node31316 = (inp[6]) ? node31324 : node31317;
														assign node31317 = (inp[13]) ? node31321 : node31318;
															assign node31318 = (inp[11]) ? 4'b0010 : 4'b1010;
															assign node31321 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node31324 = (inp[3]) ? node31328 : node31325;
															assign node31325 = (inp[13]) ? 4'b0010 : 4'b0010;
															assign node31328 = (inp[13]) ? 4'b0010 : 4'b0010;
													assign node31331 = (inp[11]) ? node31335 : node31332;
														assign node31332 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node31335 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node31338 = (inp[3]) ? node31352 : node31339;
													assign node31339 = (inp[1]) ? node31345 : node31340;
														assign node31340 = (inp[13]) ? 4'b0010 : node31341;
															assign node31341 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node31345 = (inp[6]) ? node31349 : node31346;
															assign node31346 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node31349 = (inp[11]) ? 4'b0010 : 4'b1010;
													assign node31352 = (inp[13]) ? node31358 : node31353;
														assign node31353 = (inp[6]) ? node31355 : 4'b1000;
															assign node31355 = (inp[11]) ? 4'b0000 : 4'b0000;
														assign node31358 = (inp[1]) ? node31362 : node31359;
															assign node31359 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node31362 = (inp[6]) ? 4'b0000 : 4'b0000;
											assign node31365 = (inp[5]) ? node31389 : node31366;
												assign node31366 = (inp[6]) ? node31378 : node31367;
													assign node31367 = (inp[11]) ? node31373 : node31368;
														assign node31368 = (inp[1]) ? 4'b0000 : node31369;
															assign node31369 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node31373 = (inp[13]) ? 4'b1000 : node31374;
															assign node31374 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node31378 = (inp[11]) ? node31384 : node31379;
														assign node31379 = (inp[13]) ? 4'b1000 : node31380;
															assign node31380 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node31384 = (inp[1]) ? 4'b0000 : node31385;
															assign node31385 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node31389 = (inp[3]) ? node31401 : node31390;
													assign node31390 = (inp[11]) ? node31396 : node31391;
														assign node31391 = (inp[6]) ? 4'b1000 : node31392;
															assign node31392 = (inp[1]) ? 4'b0000 : 4'b0000;
														assign node31396 = (inp[1]) ? node31398 : 4'b0000;
															assign node31398 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node31401 = (inp[11]) ? node31405 : node31402;
														assign node31402 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node31405 = (inp[6]) ? node31407 : 4'b1010;
															assign node31407 = (inp[13]) ? 4'b0010 : 4'b0010;
										assign node31410 = (inp[15]) ? node31464 : node31411;
											assign node31411 = (inp[5]) ? node31435 : node31412;
												assign node31412 = (inp[11]) ? node31424 : node31413;
													assign node31413 = (inp[6]) ? node31419 : node31414;
														assign node31414 = (inp[13]) ? 4'b0000 : node31415;
															assign node31415 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node31419 = (inp[13]) ? 4'b1000 : node31420;
															assign node31420 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node31424 = (inp[6]) ? node31430 : node31425;
														assign node31425 = (inp[13]) ? 4'b1000 : node31426;
															assign node31426 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node31430 = (inp[13]) ? 4'b0000 : node31431;
															assign node31431 = (inp[1]) ? 4'b0000 : 4'b1000;
												assign node31435 = (inp[3]) ? node31449 : node31436;
													assign node31436 = (inp[13]) ? node31442 : node31437;
														assign node31437 = (inp[11]) ? node31439 : 4'b1000;
															assign node31439 = (inp[1]) ? 4'b0000 : 4'b0000;
														assign node31442 = (inp[1]) ? node31446 : node31443;
															assign node31443 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node31446 = (inp[11]) ? 4'b0000 : 4'b0000;
													assign node31449 = (inp[11]) ? node31457 : node31450;
														assign node31450 = (inp[6]) ? node31454 : node31451;
															assign node31451 = (inp[1]) ? 4'b0010 : 4'b0010;
															assign node31454 = (inp[13]) ? 4'b1010 : 4'b0010;
														assign node31457 = (inp[6]) ? node31461 : node31458;
															assign node31458 = (inp[13]) ? 4'b1010 : 4'b0010;
															assign node31461 = (inp[1]) ? 4'b0010 : 4'b0010;
											assign node31464 = (inp[3]) ? node31488 : node31465;
												assign node31465 = (inp[11]) ? node31477 : node31466;
													assign node31466 = (inp[6]) ? node31472 : node31467;
														assign node31467 = (inp[13]) ? 4'b0010 : node31468;
															assign node31468 = (inp[1]) ? 4'b0010 : 4'b1010;
														assign node31472 = (inp[1]) ? 4'b1010 : node31473;
															assign node31473 = (inp[13]) ? 4'b1010 : 4'b0010;
													assign node31477 = (inp[6]) ? node31483 : node31478;
														assign node31478 = (inp[13]) ? 4'b1010 : node31479;
															assign node31479 = (inp[1]) ? 4'b1010 : 4'b0010;
														assign node31483 = (inp[13]) ? 4'b0010 : node31484;
															assign node31484 = (inp[1]) ? 4'b0010 : 4'b1010;
												assign node31488 = (inp[5]) ? node31502 : node31489;
													assign node31489 = (inp[6]) ? node31497 : node31490;
														assign node31490 = (inp[11]) ? node31494 : node31491;
															assign node31491 = (inp[1]) ? 4'b0010 : 4'b0010;
															assign node31494 = (inp[13]) ? 4'b1010 : 4'b0010;
														assign node31497 = (inp[11]) ? node31499 : 4'b1010;
															assign node31499 = (inp[13]) ? 4'b0010 : 4'b0010;
													assign node31502 = (inp[11]) ? node31506 : node31503;
														assign node31503 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node31506 = (inp[6]) ? node31510 : node31507;
															assign node31507 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node31510 = (inp[13]) ? 4'b0000 : 4'b0000;
								assign node31513 = (inp[5]) ? node31749 : node31514;
									assign node31514 = (inp[13]) ? node31634 : node31515;
										assign node31515 = (inp[11]) ? node31579 : node31516;
											assign node31516 = (inp[3]) ? node31548 : node31517;
												assign node31517 = (inp[6]) ? node31533 : node31518;
													assign node31518 = (inp[1]) ? node31526 : node31519;
														assign node31519 = (inp[15]) ? node31523 : node31520;
															assign node31520 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node31523 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node31526 = (inp[0]) ? node31530 : node31527;
															assign node31527 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node31530 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node31533 = (inp[1]) ? node31541 : node31534;
														assign node31534 = (inp[0]) ? node31538 : node31535;
															assign node31535 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node31538 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node31541 = (inp[15]) ? node31545 : node31542;
															assign node31542 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node31545 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node31548 = (inp[1]) ? node31564 : node31549;
													assign node31549 = (inp[6]) ? node31557 : node31550;
														assign node31550 = (inp[15]) ? node31554 : node31551;
															assign node31551 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node31554 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node31557 = (inp[2]) ? node31561 : node31558;
															assign node31558 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node31561 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node31564 = (inp[6]) ? node31572 : node31565;
														assign node31565 = (inp[0]) ? node31569 : node31566;
															assign node31566 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node31569 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node31572 = (inp[15]) ? node31576 : node31573;
															assign node31573 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node31576 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node31579 = (inp[1]) ? node31611 : node31580;
												assign node31580 = (inp[6]) ? node31596 : node31581;
													assign node31581 = (inp[3]) ? node31589 : node31582;
														assign node31582 = (inp[0]) ? node31586 : node31583;
															assign node31583 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node31586 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node31589 = (inp[0]) ? node31593 : node31590;
															assign node31590 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node31593 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node31596 = (inp[2]) ? node31604 : node31597;
														assign node31597 = (inp[0]) ? node31601 : node31598;
															assign node31598 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node31601 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node31604 = (inp[3]) ? node31608 : node31605;
															assign node31605 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node31608 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node31611 = (inp[6]) ? node31627 : node31612;
													assign node31612 = (inp[2]) ? node31620 : node31613;
														assign node31613 = (inp[3]) ? node31617 : node31614;
															assign node31614 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node31617 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node31620 = (inp[3]) ? node31624 : node31621;
															assign node31621 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node31624 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node31627 = (inp[15]) ? node31631 : node31628;
														assign node31628 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node31631 = (inp[0]) ? 4'b0010 : 4'b0000;
										assign node31634 = (inp[3]) ? node31696 : node31635;
											assign node31635 = (inp[1]) ? node31667 : node31636;
												assign node31636 = (inp[0]) ? node31652 : node31637;
													assign node31637 = (inp[15]) ? node31645 : node31638;
														assign node31638 = (inp[6]) ? node31642 : node31639;
															assign node31639 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node31642 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node31645 = (inp[11]) ? node31649 : node31646;
															assign node31646 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node31649 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node31652 = (inp[15]) ? node31660 : node31653;
														assign node31653 = (inp[2]) ? node31657 : node31654;
															assign node31654 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node31657 = (inp[11]) ? 4'b0000 : 4'b0000;
														assign node31660 = (inp[6]) ? node31664 : node31661;
															assign node31661 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node31664 = (inp[11]) ? 4'b0010 : 4'b1010;
												assign node31667 = (inp[0]) ? node31681 : node31668;
													assign node31668 = (inp[15]) ? node31674 : node31669;
														assign node31669 = (inp[11]) ? 4'b1010 : node31670;
															assign node31670 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node31674 = (inp[2]) ? node31678 : node31675;
															assign node31675 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node31678 = (inp[11]) ? 4'b0000 : 4'b0000;
													assign node31681 = (inp[15]) ? node31689 : node31682;
														assign node31682 = (inp[11]) ? node31686 : node31683;
															assign node31683 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node31686 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node31689 = (inp[11]) ? node31693 : node31690;
															assign node31690 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node31693 = (inp[6]) ? 4'b0010 : 4'b1010;
											assign node31696 = (inp[0]) ? node31720 : node31697;
												assign node31697 = (inp[15]) ? node31713 : node31698;
													assign node31698 = (inp[2]) ? node31706 : node31699;
														assign node31699 = (inp[1]) ? node31703 : node31700;
															assign node31700 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node31703 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node31706 = (inp[1]) ? node31710 : node31707;
															assign node31707 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node31710 = (inp[6]) ? 4'b0010 : 4'b0010;
													assign node31713 = (inp[6]) ? node31717 : node31714;
														assign node31714 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node31717 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node31720 = (inp[15]) ? node31736 : node31721;
													assign node31721 = (inp[2]) ? node31729 : node31722;
														assign node31722 = (inp[6]) ? node31726 : node31723;
															assign node31723 = (inp[11]) ? 4'b1000 : 4'b0000;
															assign node31726 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node31729 = (inp[1]) ? node31733 : node31730;
															assign node31730 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node31733 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node31736 = (inp[1]) ? node31744 : node31737;
														assign node31737 = (inp[11]) ? node31741 : node31738;
															assign node31738 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node31741 = (inp[6]) ? 4'b0010 : 4'b1010;
														assign node31744 = (inp[2]) ? node31746 : 4'b1010;
															assign node31746 = (inp[6]) ? 4'b0010 : 4'b0010;
									assign node31749 = (inp[13]) ? node31871 : node31750;
										assign node31750 = (inp[15]) ? node31808 : node31751;
											assign node31751 = (inp[3]) ? node31777 : node31752;
												assign node31752 = (inp[0]) ? node31768 : node31753;
													assign node31753 = (inp[2]) ? node31761 : node31754;
														assign node31754 = (inp[6]) ? node31758 : node31755;
															assign node31755 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node31758 = (inp[1]) ? 4'b0010 : 4'b0010;
														assign node31761 = (inp[11]) ? node31765 : node31762;
															assign node31762 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node31765 = (inp[1]) ? 4'b0010 : 4'b0010;
													assign node31768 = (inp[2]) ? 4'b0000 : node31769;
														assign node31769 = (inp[11]) ? node31773 : node31770;
															assign node31770 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node31773 = (inp[6]) ? 4'b0000 : 4'b0000;
												assign node31777 = (inp[0]) ? node31793 : node31778;
													assign node31778 = (inp[6]) ? node31786 : node31779;
														assign node31779 = (inp[1]) ? node31783 : node31780;
															assign node31780 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node31783 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node31786 = (inp[11]) ? node31790 : node31787;
															assign node31787 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node31790 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node31793 = (inp[2]) ? node31801 : node31794;
														assign node31794 = (inp[1]) ? node31798 : node31795;
															assign node31795 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node31798 = (inp[11]) ? 4'b0010 : 4'b0010;
														assign node31801 = (inp[11]) ? node31805 : node31802;
															assign node31802 = (inp[1]) ? 4'b0010 : 4'b0010;
															assign node31805 = (inp[6]) ? 4'b0010 : 4'b0010;
											assign node31808 = (inp[0]) ? node31840 : node31809;
												assign node31809 = (inp[3]) ? node31825 : node31810;
													assign node31810 = (inp[1]) ? node31818 : node31811;
														assign node31811 = (inp[2]) ? node31815 : node31812;
															assign node31812 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node31815 = (inp[11]) ? 4'b0000 : 4'b0000;
														assign node31818 = (inp[2]) ? node31822 : node31819;
															assign node31819 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node31822 = (inp[11]) ? 4'b0000 : 4'b0000;
													assign node31825 = (inp[1]) ? node31833 : node31826;
														assign node31826 = (inp[6]) ? node31830 : node31827;
															assign node31827 = (inp[11]) ? 4'b0010 : 4'b1010;
															assign node31830 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node31833 = (inp[11]) ? node31837 : node31834;
															assign node31834 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node31837 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node31840 = (inp[3]) ? node31856 : node31841;
													assign node31841 = (inp[1]) ? node31849 : node31842;
														assign node31842 = (inp[6]) ? node31846 : node31843;
															assign node31843 = (inp[11]) ? 4'b0010 : 4'b1010;
															assign node31846 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node31849 = (inp[11]) ? node31853 : node31850;
															assign node31850 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node31853 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node31856 = (inp[11]) ? node31864 : node31857;
														assign node31857 = (inp[2]) ? node31861 : node31858;
															assign node31858 = (inp[1]) ? 4'b0000 : 4'b0000;
															assign node31861 = (inp[1]) ? 4'b0000 : 4'b0000;
														assign node31864 = (inp[2]) ? node31868 : node31865;
															assign node31865 = (inp[1]) ? 4'b0000 : 4'b0000;
															assign node31868 = (inp[1]) ? 4'b0000 : 4'b0000;
										assign node31871 = (inp[2]) ? node31935 : node31872;
											assign node31872 = (inp[0]) ? node31904 : node31873;
												assign node31873 = (inp[1]) ? node31889 : node31874;
													assign node31874 = (inp[3]) ? node31882 : node31875;
														assign node31875 = (inp[15]) ? node31879 : node31876;
															assign node31876 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node31879 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node31882 = (inp[15]) ? node31886 : node31883;
															assign node31883 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node31886 = (inp[6]) ? 4'b0010 : 4'b0010;
													assign node31889 = (inp[3]) ? node31897 : node31890;
														assign node31890 = (inp[15]) ? node31894 : node31891;
															assign node31891 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node31894 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node31897 = (inp[15]) ? node31901 : node31898;
															assign node31898 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node31901 = (inp[11]) ? 4'b0010 : 4'b0010;
												assign node31904 = (inp[1]) ? node31920 : node31905;
													assign node31905 = (inp[11]) ? node31913 : node31906;
														assign node31906 = (inp[6]) ? node31910 : node31907;
															assign node31907 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node31910 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node31913 = (inp[6]) ? node31917 : node31914;
															assign node31914 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node31917 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node31920 = (inp[15]) ? node31928 : node31921;
														assign node31921 = (inp[3]) ? node31925 : node31922;
															assign node31922 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node31925 = (inp[11]) ? 4'b0010 : 4'b0010;
														assign node31928 = (inp[3]) ? node31932 : node31929;
															assign node31929 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node31932 = (inp[6]) ? 4'b0000 : 4'b0000;
											assign node31935 = (inp[15]) ? node31965 : node31936;
												assign node31936 = (inp[11]) ? node31952 : node31937;
													assign node31937 = (inp[6]) ? node31945 : node31938;
														assign node31938 = (inp[1]) ? node31942 : node31939;
															assign node31939 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node31942 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node31945 = (inp[0]) ? node31949 : node31946;
															assign node31946 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node31949 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node31952 = (inp[6]) ? node31960 : node31953;
														assign node31953 = (inp[1]) ? node31957 : node31954;
															assign node31954 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node31957 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node31960 = (inp[1]) ? node31962 : 4'b0010;
															assign node31962 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node31965 = (inp[6]) ? node31981 : node31966;
													assign node31966 = (inp[11]) ? node31974 : node31967;
														assign node31967 = (inp[3]) ? node31971 : node31968;
															assign node31968 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node31971 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node31974 = (inp[3]) ? node31978 : node31975;
															assign node31975 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node31978 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node31981 = (inp[11]) ? node31989 : node31982;
														assign node31982 = (inp[3]) ? node31986 : node31983;
															assign node31983 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node31986 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node31989 = (inp[1]) ? node31993 : node31990;
															assign node31990 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node31993 = (inp[0]) ? 4'b0000 : 4'b0000;
					assign node31996 = (inp[11]) ? node33822 : node31997;
						assign node31997 = (inp[6]) ? node32879 : node31998;
							assign node31998 = (inp[13]) ? node32450 : node31999;
								assign node31999 = (inp[1]) ? node32227 : node32000;
									assign node32000 = (inp[7]) ? node32110 : node32001;
										assign node32001 = (inp[8]) ? node32051 : node32002;
											assign node32002 = (inp[2]) ? node32028 : node32003;
												assign node32003 = (inp[14]) ? node32017 : node32004;
													assign node32004 = (inp[5]) ? node32012 : node32005;
														assign node32005 = (inp[0]) ? node32009 : node32006;
															assign node32006 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node32009 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node32012 = (inp[0]) ? node32014 : 4'b1001;
															assign node32014 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node32017 = (inp[15]) ? node32023 : node32018;
														assign node32018 = (inp[0]) ? 4'b1000 : node32019;
															assign node32019 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node32023 = (inp[0]) ? 4'b1010 : node32024;
															assign node32024 = (inp[3]) ? 4'b1000 : 4'b1000;
												assign node32028 = (inp[0]) ? node32040 : node32029;
													assign node32029 = (inp[15]) ? node32035 : node32030;
														assign node32030 = (inp[3]) ? node32032 : 4'b1010;
															assign node32032 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node32035 = (inp[3]) ? node32037 : 4'b1000;
															assign node32037 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node32040 = (inp[15]) ? node32046 : node32041;
														assign node32041 = (inp[3]) ? node32043 : 4'b1000;
															assign node32043 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node32046 = (inp[3]) ? node32048 : 4'b1010;
															assign node32048 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node32051 = (inp[2]) ? node32081 : node32052;
												assign node32052 = (inp[14]) ? node32068 : node32053;
													assign node32053 = (inp[3]) ? node32061 : node32054;
														assign node32054 = (inp[0]) ? node32058 : node32055;
															assign node32055 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node32058 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node32061 = (inp[5]) ? node32065 : node32062;
															assign node32062 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node32065 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node32068 = (inp[3]) ? node32076 : node32069;
														assign node32069 = (inp[5]) ? node32073 : node32070;
															assign node32070 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node32073 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node32076 = (inp[0]) ? 4'b1001 : node32077;
															assign node32077 = (inp[15]) ? 4'b1001 : 4'b1001;
												assign node32081 = (inp[3]) ? node32095 : node32082;
													assign node32082 = (inp[5]) ? node32088 : node32083;
														assign node32083 = (inp[14]) ? node32085 : 4'b1001;
															assign node32085 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node32088 = (inp[14]) ? node32092 : node32089;
															assign node32089 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node32092 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node32095 = (inp[5]) ? node32103 : node32096;
														assign node32096 = (inp[15]) ? node32100 : node32097;
															assign node32097 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node32100 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node32103 = (inp[14]) ? node32107 : node32104;
															assign node32104 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node32107 = (inp[0]) ? 4'b1001 : 4'b1001;
										assign node32110 = (inp[8]) ? node32166 : node32111;
											assign node32111 = (inp[14]) ? node32143 : node32112;
												assign node32112 = (inp[2]) ? node32128 : node32113;
													assign node32113 = (inp[0]) ? node32121 : node32114;
														assign node32114 = (inp[15]) ? node32118 : node32115;
															assign node32115 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node32118 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node32121 = (inp[15]) ? node32125 : node32122;
															assign node32122 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node32125 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node32128 = (inp[15]) ? node32136 : node32129;
														assign node32129 = (inp[0]) ? node32133 : node32130;
															assign node32130 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node32133 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node32136 = (inp[0]) ? node32140 : node32137;
															assign node32137 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node32140 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node32143 = (inp[15]) ? node32155 : node32144;
													assign node32144 = (inp[0]) ? node32150 : node32145;
														assign node32145 = (inp[5]) ? node32147 : 4'b1011;
															assign node32147 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node32150 = (inp[5]) ? node32152 : 4'b1001;
															assign node32152 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node32155 = (inp[0]) ? node32161 : node32156;
														assign node32156 = (inp[3]) ? node32158 : 4'b1001;
															assign node32158 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node32161 = (inp[5]) ? node32163 : 4'b1011;
															assign node32163 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node32166 = (inp[14]) ? node32198 : node32167;
												assign node32167 = (inp[2]) ? node32183 : node32168;
													assign node32168 = (inp[5]) ? node32176 : node32169;
														assign node32169 = (inp[15]) ? node32173 : node32170;
															assign node32170 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node32173 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node32176 = (inp[15]) ? node32180 : node32177;
															assign node32177 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node32180 = (inp[3]) ? 4'b1001 : 4'b1001;
													assign node32183 = (inp[5]) ? node32191 : node32184;
														assign node32184 = (inp[15]) ? node32188 : node32185;
															assign node32185 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node32188 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node32191 = (inp[15]) ? node32195 : node32192;
															assign node32192 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node32195 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node32198 = (inp[5]) ? node32212 : node32199;
													assign node32199 = (inp[3]) ? node32205 : node32200;
														assign node32200 = (inp[2]) ? node32202 : 4'b1000;
															assign node32202 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node32205 = (inp[2]) ? node32209 : node32206;
															assign node32206 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node32209 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node32212 = (inp[15]) ? node32220 : node32213;
														assign node32213 = (inp[3]) ? node32217 : node32214;
															assign node32214 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node32217 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node32220 = (inp[0]) ? node32224 : node32221;
															assign node32221 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node32224 = (inp[3]) ? 4'b1000 : 4'b1010;
									assign node32227 = (inp[7]) ? node32333 : node32228;
										assign node32228 = (inp[8]) ? node32280 : node32229;
											assign node32229 = (inp[14]) ? node32261 : node32230;
												assign node32230 = (inp[2]) ? node32246 : node32231;
													assign node32231 = (inp[3]) ? node32239 : node32232;
														assign node32232 = (inp[5]) ? node32236 : node32233;
															assign node32233 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node32236 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node32239 = (inp[15]) ? node32243 : node32240;
															assign node32240 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node32243 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node32246 = (inp[15]) ? node32254 : node32247;
														assign node32247 = (inp[0]) ? node32251 : node32248;
															assign node32248 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node32251 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node32254 = (inp[0]) ? node32258 : node32255;
															assign node32255 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node32258 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node32261 = (inp[15]) ? node32273 : node32262;
													assign node32262 = (inp[0]) ? node32268 : node32263;
														assign node32263 = (inp[3]) ? node32265 : 4'b1010;
															assign node32265 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node32268 = (inp[3]) ? node32270 : 4'b1000;
															assign node32270 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node32273 = (inp[0]) ? 4'b1010 : node32274;
														assign node32274 = (inp[3]) ? node32276 : 4'b1000;
															assign node32276 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node32280 = (inp[14]) ? node32310 : node32281;
												assign node32281 = (inp[2]) ? node32297 : node32282;
													assign node32282 = (inp[5]) ? node32290 : node32283;
														assign node32283 = (inp[15]) ? node32287 : node32284;
															assign node32284 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node32287 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node32290 = (inp[0]) ? node32294 : node32291;
															assign node32291 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node32294 = (inp[3]) ? 4'b1000 : 4'b1000;
													assign node32297 = (inp[15]) ? node32303 : node32298;
														assign node32298 = (inp[3]) ? node32300 : 4'b0011;
															assign node32300 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node32303 = (inp[0]) ? node32307 : node32304;
															assign node32304 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node32307 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node32310 = (inp[15]) ? node32322 : node32311;
													assign node32311 = (inp[0]) ? node32317 : node32312;
														assign node32312 = (inp[3]) ? node32314 : 4'b0011;
															assign node32314 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node32317 = (inp[5]) ? node32319 : 4'b0001;
															assign node32319 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node32322 = (inp[0]) ? node32328 : node32323;
														assign node32323 = (inp[5]) ? node32325 : 4'b0001;
															assign node32325 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node32328 = (inp[5]) ? node32330 : 4'b0011;
															assign node32330 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node32333 = (inp[8]) ? node32391 : node32334;
											assign node32334 = (inp[14]) ? node32362 : node32335;
												assign node32335 = (inp[2]) ? node32351 : node32336;
													assign node32336 = (inp[5]) ? node32344 : node32337;
														assign node32337 = (inp[3]) ? node32341 : node32338;
															assign node32338 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node32341 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node32344 = (inp[0]) ? node32348 : node32345;
															assign node32345 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node32348 = (inp[3]) ? 4'b1000 : 4'b1000;
													assign node32351 = (inp[15]) ? node32355 : node32352;
														assign node32352 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node32355 = (inp[0]) ? node32359 : node32356;
															assign node32356 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node32359 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node32362 = (inp[2]) ? node32376 : node32363;
													assign node32363 = (inp[3]) ? node32369 : node32364;
														assign node32364 = (inp[5]) ? 4'b0001 : node32365;
															assign node32365 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node32369 = (inp[5]) ? node32373 : node32370;
															assign node32370 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node32373 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node32376 = (inp[3]) ? node32384 : node32377;
														assign node32377 = (inp[0]) ? node32381 : node32378;
															assign node32378 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node32381 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node32384 = (inp[0]) ? node32388 : node32385;
															assign node32385 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node32388 = (inp[15]) ? 4'b0001 : 4'b0001;
											assign node32391 = (inp[2]) ? node32421 : node32392;
												assign node32392 = (inp[14]) ? node32408 : node32393;
													assign node32393 = (inp[5]) ? node32401 : node32394;
														assign node32394 = (inp[0]) ? node32398 : node32395;
															assign node32395 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node32398 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node32401 = (inp[3]) ? node32405 : node32402;
															assign node32402 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node32405 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node32408 = (inp[0]) ? node32414 : node32409;
														assign node32409 = (inp[15]) ? node32411 : 4'b0010;
															assign node32411 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node32414 = (inp[15]) ? node32418 : node32415;
															assign node32415 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node32418 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node32421 = (inp[3]) ? node32435 : node32422;
													assign node32422 = (inp[5]) ? node32430 : node32423;
														assign node32423 = (inp[14]) ? node32427 : node32424;
															assign node32424 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node32427 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node32430 = (inp[14]) ? 4'b0000 : node32431;
															assign node32431 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node32435 = (inp[5]) ? node32443 : node32436;
														assign node32436 = (inp[14]) ? node32440 : node32437;
															assign node32437 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node32440 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node32443 = (inp[15]) ? node32447 : node32444;
															assign node32444 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node32447 = (inp[0]) ? 4'b0000 : 4'b0010;
								assign node32450 = (inp[1]) ? node32666 : node32451;
									assign node32451 = (inp[7]) ? node32559 : node32452;
										assign node32452 = (inp[8]) ? node32506 : node32453;
											assign node32453 = (inp[2]) ? node32483 : node32454;
												assign node32454 = (inp[14]) ? node32470 : node32455;
													assign node32455 = (inp[0]) ? node32463 : node32456;
														assign node32456 = (inp[15]) ? node32460 : node32457;
															assign node32457 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node32460 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node32463 = (inp[15]) ? node32467 : node32464;
															assign node32464 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node32467 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node32470 = (inp[5]) ? node32478 : node32471;
														assign node32471 = (inp[15]) ? node32475 : node32472;
															assign node32472 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node32475 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node32478 = (inp[15]) ? 4'b1010 : node32479;
															assign node32479 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node32483 = (inp[0]) ? node32495 : node32484;
													assign node32484 = (inp[15]) ? node32490 : node32485;
														assign node32485 = (inp[5]) ? node32487 : 4'b1010;
															assign node32487 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node32490 = (inp[5]) ? node32492 : 4'b1000;
															assign node32492 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node32495 = (inp[15]) ? node32501 : node32496;
														assign node32496 = (inp[5]) ? node32498 : 4'b1000;
															assign node32498 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node32501 = (inp[3]) ? node32503 : 4'b1010;
															assign node32503 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node32506 = (inp[2]) ? node32538 : node32507;
												assign node32507 = (inp[14]) ? node32523 : node32508;
													assign node32508 = (inp[5]) ? node32516 : node32509;
														assign node32509 = (inp[3]) ? node32513 : node32510;
															assign node32510 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node32513 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node32516 = (inp[15]) ? node32520 : node32517;
															assign node32517 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node32520 = (inp[3]) ? 4'b1000 : 4'b1000;
													assign node32523 = (inp[5]) ? node32531 : node32524;
														assign node32524 = (inp[3]) ? node32528 : node32525;
															assign node32525 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node32528 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node32531 = (inp[15]) ? node32535 : node32532;
															assign node32532 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node32535 = (inp[0]) ? 4'b0001 : 4'b0001;
												assign node32538 = (inp[5]) ? node32546 : node32539;
													assign node32539 = (inp[15]) ? node32543 : node32540;
														assign node32540 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node32543 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node32546 = (inp[0]) ? node32552 : node32547;
														assign node32547 = (inp[15]) ? node32549 : 4'b0011;
															assign node32549 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node32552 = (inp[3]) ? node32556 : node32553;
															assign node32553 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node32556 = (inp[15]) ? 4'b0001 : 4'b0011;
										assign node32559 = (inp[8]) ? node32613 : node32560;
											assign node32560 = (inp[2]) ? node32590 : node32561;
												assign node32561 = (inp[14]) ? node32577 : node32562;
													assign node32562 = (inp[3]) ? node32570 : node32563;
														assign node32563 = (inp[15]) ? node32567 : node32564;
															assign node32564 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node32567 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node32570 = (inp[5]) ? node32574 : node32571;
															assign node32571 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node32574 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node32577 = (inp[3]) ? node32585 : node32578;
														assign node32578 = (inp[5]) ? node32582 : node32579;
															assign node32579 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node32582 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node32585 = (inp[5]) ? 4'b0001 : node32586;
															assign node32586 = (inp[0]) ? 4'b0001 : 4'b0001;
												assign node32590 = (inp[5]) ? node32598 : node32591;
													assign node32591 = (inp[0]) ? node32595 : node32592;
														assign node32592 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node32595 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node32598 = (inp[0]) ? node32606 : node32599;
														assign node32599 = (inp[3]) ? node32603 : node32600;
															assign node32600 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node32603 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node32606 = (inp[15]) ? node32610 : node32607;
															assign node32607 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node32610 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node32613 = (inp[14]) ? node32643 : node32614;
												assign node32614 = (inp[2]) ? node32630 : node32615;
													assign node32615 = (inp[0]) ? node32623 : node32616;
														assign node32616 = (inp[15]) ? node32620 : node32617;
															assign node32617 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node32620 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node32623 = (inp[15]) ? node32627 : node32624;
															assign node32624 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node32627 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node32630 = (inp[15]) ? node32636 : node32631;
														assign node32631 = (inp[0]) ? node32633 : 4'b0010;
															assign node32633 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node32636 = (inp[0]) ? node32640 : node32637;
															assign node32637 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node32640 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node32643 = (inp[0]) ? node32655 : node32644;
													assign node32644 = (inp[15]) ? node32650 : node32645;
														assign node32645 = (inp[5]) ? node32647 : 4'b0010;
															assign node32647 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node32650 = (inp[3]) ? node32652 : 4'b0000;
															assign node32652 = (inp[2]) ? 4'b0000 : 4'b0010;
													assign node32655 = (inp[15]) ? node32661 : node32656;
														assign node32656 = (inp[5]) ? node32658 : 4'b0000;
															assign node32658 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node32661 = (inp[5]) ? node32663 : 4'b0010;
															assign node32663 = (inp[3]) ? 4'b0000 : 4'b0010;
									assign node32666 = (inp[7]) ? node32776 : node32667;
										assign node32667 = (inp[8]) ? node32723 : node32668;
											assign node32668 = (inp[14]) ? node32700 : node32669;
												assign node32669 = (inp[2]) ? node32685 : node32670;
													assign node32670 = (inp[0]) ? node32678 : node32671;
														assign node32671 = (inp[15]) ? node32675 : node32672;
															assign node32672 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node32675 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node32678 = (inp[15]) ? node32682 : node32679;
															assign node32679 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node32682 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node32685 = (inp[15]) ? node32693 : node32686;
														assign node32686 = (inp[0]) ? node32690 : node32687;
															assign node32687 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node32690 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node32693 = (inp[0]) ? node32697 : node32694;
															assign node32694 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node32697 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node32700 = (inp[15]) ? node32712 : node32701;
													assign node32701 = (inp[0]) ? node32707 : node32702;
														assign node32702 = (inp[3]) ? node32704 : 4'b0010;
															assign node32704 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node32707 = (inp[5]) ? node32709 : 4'b0000;
															assign node32709 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node32712 = (inp[0]) ? node32718 : node32713;
														assign node32713 = (inp[3]) ? node32715 : 4'b0000;
															assign node32715 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node32718 = (inp[3]) ? node32720 : 4'b0010;
															assign node32720 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node32723 = (inp[2]) ? node32753 : node32724;
												assign node32724 = (inp[14]) ? node32740 : node32725;
													assign node32725 = (inp[3]) ? node32733 : node32726;
														assign node32726 = (inp[15]) ? node32730 : node32727;
															assign node32727 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node32730 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node32733 = (inp[0]) ? node32737 : node32734;
															assign node32734 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node32737 = (inp[5]) ? 4'b0000 : 4'b0000;
													assign node32740 = (inp[0]) ? node32746 : node32741;
														assign node32741 = (inp[15]) ? node32743 : 4'b0011;
															assign node32743 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node32746 = (inp[15]) ? node32750 : node32747;
															assign node32747 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node32750 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node32753 = (inp[5]) ? node32761 : node32754;
													assign node32754 = (inp[0]) ? node32758 : node32755;
														assign node32755 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node32758 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node32761 = (inp[15]) ? node32769 : node32762;
														assign node32762 = (inp[3]) ? node32766 : node32763;
															assign node32763 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node32766 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node32769 = (inp[0]) ? node32773 : node32770;
															assign node32770 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node32773 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node32776 = (inp[8]) ? node32830 : node32777;
											assign node32777 = (inp[2]) ? node32807 : node32778;
												assign node32778 = (inp[14]) ? node32792 : node32779;
													assign node32779 = (inp[15]) ? node32787 : node32780;
														assign node32780 = (inp[0]) ? node32784 : node32781;
															assign node32781 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node32784 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node32787 = (inp[3]) ? node32789 : 4'b0000;
															assign node32789 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node32792 = (inp[0]) ? node32800 : node32793;
														assign node32793 = (inp[15]) ? node32797 : node32794;
															assign node32794 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node32797 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node32800 = (inp[15]) ? node32804 : node32801;
															assign node32801 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node32804 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node32807 = (inp[15]) ? node32819 : node32808;
													assign node32808 = (inp[0]) ? node32814 : node32809;
														assign node32809 = (inp[5]) ? node32811 : 4'b0011;
															assign node32811 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node32814 = (inp[5]) ? node32816 : 4'b0001;
															assign node32816 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node32819 = (inp[0]) ? node32825 : node32820;
														assign node32820 = (inp[5]) ? node32822 : 4'b0001;
															assign node32822 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node32825 = (inp[3]) ? node32827 : 4'b0011;
															assign node32827 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node32830 = (inp[2]) ? node32856 : node32831;
												assign node32831 = (inp[14]) ? node32845 : node32832;
													assign node32832 = (inp[0]) ? node32838 : node32833;
														assign node32833 = (inp[15]) ? 4'b0001 : node32834;
															assign node32834 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node32838 = (inp[15]) ? node32842 : node32839;
															assign node32839 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node32842 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node32845 = (inp[15]) ? node32851 : node32846;
														assign node32846 = (inp[0]) ? 4'b0000 : node32847;
															assign node32847 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node32851 = (inp[0]) ? 4'b0010 : node32852;
															assign node32852 = (inp[3]) ? 4'b0000 : 4'b0000;
												assign node32856 = (inp[0]) ? node32868 : node32857;
													assign node32857 = (inp[15]) ? node32863 : node32858;
														assign node32858 = (inp[3]) ? node32860 : 4'b0010;
															assign node32860 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node32863 = (inp[5]) ? node32865 : 4'b0000;
															assign node32865 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node32868 = (inp[15]) ? node32874 : node32869;
														assign node32869 = (inp[3]) ? node32871 : 4'b0000;
															assign node32871 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node32874 = (inp[5]) ? node32876 : 4'b0010;
															assign node32876 = (inp[3]) ? 4'b0000 : 4'b0010;
							assign node32879 = (inp[13]) ? node33353 : node32880;
								assign node32880 = (inp[1]) ? node33122 : node32881;
									assign node32881 = (inp[5]) ? node32999 : node32882;
										assign node32882 = (inp[7]) ? node32946 : node32883;
											assign node32883 = (inp[8]) ? node32915 : node32884;
												assign node32884 = (inp[2]) ? node32900 : node32885;
													assign node32885 = (inp[14]) ? node32893 : node32886;
														assign node32886 = (inp[0]) ? node32890 : node32887;
															assign node32887 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node32890 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node32893 = (inp[0]) ? node32897 : node32894;
															assign node32894 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node32897 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node32900 = (inp[3]) ? node32908 : node32901;
														assign node32901 = (inp[15]) ? node32905 : node32902;
															assign node32902 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node32905 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node32908 = (inp[14]) ? node32912 : node32909;
															assign node32909 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node32912 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node32915 = (inp[14]) ? node32931 : node32916;
													assign node32916 = (inp[2]) ? node32924 : node32917;
														assign node32917 = (inp[15]) ? node32921 : node32918;
															assign node32918 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node32921 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node32924 = (inp[0]) ? node32928 : node32925;
															assign node32925 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node32928 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node32931 = (inp[2]) ? node32939 : node32932;
														assign node32932 = (inp[0]) ? node32936 : node32933;
															assign node32933 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node32936 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node32939 = (inp[15]) ? node32943 : node32940;
															assign node32940 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node32943 = (inp[0]) ? 4'b0011 : 4'b0001;
											assign node32946 = (inp[8]) ? node32976 : node32947;
												assign node32947 = (inp[2]) ? node32961 : node32948;
													assign node32948 = (inp[14]) ? node32956 : node32949;
														assign node32949 = (inp[3]) ? node32953 : node32950;
															assign node32950 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node32953 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node32956 = (inp[0]) ? 4'b0001 : node32957;
															assign node32957 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node32961 = (inp[3]) ? node32969 : node32962;
														assign node32962 = (inp[15]) ? node32966 : node32963;
															assign node32963 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node32966 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node32969 = (inp[15]) ? node32973 : node32970;
															assign node32970 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node32973 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node32976 = (inp[2]) ? node32992 : node32977;
													assign node32977 = (inp[14]) ? node32985 : node32978;
														assign node32978 = (inp[15]) ? node32982 : node32979;
															assign node32979 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node32982 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node32985 = (inp[15]) ? node32989 : node32986;
															assign node32986 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node32989 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node32992 = (inp[0]) ? node32996 : node32993;
														assign node32993 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node32996 = (inp[15]) ? 4'b0010 : 4'b0000;
										assign node32999 = (inp[3]) ? node33063 : node33000;
											assign node33000 = (inp[15]) ? node33032 : node33001;
												assign node33001 = (inp[0]) ? node33017 : node33002;
													assign node33002 = (inp[8]) ? node33010 : node33003;
														assign node33003 = (inp[7]) ? node33007 : node33004;
															assign node33004 = (inp[14]) ? 4'b0010 : 4'b0010;
															assign node33007 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node33010 = (inp[7]) ? node33014 : node33011;
															assign node33011 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node33014 = (inp[2]) ? 4'b0010 : 4'b0010;
													assign node33017 = (inp[8]) ? node33025 : node33018;
														assign node33018 = (inp[7]) ? node33022 : node33019;
															assign node33019 = (inp[2]) ? 4'b0000 : 4'b0000;
															assign node33022 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node33025 = (inp[7]) ? node33029 : node33026;
															assign node33026 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node33029 = (inp[2]) ? 4'b0000 : 4'b0000;
												assign node33032 = (inp[0]) ? node33048 : node33033;
													assign node33033 = (inp[2]) ? node33041 : node33034;
														assign node33034 = (inp[8]) ? node33038 : node33035;
															assign node33035 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node33038 = (inp[7]) ? 4'b0000 : 4'b0000;
														assign node33041 = (inp[14]) ? node33045 : node33042;
															assign node33042 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node33045 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node33048 = (inp[2]) ? node33056 : node33049;
														assign node33049 = (inp[8]) ? node33053 : node33050;
															assign node33050 = (inp[14]) ? 4'b0010 : 4'b0010;
															assign node33053 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node33056 = (inp[7]) ? node33060 : node33057;
															assign node33057 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node33060 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node33063 = (inp[2]) ? node33095 : node33064;
												assign node33064 = (inp[14]) ? node33080 : node33065;
													assign node33065 = (inp[15]) ? node33073 : node33066;
														assign node33066 = (inp[0]) ? node33070 : node33067;
															assign node33067 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node33070 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node33073 = (inp[0]) ? node33077 : node33074;
															assign node33074 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node33077 = (inp[8]) ? 4'b0000 : 4'b0000;
													assign node33080 = (inp[0]) ? node33088 : node33081;
														assign node33081 = (inp[15]) ? node33085 : node33082;
															assign node33082 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node33085 = (inp[8]) ? 4'b0010 : 4'b0010;
														assign node33088 = (inp[15]) ? node33092 : node33089;
															assign node33089 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node33092 = (inp[8]) ? 4'b0000 : 4'b0000;
												assign node33095 = (inp[0]) ? node33109 : node33096;
													assign node33096 = (inp[15]) ? node33102 : node33097;
														assign node33097 = (inp[8]) ? node33099 : 4'b0000;
															assign node33099 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node33102 = (inp[7]) ? node33106 : node33103;
															assign node33103 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node33106 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node33109 = (inp[15]) ? node33117 : node33110;
														assign node33110 = (inp[14]) ? node33114 : node33111;
															assign node33111 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node33114 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node33117 = (inp[8]) ? node33119 : 4'b0001;
															assign node33119 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node33122 = (inp[8]) ? node33244 : node33123;
										assign node33123 = (inp[7]) ? node33185 : node33124;
											assign node33124 = (inp[14]) ? node33154 : node33125;
												assign node33125 = (inp[2]) ? node33139 : node33126;
													assign node33126 = (inp[0]) ? node33134 : node33127;
														assign node33127 = (inp[15]) ? node33131 : node33128;
															assign node33128 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node33131 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node33134 = (inp[15]) ? node33136 : 4'b0001;
															assign node33136 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node33139 = (inp[15]) ? node33147 : node33140;
														assign node33140 = (inp[0]) ? node33144 : node33141;
															assign node33141 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node33144 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node33147 = (inp[0]) ? node33151 : node33148;
															assign node33148 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node33151 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node33154 = (inp[2]) ? node33170 : node33155;
													assign node33155 = (inp[3]) ? node33163 : node33156;
														assign node33156 = (inp[5]) ? node33160 : node33157;
															assign node33157 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node33160 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node33163 = (inp[5]) ? node33167 : node33164;
															assign node33164 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node33167 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node33170 = (inp[0]) ? node33178 : node33171;
														assign node33171 = (inp[15]) ? node33175 : node33172;
															assign node33172 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node33175 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node33178 = (inp[15]) ? node33182 : node33179;
															assign node33179 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node33182 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node33185 = (inp[14]) ? node33215 : node33186;
												assign node33186 = (inp[2]) ? node33202 : node33187;
													assign node33187 = (inp[3]) ? node33195 : node33188;
														assign node33188 = (inp[15]) ? node33192 : node33189;
															assign node33189 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node33192 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node33195 = (inp[15]) ? node33199 : node33196;
															assign node33196 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node33199 = (inp[5]) ? 4'b0000 : 4'b0000;
													assign node33202 = (inp[0]) ? node33208 : node33203;
														assign node33203 = (inp[15]) ? 4'b1111 : node33204;
															assign node33204 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node33208 = (inp[15]) ? node33212 : node33209;
															assign node33209 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node33212 = (inp[3]) ? 4'b1101 : 4'b1101;
												assign node33215 = (inp[2]) ? node33231 : node33216;
													assign node33216 = (inp[15]) ? node33224 : node33217;
														assign node33217 = (inp[0]) ? node33221 : node33218;
															assign node33218 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node33221 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node33224 = (inp[0]) ? node33228 : node33225;
															assign node33225 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node33228 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node33231 = (inp[0]) ? node33237 : node33232;
														assign node33232 = (inp[3]) ? 4'b1111 : node33233;
															assign node33233 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node33237 = (inp[15]) ? node33241 : node33238;
															assign node33238 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node33241 = (inp[5]) ? 4'b1101 : 4'b1101;
										assign node33244 = (inp[7]) ? node33302 : node33245;
											assign node33245 = (inp[2]) ? node33273 : node33246;
												assign node33246 = (inp[14]) ? node33260 : node33247;
													assign node33247 = (inp[15]) ? node33253 : node33248;
														assign node33248 = (inp[0]) ? 4'b0000 : node33249;
															assign node33249 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node33253 = (inp[0]) ? node33257 : node33254;
															assign node33254 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node33257 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node33260 = (inp[15]) ? node33268 : node33261;
														assign node33261 = (inp[0]) ? node33265 : node33262;
															assign node33262 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node33265 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node33268 = (inp[0]) ? 4'b1101 : node33269;
															assign node33269 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node33273 = (inp[3]) ? node33287 : node33274;
													assign node33274 = (inp[5]) ? node33280 : node33275;
														assign node33275 = (inp[14]) ? 4'b1111 : node33276;
															assign node33276 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node33280 = (inp[14]) ? node33284 : node33281;
															assign node33281 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node33284 = (inp[0]) ? 4'b1101 : 4'b1101;
													assign node33287 = (inp[14]) ? node33295 : node33288;
														assign node33288 = (inp[0]) ? node33292 : node33289;
															assign node33289 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node33292 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node33295 = (inp[5]) ? node33299 : node33296;
															assign node33296 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node33299 = (inp[0]) ? 4'b1101 : 4'b1101;
											assign node33302 = (inp[14]) ? node33330 : node33303;
												assign node33303 = (inp[2]) ? node33317 : node33304;
													assign node33304 = (inp[5]) ? node33310 : node33305;
														assign node33305 = (inp[3]) ? 4'b1111 : node33306;
															assign node33306 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node33310 = (inp[0]) ? node33314 : node33311;
															assign node33311 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node33314 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node33317 = (inp[3]) ? node33323 : node33318;
														assign node33318 = (inp[15]) ? node33320 : 4'b1100;
															assign node33320 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node33323 = (inp[5]) ? node33327 : node33324;
															assign node33324 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node33327 = (inp[0]) ? 4'b1100 : 4'b1100;
												assign node33330 = (inp[0]) ? node33342 : node33331;
													assign node33331 = (inp[15]) ? node33337 : node33332;
														assign node33332 = (inp[5]) ? 4'b1100 : node33333;
															assign node33333 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node33337 = (inp[5]) ? 4'b1110 : node33338;
															assign node33338 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node33342 = (inp[15]) ? node33348 : node33343;
														assign node33343 = (inp[3]) ? 4'b1110 : node33344;
															assign node33344 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node33348 = (inp[3]) ? 4'b1100 : node33349;
															assign node33349 = (inp[5]) ? 4'b1100 : 4'b1110;
								assign node33353 = (inp[1]) ? node33591 : node33354;
									assign node33354 = (inp[7]) ? node33470 : node33355;
										assign node33355 = (inp[8]) ? node33407 : node33356;
											assign node33356 = (inp[14]) ? node33384 : node33357;
												assign node33357 = (inp[2]) ? node33373 : node33358;
													assign node33358 = (inp[3]) ? node33366 : node33359;
														assign node33359 = (inp[5]) ? node33363 : node33360;
															assign node33360 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node33363 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node33366 = (inp[15]) ? node33370 : node33367;
															assign node33367 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node33370 = (inp[5]) ? 4'b0001 : 4'b0001;
													assign node33373 = (inp[0]) ? node33379 : node33374;
														assign node33374 = (inp[15]) ? node33376 : 4'b0010;
															assign node33376 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node33379 = (inp[5]) ? node33381 : 4'b0000;
															assign node33381 = (inp[3]) ? 4'b0000 : 4'b0000;
												assign node33384 = (inp[15]) ? node33396 : node33385;
													assign node33385 = (inp[0]) ? node33391 : node33386;
														assign node33386 = (inp[3]) ? node33388 : 4'b0010;
															assign node33388 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node33391 = (inp[3]) ? node33393 : 4'b0000;
															assign node33393 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node33396 = (inp[0]) ? node33402 : node33397;
														assign node33397 = (inp[5]) ? node33399 : 4'b0000;
															assign node33399 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node33402 = (inp[3]) ? node33404 : 4'b0010;
															assign node33404 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node33407 = (inp[14]) ? node33439 : node33408;
												assign node33408 = (inp[2]) ? node33424 : node33409;
													assign node33409 = (inp[3]) ? node33417 : node33410;
														assign node33410 = (inp[15]) ? node33414 : node33411;
															assign node33411 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node33414 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node33417 = (inp[5]) ? node33421 : node33418;
															assign node33418 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node33421 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node33424 = (inp[5]) ? node33432 : node33425;
														assign node33425 = (inp[3]) ? node33429 : node33426;
															assign node33426 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node33429 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node33432 = (inp[3]) ? node33436 : node33433;
															assign node33433 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node33436 = (inp[15]) ? 4'b1101 : 4'b1101;
												assign node33439 = (inp[2]) ? node33455 : node33440;
													assign node33440 = (inp[15]) ? node33448 : node33441;
														assign node33441 = (inp[0]) ? node33445 : node33442;
															assign node33442 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node33445 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node33448 = (inp[0]) ? node33452 : node33449;
															assign node33449 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node33452 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node33455 = (inp[5]) ? node33463 : node33456;
														assign node33456 = (inp[0]) ? node33460 : node33457;
															assign node33457 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node33460 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node33463 = (inp[0]) ? node33467 : node33464;
															assign node33464 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node33467 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node33470 = (inp[8]) ? node33528 : node33471;
											assign node33471 = (inp[14]) ? node33497 : node33472;
												assign node33472 = (inp[2]) ? node33484 : node33473;
													assign node33473 = (inp[15]) ? node33479 : node33474;
														assign node33474 = (inp[0]) ? node33476 : 4'b0010;
															assign node33476 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node33479 = (inp[0]) ? node33481 : 4'b0000;
															assign node33481 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node33484 = (inp[0]) ? node33490 : node33485;
														assign node33485 = (inp[15]) ? 4'b1111 : node33486;
															assign node33486 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node33490 = (inp[15]) ? node33494 : node33491;
															assign node33491 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node33494 = (inp[3]) ? 4'b1101 : 4'b1101;
												assign node33497 = (inp[5]) ? node33513 : node33498;
													assign node33498 = (inp[2]) ? node33506 : node33499;
														assign node33499 = (inp[15]) ? node33503 : node33500;
															assign node33500 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node33503 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node33506 = (inp[0]) ? node33510 : node33507;
															assign node33507 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node33510 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node33513 = (inp[3]) ? node33521 : node33514;
														assign node33514 = (inp[0]) ? node33518 : node33515;
															assign node33515 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node33518 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node33521 = (inp[0]) ? node33525 : node33522;
															assign node33522 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node33525 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node33528 = (inp[14]) ? node33560 : node33529;
												assign node33529 = (inp[2]) ? node33545 : node33530;
													assign node33530 = (inp[5]) ? node33538 : node33531;
														assign node33531 = (inp[0]) ? node33535 : node33532;
															assign node33532 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node33535 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node33538 = (inp[0]) ? node33542 : node33539;
															assign node33539 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node33542 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node33545 = (inp[0]) ? node33553 : node33546;
														assign node33546 = (inp[15]) ? node33550 : node33547;
															assign node33547 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node33550 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node33553 = (inp[15]) ? node33557 : node33554;
															assign node33554 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node33557 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node33560 = (inp[3]) ? node33576 : node33561;
													assign node33561 = (inp[0]) ? node33569 : node33562;
														assign node33562 = (inp[2]) ? node33566 : node33563;
															assign node33563 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node33566 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node33569 = (inp[15]) ? node33573 : node33570;
															assign node33570 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node33573 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node33576 = (inp[2]) ? node33584 : node33577;
														assign node33577 = (inp[15]) ? node33581 : node33578;
															assign node33578 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node33581 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node33584 = (inp[0]) ? node33588 : node33585;
															assign node33585 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node33588 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node33591 = (inp[8]) ? node33711 : node33592;
										assign node33592 = (inp[7]) ? node33652 : node33593;
											assign node33593 = (inp[14]) ? node33623 : node33594;
												assign node33594 = (inp[2]) ? node33608 : node33595;
													assign node33595 = (inp[3]) ? node33603 : node33596;
														assign node33596 = (inp[15]) ? node33600 : node33597;
															assign node33597 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node33600 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node33603 = (inp[15]) ? node33605 : 4'b1101;
															assign node33605 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node33608 = (inp[3]) ? node33616 : node33609;
														assign node33609 = (inp[15]) ? node33613 : node33610;
															assign node33610 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node33613 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node33616 = (inp[0]) ? node33620 : node33617;
															assign node33617 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node33620 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node33623 = (inp[2]) ? node33639 : node33624;
													assign node33624 = (inp[3]) ? node33632 : node33625;
														assign node33625 = (inp[0]) ? node33629 : node33626;
															assign node33626 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node33629 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node33632 = (inp[5]) ? node33636 : node33633;
															assign node33633 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node33636 = (inp[0]) ? 4'b1100 : 4'b1100;
													assign node33639 = (inp[15]) ? node33647 : node33640;
														assign node33640 = (inp[0]) ? node33644 : node33641;
															assign node33641 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node33644 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node33647 = (inp[5]) ? 4'b1110 : node33648;
															assign node33648 = (inp[3]) ? 4'b1110 : 4'b1100;
											assign node33652 = (inp[14]) ? node33680 : node33653;
												assign node33653 = (inp[2]) ? node33667 : node33654;
													assign node33654 = (inp[3]) ? node33662 : node33655;
														assign node33655 = (inp[5]) ? node33659 : node33656;
															assign node33656 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node33659 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node33662 = (inp[15]) ? 4'b1100 : node33663;
															assign node33663 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node33667 = (inp[15]) ? node33673 : node33668;
														assign node33668 = (inp[3]) ? 4'b1101 : node33669;
															assign node33669 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node33673 = (inp[0]) ? node33677 : node33674;
															assign node33674 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node33677 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node33680 = (inp[5]) ? node33696 : node33681;
													assign node33681 = (inp[15]) ? node33689 : node33682;
														assign node33682 = (inp[3]) ? node33686 : node33683;
															assign node33683 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node33686 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node33689 = (inp[2]) ? node33693 : node33690;
															assign node33690 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node33693 = (inp[0]) ? 4'b1101 : 4'b1101;
													assign node33696 = (inp[2]) ? node33704 : node33697;
														assign node33697 = (inp[0]) ? node33701 : node33698;
															assign node33698 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node33701 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node33704 = (inp[3]) ? node33708 : node33705;
															assign node33705 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node33708 = (inp[15]) ? 4'b1101 : 4'b1101;
										assign node33711 = (inp[7]) ? node33769 : node33712;
											assign node33712 = (inp[14]) ? node33742 : node33713;
												assign node33713 = (inp[2]) ? node33727 : node33714;
													assign node33714 = (inp[15]) ? node33722 : node33715;
														assign node33715 = (inp[0]) ? node33719 : node33716;
															assign node33716 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node33719 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node33722 = (inp[0]) ? node33724 : 4'b1110;
															assign node33724 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node33727 = (inp[5]) ? node33735 : node33728;
														assign node33728 = (inp[3]) ? node33732 : node33729;
															assign node33729 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node33732 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node33735 = (inp[3]) ? node33739 : node33736;
															assign node33736 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node33739 = (inp[0]) ? 4'b1101 : 4'b1101;
												assign node33742 = (inp[2]) ? node33756 : node33743;
													assign node33743 = (inp[0]) ? node33751 : node33744;
														assign node33744 = (inp[15]) ? node33748 : node33745;
															assign node33745 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node33748 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node33751 = (inp[15]) ? node33753 : 4'b1111;
															assign node33753 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node33756 = (inp[0]) ? node33764 : node33757;
														assign node33757 = (inp[15]) ? node33761 : node33758;
															assign node33758 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node33761 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node33764 = (inp[15]) ? node33766 : 4'b1111;
															assign node33766 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node33769 = (inp[14]) ? node33799 : node33770;
												assign node33770 = (inp[2]) ? node33786 : node33771;
													assign node33771 = (inp[0]) ? node33779 : node33772;
														assign node33772 = (inp[15]) ? node33776 : node33773;
															assign node33773 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node33776 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node33779 = (inp[15]) ? node33783 : node33780;
															assign node33780 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node33783 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node33786 = (inp[5]) ? node33792 : node33787;
														assign node33787 = (inp[15]) ? 4'b1110 : node33788;
															assign node33788 = (inp[3]) ? 4'b1100 : 4'b1100;
														assign node33792 = (inp[15]) ? node33796 : node33793;
															assign node33793 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node33796 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node33799 = (inp[3]) ? node33815 : node33800;
													assign node33800 = (inp[15]) ? node33808 : node33801;
														assign node33801 = (inp[0]) ? node33805 : node33802;
															assign node33802 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node33805 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node33808 = (inp[5]) ? node33812 : node33809;
															assign node33809 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node33812 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node33815 = (inp[15]) ? node33819 : node33816;
														assign node33816 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node33819 = (inp[0]) ? 4'b1100 : 4'b1110;
						assign node33822 = (inp[6]) ? node34712 : node33823;
							assign node33823 = (inp[1]) ? node34263 : node33824;
								assign node33824 = (inp[13]) ? node34054 : node33825;
									assign node33825 = (inp[2]) ? node33945 : node33826;
										assign node33826 = (inp[8]) ? node33888 : node33827;
											assign node33827 = (inp[5]) ? node33857 : node33828;
												assign node33828 = (inp[15]) ? node33844 : node33829;
													assign node33829 = (inp[0]) ? node33837 : node33830;
														assign node33830 = (inp[3]) ? node33834 : node33831;
															assign node33831 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node33834 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node33837 = (inp[7]) ? node33841 : node33838;
															assign node33838 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node33841 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node33844 = (inp[0]) ? node33852 : node33845;
														assign node33845 = (inp[3]) ? node33849 : node33846;
															assign node33846 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node33849 = (inp[14]) ? 4'b0000 : 4'b0000;
														assign node33852 = (inp[3]) ? 4'b0010 : node33853;
															assign node33853 = (inp[7]) ? 4'b0010 : 4'b0010;
												assign node33857 = (inp[15]) ? node33873 : node33858;
													assign node33858 = (inp[7]) ? node33866 : node33859;
														assign node33859 = (inp[14]) ? node33863 : node33860;
															assign node33860 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node33863 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node33866 = (inp[14]) ? node33870 : node33867;
															assign node33867 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node33870 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node33873 = (inp[0]) ? node33881 : node33874;
														assign node33874 = (inp[3]) ? node33878 : node33875;
															assign node33875 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node33878 = (inp[14]) ? 4'b0010 : 4'b0010;
														assign node33881 = (inp[3]) ? node33885 : node33882;
															assign node33882 = (inp[14]) ? 4'b0010 : 4'b0010;
															assign node33885 = (inp[14]) ? 4'b0000 : 4'b0001;
											assign node33888 = (inp[15]) ? node33920 : node33889;
												assign node33889 = (inp[0]) ? node33905 : node33890;
													assign node33890 = (inp[5]) ? node33898 : node33891;
														assign node33891 = (inp[3]) ? node33895 : node33892;
															assign node33892 = (inp[14]) ? 4'b0010 : 4'b0010;
															assign node33895 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node33898 = (inp[3]) ? node33902 : node33899;
															assign node33899 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node33902 = (inp[14]) ? 4'b0000 : 4'b0000;
													assign node33905 = (inp[3]) ? node33913 : node33906;
														assign node33906 = (inp[7]) ? node33910 : node33907;
															assign node33907 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node33910 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node33913 = (inp[5]) ? node33917 : node33914;
															assign node33914 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node33917 = (inp[14]) ? 4'b0010 : 4'b0010;
												assign node33920 = (inp[0]) ? node33934 : node33921;
													assign node33921 = (inp[5]) ? node33929 : node33922;
														assign node33922 = (inp[14]) ? node33926 : node33923;
															assign node33923 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node33926 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node33929 = (inp[3]) ? 4'b0011 : node33930;
															assign node33930 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node33934 = (inp[3]) ? node33940 : node33935;
														assign node33935 = (inp[5]) ? 4'b0011 : node33936;
															assign node33936 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node33940 = (inp[5]) ? node33942 : 4'b0010;
															assign node33942 = (inp[7]) ? 4'b0000 : 4'b0000;
										assign node33945 = (inp[15]) ? node34007 : node33946;
											assign node33946 = (inp[0]) ? node33978 : node33947;
												assign node33947 = (inp[5]) ? node33963 : node33948;
													assign node33948 = (inp[3]) ? node33956 : node33949;
														assign node33949 = (inp[7]) ? node33953 : node33950;
															assign node33950 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node33953 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node33956 = (inp[8]) ? node33960 : node33957;
															assign node33957 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node33960 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node33963 = (inp[3]) ? node33971 : node33964;
														assign node33964 = (inp[7]) ? node33968 : node33965;
															assign node33965 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node33968 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node33971 = (inp[7]) ? node33975 : node33972;
															assign node33972 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node33975 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node33978 = (inp[5]) ? node33992 : node33979;
													assign node33979 = (inp[3]) ? node33985 : node33980;
														assign node33980 = (inp[8]) ? 4'b0001 : node33981;
															assign node33981 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node33985 = (inp[7]) ? node33989 : node33986;
															assign node33986 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node33989 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node33992 = (inp[3]) ? node34000 : node33993;
														assign node33993 = (inp[14]) ? node33997 : node33994;
															assign node33994 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node33997 = (inp[7]) ? 4'b0000 : 4'b0000;
														assign node34000 = (inp[14]) ? node34004 : node34001;
															assign node34001 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node34004 = (inp[8]) ? 4'b0010 : 4'b0010;
											assign node34007 = (inp[0]) ? node34031 : node34008;
												assign node34008 = (inp[3]) ? node34016 : node34009;
													assign node34009 = (inp[8]) ? node34013 : node34010;
														assign node34010 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node34013 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node34016 = (inp[5]) ? node34024 : node34017;
														assign node34017 = (inp[8]) ? node34021 : node34018;
															assign node34018 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node34021 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node34024 = (inp[7]) ? node34028 : node34025;
															assign node34025 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node34028 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node34031 = (inp[5]) ? node34039 : node34032;
													assign node34032 = (inp[7]) ? node34036 : node34033;
														assign node34033 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node34036 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node34039 = (inp[3]) ? node34047 : node34040;
														assign node34040 = (inp[7]) ? node34044 : node34041;
															assign node34041 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node34044 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node34047 = (inp[7]) ? node34051 : node34048;
															assign node34048 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node34051 = (inp[8]) ? 4'b0000 : 4'b0001;
									assign node34054 = (inp[7]) ? node34162 : node34055;
										assign node34055 = (inp[8]) ? node34115 : node34056;
											assign node34056 = (inp[2]) ? node34084 : node34057;
												assign node34057 = (inp[14]) ? node34071 : node34058;
													assign node34058 = (inp[0]) ? node34064 : node34059;
														assign node34059 = (inp[15]) ? node34061 : 4'b0011;
															assign node34061 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node34064 = (inp[15]) ? node34068 : node34065;
															assign node34065 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node34068 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node34071 = (inp[3]) ? node34077 : node34072;
														assign node34072 = (inp[5]) ? node34074 : 4'b0010;
															assign node34074 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node34077 = (inp[0]) ? node34081 : node34078;
															assign node34078 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node34081 = (inp[5]) ? 4'b0000 : 4'b0000;
												assign node34084 = (inp[5]) ? node34100 : node34085;
													assign node34085 = (inp[3]) ? node34093 : node34086;
														assign node34086 = (inp[15]) ? node34090 : node34087;
															assign node34087 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node34090 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node34093 = (inp[0]) ? node34097 : node34094;
															assign node34094 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node34097 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node34100 = (inp[15]) ? node34108 : node34101;
														assign node34101 = (inp[14]) ? node34105 : node34102;
															assign node34102 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node34105 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node34108 = (inp[3]) ? node34112 : node34109;
															assign node34109 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node34112 = (inp[0]) ? 4'b0000 : 4'b0010;
											assign node34115 = (inp[2]) ? node34141 : node34116;
												assign node34116 = (inp[14]) ? node34130 : node34117;
													assign node34117 = (inp[5]) ? node34125 : node34118;
														assign node34118 = (inp[15]) ? node34122 : node34119;
															assign node34119 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node34122 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node34125 = (inp[3]) ? 4'b0000 : node34126;
															assign node34126 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node34130 = (inp[0]) ? node34134 : node34131;
														assign node34131 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node34134 = (inp[15]) ? node34138 : node34135;
															assign node34135 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node34138 = (inp[5]) ? 4'b1101 : 4'b1101;
												assign node34141 = (inp[5]) ? node34155 : node34142;
													assign node34142 = (inp[15]) ? node34150 : node34143;
														assign node34143 = (inp[0]) ? node34147 : node34144;
															assign node34144 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node34147 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node34150 = (inp[3]) ? node34152 : 4'b1111;
															assign node34152 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node34155 = (inp[0]) ? node34159 : node34156;
														assign node34156 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node34159 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node34162 = (inp[8]) ? node34212 : node34163;
											assign node34163 = (inp[14]) ? node34189 : node34164;
												assign node34164 = (inp[2]) ? node34178 : node34165;
													assign node34165 = (inp[0]) ? node34173 : node34166;
														assign node34166 = (inp[15]) ? node34170 : node34167;
															assign node34167 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node34170 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node34173 = (inp[15]) ? node34175 : 4'b0000;
															assign node34175 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node34178 = (inp[0]) ? node34184 : node34179;
														assign node34179 = (inp[15]) ? node34181 : 4'b1101;
															assign node34181 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node34184 = (inp[15]) ? node34186 : 4'b1111;
															assign node34186 = (inp[5]) ? 4'b1101 : 4'b1101;
												assign node34189 = (inp[3]) ? node34205 : node34190;
													assign node34190 = (inp[15]) ? node34198 : node34191;
														assign node34191 = (inp[5]) ? node34195 : node34192;
															assign node34192 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node34195 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node34198 = (inp[5]) ? node34202 : node34199;
															assign node34199 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node34202 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node34205 = (inp[0]) ? node34209 : node34206;
														assign node34206 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node34209 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node34212 = (inp[14]) ? node34240 : node34213;
												assign node34213 = (inp[2]) ? node34227 : node34214;
													assign node34214 = (inp[5]) ? node34220 : node34215;
														assign node34215 = (inp[15]) ? 4'b1101 : node34216;
															assign node34216 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node34220 = (inp[0]) ? node34224 : node34221;
															assign node34221 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node34224 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node34227 = (inp[5]) ? node34235 : node34228;
														assign node34228 = (inp[3]) ? node34232 : node34229;
															assign node34229 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node34232 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node34235 = (inp[3]) ? node34237 : 4'b1110;
															assign node34237 = (inp[0]) ? 4'b1100 : 4'b1100;
												assign node34240 = (inp[0]) ? node34252 : node34241;
													assign node34241 = (inp[15]) ? node34247 : node34242;
														assign node34242 = (inp[3]) ? 4'b1100 : node34243;
															assign node34243 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node34247 = (inp[3]) ? 4'b1110 : node34248;
															assign node34248 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node34252 = (inp[15]) ? node34258 : node34253;
														assign node34253 = (inp[5]) ? 4'b1110 : node34254;
															assign node34254 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node34258 = (inp[5]) ? 4'b1100 : node34259;
															assign node34259 = (inp[3]) ? 4'b1100 : 4'b1110;
								assign node34263 = (inp[13]) ? node34489 : node34264;
									assign node34264 = (inp[8]) ? node34376 : node34265;
										assign node34265 = (inp[7]) ? node34321 : node34266;
											assign node34266 = (inp[14]) ? node34294 : node34267;
												assign node34267 = (inp[2]) ? node34283 : node34268;
													assign node34268 = (inp[3]) ? node34276 : node34269;
														assign node34269 = (inp[5]) ? node34273 : node34270;
															assign node34270 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node34273 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node34276 = (inp[0]) ? node34280 : node34277;
															assign node34277 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node34280 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node34283 = (inp[0]) ? node34291 : node34284;
														assign node34284 = (inp[15]) ? node34288 : node34285;
															assign node34285 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node34288 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node34291 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node34294 = (inp[3]) ? node34308 : node34295;
													assign node34295 = (inp[2]) ? node34303 : node34296;
														assign node34296 = (inp[0]) ? node34300 : node34297;
															assign node34297 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node34300 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node34303 = (inp[15]) ? node34305 : 4'b0010;
															assign node34305 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node34308 = (inp[0]) ? node34314 : node34309;
														assign node34309 = (inp[2]) ? node34311 : 4'b0000;
															assign node34311 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node34314 = (inp[2]) ? node34318 : node34315;
															assign node34315 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node34318 = (inp[15]) ? 4'b0000 : 4'b0000;
											assign node34321 = (inp[2]) ? node34353 : node34322;
												assign node34322 = (inp[14]) ? node34338 : node34323;
													assign node34323 = (inp[3]) ? node34331 : node34324;
														assign node34324 = (inp[5]) ? node34328 : node34325;
															assign node34325 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node34328 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node34331 = (inp[0]) ? node34335 : node34332;
															assign node34332 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node34335 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node34338 = (inp[5]) ? node34346 : node34339;
														assign node34339 = (inp[3]) ? node34343 : node34340;
															assign node34340 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node34343 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node34346 = (inp[3]) ? node34350 : node34347;
															assign node34347 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node34350 = (inp[0]) ? 4'b1101 : 4'b1101;
												assign node34353 = (inp[15]) ? node34365 : node34354;
													assign node34354 = (inp[0]) ? node34360 : node34355;
														assign node34355 = (inp[5]) ? 4'b1101 : node34356;
															assign node34356 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node34360 = (inp[3]) ? 4'b1111 : node34361;
															assign node34361 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node34365 = (inp[0]) ? node34371 : node34366;
														assign node34366 = (inp[5]) ? 4'b1111 : node34367;
															assign node34367 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node34371 = (inp[3]) ? 4'b1101 : node34372;
															assign node34372 = (inp[5]) ? 4'b1101 : 4'b1111;
										assign node34376 = (inp[7]) ? node34436 : node34377;
											assign node34377 = (inp[14]) ? node34407 : node34378;
												assign node34378 = (inp[2]) ? node34392 : node34379;
													assign node34379 = (inp[15]) ? node34385 : node34380;
														assign node34380 = (inp[5]) ? node34382 : 4'b0010;
															assign node34382 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node34385 = (inp[0]) ? node34389 : node34386;
															assign node34386 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node34389 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node34392 = (inp[0]) ? node34400 : node34393;
														assign node34393 = (inp[15]) ? node34397 : node34394;
															assign node34394 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node34397 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node34400 = (inp[15]) ? node34404 : node34401;
															assign node34401 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node34404 = (inp[5]) ? 4'b1101 : 4'b1101;
												assign node34407 = (inp[2]) ? node34421 : node34408;
													assign node34408 = (inp[15]) ? node34414 : node34409;
														assign node34409 = (inp[0]) ? node34411 : 4'b1101;
															assign node34411 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node34414 = (inp[0]) ? node34418 : node34415;
															assign node34415 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node34418 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node34421 = (inp[0]) ? node34429 : node34422;
														assign node34422 = (inp[15]) ? node34426 : node34423;
															assign node34423 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node34426 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node34429 = (inp[15]) ? node34433 : node34430;
															assign node34430 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node34433 = (inp[5]) ? 4'b1101 : 4'b1101;
											assign node34436 = (inp[14]) ? node34466 : node34437;
												assign node34437 = (inp[2]) ? node34453 : node34438;
													assign node34438 = (inp[0]) ? node34446 : node34439;
														assign node34439 = (inp[15]) ? node34443 : node34440;
															assign node34440 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node34443 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node34446 = (inp[15]) ? node34450 : node34447;
															assign node34447 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node34450 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node34453 = (inp[0]) ? node34461 : node34454;
														assign node34454 = (inp[15]) ? node34458 : node34455;
															assign node34455 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node34458 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node34461 = (inp[15]) ? node34463 : 4'b1110;
															assign node34463 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node34466 = (inp[15]) ? node34478 : node34467;
													assign node34467 = (inp[0]) ? node34473 : node34468;
														assign node34468 = (inp[3]) ? 4'b1100 : node34469;
															assign node34469 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node34473 = (inp[3]) ? 4'b1110 : node34474;
															assign node34474 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node34478 = (inp[0]) ? node34484 : node34479;
														assign node34479 = (inp[3]) ? 4'b1110 : node34480;
															assign node34480 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node34484 = (inp[5]) ? 4'b1100 : node34485;
															assign node34485 = (inp[3]) ? 4'b1100 : 4'b1110;
									assign node34489 = (inp[2]) ? node34611 : node34490;
										assign node34490 = (inp[14]) ? node34552 : node34491;
											assign node34491 = (inp[15]) ? node34523 : node34492;
												assign node34492 = (inp[0]) ? node34508 : node34493;
													assign node34493 = (inp[5]) ? node34501 : node34494;
														assign node34494 = (inp[3]) ? node34498 : node34495;
															assign node34495 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node34498 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node34501 = (inp[7]) ? node34505 : node34502;
															assign node34502 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node34505 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node34508 = (inp[5]) ? node34516 : node34509;
														assign node34509 = (inp[3]) ? node34513 : node34510;
															assign node34510 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node34513 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node34516 = (inp[7]) ? node34520 : node34517;
															assign node34517 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node34520 = (inp[8]) ? 4'b1111 : 4'b1110;
												assign node34523 = (inp[0]) ? node34537 : node34524;
													assign node34524 = (inp[3]) ? node34532 : node34525;
														assign node34525 = (inp[5]) ? node34529 : node34526;
															assign node34526 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node34529 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node34532 = (inp[5]) ? 4'b1111 : node34533;
															assign node34533 = (inp[8]) ? 4'b1110 : 4'b1110;
													assign node34537 = (inp[5]) ? node34545 : node34538;
														assign node34538 = (inp[3]) ? node34542 : node34539;
															assign node34539 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node34542 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node34545 = (inp[3]) ? node34549 : node34546;
															assign node34546 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node34549 = (inp[7]) ? 4'b1100 : 4'b1100;
											assign node34552 = (inp[8]) ? node34584 : node34553;
												assign node34553 = (inp[7]) ? node34569 : node34554;
													assign node34554 = (inp[3]) ? node34562 : node34555;
														assign node34555 = (inp[15]) ? node34559 : node34556;
															assign node34556 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node34559 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node34562 = (inp[15]) ? node34566 : node34563;
															assign node34563 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node34566 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node34569 = (inp[3]) ? node34577 : node34570;
														assign node34570 = (inp[5]) ? node34574 : node34571;
															assign node34571 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node34574 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node34577 = (inp[15]) ? node34581 : node34578;
															assign node34578 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node34581 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node34584 = (inp[7]) ? node34600 : node34585;
													assign node34585 = (inp[0]) ? node34593 : node34586;
														assign node34586 = (inp[15]) ? node34590 : node34587;
															assign node34587 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node34590 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node34593 = (inp[15]) ? node34597 : node34594;
															assign node34594 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node34597 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node34600 = (inp[0]) ? node34606 : node34601;
														assign node34601 = (inp[15]) ? 4'b1110 : node34602;
															assign node34602 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node34606 = (inp[15]) ? node34608 : 4'b1110;
															assign node34608 = (inp[3]) ? 4'b1100 : 4'b1100;
										assign node34611 = (inp[8]) ? node34659 : node34612;
											assign node34612 = (inp[7]) ? node34636 : node34613;
												assign node34613 = (inp[15]) ? node34625 : node34614;
													assign node34614 = (inp[0]) ? node34620 : node34615;
														assign node34615 = (inp[3]) ? 4'b1100 : node34616;
															assign node34616 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node34620 = (inp[3]) ? 4'b1110 : node34621;
															assign node34621 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node34625 = (inp[0]) ? node34631 : node34626;
														assign node34626 = (inp[3]) ? 4'b1110 : node34627;
															assign node34627 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node34631 = (inp[3]) ? 4'b1100 : node34632;
															assign node34632 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node34636 = (inp[15]) ? node34648 : node34637;
													assign node34637 = (inp[0]) ? node34643 : node34638;
														assign node34638 = (inp[3]) ? 4'b1101 : node34639;
															assign node34639 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node34643 = (inp[5]) ? 4'b1111 : node34644;
															assign node34644 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node34648 = (inp[0]) ? node34654 : node34649;
														assign node34649 = (inp[5]) ? 4'b1111 : node34650;
															assign node34650 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node34654 = (inp[5]) ? 4'b1101 : node34655;
															assign node34655 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node34659 = (inp[7]) ? node34681 : node34660;
												assign node34660 = (inp[3]) ? node34674 : node34661;
													assign node34661 = (inp[14]) ? node34669 : node34662;
														assign node34662 = (inp[5]) ? node34666 : node34663;
															assign node34663 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node34666 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node34669 = (inp[15]) ? node34671 : 4'b1101;
															assign node34671 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node34674 = (inp[15]) ? node34678 : node34675;
														assign node34675 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node34678 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node34681 = (inp[14]) ? node34697 : node34682;
													assign node34682 = (inp[0]) ? node34690 : node34683;
														assign node34683 = (inp[15]) ? node34687 : node34684;
															assign node34684 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node34687 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node34690 = (inp[15]) ? node34694 : node34691;
															assign node34691 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node34694 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node34697 = (inp[0]) ? node34705 : node34698;
														assign node34698 = (inp[15]) ? node34702 : node34699;
															assign node34699 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node34702 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node34705 = (inp[15]) ? node34709 : node34706;
															assign node34706 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node34709 = (inp[3]) ? 4'b1100 : 4'b1100;
							assign node34712 = (inp[13]) ? node35180 : node34713;
								assign node34713 = (inp[1]) ? node34951 : node34714;
									assign node34714 = (inp[5]) ? node34836 : node34715;
										assign node34715 = (inp[14]) ? node34775 : node34716;
											assign node34716 = (inp[8]) ? node34748 : node34717;
												assign node34717 = (inp[15]) ? node34733 : node34718;
													assign node34718 = (inp[3]) ? node34726 : node34719;
														assign node34719 = (inp[0]) ? node34723 : node34720;
															assign node34720 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node34723 = (inp[2]) ? 4'b1100 : 4'b1100;
														assign node34726 = (inp[0]) ? node34730 : node34727;
															assign node34727 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node34730 = (inp[7]) ? 4'b1110 : 4'b1110;
													assign node34733 = (inp[3]) ? node34741 : node34734;
														assign node34734 = (inp[0]) ? node34738 : node34735;
															assign node34735 = (inp[2]) ? 4'b1100 : 4'b1100;
															assign node34738 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node34741 = (inp[0]) ? node34745 : node34742;
															assign node34742 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node34745 = (inp[2]) ? 4'b1100 : 4'b1100;
												assign node34748 = (inp[3]) ? node34762 : node34749;
													assign node34749 = (inp[2]) ? node34757 : node34750;
														assign node34750 = (inp[7]) ? node34754 : node34751;
															assign node34751 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node34754 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node34757 = (inp[7]) ? node34759 : 4'b1101;
															assign node34759 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node34762 = (inp[7]) ? node34770 : node34763;
														assign node34763 = (inp[2]) ? node34767 : node34764;
															assign node34764 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node34767 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node34770 = (inp[2]) ? node34772 : 4'b1101;
															assign node34772 = (inp[0]) ? 4'b1100 : 4'b1100;
											assign node34775 = (inp[8]) ? node34807 : node34776;
												assign node34776 = (inp[7]) ? node34792 : node34777;
													assign node34777 = (inp[0]) ? node34785 : node34778;
														assign node34778 = (inp[2]) ? node34782 : node34779;
															assign node34779 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node34782 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node34785 = (inp[15]) ? node34789 : node34786;
															assign node34786 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node34789 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node34792 = (inp[2]) ? node34800 : node34793;
														assign node34793 = (inp[3]) ? node34797 : node34794;
															assign node34794 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node34797 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node34800 = (inp[15]) ? node34804 : node34801;
															assign node34801 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node34804 = (inp[3]) ? 4'b1101 : 4'b1101;
												assign node34807 = (inp[7]) ? node34821 : node34808;
													assign node34808 = (inp[0]) ? node34814 : node34809;
														assign node34809 = (inp[2]) ? node34811 : 4'b1111;
															assign node34811 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node34814 = (inp[15]) ? node34818 : node34815;
															assign node34815 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node34818 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node34821 = (inp[3]) ? node34829 : node34822;
														assign node34822 = (inp[15]) ? node34826 : node34823;
															assign node34823 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node34826 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node34829 = (inp[2]) ? node34833 : node34830;
															assign node34830 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node34833 = (inp[15]) ? 4'b1100 : 4'b1100;
										assign node34836 = (inp[14]) ? node34898 : node34837;
											assign node34837 = (inp[15]) ? node34867 : node34838;
												assign node34838 = (inp[0]) ? node34854 : node34839;
													assign node34839 = (inp[2]) ? node34847 : node34840;
														assign node34840 = (inp[7]) ? node34844 : node34841;
															assign node34841 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node34844 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node34847 = (inp[8]) ? node34851 : node34848;
															assign node34848 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node34851 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node34854 = (inp[3]) ? node34860 : node34855;
														assign node34855 = (inp[8]) ? 4'b1111 : node34856;
															assign node34856 = (inp[2]) ? 4'b1110 : 4'b1110;
														assign node34860 = (inp[7]) ? node34864 : node34861;
															assign node34861 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node34864 = (inp[2]) ? 4'b1110 : 4'b1110;
												assign node34867 = (inp[0]) ? node34883 : node34868;
													assign node34868 = (inp[7]) ? node34876 : node34869;
														assign node34869 = (inp[3]) ? node34873 : node34870;
															assign node34870 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node34873 = (inp[2]) ? 4'b1110 : 4'b1110;
														assign node34876 = (inp[2]) ? node34880 : node34877;
															assign node34877 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node34880 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node34883 = (inp[8]) ? node34891 : node34884;
														assign node34884 = (inp[2]) ? node34888 : node34885;
															assign node34885 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node34888 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node34891 = (inp[2]) ? node34895 : node34892;
															assign node34892 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node34895 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node34898 = (inp[7]) ? node34928 : node34899;
												assign node34899 = (inp[8]) ? node34915 : node34900;
													assign node34900 = (inp[3]) ? node34908 : node34901;
														assign node34901 = (inp[0]) ? node34905 : node34902;
															assign node34902 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node34905 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node34908 = (inp[15]) ? node34912 : node34909;
															assign node34909 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node34912 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node34915 = (inp[3]) ? node34921 : node34916;
														assign node34916 = (inp[0]) ? 4'b1101 : node34917;
															assign node34917 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node34921 = (inp[0]) ? node34925 : node34922;
															assign node34922 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node34925 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node34928 = (inp[8]) ? node34936 : node34929;
													assign node34929 = (inp[0]) ? node34933 : node34930;
														assign node34930 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node34933 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node34936 = (inp[3]) ? node34944 : node34937;
														assign node34937 = (inp[2]) ? node34941 : node34938;
															assign node34938 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node34941 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node34944 = (inp[2]) ? node34948 : node34945;
															assign node34945 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node34948 = (inp[0]) ? 4'b1100 : 4'b1110;
									assign node34951 = (inp[8]) ? node35065 : node34952;
										assign node34952 = (inp[7]) ? node35006 : node34953;
											assign node34953 = (inp[14]) ? node34983 : node34954;
												assign node34954 = (inp[2]) ? node34970 : node34955;
													assign node34955 = (inp[15]) ? node34963 : node34956;
														assign node34956 = (inp[0]) ? node34960 : node34957;
															assign node34957 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node34960 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node34963 = (inp[0]) ? node34967 : node34964;
															assign node34964 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node34967 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node34970 = (inp[15]) ? node34978 : node34971;
														assign node34971 = (inp[0]) ? node34975 : node34972;
															assign node34972 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node34975 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node34978 = (inp[0]) ? node34980 : 4'b1110;
															assign node34980 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node34983 = (inp[15]) ? node34995 : node34984;
													assign node34984 = (inp[0]) ? node34990 : node34985;
														assign node34985 = (inp[5]) ? 4'b1100 : node34986;
															assign node34986 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node34990 = (inp[5]) ? 4'b1110 : node34991;
															assign node34991 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node34995 = (inp[0]) ? node35001 : node34996;
														assign node34996 = (inp[3]) ? 4'b1110 : node34997;
															assign node34997 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node35001 = (inp[5]) ? 4'b1100 : node35002;
															assign node35002 = (inp[3]) ? 4'b1100 : 4'b1110;
											assign node35006 = (inp[2]) ? node35036 : node35007;
												assign node35007 = (inp[14]) ? node35023 : node35008;
													assign node35008 = (inp[5]) ? node35016 : node35009;
														assign node35009 = (inp[15]) ? node35013 : node35010;
															assign node35010 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node35013 = (inp[3]) ? 4'b1100 : 4'b1100;
														assign node35016 = (inp[0]) ? node35020 : node35017;
															assign node35017 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node35020 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node35023 = (inp[15]) ? node35029 : node35024;
														assign node35024 = (inp[0]) ? 4'b0111 : node35025;
															assign node35025 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node35029 = (inp[0]) ? node35033 : node35030;
															assign node35030 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node35033 = (inp[3]) ? 4'b0101 : 4'b0101;
												assign node35036 = (inp[5]) ? node35052 : node35037;
													assign node35037 = (inp[0]) ? node35045 : node35038;
														assign node35038 = (inp[14]) ? node35042 : node35039;
															assign node35039 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node35042 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node35045 = (inp[15]) ? node35049 : node35046;
															assign node35046 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node35049 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node35052 = (inp[3]) ? node35060 : node35053;
														assign node35053 = (inp[15]) ? node35057 : node35054;
															assign node35054 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node35057 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node35060 = (inp[14]) ? node35062 : 4'b0101;
															assign node35062 = (inp[15]) ? 4'b0101 : 4'b0101;
										assign node35065 = (inp[7]) ? node35121 : node35066;
											assign node35066 = (inp[2]) ? node35098 : node35067;
												assign node35067 = (inp[14]) ? node35083 : node35068;
													assign node35068 = (inp[3]) ? node35076 : node35069;
														assign node35069 = (inp[5]) ? node35073 : node35070;
															assign node35070 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node35073 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node35076 = (inp[5]) ? node35080 : node35077;
															assign node35077 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node35080 = (inp[0]) ? 4'b1100 : 4'b1100;
													assign node35083 = (inp[3]) ? node35091 : node35084;
														assign node35084 = (inp[15]) ? node35088 : node35085;
															assign node35085 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node35088 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node35091 = (inp[0]) ? node35095 : node35092;
															assign node35092 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node35095 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node35098 = (inp[0]) ? node35110 : node35099;
													assign node35099 = (inp[15]) ? node35105 : node35100;
														assign node35100 = (inp[5]) ? 4'b0101 : node35101;
															assign node35101 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node35105 = (inp[5]) ? 4'b0111 : node35106;
															assign node35106 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node35110 = (inp[15]) ? node35116 : node35111;
														assign node35111 = (inp[3]) ? 4'b0111 : node35112;
															assign node35112 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node35116 = (inp[5]) ? 4'b0101 : node35117;
															assign node35117 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node35121 = (inp[14]) ? node35149 : node35122;
												assign node35122 = (inp[2]) ? node35136 : node35123;
													assign node35123 = (inp[5]) ? node35129 : node35124;
														assign node35124 = (inp[15]) ? node35126 : 4'b0101;
															assign node35126 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node35129 = (inp[3]) ? node35133 : node35130;
															assign node35130 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node35133 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node35136 = (inp[5]) ? node35144 : node35137;
														assign node35137 = (inp[15]) ? node35141 : node35138;
															assign node35138 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node35141 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node35144 = (inp[15]) ? 4'b0110 : node35145;
															assign node35145 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node35149 = (inp[3]) ? node35165 : node35150;
													assign node35150 = (inp[15]) ? node35158 : node35151;
														assign node35151 = (inp[5]) ? node35155 : node35152;
															assign node35152 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node35155 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node35158 = (inp[0]) ? node35162 : node35159;
															assign node35159 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node35162 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node35165 = (inp[5]) ? node35173 : node35166;
														assign node35166 = (inp[15]) ? node35170 : node35167;
															assign node35167 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node35170 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node35173 = (inp[0]) ? node35177 : node35174;
															assign node35174 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node35177 = (inp[15]) ? 4'b0100 : 4'b0110;
								assign node35180 = (inp[1]) ? node35408 : node35181;
									assign node35181 = (inp[7]) ? node35293 : node35182;
										assign node35182 = (inp[8]) ? node35240 : node35183;
											assign node35183 = (inp[14]) ? node35213 : node35184;
												assign node35184 = (inp[2]) ? node35200 : node35185;
													assign node35185 = (inp[15]) ? node35193 : node35186;
														assign node35186 = (inp[0]) ? node35190 : node35187;
															assign node35187 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node35190 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node35193 = (inp[0]) ? node35197 : node35194;
															assign node35194 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node35197 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node35200 = (inp[15]) ? node35206 : node35201;
														assign node35201 = (inp[5]) ? 4'b1110 : node35202;
															assign node35202 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node35206 = (inp[0]) ? node35210 : node35207;
															assign node35207 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node35210 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node35213 = (inp[2]) ? node35227 : node35214;
													assign node35214 = (inp[15]) ? node35220 : node35215;
														assign node35215 = (inp[0]) ? 4'b1110 : node35216;
															assign node35216 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node35220 = (inp[0]) ? node35224 : node35221;
															assign node35221 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node35224 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node35227 = (inp[0]) ? node35235 : node35228;
														assign node35228 = (inp[15]) ? node35232 : node35229;
															assign node35229 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node35232 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node35235 = (inp[15]) ? 4'b1100 : node35236;
															assign node35236 = (inp[3]) ? 4'b1110 : 4'b1100;
											assign node35240 = (inp[2]) ? node35270 : node35241;
												assign node35241 = (inp[14]) ? node35257 : node35242;
													assign node35242 = (inp[5]) ? node35250 : node35243;
														assign node35243 = (inp[15]) ? node35247 : node35244;
															assign node35244 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node35247 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node35250 = (inp[3]) ? node35254 : node35251;
															assign node35251 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node35254 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node35257 = (inp[5]) ? node35265 : node35258;
														assign node35258 = (inp[3]) ? node35262 : node35259;
															assign node35259 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node35262 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node35265 = (inp[3]) ? node35267 : 4'b0101;
															assign node35267 = (inp[15]) ? 4'b0101 : 4'b0101;
												assign node35270 = (inp[15]) ? node35282 : node35271;
													assign node35271 = (inp[0]) ? node35277 : node35272;
														assign node35272 = (inp[5]) ? 4'b0101 : node35273;
															assign node35273 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node35277 = (inp[5]) ? 4'b0111 : node35278;
															assign node35278 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node35282 = (inp[0]) ? node35288 : node35283;
														assign node35283 = (inp[5]) ? 4'b0111 : node35284;
															assign node35284 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node35288 = (inp[3]) ? 4'b0101 : node35289;
															assign node35289 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node35293 = (inp[8]) ? node35347 : node35294;
											assign node35294 = (inp[2]) ? node35324 : node35295;
												assign node35295 = (inp[14]) ? node35311 : node35296;
													assign node35296 = (inp[3]) ? node35304 : node35297;
														assign node35297 = (inp[5]) ? node35301 : node35298;
															assign node35298 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node35301 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node35304 = (inp[15]) ? node35308 : node35305;
															assign node35305 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node35308 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node35311 = (inp[0]) ? node35319 : node35312;
														assign node35312 = (inp[15]) ? node35316 : node35313;
															assign node35313 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node35316 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node35319 = (inp[15]) ? node35321 : 4'b0111;
															assign node35321 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node35324 = (inp[15]) ? node35336 : node35325;
													assign node35325 = (inp[0]) ? node35331 : node35326;
														assign node35326 = (inp[3]) ? 4'b0101 : node35327;
															assign node35327 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node35331 = (inp[3]) ? 4'b0111 : node35332;
															assign node35332 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node35336 = (inp[0]) ? node35342 : node35337;
														assign node35337 = (inp[5]) ? 4'b0111 : node35338;
															assign node35338 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node35342 = (inp[3]) ? 4'b0101 : node35343;
															assign node35343 = (inp[5]) ? 4'b0101 : 4'b0111;
											assign node35347 = (inp[2]) ? node35377 : node35348;
												assign node35348 = (inp[14]) ? node35364 : node35349;
													assign node35349 = (inp[0]) ? node35357 : node35350;
														assign node35350 = (inp[15]) ? node35354 : node35351;
															assign node35351 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node35354 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node35357 = (inp[15]) ? node35361 : node35358;
															assign node35358 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node35361 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node35364 = (inp[3]) ? node35370 : node35365;
														assign node35365 = (inp[0]) ? 4'b0100 : node35366;
															assign node35366 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node35370 = (inp[15]) ? node35374 : node35371;
															assign node35371 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node35374 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node35377 = (inp[3]) ? node35393 : node35378;
													assign node35378 = (inp[14]) ? node35386 : node35379;
														assign node35379 = (inp[15]) ? node35383 : node35380;
															assign node35380 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node35383 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node35386 = (inp[15]) ? node35390 : node35387;
															assign node35387 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node35390 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node35393 = (inp[5]) ? node35401 : node35394;
														assign node35394 = (inp[14]) ? node35398 : node35395;
															assign node35395 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node35398 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node35401 = (inp[15]) ? node35405 : node35402;
															assign node35402 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node35405 = (inp[0]) ? 4'b0100 : 4'b0110;
									assign node35408 = (inp[2]) ? node35532 : node35409;
										assign node35409 = (inp[0]) ? node35473 : node35410;
											assign node35410 = (inp[15]) ? node35442 : node35411;
												assign node35411 = (inp[3]) ? node35427 : node35412;
													assign node35412 = (inp[5]) ? node35420 : node35413;
														assign node35413 = (inp[8]) ? node35417 : node35414;
															assign node35414 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node35417 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node35420 = (inp[14]) ? node35424 : node35421;
															assign node35421 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node35424 = (inp[7]) ? 4'b0100 : 4'b0100;
													assign node35427 = (inp[14]) ? node35435 : node35428;
														assign node35428 = (inp[7]) ? node35432 : node35429;
															assign node35429 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node35432 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node35435 = (inp[7]) ? node35439 : node35436;
															assign node35436 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node35439 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node35442 = (inp[5]) ? node35458 : node35443;
													assign node35443 = (inp[3]) ? node35451 : node35444;
														assign node35444 = (inp[8]) ? node35448 : node35445;
															assign node35445 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node35448 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node35451 = (inp[8]) ? node35455 : node35452;
															assign node35452 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node35455 = (inp[14]) ? 4'b0110 : 4'b0110;
													assign node35458 = (inp[8]) ? node35466 : node35459;
														assign node35459 = (inp[7]) ? node35463 : node35460;
															assign node35460 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node35463 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node35466 = (inp[3]) ? node35470 : node35467;
															assign node35467 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node35470 = (inp[7]) ? 4'b0110 : 4'b0110;
											assign node35473 = (inp[15]) ? node35503 : node35474;
												assign node35474 = (inp[5]) ? node35490 : node35475;
													assign node35475 = (inp[3]) ? node35483 : node35476;
														assign node35476 = (inp[7]) ? node35480 : node35477;
															assign node35477 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node35480 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node35483 = (inp[14]) ? node35487 : node35484;
															assign node35484 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node35487 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node35490 = (inp[3]) ? node35498 : node35491;
														assign node35491 = (inp[7]) ? node35495 : node35492;
															assign node35492 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node35495 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node35498 = (inp[14]) ? 4'b0111 : node35499;
															assign node35499 = (inp[7]) ? 4'b0110 : 4'b0110;
												assign node35503 = (inp[3]) ? node35517 : node35504;
													assign node35504 = (inp[5]) ? node35510 : node35505;
														assign node35505 = (inp[7]) ? node35507 : 4'b0111;
															assign node35507 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node35510 = (inp[8]) ? node35514 : node35511;
															assign node35511 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node35514 = (inp[7]) ? 4'b0100 : 4'b0100;
													assign node35517 = (inp[8]) ? node35525 : node35518;
														assign node35518 = (inp[7]) ? node35522 : node35519;
															assign node35519 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node35522 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node35525 = (inp[5]) ? node35529 : node35526;
															assign node35526 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node35529 = (inp[14]) ? 4'b0100 : 4'b0100;
										assign node35532 = (inp[15]) ? node35594 : node35533;
											assign node35533 = (inp[0]) ? node35563 : node35534;
												assign node35534 = (inp[3]) ? node35550 : node35535;
													assign node35535 = (inp[5]) ? node35543 : node35536;
														assign node35536 = (inp[7]) ? node35540 : node35537;
															assign node35537 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node35540 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node35543 = (inp[7]) ? node35547 : node35544;
															assign node35544 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node35547 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node35550 = (inp[14]) ? node35556 : node35551;
														assign node35551 = (inp[5]) ? 4'b0100 : node35552;
															assign node35552 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node35556 = (inp[8]) ? node35560 : node35557;
															assign node35557 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node35560 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node35563 = (inp[3]) ? node35579 : node35564;
													assign node35564 = (inp[5]) ? node35572 : node35565;
														assign node35565 = (inp[8]) ? node35569 : node35566;
															assign node35566 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node35569 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node35572 = (inp[8]) ? node35576 : node35573;
															assign node35573 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node35576 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node35579 = (inp[14]) ? node35587 : node35580;
														assign node35580 = (inp[7]) ? node35584 : node35581;
															assign node35581 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node35584 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node35587 = (inp[8]) ? node35591 : node35588;
															assign node35588 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node35591 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node35594 = (inp[0]) ? node35626 : node35595;
												assign node35595 = (inp[5]) ? node35611 : node35596;
													assign node35596 = (inp[3]) ? node35604 : node35597;
														assign node35597 = (inp[7]) ? node35601 : node35598;
															assign node35598 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node35601 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node35604 = (inp[8]) ? node35608 : node35605;
															assign node35605 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node35608 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node35611 = (inp[14]) ? node35619 : node35612;
														assign node35612 = (inp[7]) ? node35616 : node35613;
															assign node35613 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node35616 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node35619 = (inp[3]) ? node35623 : node35620;
															assign node35620 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node35623 = (inp[8]) ? 4'b0110 : 4'b0110;
												assign node35626 = (inp[3]) ? node35642 : node35627;
													assign node35627 = (inp[5]) ? node35635 : node35628;
														assign node35628 = (inp[14]) ? node35632 : node35629;
															assign node35629 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node35632 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node35635 = (inp[7]) ? node35639 : node35636;
															assign node35636 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node35639 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node35642 = (inp[14]) ? node35650 : node35643;
														assign node35643 = (inp[8]) ? node35647 : node35644;
															assign node35644 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node35647 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node35650 = (inp[7]) ? node35654 : node35651;
															assign node35651 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node35654 = (inp[8]) ? 4'b0100 : 4'b0101;
				assign node35657 = (inp[12]) ? node39223 : node35658;
					assign node35658 = (inp[11]) ? node37436 : node35659;
						assign node35659 = (inp[6]) ? node36545 : node35660;
							assign node35660 = (inp[13]) ? node36086 : node35661;
								assign node35661 = (inp[1]) ? node35873 : node35662;
									assign node35662 = (inp[15]) ? node35770 : node35663;
										assign node35663 = (inp[0]) ? node35719 : node35664;
											assign node35664 = (inp[5]) ? node35688 : node35665;
												assign node35665 = (inp[8]) ? node35677 : node35666;
													assign node35666 = (inp[7]) ? node35672 : node35667;
														assign node35667 = (inp[14]) ? 4'b1010 : node35668;
															assign node35668 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node35672 = (inp[14]) ? 4'b1011 : node35673;
															assign node35673 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node35677 = (inp[7]) ? node35683 : node35678;
														assign node35678 = (inp[2]) ? 4'b1011 : node35679;
															assign node35679 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node35683 = (inp[14]) ? 4'b1010 : node35684;
															assign node35684 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node35688 = (inp[3]) ? node35704 : node35689;
													assign node35689 = (inp[2]) ? node35697 : node35690;
														assign node35690 = (inp[7]) ? node35694 : node35691;
															assign node35691 = (inp[8]) ? 4'b1010 : 4'b1010;
															assign node35694 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node35697 = (inp[8]) ? node35701 : node35698;
															assign node35698 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node35701 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node35704 = (inp[8]) ? node35712 : node35705;
														assign node35705 = (inp[7]) ? node35709 : node35706;
															assign node35706 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node35709 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node35712 = (inp[7]) ? node35716 : node35713;
															assign node35713 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node35716 = (inp[14]) ? 4'b1000 : 4'b1000;
											assign node35719 = (inp[3]) ? node35743 : node35720;
												assign node35720 = (inp[2]) ? node35736 : node35721;
													assign node35721 = (inp[7]) ? node35729 : node35722;
														assign node35722 = (inp[14]) ? node35726 : node35723;
															assign node35723 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node35726 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node35729 = (inp[5]) ? node35733 : node35730;
															assign node35730 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node35733 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node35736 = (inp[8]) ? node35740 : node35737;
														assign node35737 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node35740 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node35743 = (inp[5]) ? node35757 : node35744;
													assign node35744 = (inp[7]) ? node35752 : node35745;
														assign node35745 = (inp[8]) ? node35749 : node35746;
															assign node35746 = (inp[2]) ? 4'b1000 : 4'b1000;
															assign node35749 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node35752 = (inp[8]) ? node35754 : 4'b1001;
															assign node35754 = (inp[2]) ? 4'b1000 : 4'b1000;
													assign node35757 = (inp[14]) ? node35763 : node35758;
														assign node35758 = (inp[7]) ? 4'b1011 : node35759;
															assign node35759 = (inp[2]) ? 4'b1010 : 4'b1010;
														assign node35763 = (inp[8]) ? node35767 : node35764;
															assign node35764 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node35767 = (inp[7]) ? 4'b1010 : 4'b1011;
										assign node35770 = (inp[0]) ? node35820 : node35771;
											assign node35771 = (inp[3]) ? node35795 : node35772;
												assign node35772 = (inp[8]) ? node35784 : node35773;
													assign node35773 = (inp[7]) ? node35779 : node35774;
														assign node35774 = (inp[2]) ? 4'b1000 : node35775;
															assign node35775 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node35779 = (inp[2]) ? 4'b1001 : node35780;
															assign node35780 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node35784 = (inp[7]) ? node35790 : node35785;
														assign node35785 = (inp[2]) ? 4'b1001 : node35786;
															assign node35786 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node35790 = (inp[2]) ? 4'b1000 : node35791;
															assign node35791 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node35795 = (inp[5]) ? node35809 : node35796;
													assign node35796 = (inp[7]) ? node35804 : node35797;
														assign node35797 = (inp[8]) ? node35801 : node35798;
															assign node35798 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node35801 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node35804 = (inp[8]) ? node35806 : 4'b1001;
															assign node35806 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node35809 = (inp[2]) ? node35815 : node35810;
														assign node35810 = (inp[14]) ? 4'b1010 : node35811;
															assign node35811 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node35815 = (inp[7]) ? 4'b1011 : node35816;
															assign node35816 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node35820 = (inp[3]) ? node35844 : node35821;
												assign node35821 = (inp[7]) ? node35833 : node35822;
													assign node35822 = (inp[8]) ? node35828 : node35823;
														assign node35823 = (inp[2]) ? 4'b1010 : node35824;
															assign node35824 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node35828 = (inp[14]) ? 4'b1011 : node35829;
															assign node35829 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node35833 = (inp[8]) ? node35839 : node35834;
														assign node35834 = (inp[14]) ? 4'b1011 : node35835;
															assign node35835 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node35839 = (inp[14]) ? 4'b1010 : node35840;
															assign node35840 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node35844 = (inp[5]) ? node35858 : node35845;
													assign node35845 = (inp[14]) ? node35853 : node35846;
														assign node35846 = (inp[2]) ? node35850 : node35847;
															assign node35847 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node35850 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node35853 = (inp[8]) ? 4'b1011 : node35854;
															assign node35854 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node35858 = (inp[8]) ? node35866 : node35859;
														assign node35859 = (inp[7]) ? node35863 : node35860;
															assign node35860 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node35863 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node35866 = (inp[7]) ? node35870 : node35867;
															assign node35867 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node35870 = (inp[2]) ? 4'b1000 : 4'b1001;
									assign node35873 = (inp[8]) ? node35977 : node35874;
										assign node35874 = (inp[7]) ? node35924 : node35875;
											assign node35875 = (inp[14]) ? node35903 : node35876;
												assign node35876 = (inp[2]) ? node35890 : node35877;
													assign node35877 = (inp[0]) ? node35885 : node35878;
														assign node35878 = (inp[15]) ? node35882 : node35879;
															assign node35879 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node35882 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node35885 = (inp[5]) ? node35887 : 4'b1011;
															assign node35887 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node35890 = (inp[15]) ? node35896 : node35891;
														assign node35891 = (inp[0]) ? 4'b1000 : node35892;
															assign node35892 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node35896 = (inp[0]) ? node35900 : node35897;
															assign node35897 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node35900 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node35903 = (inp[5]) ? node35911 : node35904;
													assign node35904 = (inp[15]) ? node35908 : node35905;
														assign node35905 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node35908 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node35911 = (inp[2]) ? node35917 : node35912;
														assign node35912 = (inp[3]) ? node35914 : 4'b1010;
															assign node35914 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node35917 = (inp[0]) ? node35921 : node35918;
															assign node35918 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node35921 = (inp[15]) ? 4'b1000 : 4'b1000;
											assign node35924 = (inp[14]) ? node35954 : node35925;
												assign node35925 = (inp[2]) ? node35941 : node35926;
													assign node35926 = (inp[0]) ? node35934 : node35927;
														assign node35927 = (inp[15]) ? node35931 : node35928;
															assign node35928 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node35931 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node35934 = (inp[15]) ? node35938 : node35935;
															assign node35935 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node35938 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node35941 = (inp[5]) ? node35949 : node35942;
														assign node35942 = (inp[0]) ? node35946 : node35943;
															assign node35943 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node35946 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node35949 = (inp[0]) ? 4'b0001 : node35950;
															assign node35950 = (inp[15]) ? 4'b0001 : 4'b0001;
												assign node35954 = (inp[0]) ? node35966 : node35955;
													assign node35955 = (inp[15]) ? node35961 : node35956;
														assign node35956 = (inp[5]) ? node35958 : 4'b0011;
															assign node35958 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node35961 = (inp[3]) ? node35963 : 4'b0001;
															assign node35963 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node35966 = (inp[15]) ? node35972 : node35967;
														assign node35967 = (inp[5]) ? node35969 : 4'b0001;
															assign node35969 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node35972 = (inp[5]) ? node35974 : 4'b0011;
															assign node35974 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node35977 = (inp[7]) ? node36031 : node35978;
											assign node35978 = (inp[2]) ? node36008 : node35979;
												assign node35979 = (inp[14]) ? node35993 : node35980;
													assign node35980 = (inp[0]) ? node35988 : node35981;
														assign node35981 = (inp[15]) ? node35985 : node35982;
															assign node35982 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node35985 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node35988 = (inp[15]) ? node35990 : 4'b1000;
															assign node35990 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node35993 = (inp[15]) ? node36001 : node35994;
														assign node35994 = (inp[0]) ? node35998 : node35995;
															assign node35995 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node35998 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node36001 = (inp[0]) ? node36005 : node36002;
															assign node36002 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node36005 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node36008 = (inp[15]) ? node36020 : node36009;
													assign node36009 = (inp[0]) ? node36015 : node36010;
														assign node36010 = (inp[5]) ? node36012 : 4'b0011;
															assign node36012 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node36015 = (inp[3]) ? node36017 : 4'b0001;
															assign node36017 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node36020 = (inp[0]) ? node36026 : node36021;
														assign node36021 = (inp[5]) ? node36023 : 4'b0001;
															assign node36023 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node36026 = (inp[3]) ? node36028 : 4'b0011;
															assign node36028 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node36031 = (inp[14]) ? node36063 : node36032;
												assign node36032 = (inp[2]) ? node36048 : node36033;
													assign node36033 = (inp[15]) ? node36041 : node36034;
														assign node36034 = (inp[0]) ? node36038 : node36035;
															assign node36035 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node36038 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node36041 = (inp[0]) ? node36045 : node36042;
															assign node36042 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node36045 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node36048 = (inp[0]) ? node36056 : node36049;
														assign node36049 = (inp[15]) ? node36053 : node36050;
															assign node36050 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node36053 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node36056 = (inp[15]) ? node36060 : node36057;
															assign node36057 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node36060 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node36063 = (inp[0]) ? node36075 : node36064;
													assign node36064 = (inp[15]) ? node36070 : node36065;
														assign node36065 = (inp[5]) ? node36067 : 4'b0010;
															assign node36067 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node36070 = (inp[5]) ? node36072 : 4'b0000;
															assign node36072 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node36075 = (inp[15]) ? node36081 : node36076;
														assign node36076 = (inp[5]) ? node36078 : 4'b0000;
															assign node36078 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node36081 = (inp[5]) ? node36083 : 4'b0010;
															assign node36083 = (inp[3]) ? 4'b0000 : 4'b0010;
								assign node36086 = (inp[1]) ? node36312 : node36087;
									assign node36087 = (inp[7]) ? node36205 : node36088;
										assign node36088 = (inp[8]) ? node36142 : node36089;
											assign node36089 = (inp[2]) ? node36119 : node36090;
												assign node36090 = (inp[14]) ? node36106 : node36091;
													assign node36091 = (inp[3]) ? node36099 : node36092;
														assign node36092 = (inp[5]) ? node36096 : node36093;
															assign node36093 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node36096 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node36099 = (inp[0]) ? node36103 : node36100;
															assign node36100 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node36103 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node36106 = (inp[5]) ? node36114 : node36107;
														assign node36107 = (inp[15]) ? node36111 : node36108;
															assign node36108 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node36111 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node36114 = (inp[3]) ? 4'b1010 : node36115;
															assign node36115 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node36119 = (inp[15]) ? node36131 : node36120;
													assign node36120 = (inp[0]) ? node36126 : node36121;
														assign node36121 = (inp[5]) ? node36123 : 4'b1010;
															assign node36123 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node36126 = (inp[5]) ? node36128 : 4'b1000;
															assign node36128 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node36131 = (inp[0]) ? node36137 : node36132;
														assign node36132 = (inp[3]) ? node36134 : 4'b1000;
															assign node36134 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node36137 = (inp[5]) ? node36139 : 4'b1010;
															assign node36139 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node36142 = (inp[14]) ? node36174 : node36143;
												assign node36143 = (inp[2]) ? node36159 : node36144;
													assign node36144 = (inp[0]) ? node36152 : node36145;
														assign node36145 = (inp[15]) ? node36149 : node36146;
															assign node36146 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node36149 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node36152 = (inp[15]) ? node36156 : node36153;
															assign node36153 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node36156 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node36159 = (inp[15]) ? node36167 : node36160;
														assign node36160 = (inp[0]) ? node36164 : node36161;
															assign node36161 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node36164 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node36167 = (inp[0]) ? node36171 : node36168;
															assign node36168 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node36171 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node36174 = (inp[3]) ? node36190 : node36175;
													assign node36175 = (inp[5]) ? node36183 : node36176;
														assign node36176 = (inp[0]) ? node36180 : node36177;
															assign node36177 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node36180 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node36183 = (inp[2]) ? node36187 : node36184;
															assign node36184 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node36187 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node36190 = (inp[0]) ? node36198 : node36191;
														assign node36191 = (inp[15]) ? node36195 : node36192;
															assign node36192 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node36195 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node36198 = (inp[2]) ? node36202 : node36199;
															assign node36199 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node36202 = (inp[5]) ? 4'b0001 : 4'b0001;
										assign node36205 = (inp[8]) ? node36261 : node36206;
											assign node36206 = (inp[2]) ? node36238 : node36207;
												assign node36207 = (inp[14]) ? node36223 : node36208;
													assign node36208 = (inp[5]) ? node36216 : node36209;
														assign node36209 = (inp[3]) ? node36213 : node36210;
															assign node36210 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node36213 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node36216 = (inp[15]) ? node36220 : node36217;
															assign node36217 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node36220 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node36223 = (inp[3]) ? node36231 : node36224;
														assign node36224 = (inp[0]) ? node36228 : node36225;
															assign node36225 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node36228 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node36231 = (inp[5]) ? node36235 : node36232;
															assign node36232 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node36235 = (inp[15]) ? 4'b0001 : 4'b0001;
												assign node36238 = (inp[5]) ? node36246 : node36239;
													assign node36239 = (inp[0]) ? node36243 : node36240;
														assign node36240 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node36243 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node36246 = (inp[3]) ? node36254 : node36247;
														assign node36247 = (inp[14]) ? node36251 : node36248;
															assign node36248 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node36251 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node36254 = (inp[15]) ? node36258 : node36255;
															assign node36255 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node36258 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node36261 = (inp[2]) ? node36289 : node36262;
												assign node36262 = (inp[14]) ? node36276 : node36263;
													assign node36263 = (inp[3]) ? node36271 : node36264;
														assign node36264 = (inp[5]) ? node36268 : node36265;
															assign node36265 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node36268 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node36271 = (inp[5]) ? 4'b0001 : node36272;
															assign node36272 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node36276 = (inp[3]) ? node36282 : node36277;
														assign node36277 = (inp[15]) ? node36279 : 4'b0010;
															assign node36279 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node36282 = (inp[5]) ? node36286 : node36283;
															assign node36283 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node36286 = (inp[0]) ? 4'b0000 : 4'b0000;
												assign node36289 = (inp[0]) ? node36301 : node36290;
													assign node36290 = (inp[15]) ? node36296 : node36291;
														assign node36291 = (inp[5]) ? node36293 : 4'b0010;
															assign node36293 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node36296 = (inp[5]) ? node36298 : 4'b0000;
															assign node36298 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node36301 = (inp[15]) ? node36307 : node36302;
														assign node36302 = (inp[3]) ? node36304 : 4'b0000;
															assign node36304 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node36307 = (inp[3]) ? node36309 : 4'b0010;
															assign node36309 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node36312 = (inp[0]) ? node36434 : node36313;
										assign node36313 = (inp[15]) ? node36375 : node36314;
											assign node36314 = (inp[5]) ? node36346 : node36315;
												assign node36315 = (inp[3]) ? node36331 : node36316;
													assign node36316 = (inp[14]) ? node36324 : node36317;
														assign node36317 = (inp[2]) ? node36321 : node36318;
															assign node36318 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node36321 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node36324 = (inp[8]) ? node36328 : node36325;
															assign node36325 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node36328 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node36331 = (inp[8]) ? node36339 : node36332;
														assign node36332 = (inp[7]) ? node36336 : node36333;
															assign node36333 = (inp[2]) ? 4'b0010 : 4'b0010;
															assign node36336 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node36339 = (inp[7]) ? node36343 : node36340;
															assign node36340 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node36343 = (inp[14]) ? 4'b0010 : 4'b0010;
												assign node36346 = (inp[3]) ? node36360 : node36347;
													assign node36347 = (inp[2]) ? node36355 : node36348;
														assign node36348 = (inp[14]) ? node36352 : node36349;
															assign node36349 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node36352 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node36355 = (inp[14]) ? 4'b0011 : node36356;
															assign node36356 = (inp[7]) ? 4'b0010 : 4'b0010;
													assign node36360 = (inp[2]) ? node36368 : node36361;
														assign node36361 = (inp[7]) ? node36365 : node36362;
															assign node36362 = (inp[14]) ? 4'b0000 : 4'b0000;
															assign node36365 = (inp[14]) ? 4'b0000 : 4'b0000;
														assign node36368 = (inp[14]) ? node36372 : node36369;
															assign node36369 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node36372 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node36375 = (inp[5]) ? node36407 : node36376;
												assign node36376 = (inp[3]) ? node36392 : node36377;
													assign node36377 = (inp[14]) ? node36385 : node36378;
														assign node36378 = (inp[8]) ? node36382 : node36379;
															assign node36379 = (inp[2]) ? 4'b0000 : 4'b0000;
															assign node36382 = (inp[7]) ? 4'b0000 : 4'b0000;
														assign node36385 = (inp[7]) ? node36389 : node36386;
															assign node36386 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node36389 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node36392 = (inp[8]) ? node36400 : node36393;
														assign node36393 = (inp[7]) ? node36397 : node36394;
															assign node36394 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node36397 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node36400 = (inp[7]) ? node36404 : node36401;
															assign node36401 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node36404 = (inp[2]) ? 4'b0000 : 4'b0000;
												assign node36407 = (inp[3]) ? node36421 : node36408;
													assign node36408 = (inp[14]) ? node36416 : node36409;
														assign node36409 = (inp[2]) ? node36413 : node36410;
															assign node36410 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node36413 = (inp[7]) ? 4'b0000 : 4'b0000;
														assign node36416 = (inp[2]) ? node36418 : 4'b0001;
															assign node36418 = (inp[7]) ? 4'b0000 : 4'b0000;
													assign node36421 = (inp[7]) ? node36427 : node36422;
														assign node36422 = (inp[8]) ? 4'b0011 : node36423;
															assign node36423 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node36427 = (inp[8]) ? node36431 : node36428;
															assign node36428 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node36431 = (inp[14]) ? 4'b0010 : 4'b0010;
										assign node36434 = (inp[15]) ? node36490 : node36435;
											assign node36435 = (inp[3]) ? node36459 : node36436;
												assign node36436 = (inp[7]) ? node36448 : node36437;
													assign node36437 = (inp[8]) ? node36443 : node36438;
														assign node36438 = (inp[14]) ? 4'b0000 : node36439;
															assign node36439 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node36443 = (inp[2]) ? 4'b0001 : node36444;
															assign node36444 = (inp[14]) ? 4'b0001 : 4'b0000;
													assign node36448 = (inp[8]) ? node36454 : node36449;
														assign node36449 = (inp[14]) ? 4'b0001 : node36450;
															assign node36450 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node36454 = (inp[2]) ? 4'b0000 : node36455;
															assign node36455 = (inp[14]) ? 4'b0000 : 4'b0001;
												assign node36459 = (inp[5]) ? node36475 : node36460;
													assign node36460 = (inp[8]) ? node36468 : node36461;
														assign node36461 = (inp[7]) ? node36465 : node36462;
															assign node36462 = (inp[2]) ? 4'b0000 : 4'b0000;
															assign node36465 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node36468 = (inp[7]) ? node36472 : node36469;
															assign node36469 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node36472 = (inp[14]) ? 4'b0000 : 4'b0000;
													assign node36475 = (inp[8]) ? node36483 : node36476;
														assign node36476 = (inp[7]) ? node36480 : node36477;
															assign node36477 = (inp[2]) ? 4'b0010 : 4'b0010;
															assign node36480 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node36483 = (inp[7]) ? node36487 : node36484;
															assign node36484 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node36487 = (inp[14]) ? 4'b0010 : 4'b0010;
											assign node36490 = (inp[5]) ? node36514 : node36491;
												assign node36491 = (inp[7]) ? node36503 : node36492;
													assign node36492 = (inp[8]) ? node36498 : node36493;
														assign node36493 = (inp[2]) ? 4'b0010 : node36494;
															assign node36494 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node36498 = (inp[14]) ? 4'b0011 : node36499;
															assign node36499 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node36503 = (inp[8]) ? node36509 : node36504;
														assign node36504 = (inp[2]) ? 4'b0011 : node36505;
															assign node36505 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node36509 = (inp[14]) ? 4'b0010 : node36510;
															assign node36510 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node36514 = (inp[3]) ? node36530 : node36515;
													assign node36515 = (inp[2]) ? node36523 : node36516;
														assign node36516 = (inp[7]) ? node36520 : node36517;
															assign node36517 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node36520 = (inp[14]) ? 4'b0010 : 4'b0010;
														assign node36523 = (inp[14]) ? node36527 : node36524;
															assign node36524 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node36527 = (inp[8]) ? 4'b0010 : 4'b0010;
													assign node36530 = (inp[2]) ? node36538 : node36531;
														assign node36531 = (inp[7]) ? node36535 : node36532;
															assign node36532 = (inp[14]) ? 4'b0000 : 4'b0000;
															assign node36535 = (inp[14]) ? 4'b0000 : 4'b0000;
														assign node36538 = (inp[14]) ? node36542 : node36539;
															assign node36539 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node36542 = (inp[8]) ? 4'b0000 : 4'b0000;
							assign node36545 = (inp[13]) ? node36979 : node36546;
								assign node36546 = (inp[1]) ? node36766 : node36547;
									assign node36547 = (inp[7]) ? node36653 : node36548;
										assign node36548 = (inp[8]) ? node36600 : node36549;
											assign node36549 = (inp[2]) ? node36577 : node36550;
												assign node36550 = (inp[14]) ? node36564 : node36551;
													assign node36551 = (inp[15]) ? node36557 : node36552;
														assign node36552 = (inp[0]) ? 4'b0001 : node36553;
															assign node36553 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node36557 = (inp[0]) ? node36561 : node36558;
															assign node36558 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node36561 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node36564 = (inp[15]) ? node36572 : node36565;
														assign node36565 = (inp[0]) ? node36569 : node36566;
															assign node36566 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node36569 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node36572 = (inp[0]) ? node36574 : 4'b0000;
															assign node36574 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node36577 = (inp[0]) ? node36589 : node36578;
													assign node36578 = (inp[15]) ? node36584 : node36579;
														assign node36579 = (inp[5]) ? node36581 : 4'b0010;
															assign node36581 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node36584 = (inp[3]) ? node36586 : 4'b0000;
															assign node36586 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node36589 = (inp[15]) ? node36595 : node36590;
														assign node36590 = (inp[5]) ? node36592 : 4'b0000;
															assign node36592 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node36595 = (inp[5]) ? node36597 : 4'b0010;
															assign node36597 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node36600 = (inp[2]) ? node36630 : node36601;
												assign node36601 = (inp[14]) ? node36617 : node36602;
													assign node36602 = (inp[0]) ? node36610 : node36603;
														assign node36603 = (inp[15]) ? node36607 : node36604;
															assign node36604 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node36607 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node36610 = (inp[15]) ? node36614 : node36611;
															assign node36611 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node36614 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node36617 = (inp[3]) ? node36623 : node36618;
														assign node36618 = (inp[15]) ? node36620 : 4'b0001;
															assign node36620 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node36623 = (inp[0]) ? node36627 : node36624;
															assign node36624 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node36627 = (inp[5]) ? 4'b0001 : 4'b0001;
												assign node36630 = (inp[0]) ? node36642 : node36631;
													assign node36631 = (inp[15]) ? node36637 : node36632;
														assign node36632 = (inp[5]) ? node36634 : 4'b0011;
															assign node36634 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node36637 = (inp[5]) ? node36639 : 4'b0001;
															assign node36639 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node36642 = (inp[15]) ? node36648 : node36643;
														assign node36643 = (inp[5]) ? node36645 : 4'b0001;
															assign node36645 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node36648 = (inp[3]) ? node36650 : 4'b0011;
															assign node36650 = (inp[5]) ? 4'b0001 : 4'b0011;
										assign node36653 = (inp[8]) ? node36711 : node36654;
											assign node36654 = (inp[2]) ? node36682 : node36655;
												assign node36655 = (inp[14]) ? node36671 : node36656;
													assign node36656 = (inp[15]) ? node36664 : node36657;
														assign node36657 = (inp[0]) ? node36661 : node36658;
															assign node36658 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node36661 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node36664 = (inp[0]) ? node36668 : node36665;
															assign node36665 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node36668 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node36671 = (inp[15]) ? node36677 : node36672;
														assign node36672 = (inp[0]) ? node36674 : 4'b0011;
															assign node36674 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node36677 = (inp[0]) ? node36679 : 4'b0001;
															assign node36679 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node36682 = (inp[14]) ? node36698 : node36683;
													assign node36683 = (inp[3]) ? node36691 : node36684;
														assign node36684 = (inp[5]) ? node36688 : node36685;
															assign node36685 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node36688 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node36691 = (inp[0]) ? node36695 : node36692;
															assign node36692 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node36695 = (inp[5]) ? 4'b0001 : 4'b0001;
													assign node36698 = (inp[0]) ? node36706 : node36699;
														assign node36699 = (inp[15]) ? node36703 : node36700;
															assign node36700 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node36703 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node36706 = (inp[15]) ? 4'b0011 : node36707;
															assign node36707 = (inp[3]) ? 4'b0011 : 4'b0001;
											assign node36711 = (inp[14]) ? node36743 : node36712;
												assign node36712 = (inp[2]) ? node36728 : node36713;
													assign node36713 = (inp[5]) ? node36721 : node36714;
														assign node36714 = (inp[15]) ? node36718 : node36715;
															assign node36715 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node36718 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node36721 = (inp[15]) ? node36725 : node36722;
															assign node36722 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node36725 = (inp[3]) ? 4'b0001 : 4'b0001;
													assign node36728 = (inp[3]) ? node36736 : node36729;
														assign node36729 = (inp[5]) ? node36733 : node36730;
															assign node36730 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node36733 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node36736 = (inp[5]) ? node36740 : node36737;
															assign node36737 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node36740 = (inp[0]) ? 4'b0000 : 4'b0000;
												assign node36743 = (inp[5]) ? node36751 : node36744;
													assign node36744 = (inp[15]) ? node36748 : node36745;
														assign node36745 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node36748 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node36751 = (inp[3]) ? node36759 : node36752;
														assign node36752 = (inp[15]) ? node36756 : node36753;
															assign node36753 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node36756 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node36759 = (inp[15]) ? node36763 : node36760;
															assign node36760 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node36763 = (inp[0]) ? 4'b0000 : 4'b0010;
									assign node36766 = (inp[7]) ? node36874 : node36767;
										assign node36767 = (inp[8]) ? node36821 : node36768;
											assign node36768 = (inp[2]) ? node36798 : node36769;
												assign node36769 = (inp[14]) ? node36783 : node36770;
													assign node36770 = (inp[5]) ? node36778 : node36771;
														assign node36771 = (inp[3]) ? node36775 : node36772;
															assign node36772 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node36775 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node36778 = (inp[3]) ? node36780 : 4'b0001;
															assign node36780 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node36783 = (inp[5]) ? node36791 : node36784;
														assign node36784 = (inp[0]) ? node36788 : node36785;
															assign node36785 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node36788 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node36791 = (inp[3]) ? node36795 : node36792;
															assign node36792 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node36795 = (inp[0]) ? 4'b0000 : 4'b0000;
												assign node36798 = (inp[15]) ? node36810 : node36799;
													assign node36799 = (inp[0]) ? node36805 : node36800;
														assign node36800 = (inp[5]) ? node36802 : 4'b0010;
															assign node36802 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node36805 = (inp[5]) ? node36807 : 4'b0000;
															assign node36807 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node36810 = (inp[0]) ? node36816 : node36811;
														assign node36811 = (inp[5]) ? node36813 : 4'b0000;
															assign node36813 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node36816 = (inp[3]) ? node36818 : 4'b0010;
															assign node36818 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node36821 = (inp[2]) ? node36851 : node36822;
												assign node36822 = (inp[14]) ? node36838 : node36823;
													assign node36823 = (inp[15]) ? node36831 : node36824;
														assign node36824 = (inp[0]) ? node36828 : node36825;
															assign node36825 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node36828 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node36831 = (inp[0]) ? node36835 : node36832;
															assign node36832 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node36835 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node36838 = (inp[0]) ? node36844 : node36839;
														assign node36839 = (inp[15]) ? node36841 : 4'b1101;
															assign node36841 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node36844 = (inp[15]) ? node36848 : node36845;
															assign node36845 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node36848 = (inp[3]) ? 4'b1101 : 4'b1101;
												assign node36851 = (inp[3]) ? node36867 : node36852;
													assign node36852 = (inp[0]) ? node36860 : node36853;
														assign node36853 = (inp[14]) ? node36857 : node36854;
															assign node36854 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node36857 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node36860 = (inp[14]) ? node36864 : node36861;
															assign node36861 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node36864 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node36867 = (inp[0]) ? node36871 : node36868;
														assign node36868 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node36871 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node36874 = (inp[8]) ? node36924 : node36875;
											assign node36875 = (inp[14]) ? node36901 : node36876;
												assign node36876 = (inp[2]) ? node36890 : node36877;
													assign node36877 = (inp[5]) ? node36883 : node36878;
														assign node36878 = (inp[0]) ? 4'b0010 : node36879;
															assign node36879 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node36883 = (inp[0]) ? node36887 : node36884;
															assign node36884 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node36887 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node36890 = (inp[15]) ? node36896 : node36891;
														assign node36891 = (inp[0]) ? 4'b1111 : node36892;
															assign node36892 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node36896 = (inp[0]) ? 4'b1101 : node36897;
															assign node36897 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node36901 = (inp[15]) ? node36913 : node36902;
													assign node36902 = (inp[0]) ? node36908 : node36903;
														assign node36903 = (inp[5]) ? 4'b1101 : node36904;
															assign node36904 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node36908 = (inp[5]) ? 4'b1111 : node36909;
															assign node36909 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node36913 = (inp[0]) ? node36919 : node36914;
														assign node36914 = (inp[5]) ? 4'b1111 : node36915;
															assign node36915 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node36919 = (inp[3]) ? 4'b1101 : node36920;
															assign node36920 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node36924 = (inp[14]) ? node36948 : node36925;
												assign node36925 = (inp[2]) ? node36937 : node36926;
													assign node36926 = (inp[0]) ? node36932 : node36927;
														assign node36927 = (inp[15]) ? 4'b1111 : node36928;
															assign node36928 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node36932 = (inp[5]) ? 4'b1101 : node36933;
															assign node36933 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node36937 = (inp[15]) ? node36943 : node36938;
														assign node36938 = (inp[0]) ? node36940 : 4'b1100;
															assign node36940 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node36943 = (inp[0]) ? node36945 : 4'b1110;
															assign node36945 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node36948 = (inp[3]) ? node36964 : node36949;
													assign node36949 = (inp[0]) ? node36957 : node36950;
														assign node36950 = (inp[2]) ? node36954 : node36951;
															assign node36951 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node36954 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node36957 = (inp[15]) ? node36961 : node36958;
															assign node36958 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node36961 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node36964 = (inp[5]) ? node36972 : node36965;
														assign node36965 = (inp[2]) ? node36969 : node36966;
															assign node36966 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node36969 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node36972 = (inp[15]) ? node36976 : node36973;
															assign node36973 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node36976 = (inp[0]) ? 4'b1100 : 4'b1110;
								assign node36979 = (inp[1]) ? node37209 : node36980;
									assign node36980 = (inp[7]) ? node37092 : node36981;
										assign node36981 = (inp[8]) ? node37031 : node36982;
											assign node36982 = (inp[14]) ? node37014 : node36983;
												assign node36983 = (inp[2]) ? node36999 : node36984;
													assign node36984 = (inp[5]) ? node36992 : node36985;
														assign node36985 = (inp[15]) ? node36989 : node36986;
															assign node36986 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node36989 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node36992 = (inp[3]) ? node36996 : node36993;
															assign node36993 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node36996 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node36999 = (inp[5]) ? node37007 : node37000;
														assign node37000 = (inp[3]) ? node37004 : node37001;
															assign node37001 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node37004 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node37007 = (inp[3]) ? node37011 : node37008;
															assign node37008 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node37011 = (inp[15]) ? 4'b0000 : 4'b0000;
												assign node37014 = (inp[0]) ? node37020 : node37015;
													assign node37015 = (inp[3]) ? 4'b0010 : node37016;
														assign node37016 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node37020 = (inp[15]) ? node37026 : node37021;
														assign node37021 = (inp[3]) ? node37023 : 4'b0000;
															assign node37023 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node37026 = (inp[5]) ? node37028 : 4'b0010;
															assign node37028 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node37031 = (inp[2]) ? node37063 : node37032;
												assign node37032 = (inp[14]) ? node37048 : node37033;
													assign node37033 = (inp[3]) ? node37041 : node37034;
														assign node37034 = (inp[15]) ? node37038 : node37035;
															assign node37035 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node37038 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node37041 = (inp[0]) ? node37045 : node37042;
															assign node37042 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node37045 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node37048 = (inp[15]) ? node37056 : node37049;
														assign node37049 = (inp[0]) ? node37053 : node37050;
															assign node37050 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node37053 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node37056 = (inp[0]) ? node37060 : node37057;
															assign node37057 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node37060 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node37063 = (inp[14]) ? node37077 : node37064;
													assign node37064 = (inp[0]) ? node37072 : node37065;
														assign node37065 = (inp[15]) ? node37069 : node37066;
															assign node37066 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node37069 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node37072 = (inp[15]) ? node37074 : 4'b1111;
															assign node37074 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node37077 = (inp[5]) ? node37085 : node37078;
														assign node37078 = (inp[15]) ? node37082 : node37079;
															assign node37079 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node37082 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node37085 = (inp[15]) ? node37089 : node37086;
															assign node37086 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node37089 = (inp[0]) ? 4'b1101 : 4'b1111;
										assign node37092 = (inp[8]) ? node37156 : node37093;
											assign node37093 = (inp[14]) ? node37125 : node37094;
												assign node37094 = (inp[2]) ? node37110 : node37095;
													assign node37095 = (inp[3]) ? node37103 : node37096;
														assign node37096 = (inp[5]) ? node37100 : node37097;
															assign node37097 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node37100 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node37103 = (inp[5]) ? node37107 : node37104;
															assign node37104 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node37107 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node37110 = (inp[5]) ? node37118 : node37111;
														assign node37111 = (inp[3]) ? node37115 : node37112;
															assign node37112 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node37115 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node37118 = (inp[15]) ? node37122 : node37119;
															assign node37119 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node37122 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node37125 = (inp[5]) ? node37141 : node37126;
													assign node37126 = (inp[15]) ? node37134 : node37127;
														assign node37127 = (inp[3]) ? node37131 : node37128;
															assign node37128 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node37131 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node37134 = (inp[3]) ? node37138 : node37135;
															assign node37135 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node37138 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node37141 = (inp[3]) ? node37149 : node37142;
														assign node37142 = (inp[2]) ? node37146 : node37143;
															assign node37143 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node37146 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node37149 = (inp[0]) ? node37153 : node37150;
															assign node37150 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node37153 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node37156 = (inp[2]) ? node37186 : node37157;
												assign node37157 = (inp[14]) ? node37171 : node37158;
													assign node37158 = (inp[3]) ? node37164 : node37159;
														assign node37159 = (inp[5]) ? node37161 : 4'b1101;
															assign node37161 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node37164 = (inp[5]) ? node37168 : node37165;
															assign node37165 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node37168 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node37171 = (inp[15]) ? node37179 : node37172;
														assign node37172 = (inp[0]) ? node37176 : node37173;
															assign node37173 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node37176 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node37179 = (inp[0]) ? node37183 : node37180;
															assign node37180 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node37183 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node37186 = (inp[5]) ? node37202 : node37187;
													assign node37187 = (inp[14]) ? node37195 : node37188;
														assign node37188 = (inp[0]) ? node37192 : node37189;
															assign node37189 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node37192 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node37195 = (inp[3]) ? node37199 : node37196;
															assign node37196 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node37199 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node37202 = (inp[0]) ? node37206 : node37203;
														assign node37203 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node37206 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node37209 = (inp[3]) ? node37329 : node37210;
										assign node37210 = (inp[7]) ? node37270 : node37211;
											assign node37211 = (inp[8]) ? node37241 : node37212;
												assign node37212 = (inp[14]) ? node37226 : node37213;
													assign node37213 = (inp[2]) ? node37221 : node37214;
														assign node37214 = (inp[0]) ? node37218 : node37215;
															assign node37215 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node37218 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node37221 = (inp[5]) ? 4'b1110 : node37222;
															assign node37222 = (inp[0]) ? 4'b1100 : 4'b1100;
													assign node37226 = (inp[2]) ? node37234 : node37227;
														assign node37227 = (inp[0]) ? node37231 : node37228;
															assign node37228 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node37231 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node37234 = (inp[5]) ? node37238 : node37235;
															assign node37235 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node37238 = (inp[15]) ? 4'b1100 : 4'b1100;
												assign node37241 = (inp[14]) ? node37255 : node37242;
													assign node37242 = (inp[2]) ? node37250 : node37243;
														assign node37243 = (inp[15]) ? node37247 : node37244;
															assign node37244 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node37247 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node37250 = (inp[5]) ? 4'b1111 : node37251;
															assign node37251 = (inp[0]) ? 4'b1101 : 4'b1101;
													assign node37255 = (inp[0]) ? node37263 : node37256;
														assign node37256 = (inp[15]) ? node37260 : node37257;
															assign node37257 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node37260 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node37263 = (inp[15]) ? node37267 : node37264;
															assign node37264 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node37267 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node37270 = (inp[8]) ? node37298 : node37271;
												assign node37271 = (inp[14]) ? node37285 : node37272;
													assign node37272 = (inp[2]) ? node37280 : node37273;
														assign node37273 = (inp[15]) ? node37277 : node37274;
															assign node37274 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node37277 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node37280 = (inp[0]) ? 4'b1101 : node37281;
															assign node37281 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node37285 = (inp[2]) ? node37293 : node37286;
														assign node37286 = (inp[0]) ? node37290 : node37287;
															assign node37287 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node37290 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node37293 = (inp[15]) ? node37295 : 4'b1101;
															assign node37295 = (inp[5]) ? 4'b1101 : 4'b1101;
												assign node37298 = (inp[14]) ? node37314 : node37299;
													assign node37299 = (inp[2]) ? node37307 : node37300;
														assign node37300 = (inp[15]) ? node37304 : node37301;
															assign node37301 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node37304 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node37307 = (inp[0]) ? node37311 : node37308;
															assign node37308 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node37311 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node37314 = (inp[15]) ? node37322 : node37315;
														assign node37315 = (inp[0]) ? node37319 : node37316;
															assign node37316 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node37319 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node37322 = (inp[0]) ? node37326 : node37323;
															assign node37323 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node37326 = (inp[5]) ? 4'b1100 : 4'b1110;
										assign node37329 = (inp[2]) ? node37389 : node37330;
											assign node37330 = (inp[8]) ? node37358 : node37331;
												assign node37331 = (inp[5]) ? node37345 : node37332;
													assign node37332 = (inp[0]) ? node37340 : node37333;
														assign node37333 = (inp[15]) ? node37337 : node37334;
															assign node37334 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node37337 = (inp[7]) ? 4'b1110 : 4'b1110;
														assign node37340 = (inp[15]) ? 4'b1101 : node37341;
															assign node37341 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node37345 = (inp[0]) ? node37351 : node37346;
														assign node37346 = (inp[15]) ? 4'b1111 : node37347;
															assign node37347 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node37351 = (inp[15]) ? node37355 : node37352;
															assign node37352 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node37355 = (inp[14]) ? 4'b1100 : 4'b1100;
												assign node37358 = (inp[15]) ? node37374 : node37359;
													assign node37359 = (inp[0]) ? node37367 : node37360;
														assign node37360 = (inp[14]) ? node37364 : node37361;
															assign node37361 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node37364 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node37367 = (inp[14]) ? node37371 : node37368;
															assign node37368 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node37371 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node37374 = (inp[0]) ? node37382 : node37375;
														assign node37375 = (inp[14]) ? node37379 : node37376;
															assign node37376 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node37379 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node37382 = (inp[7]) ? node37386 : node37383;
															assign node37383 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node37386 = (inp[14]) ? 4'b1100 : 4'b1101;
											assign node37389 = (inp[0]) ? node37421 : node37390;
												assign node37390 = (inp[15]) ? node37406 : node37391;
													assign node37391 = (inp[14]) ? node37399 : node37392;
														assign node37392 = (inp[5]) ? node37396 : node37393;
															assign node37393 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node37396 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node37399 = (inp[7]) ? node37403 : node37400;
															assign node37400 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node37403 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node37406 = (inp[14]) ? node37414 : node37407;
														assign node37407 = (inp[5]) ? node37411 : node37408;
															assign node37408 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node37411 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node37414 = (inp[8]) ? node37418 : node37415;
															assign node37415 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node37418 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node37421 = (inp[15]) ? node37429 : node37422;
													assign node37422 = (inp[7]) ? node37426 : node37423;
														assign node37423 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node37426 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node37429 = (inp[8]) ? node37433 : node37430;
														assign node37430 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node37433 = (inp[7]) ? 4'b1100 : 4'b1101;
						assign node37436 = (inp[6]) ? node38326 : node37437;
							assign node37437 = (inp[13]) ? node37889 : node37438;
								assign node37438 = (inp[1]) ? node37668 : node37439;
									assign node37439 = (inp[5]) ? node37545 : node37440;
										assign node37440 = (inp[8]) ? node37494 : node37441;
											assign node37441 = (inp[7]) ? node37465 : node37442;
												assign node37442 = (inp[14]) ? node37458 : node37443;
													assign node37443 = (inp[2]) ? node37451 : node37444;
														assign node37444 = (inp[3]) ? node37448 : node37445;
															assign node37445 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node37448 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node37451 = (inp[0]) ? node37455 : node37452;
															assign node37452 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node37455 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node37458 = (inp[0]) ? node37462 : node37459;
														assign node37459 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node37462 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node37465 = (inp[14]) ? node37481 : node37466;
													assign node37466 = (inp[2]) ? node37474 : node37467;
														assign node37467 = (inp[0]) ? node37471 : node37468;
															assign node37468 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node37471 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node37474 = (inp[3]) ? node37478 : node37475;
															assign node37475 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node37478 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node37481 = (inp[2]) ? node37489 : node37482;
														assign node37482 = (inp[15]) ? node37486 : node37483;
															assign node37483 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node37486 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node37489 = (inp[3]) ? node37491 : 4'b0001;
															assign node37491 = (inp[15]) ? 4'b0001 : 4'b0001;
											assign node37494 = (inp[7]) ? node37518 : node37495;
												assign node37495 = (inp[2]) ? node37511 : node37496;
													assign node37496 = (inp[14]) ? node37504 : node37497;
														assign node37497 = (inp[0]) ? node37501 : node37498;
															assign node37498 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node37501 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node37504 = (inp[15]) ? node37508 : node37505;
															assign node37505 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node37508 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node37511 = (inp[0]) ? node37515 : node37512;
														assign node37512 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node37515 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node37518 = (inp[2]) ? node37532 : node37519;
													assign node37519 = (inp[14]) ? node37527 : node37520;
														assign node37520 = (inp[15]) ? node37524 : node37521;
															assign node37521 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node37524 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node37527 = (inp[15]) ? 4'b0010 : node37528;
															assign node37528 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node37532 = (inp[3]) ? node37538 : node37533;
														assign node37533 = (inp[14]) ? node37535 : 4'b0010;
															assign node37535 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node37538 = (inp[0]) ? node37542 : node37539;
															assign node37539 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node37542 = (inp[15]) ? 4'b0010 : 4'b0000;
										assign node37545 = (inp[0]) ? node37607 : node37546;
											assign node37546 = (inp[14]) ? node37576 : node37547;
												assign node37547 = (inp[3]) ? node37561 : node37548;
													assign node37548 = (inp[15]) ? node37554 : node37549;
														assign node37549 = (inp[8]) ? 4'b0010 : node37550;
															assign node37550 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node37554 = (inp[8]) ? node37558 : node37555;
															assign node37555 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node37558 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node37561 = (inp[15]) ? node37569 : node37562;
														assign node37562 = (inp[8]) ? node37566 : node37563;
															assign node37563 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node37566 = (inp[7]) ? 4'b0000 : 4'b0000;
														assign node37569 = (inp[8]) ? node37573 : node37570;
															assign node37570 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node37573 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node37576 = (inp[7]) ? node37592 : node37577;
													assign node37577 = (inp[8]) ? node37585 : node37578;
														assign node37578 = (inp[3]) ? node37582 : node37579;
															assign node37579 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node37582 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node37585 = (inp[15]) ? node37589 : node37586;
															assign node37586 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node37589 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node37592 = (inp[8]) ? node37600 : node37593;
														assign node37593 = (inp[15]) ? node37597 : node37594;
															assign node37594 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node37597 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node37600 = (inp[2]) ? node37604 : node37601;
															assign node37601 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node37604 = (inp[3]) ? 4'b0000 : 4'b0000;
											assign node37607 = (inp[2]) ? node37639 : node37608;
												assign node37608 = (inp[7]) ? node37624 : node37609;
													assign node37609 = (inp[14]) ? node37617 : node37610;
														assign node37610 = (inp[8]) ? node37614 : node37611;
															assign node37611 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node37614 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node37617 = (inp[8]) ? node37621 : node37618;
															assign node37618 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node37621 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node37624 = (inp[15]) ? node37632 : node37625;
														assign node37625 = (inp[3]) ? node37629 : node37626;
															assign node37626 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node37629 = (inp[14]) ? 4'b0010 : 4'b0010;
														assign node37632 = (inp[3]) ? node37636 : node37633;
															assign node37633 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node37636 = (inp[14]) ? 4'b0000 : 4'b0000;
												assign node37639 = (inp[3]) ? node37655 : node37640;
													assign node37640 = (inp[15]) ? node37648 : node37641;
														assign node37641 = (inp[14]) ? node37645 : node37642;
															assign node37642 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node37645 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node37648 = (inp[7]) ? node37652 : node37649;
															assign node37649 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node37652 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node37655 = (inp[15]) ? node37663 : node37656;
														assign node37656 = (inp[8]) ? node37660 : node37657;
															assign node37657 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node37660 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node37663 = (inp[14]) ? 4'b0000 : node37664;
															assign node37664 = (inp[8]) ? 4'b0000 : 4'b0000;
									assign node37668 = (inp[8]) ? node37780 : node37669;
										assign node37669 = (inp[7]) ? node37729 : node37670;
											assign node37670 = (inp[2]) ? node37698 : node37671;
												assign node37671 = (inp[14]) ? node37685 : node37672;
													assign node37672 = (inp[5]) ? node37680 : node37673;
														assign node37673 = (inp[0]) ? node37677 : node37674;
															assign node37674 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node37677 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node37680 = (inp[15]) ? 4'b0011 : node37681;
															assign node37681 = (inp[3]) ? 4'b0001 : 4'b0001;
													assign node37685 = (inp[15]) ? node37693 : node37686;
														assign node37686 = (inp[0]) ? node37690 : node37687;
															assign node37687 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node37690 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node37693 = (inp[5]) ? node37695 : 4'b0000;
															assign node37695 = (inp[0]) ? 4'b0000 : 4'b0000;
												assign node37698 = (inp[3]) ? node37714 : node37699;
													assign node37699 = (inp[14]) ? node37707 : node37700;
														assign node37700 = (inp[5]) ? node37704 : node37701;
															assign node37701 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node37704 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node37707 = (inp[15]) ? node37711 : node37708;
															assign node37708 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node37711 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node37714 = (inp[15]) ? node37722 : node37715;
														assign node37715 = (inp[0]) ? node37719 : node37716;
															assign node37716 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node37719 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node37722 = (inp[5]) ? node37726 : node37723;
															assign node37723 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node37726 = (inp[0]) ? 4'b0000 : 4'b0010;
											assign node37729 = (inp[2]) ? node37759 : node37730;
												assign node37730 = (inp[14]) ? node37746 : node37731;
													assign node37731 = (inp[0]) ? node37739 : node37732;
														assign node37732 = (inp[15]) ? node37736 : node37733;
															assign node37733 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node37736 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node37739 = (inp[15]) ? node37743 : node37740;
															assign node37740 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node37743 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node37746 = (inp[5]) ? node37754 : node37747;
														assign node37747 = (inp[15]) ? node37751 : node37748;
															assign node37748 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node37751 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node37754 = (inp[0]) ? 4'b1111 : node37755;
															assign node37755 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node37759 = (inp[3]) ? node37773 : node37760;
													assign node37760 = (inp[5]) ? node37766 : node37761;
														assign node37761 = (inp[15]) ? 4'b1101 : node37762;
															assign node37762 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node37766 = (inp[0]) ? node37770 : node37767;
															assign node37767 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node37770 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node37773 = (inp[15]) ? node37777 : node37774;
														assign node37774 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node37777 = (inp[0]) ? 4'b1101 : 4'b1111;
										assign node37780 = (inp[7]) ? node37834 : node37781;
											assign node37781 = (inp[14]) ? node37811 : node37782;
												assign node37782 = (inp[2]) ? node37798 : node37783;
													assign node37783 = (inp[0]) ? node37791 : node37784;
														assign node37784 = (inp[15]) ? node37788 : node37785;
															assign node37785 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node37788 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node37791 = (inp[15]) ? node37795 : node37792;
															assign node37792 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node37795 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node37798 = (inp[5]) ? node37804 : node37799;
														assign node37799 = (inp[3]) ? 4'b1111 : node37800;
															assign node37800 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node37804 = (inp[15]) ? node37808 : node37805;
															assign node37805 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node37808 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node37811 = (inp[15]) ? node37823 : node37812;
													assign node37812 = (inp[0]) ? node37818 : node37813;
														assign node37813 = (inp[5]) ? 4'b1101 : node37814;
															assign node37814 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node37818 = (inp[5]) ? 4'b1111 : node37819;
															assign node37819 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node37823 = (inp[0]) ? node37829 : node37824;
														assign node37824 = (inp[3]) ? 4'b1111 : node37825;
															assign node37825 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node37829 = (inp[5]) ? 4'b1101 : node37830;
															assign node37830 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node37834 = (inp[2]) ? node37866 : node37835;
												assign node37835 = (inp[14]) ? node37851 : node37836;
													assign node37836 = (inp[3]) ? node37844 : node37837;
														assign node37837 = (inp[5]) ? node37841 : node37838;
															assign node37838 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node37841 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node37844 = (inp[5]) ? node37848 : node37845;
															assign node37845 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node37848 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node37851 = (inp[15]) ? node37859 : node37852;
														assign node37852 = (inp[0]) ? node37856 : node37853;
															assign node37853 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node37856 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node37859 = (inp[0]) ? node37863 : node37860;
															assign node37860 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node37863 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node37866 = (inp[0]) ? node37878 : node37867;
													assign node37867 = (inp[15]) ? node37873 : node37868;
														assign node37868 = (inp[5]) ? 4'b1100 : node37869;
															assign node37869 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node37873 = (inp[5]) ? 4'b1110 : node37874;
															assign node37874 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node37878 = (inp[15]) ? node37884 : node37879;
														assign node37879 = (inp[5]) ? 4'b1110 : node37880;
															assign node37880 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node37884 = (inp[3]) ? 4'b1100 : node37885;
															assign node37885 = (inp[5]) ? 4'b1100 : 4'b1110;
								assign node37889 = (inp[1]) ? node38113 : node37890;
									assign node37890 = (inp[8]) ? node37998 : node37891;
										assign node37891 = (inp[7]) ? node37947 : node37892;
											assign node37892 = (inp[14]) ? node37918 : node37893;
												assign node37893 = (inp[2]) ? node37907 : node37894;
													assign node37894 = (inp[3]) ? node37902 : node37895;
														assign node37895 = (inp[5]) ? node37899 : node37896;
															assign node37896 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node37899 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node37902 = (inp[5]) ? 4'b0001 : node37903;
															assign node37903 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node37907 = (inp[0]) ? node37911 : node37908;
														assign node37908 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node37911 = (inp[15]) ? node37915 : node37912;
															assign node37912 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node37915 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node37918 = (inp[2]) ? node37934 : node37919;
													assign node37919 = (inp[0]) ? node37927 : node37920;
														assign node37920 = (inp[15]) ? node37924 : node37921;
															assign node37921 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node37924 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node37927 = (inp[15]) ? node37931 : node37928;
															assign node37928 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node37931 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node37934 = (inp[5]) ? node37942 : node37935;
														assign node37935 = (inp[3]) ? node37939 : node37936;
															assign node37936 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node37939 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node37942 = (inp[15]) ? 4'b0000 : node37943;
															assign node37943 = (inp[0]) ? 4'b0000 : 4'b0000;
											assign node37947 = (inp[14]) ? node37975 : node37948;
												assign node37948 = (inp[2]) ? node37964 : node37949;
													assign node37949 = (inp[5]) ? node37957 : node37950;
														assign node37950 = (inp[0]) ? node37954 : node37951;
															assign node37951 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node37954 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node37957 = (inp[3]) ? node37961 : node37958;
															assign node37958 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node37961 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node37964 = (inp[0]) ? node37970 : node37965;
														assign node37965 = (inp[15]) ? 4'b1111 : node37966;
															assign node37966 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node37970 = (inp[5]) ? 4'b1101 : node37971;
															assign node37971 = (inp[15]) ? 4'b1101 : 4'b1101;
												assign node37975 = (inp[0]) ? node37987 : node37976;
													assign node37976 = (inp[15]) ? node37982 : node37977;
														assign node37977 = (inp[3]) ? 4'b1101 : node37978;
															assign node37978 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node37982 = (inp[3]) ? 4'b1111 : node37983;
															assign node37983 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node37987 = (inp[15]) ? node37993 : node37988;
														assign node37988 = (inp[5]) ? 4'b1111 : node37989;
															assign node37989 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node37993 = (inp[5]) ? 4'b1101 : node37994;
															assign node37994 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node37998 = (inp[7]) ? node38050 : node37999;
											assign node37999 = (inp[2]) ? node38027 : node38000;
												assign node38000 = (inp[14]) ? node38014 : node38001;
													assign node38001 = (inp[0]) ? node38009 : node38002;
														assign node38002 = (inp[15]) ? node38006 : node38003;
															assign node38003 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node38006 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node38009 = (inp[15]) ? node38011 : 4'b0000;
															assign node38011 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node38014 = (inp[0]) ? node38022 : node38015;
														assign node38015 = (inp[15]) ? node38019 : node38016;
															assign node38016 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node38019 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node38022 = (inp[15]) ? node38024 : 4'b1111;
															assign node38024 = (inp[3]) ? 4'b1101 : 4'b1101;
												assign node38027 = (inp[15]) ? node38039 : node38028;
													assign node38028 = (inp[0]) ? node38034 : node38029;
														assign node38029 = (inp[5]) ? 4'b1101 : node38030;
															assign node38030 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node38034 = (inp[3]) ? 4'b1111 : node38035;
															assign node38035 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node38039 = (inp[0]) ? node38045 : node38040;
														assign node38040 = (inp[3]) ? 4'b1111 : node38041;
															assign node38041 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node38045 = (inp[5]) ? 4'b1101 : node38046;
															assign node38046 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node38050 = (inp[14]) ? node38082 : node38051;
												assign node38051 = (inp[2]) ? node38067 : node38052;
													assign node38052 = (inp[5]) ? node38060 : node38053;
														assign node38053 = (inp[15]) ? node38057 : node38054;
															assign node38054 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node38057 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node38060 = (inp[3]) ? node38064 : node38061;
															assign node38061 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node38064 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node38067 = (inp[0]) ? node38075 : node38068;
														assign node38068 = (inp[15]) ? node38072 : node38069;
															assign node38069 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node38072 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node38075 = (inp[15]) ? node38079 : node38076;
															assign node38076 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node38079 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node38082 = (inp[5]) ? node38098 : node38083;
													assign node38083 = (inp[3]) ? node38091 : node38084;
														assign node38084 = (inp[0]) ? node38088 : node38085;
															assign node38085 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node38088 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node38091 = (inp[2]) ? node38095 : node38092;
															assign node38092 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node38095 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node38098 = (inp[2]) ? node38106 : node38099;
														assign node38099 = (inp[3]) ? node38103 : node38100;
															assign node38100 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node38103 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node38106 = (inp[3]) ? node38110 : node38107;
															assign node38107 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node38110 = (inp[0]) ? 4'b1110 : 4'b1100;
									assign node38113 = (inp[8]) ? node38219 : node38114;
										assign node38114 = (inp[7]) ? node38168 : node38115;
											assign node38115 = (inp[2]) ? node38145 : node38116;
												assign node38116 = (inp[14]) ? node38132 : node38117;
													assign node38117 = (inp[0]) ? node38125 : node38118;
														assign node38118 = (inp[15]) ? node38122 : node38119;
															assign node38119 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node38122 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node38125 = (inp[15]) ? node38129 : node38126;
															assign node38126 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node38129 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node38132 = (inp[15]) ? node38140 : node38133;
														assign node38133 = (inp[0]) ? node38137 : node38134;
															assign node38134 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node38137 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node38140 = (inp[3]) ? 4'b1100 : node38141;
															assign node38141 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node38145 = (inp[0]) ? node38157 : node38146;
													assign node38146 = (inp[15]) ? node38152 : node38147;
														assign node38147 = (inp[3]) ? 4'b1100 : node38148;
															assign node38148 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node38152 = (inp[3]) ? 4'b1110 : node38153;
															assign node38153 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node38157 = (inp[15]) ? node38163 : node38158;
														assign node38158 = (inp[5]) ? 4'b1110 : node38159;
															assign node38159 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node38163 = (inp[5]) ? 4'b1100 : node38164;
															assign node38164 = (inp[3]) ? 4'b1100 : 4'b1110;
											assign node38168 = (inp[2]) ? node38196 : node38169;
												assign node38169 = (inp[14]) ? node38181 : node38170;
													assign node38170 = (inp[15]) ? node38176 : node38171;
														assign node38171 = (inp[0]) ? 4'b1110 : node38172;
															assign node38172 = (inp[3]) ? 4'b1100 : 4'b1100;
														assign node38176 = (inp[0]) ? 4'b1100 : node38177;
															assign node38177 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node38181 = (inp[0]) ? node38189 : node38182;
														assign node38182 = (inp[15]) ? node38186 : node38183;
															assign node38183 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node38186 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node38189 = (inp[15]) ? node38193 : node38190;
															assign node38190 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node38193 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node38196 = (inp[15]) ? node38208 : node38197;
													assign node38197 = (inp[0]) ? node38203 : node38198;
														assign node38198 = (inp[5]) ? 4'b1101 : node38199;
															assign node38199 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node38203 = (inp[5]) ? 4'b1111 : node38204;
															assign node38204 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node38208 = (inp[0]) ? node38214 : node38209;
														assign node38209 = (inp[5]) ? 4'b1111 : node38210;
															assign node38210 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node38214 = (inp[14]) ? node38216 : 4'b1101;
															assign node38216 = (inp[5]) ? 4'b1101 : 4'b1101;
										assign node38219 = (inp[7]) ? node38273 : node38220;
											assign node38220 = (inp[14]) ? node38250 : node38221;
												assign node38221 = (inp[2]) ? node38237 : node38222;
													assign node38222 = (inp[5]) ? node38230 : node38223;
														assign node38223 = (inp[15]) ? node38227 : node38224;
															assign node38224 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node38227 = (inp[3]) ? 4'b1100 : 4'b1100;
														assign node38230 = (inp[0]) ? node38234 : node38231;
															assign node38231 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node38234 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node38237 = (inp[5]) ? node38245 : node38238;
														assign node38238 = (inp[15]) ? node38242 : node38239;
															assign node38239 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node38242 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node38245 = (inp[3]) ? 4'b1111 : node38246;
															assign node38246 = (inp[15]) ? 4'b1101 : 4'b1101;
												assign node38250 = (inp[5]) ? node38266 : node38251;
													assign node38251 = (inp[15]) ? node38259 : node38252;
														assign node38252 = (inp[2]) ? node38256 : node38253;
															assign node38253 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node38256 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node38259 = (inp[0]) ? node38263 : node38260;
															assign node38260 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node38263 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node38266 = (inp[0]) ? node38270 : node38267;
														assign node38267 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node38270 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node38273 = (inp[2]) ? node38303 : node38274;
												assign node38274 = (inp[14]) ? node38288 : node38275;
													assign node38275 = (inp[5]) ? node38283 : node38276;
														assign node38276 = (inp[3]) ? node38280 : node38277;
															assign node38277 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node38280 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node38283 = (inp[3]) ? 4'b1111 : node38284;
															assign node38284 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node38288 = (inp[15]) ? node38296 : node38289;
														assign node38289 = (inp[0]) ? node38293 : node38290;
															assign node38290 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node38293 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node38296 = (inp[0]) ? node38300 : node38297;
															assign node38297 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node38300 = (inp[3]) ? 4'b1100 : 4'b1100;
												assign node38303 = (inp[0]) ? node38315 : node38304;
													assign node38304 = (inp[15]) ? node38310 : node38305;
														assign node38305 = (inp[3]) ? 4'b1100 : node38306;
															assign node38306 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node38310 = (inp[5]) ? 4'b1110 : node38311;
															assign node38311 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node38315 = (inp[15]) ? node38321 : node38316;
														assign node38316 = (inp[3]) ? 4'b1110 : node38317;
															assign node38317 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node38321 = (inp[5]) ? 4'b1100 : node38322;
															assign node38322 = (inp[3]) ? 4'b1100 : 4'b1110;
							assign node38326 = (inp[1]) ? node38772 : node38327;
								assign node38327 = (inp[13]) ? node38549 : node38328;
									assign node38328 = (inp[7]) ? node38434 : node38329;
										assign node38329 = (inp[8]) ? node38383 : node38330;
											assign node38330 = (inp[14]) ? node38360 : node38331;
												assign node38331 = (inp[2]) ? node38347 : node38332;
													assign node38332 = (inp[3]) ? node38340 : node38333;
														assign node38333 = (inp[0]) ? node38337 : node38334;
															assign node38334 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node38337 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node38340 = (inp[15]) ? node38344 : node38341;
															assign node38341 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node38344 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node38347 = (inp[15]) ? node38353 : node38348;
														assign node38348 = (inp[0]) ? 4'b1110 : node38349;
															assign node38349 = (inp[3]) ? 4'b1100 : 4'b1100;
														assign node38353 = (inp[0]) ? node38357 : node38354;
															assign node38354 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node38357 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node38360 = (inp[3]) ? node38376 : node38361;
													assign node38361 = (inp[15]) ? node38369 : node38362;
														assign node38362 = (inp[0]) ? node38366 : node38363;
															assign node38363 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node38366 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node38369 = (inp[0]) ? node38373 : node38370;
															assign node38370 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node38373 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node38376 = (inp[0]) ? node38380 : node38377;
														assign node38377 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node38380 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node38383 = (inp[14]) ? node38411 : node38384;
												assign node38384 = (inp[2]) ? node38398 : node38385;
													assign node38385 = (inp[3]) ? node38393 : node38386;
														assign node38386 = (inp[5]) ? node38390 : node38387;
															assign node38387 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node38390 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node38393 = (inp[15]) ? node38395 : 4'b1100;
															assign node38395 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node38398 = (inp[3]) ? node38404 : node38399;
														assign node38399 = (inp[0]) ? 4'b1111 : node38400;
															assign node38400 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node38404 = (inp[15]) ? node38408 : node38405;
															assign node38405 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node38408 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node38411 = (inp[3]) ? node38427 : node38412;
													assign node38412 = (inp[2]) ? node38420 : node38413;
														assign node38413 = (inp[0]) ? node38417 : node38414;
															assign node38414 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node38417 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node38420 = (inp[15]) ? node38424 : node38421;
															assign node38421 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node38424 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node38427 = (inp[0]) ? node38431 : node38428;
														assign node38428 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node38431 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node38434 = (inp[8]) ? node38490 : node38435;
											assign node38435 = (inp[2]) ? node38467 : node38436;
												assign node38436 = (inp[14]) ? node38452 : node38437;
													assign node38437 = (inp[5]) ? node38445 : node38438;
														assign node38438 = (inp[0]) ? node38442 : node38439;
															assign node38439 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node38442 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node38445 = (inp[3]) ? node38449 : node38446;
															assign node38446 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node38449 = (inp[0]) ? 4'b1100 : 4'b1100;
													assign node38452 = (inp[15]) ? node38460 : node38453;
														assign node38453 = (inp[0]) ? node38457 : node38454;
															assign node38454 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node38457 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node38460 = (inp[0]) ? node38464 : node38461;
															assign node38461 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node38464 = (inp[3]) ? 4'b1101 : 4'b1101;
												assign node38467 = (inp[0]) ? node38479 : node38468;
													assign node38468 = (inp[15]) ? node38474 : node38469;
														assign node38469 = (inp[5]) ? 4'b1101 : node38470;
															assign node38470 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node38474 = (inp[3]) ? 4'b1111 : node38475;
															assign node38475 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node38479 = (inp[15]) ? node38485 : node38480;
														assign node38480 = (inp[5]) ? 4'b1111 : node38481;
															assign node38481 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node38485 = (inp[5]) ? 4'b1101 : node38486;
															assign node38486 = (inp[14]) ? 4'b1111 : 4'b1101;
											assign node38490 = (inp[14]) ? node38520 : node38491;
												assign node38491 = (inp[2]) ? node38505 : node38492;
													assign node38492 = (inp[15]) ? node38500 : node38493;
														assign node38493 = (inp[0]) ? node38497 : node38494;
															assign node38494 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node38497 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node38500 = (inp[0]) ? node38502 : 4'b1111;
															assign node38502 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node38505 = (inp[3]) ? node38513 : node38506;
														assign node38506 = (inp[0]) ? node38510 : node38507;
															assign node38507 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node38510 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node38513 = (inp[0]) ? node38517 : node38514;
															assign node38514 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node38517 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node38520 = (inp[3]) ? node38534 : node38521;
													assign node38521 = (inp[0]) ? node38529 : node38522;
														assign node38522 = (inp[15]) ? node38526 : node38523;
															assign node38523 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node38526 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node38529 = (inp[2]) ? 4'b1100 : node38530;
															assign node38530 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node38534 = (inp[2]) ? node38542 : node38535;
														assign node38535 = (inp[0]) ? node38539 : node38536;
															assign node38536 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node38539 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node38542 = (inp[5]) ? node38546 : node38543;
															assign node38543 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node38546 = (inp[0]) ? 4'b1110 : 4'b1100;
									assign node38549 = (inp[7]) ? node38661 : node38550;
										assign node38550 = (inp[8]) ? node38602 : node38551;
											assign node38551 = (inp[14]) ? node38579 : node38552;
												assign node38552 = (inp[2]) ? node38566 : node38553;
													assign node38553 = (inp[15]) ? node38559 : node38554;
														assign node38554 = (inp[0]) ? node38556 : 4'b1101;
															assign node38556 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node38559 = (inp[0]) ? node38563 : node38560;
															assign node38560 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node38563 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node38566 = (inp[3]) ? node38574 : node38567;
														assign node38567 = (inp[5]) ? node38571 : node38568;
															assign node38568 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node38571 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node38574 = (inp[0]) ? 4'b1110 : node38575;
															assign node38575 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node38579 = (inp[0]) ? node38591 : node38580;
													assign node38580 = (inp[15]) ? node38586 : node38581;
														assign node38581 = (inp[5]) ? 4'b1100 : node38582;
															assign node38582 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node38586 = (inp[3]) ? 4'b1110 : node38587;
															assign node38587 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node38591 = (inp[15]) ? node38597 : node38592;
														assign node38592 = (inp[3]) ? 4'b1110 : node38593;
															assign node38593 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node38597 = (inp[5]) ? 4'b1100 : node38598;
															assign node38598 = (inp[3]) ? 4'b1100 : 4'b1110;
											assign node38602 = (inp[14]) ? node38630 : node38603;
												assign node38603 = (inp[2]) ? node38619 : node38604;
													assign node38604 = (inp[0]) ? node38612 : node38605;
														assign node38605 = (inp[15]) ? node38609 : node38606;
															assign node38606 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node38609 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node38612 = (inp[15]) ? node38616 : node38613;
															assign node38613 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node38616 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node38619 = (inp[0]) ? node38625 : node38620;
														assign node38620 = (inp[15]) ? node38622 : 4'b0101;
															assign node38622 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node38625 = (inp[3]) ? 4'b0101 : node38626;
															assign node38626 = (inp[15]) ? 4'b0101 : 4'b0101;
												assign node38630 = (inp[3]) ? node38646 : node38631;
													assign node38631 = (inp[5]) ? node38639 : node38632;
														assign node38632 = (inp[0]) ? node38636 : node38633;
															assign node38633 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node38636 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node38639 = (inp[2]) ? node38643 : node38640;
															assign node38640 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node38643 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node38646 = (inp[5]) ? node38654 : node38647;
														assign node38647 = (inp[15]) ? node38651 : node38648;
															assign node38648 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node38651 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node38654 = (inp[15]) ? node38658 : node38655;
															assign node38655 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node38658 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node38661 = (inp[8]) ? node38721 : node38662;
											assign node38662 = (inp[14]) ? node38690 : node38663;
												assign node38663 = (inp[2]) ? node38677 : node38664;
													assign node38664 = (inp[0]) ? node38670 : node38665;
														assign node38665 = (inp[15]) ? node38667 : 4'b1100;
															assign node38667 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node38670 = (inp[15]) ? node38674 : node38671;
															assign node38671 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node38674 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node38677 = (inp[5]) ? node38685 : node38678;
														assign node38678 = (inp[0]) ? node38682 : node38679;
															assign node38679 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node38682 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node38685 = (inp[3]) ? 4'b0101 : node38686;
															assign node38686 = (inp[0]) ? 4'b0101 : 4'b0101;
												assign node38690 = (inp[5]) ? node38706 : node38691;
													assign node38691 = (inp[15]) ? node38699 : node38692;
														assign node38692 = (inp[2]) ? node38696 : node38693;
															assign node38693 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node38696 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node38699 = (inp[3]) ? node38703 : node38700;
															assign node38700 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node38703 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node38706 = (inp[2]) ? node38714 : node38707;
														assign node38707 = (inp[0]) ? node38711 : node38708;
															assign node38708 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node38711 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node38714 = (inp[0]) ? node38718 : node38715;
															assign node38715 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node38718 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node38721 = (inp[14]) ? node38749 : node38722;
												assign node38722 = (inp[2]) ? node38738 : node38723;
													assign node38723 = (inp[3]) ? node38731 : node38724;
														assign node38724 = (inp[15]) ? node38728 : node38725;
															assign node38725 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node38728 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node38731 = (inp[0]) ? node38735 : node38732;
															assign node38732 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node38735 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node38738 = (inp[0]) ? node38744 : node38739;
														assign node38739 = (inp[5]) ? 4'b0110 : node38740;
															assign node38740 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node38744 = (inp[3]) ? 4'b0100 : node38745;
															assign node38745 = (inp[15]) ? 4'b0100 : 4'b0100;
												assign node38749 = (inp[5]) ? node38765 : node38750;
													assign node38750 = (inp[2]) ? node38758 : node38751;
														assign node38751 = (inp[0]) ? node38755 : node38752;
															assign node38752 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node38755 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node38758 = (inp[15]) ? node38762 : node38759;
															assign node38759 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node38762 = (inp[0]) ? 4'b0100 : 4'b0100;
													assign node38765 = (inp[15]) ? node38769 : node38766;
														assign node38766 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node38769 = (inp[0]) ? 4'b0100 : 4'b0110;
								assign node38772 = (inp[13]) ? node38998 : node38773;
									assign node38773 = (inp[7]) ? node38887 : node38774;
										assign node38774 = (inp[8]) ? node38830 : node38775;
											assign node38775 = (inp[2]) ? node38807 : node38776;
												assign node38776 = (inp[14]) ? node38792 : node38777;
													assign node38777 = (inp[3]) ? node38785 : node38778;
														assign node38778 = (inp[15]) ? node38782 : node38779;
															assign node38779 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node38782 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node38785 = (inp[5]) ? node38789 : node38786;
															assign node38786 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node38789 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node38792 = (inp[3]) ? node38800 : node38793;
														assign node38793 = (inp[0]) ? node38797 : node38794;
															assign node38794 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node38797 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node38800 = (inp[0]) ? node38804 : node38801;
															assign node38801 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node38804 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node38807 = (inp[0]) ? node38819 : node38808;
													assign node38808 = (inp[15]) ? node38814 : node38809;
														assign node38809 = (inp[5]) ? 4'b1100 : node38810;
															assign node38810 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node38814 = (inp[5]) ? 4'b1110 : node38815;
															assign node38815 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node38819 = (inp[15]) ? node38825 : node38820;
														assign node38820 = (inp[3]) ? 4'b1110 : node38821;
															assign node38821 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node38825 = (inp[3]) ? 4'b1100 : node38826;
															assign node38826 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node38830 = (inp[14]) ? node38860 : node38831;
												assign node38831 = (inp[2]) ? node38847 : node38832;
													assign node38832 = (inp[15]) ? node38840 : node38833;
														assign node38833 = (inp[0]) ? node38837 : node38834;
															assign node38834 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node38837 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node38840 = (inp[0]) ? node38844 : node38841;
															assign node38841 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node38844 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node38847 = (inp[0]) ? node38855 : node38848;
														assign node38848 = (inp[15]) ? node38852 : node38849;
															assign node38849 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node38852 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node38855 = (inp[15]) ? 4'b0101 : node38856;
															assign node38856 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node38860 = (inp[2]) ? node38876 : node38861;
													assign node38861 = (inp[15]) ? node38869 : node38862;
														assign node38862 = (inp[0]) ? node38866 : node38863;
															assign node38863 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node38866 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node38869 = (inp[0]) ? node38873 : node38870;
															assign node38870 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node38873 = (inp[3]) ? 4'b0101 : 4'b0101;
													assign node38876 = (inp[15]) ? node38882 : node38877;
														assign node38877 = (inp[0]) ? 4'b0111 : node38878;
															assign node38878 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node38882 = (inp[0]) ? node38884 : 4'b0111;
															assign node38884 = (inp[3]) ? 4'b0101 : 4'b0101;
										assign node38887 = (inp[8]) ? node38947 : node38888;
											assign node38888 = (inp[14]) ? node38918 : node38889;
												assign node38889 = (inp[2]) ? node38905 : node38890;
													assign node38890 = (inp[3]) ? node38898 : node38891;
														assign node38891 = (inp[0]) ? node38895 : node38892;
															assign node38892 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node38895 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node38898 = (inp[5]) ? node38902 : node38899;
															assign node38899 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node38902 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node38905 = (inp[15]) ? node38911 : node38906;
														assign node38906 = (inp[0]) ? 4'b0111 : node38907;
															assign node38907 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node38911 = (inp[0]) ? node38915 : node38912;
															assign node38912 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node38915 = (inp[5]) ? 4'b0101 : 4'b0101;
												assign node38918 = (inp[2]) ? node38932 : node38919;
													assign node38919 = (inp[0]) ? node38925 : node38920;
														assign node38920 = (inp[15]) ? node38922 : 4'b0101;
															assign node38922 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node38925 = (inp[15]) ? node38929 : node38926;
															assign node38926 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node38929 = (inp[3]) ? 4'b0101 : 4'b0101;
													assign node38932 = (inp[0]) ? node38940 : node38933;
														assign node38933 = (inp[15]) ? node38937 : node38934;
															assign node38934 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node38937 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node38940 = (inp[15]) ? node38944 : node38941;
															assign node38941 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node38944 = (inp[3]) ? 4'b0101 : 4'b0101;
											assign node38947 = (inp[2]) ? node38977 : node38948;
												assign node38948 = (inp[14]) ? node38964 : node38949;
													assign node38949 = (inp[5]) ? node38957 : node38950;
														assign node38950 = (inp[0]) ? node38954 : node38951;
															assign node38951 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node38954 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node38957 = (inp[3]) ? node38961 : node38958;
															assign node38958 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node38961 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node38964 = (inp[0]) ? node38972 : node38965;
														assign node38965 = (inp[15]) ? node38969 : node38966;
															assign node38966 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node38969 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node38972 = (inp[15]) ? node38974 : 4'b0110;
															assign node38974 = (inp[3]) ? 4'b0100 : 4'b0100;
												assign node38977 = (inp[3]) ? node38991 : node38978;
													assign node38978 = (inp[0]) ? node38986 : node38979;
														assign node38979 = (inp[14]) ? node38983 : node38980;
															assign node38980 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node38983 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node38986 = (inp[5]) ? node38988 : 4'b0110;
															assign node38988 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node38991 = (inp[0]) ? node38995 : node38992;
														assign node38992 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node38995 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node38998 = (inp[0]) ? node39110 : node38999;
										assign node38999 = (inp[15]) ? node39053 : node39000;
											assign node39000 = (inp[5]) ? node39030 : node39001;
												assign node39001 = (inp[3]) ? node39017 : node39002;
													assign node39002 = (inp[14]) ? node39010 : node39003;
														assign node39003 = (inp[2]) ? node39007 : node39004;
															assign node39004 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node39007 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node39010 = (inp[7]) ? node39014 : node39011;
															assign node39011 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node39014 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node39017 = (inp[2]) ? node39025 : node39018;
														assign node39018 = (inp[7]) ? node39022 : node39019;
															assign node39019 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node39022 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node39025 = (inp[14]) ? 4'b0101 : node39026;
															assign node39026 = (inp[7]) ? 4'b0100 : 4'b0100;
												assign node39030 = (inp[7]) ? node39042 : node39031;
													assign node39031 = (inp[8]) ? node39037 : node39032;
														assign node39032 = (inp[2]) ? 4'b0100 : node39033;
															assign node39033 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node39037 = (inp[2]) ? 4'b0101 : node39038;
															assign node39038 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node39042 = (inp[8]) ? node39048 : node39043;
														assign node39043 = (inp[14]) ? 4'b0101 : node39044;
															assign node39044 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node39048 = (inp[2]) ? 4'b0100 : node39049;
															assign node39049 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node39053 = (inp[5]) ? node39081 : node39054;
												assign node39054 = (inp[3]) ? node39068 : node39055;
													assign node39055 = (inp[7]) ? node39063 : node39056;
														assign node39056 = (inp[8]) ? node39060 : node39057;
															assign node39057 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node39060 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node39063 = (inp[8]) ? node39065 : 4'b0101;
															assign node39065 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node39068 = (inp[7]) ? node39076 : node39069;
														assign node39069 = (inp[8]) ? node39073 : node39070;
															assign node39070 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node39073 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node39076 = (inp[2]) ? 4'b0110 : node39077;
															assign node39077 = (inp[14]) ? 4'b0110 : 4'b0110;
												assign node39081 = (inp[3]) ? node39095 : node39082;
													assign node39082 = (inp[14]) ? node39090 : node39083;
														assign node39083 = (inp[7]) ? node39087 : node39084;
															assign node39084 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node39087 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node39090 = (inp[2]) ? 4'b0110 : node39091;
															assign node39091 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node39095 = (inp[2]) ? node39103 : node39096;
														assign node39096 = (inp[7]) ? node39100 : node39097;
															assign node39097 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node39100 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node39103 = (inp[8]) ? node39107 : node39104;
															assign node39104 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node39107 = (inp[7]) ? 4'b0110 : 4'b0111;
										assign node39110 = (inp[15]) ? node39162 : node39111;
											assign node39111 = (inp[3]) ? node39139 : node39112;
												assign node39112 = (inp[5]) ? node39126 : node39113;
													assign node39113 = (inp[14]) ? node39121 : node39114;
														assign node39114 = (inp[8]) ? node39118 : node39115;
															assign node39115 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node39118 = (inp[2]) ? 4'b0100 : 4'b0100;
														assign node39121 = (inp[7]) ? 4'b0101 : node39122;
															assign node39122 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node39126 = (inp[2]) ? node39132 : node39127;
														assign node39127 = (inp[14]) ? node39129 : 4'b0110;
															assign node39129 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node39132 = (inp[8]) ? node39136 : node39133;
															assign node39133 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node39136 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node39139 = (inp[7]) ? node39151 : node39140;
													assign node39140 = (inp[8]) ? node39146 : node39141;
														assign node39141 = (inp[14]) ? 4'b0110 : node39142;
															assign node39142 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node39146 = (inp[2]) ? 4'b0111 : node39147;
															assign node39147 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node39151 = (inp[8]) ? node39157 : node39152;
														assign node39152 = (inp[14]) ? 4'b0111 : node39153;
															assign node39153 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node39157 = (inp[14]) ? 4'b0110 : node39158;
															assign node39158 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node39162 = (inp[5]) ? node39192 : node39163;
												assign node39163 = (inp[3]) ? node39177 : node39164;
													assign node39164 = (inp[14]) ? node39172 : node39165;
														assign node39165 = (inp[8]) ? node39169 : node39166;
															assign node39166 = (inp[2]) ? 4'b0110 : 4'b0110;
															assign node39169 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node39172 = (inp[8]) ? node39174 : 4'b0110;
															assign node39174 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node39177 = (inp[8]) ? node39185 : node39178;
														assign node39178 = (inp[7]) ? node39182 : node39179;
															assign node39179 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node39182 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node39185 = (inp[7]) ? node39189 : node39186;
															assign node39186 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node39189 = (inp[14]) ? 4'b0100 : 4'b0100;
												assign node39192 = (inp[3]) ? node39208 : node39193;
													assign node39193 = (inp[8]) ? node39201 : node39194;
														assign node39194 = (inp[7]) ? node39198 : node39195;
															assign node39195 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node39198 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node39201 = (inp[7]) ? node39205 : node39202;
															assign node39202 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node39205 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node39208 = (inp[2]) ? node39216 : node39209;
														assign node39209 = (inp[7]) ? node39213 : node39210;
															assign node39210 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node39213 = (inp[14]) ? 4'b0100 : 4'b0100;
														assign node39216 = (inp[8]) ? node39220 : node39217;
															assign node39217 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node39220 = (inp[7]) ? 4'b0100 : 4'b0101;
					assign node39223 = (inp[2]) ? node41201 : node39224;
						assign node39224 = (inp[3]) ? node40218 : node39225;
							assign node39225 = (inp[11]) ? node39719 : node39226;
								assign node39226 = (inp[0]) ? node39472 : node39227;
									assign node39227 = (inp[15]) ? node39351 : node39228;
										assign node39228 = (inp[5]) ? node39290 : node39229;
											assign node39229 = (inp[13]) ? node39259 : node39230;
												assign node39230 = (inp[6]) ? node39246 : node39231;
													assign node39231 = (inp[1]) ? node39239 : node39232;
														assign node39232 = (inp[7]) ? node39236 : node39233;
															assign node39233 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node39236 = (inp[14]) ? 4'b1110 : 4'b1110;
														assign node39239 = (inp[14]) ? node39243 : node39240;
															assign node39240 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node39243 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node39246 = (inp[1]) ? node39252 : node39247;
														assign node39247 = (inp[14]) ? 4'b0110 : node39248;
															assign node39248 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node39252 = (inp[14]) ? node39256 : node39253;
															assign node39253 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node39256 = (inp[8]) ? 4'b1110 : 4'b0110;
												assign node39259 = (inp[6]) ? node39275 : node39260;
													assign node39260 = (inp[14]) ? node39268 : node39261;
														assign node39261 = (inp[1]) ? node39265 : node39262;
															assign node39262 = (inp[8]) ? 4'b0110 : 4'b1110;
															assign node39265 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node39268 = (inp[7]) ? node39272 : node39269;
															assign node39269 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node39272 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node39275 = (inp[8]) ? node39283 : node39276;
														assign node39276 = (inp[1]) ? node39280 : node39277;
															assign node39277 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node39280 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node39283 = (inp[7]) ? node39287 : node39284;
															assign node39284 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node39287 = (inp[14]) ? 4'b1110 : 4'b1111;
											assign node39290 = (inp[6]) ? node39320 : node39291;
												assign node39291 = (inp[13]) ? node39307 : node39292;
													assign node39292 = (inp[1]) ? node39300 : node39293;
														assign node39293 = (inp[14]) ? node39297 : node39294;
															assign node39294 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node39297 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node39300 = (inp[14]) ? node39304 : node39301;
															assign node39301 = (inp[8]) ? 4'b0100 : 4'b1100;
															assign node39304 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node39307 = (inp[8]) ? node39313 : node39308;
														assign node39308 = (inp[7]) ? 4'b0101 : node39309;
															assign node39309 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node39313 = (inp[14]) ? node39317 : node39314;
															assign node39314 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node39317 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node39320 = (inp[13]) ? node39336 : node39321;
													assign node39321 = (inp[1]) ? node39329 : node39322;
														assign node39322 = (inp[14]) ? node39326 : node39323;
															assign node39323 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node39326 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node39329 = (inp[14]) ? node39333 : node39330;
															assign node39330 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node39333 = (inp[7]) ? 4'b1100 : 4'b0100;
													assign node39336 = (inp[1]) ? node39344 : node39337;
														assign node39337 = (inp[7]) ? node39341 : node39338;
															assign node39338 = (inp[8]) ? 4'b1101 : 4'b0100;
															assign node39341 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node39344 = (inp[8]) ? node39348 : node39345;
															assign node39345 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node39348 = (inp[7]) ? 4'b1100 : 4'b1100;
										assign node39351 = (inp[5]) ? node39413 : node39352;
											assign node39352 = (inp[6]) ? node39384 : node39353;
												assign node39353 = (inp[13]) ? node39369 : node39354;
													assign node39354 = (inp[1]) ? node39362 : node39355;
														assign node39355 = (inp[14]) ? node39359 : node39356;
															assign node39356 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node39359 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node39362 = (inp[14]) ? node39366 : node39363;
															assign node39363 = (inp[8]) ? 4'b0100 : 4'b1100;
															assign node39366 = (inp[8]) ? 4'b0100 : 4'b0100;
													assign node39369 = (inp[1]) ? node39377 : node39370;
														assign node39370 = (inp[14]) ? node39374 : node39371;
															assign node39371 = (inp[8]) ? 4'b0100 : 4'b1100;
															assign node39374 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node39377 = (inp[8]) ? node39381 : node39378;
															assign node39378 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node39381 = (inp[7]) ? 4'b0100 : 4'b0100;
												assign node39384 = (inp[1]) ? node39400 : node39385;
													assign node39385 = (inp[13]) ? node39393 : node39386;
														assign node39386 = (inp[7]) ? node39390 : node39387;
															assign node39387 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node39390 = (inp[14]) ? 4'b0100 : 4'b0100;
														assign node39393 = (inp[8]) ? node39397 : node39394;
															assign node39394 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node39397 = (inp[7]) ? 4'b1101 : 4'b0100;
													assign node39400 = (inp[14]) ? node39408 : node39401;
														assign node39401 = (inp[13]) ? node39405 : node39402;
															assign node39402 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node39405 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node39408 = (inp[7]) ? node39410 : 4'b1101;
															assign node39410 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node39413 = (inp[14]) ? node39445 : node39414;
												assign node39414 = (inp[6]) ? node39430 : node39415;
													assign node39415 = (inp[1]) ? node39423 : node39416;
														assign node39416 = (inp[13]) ? node39420 : node39417;
															assign node39417 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node39420 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node39423 = (inp[13]) ? node39427 : node39424;
															assign node39424 = (inp[7]) ? 4'b0110 : 4'b1110;
															assign node39427 = (inp[8]) ? 4'b0110 : 4'b0110;
													assign node39430 = (inp[13]) ? node39438 : node39431;
														assign node39431 = (inp[8]) ? node39435 : node39432;
															assign node39432 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node39435 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node39438 = (inp[1]) ? node39442 : node39439;
															assign node39439 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node39442 = (inp[8]) ? 4'b1110 : 4'b1110;
												assign node39445 = (inp[6]) ? node39459 : node39446;
													assign node39446 = (inp[13]) ? node39454 : node39447;
														assign node39447 = (inp[1]) ? node39451 : node39448;
															assign node39448 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node39451 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node39454 = (inp[1]) ? node39456 : 4'b0111;
															assign node39456 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node39459 = (inp[1]) ? node39467 : node39460;
														assign node39460 = (inp[8]) ? node39464 : node39461;
															assign node39461 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node39464 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node39467 = (inp[13]) ? node39469 : 4'b1111;
															assign node39469 = (inp[7]) ? 4'b1110 : 4'b1110;
									assign node39472 = (inp[13]) ? node39596 : node39473;
										assign node39473 = (inp[6]) ? node39535 : node39474;
											assign node39474 = (inp[1]) ? node39504 : node39475;
												assign node39475 = (inp[5]) ? node39489 : node39476;
													assign node39476 = (inp[15]) ? node39482 : node39477;
														assign node39477 = (inp[14]) ? 4'b1100 : node39478;
															assign node39478 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node39482 = (inp[14]) ? node39486 : node39483;
															assign node39483 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node39486 = (inp[7]) ? 4'b1110 : 4'b1110;
													assign node39489 = (inp[15]) ? node39497 : node39490;
														assign node39490 = (inp[14]) ? node39494 : node39491;
															assign node39491 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node39494 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node39497 = (inp[14]) ? node39501 : node39498;
															assign node39498 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node39501 = (inp[7]) ? 4'b1100 : 4'b1100;
												assign node39504 = (inp[7]) ? node39520 : node39505;
													assign node39505 = (inp[14]) ? node39513 : node39506;
														assign node39506 = (inp[8]) ? node39510 : node39507;
															assign node39507 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node39510 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node39513 = (inp[8]) ? node39517 : node39514;
															assign node39514 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node39517 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node39520 = (inp[14]) ? node39528 : node39521;
														assign node39521 = (inp[8]) ? node39525 : node39522;
															assign node39522 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node39525 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node39528 = (inp[8]) ? node39532 : node39529;
															assign node39529 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node39532 = (inp[5]) ? 4'b0100 : 4'b0100;
											assign node39535 = (inp[1]) ? node39565 : node39536;
												assign node39536 = (inp[15]) ? node39552 : node39537;
													assign node39537 = (inp[5]) ? node39545 : node39538;
														assign node39538 = (inp[8]) ? node39542 : node39539;
															assign node39539 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node39542 = (inp[14]) ? 4'b0100 : 4'b0100;
														assign node39545 = (inp[14]) ? node39549 : node39546;
															assign node39546 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node39549 = (inp[8]) ? 4'b0110 : 4'b0110;
													assign node39552 = (inp[5]) ? node39560 : node39553;
														assign node39553 = (inp[8]) ? node39557 : node39554;
															assign node39554 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node39557 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node39560 = (inp[7]) ? 4'b0100 : node39561;
															assign node39561 = (inp[14]) ? 4'b0100 : 4'b0100;
												assign node39565 = (inp[14]) ? node39581 : node39566;
													assign node39566 = (inp[8]) ? node39574 : node39567;
														assign node39567 = (inp[7]) ? node39571 : node39568;
															assign node39568 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node39571 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node39574 = (inp[7]) ? node39578 : node39575;
															assign node39575 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node39578 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node39581 = (inp[7]) ? node39589 : node39582;
														assign node39582 = (inp[8]) ? node39586 : node39583;
															assign node39583 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node39586 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node39589 = (inp[8]) ? node39593 : node39590;
															assign node39590 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node39593 = (inp[5]) ? 4'b1110 : 4'b1100;
										assign node39596 = (inp[6]) ? node39660 : node39597;
											assign node39597 = (inp[1]) ? node39629 : node39598;
												assign node39598 = (inp[14]) ? node39614 : node39599;
													assign node39599 = (inp[8]) ? node39607 : node39600;
														assign node39600 = (inp[7]) ? node39604 : node39601;
															assign node39601 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node39604 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node39607 = (inp[7]) ? node39611 : node39608;
															assign node39608 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node39611 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node39614 = (inp[8]) ? node39622 : node39615;
														assign node39615 = (inp[7]) ? node39619 : node39616;
															assign node39616 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node39619 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node39622 = (inp[7]) ? node39626 : node39623;
															assign node39623 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node39626 = (inp[5]) ? 4'b0100 : 4'b0100;
												assign node39629 = (inp[7]) ? node39645 : node39630;
													assign node39630 = (inp[14]) ? node39638 : node39631;
														assign node39631 = (inp[8]) ? node39635 : node39632;
															assign node39632 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node39635 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node39638 = (inp[8]) ? node39642 : node39639;
															assign node39639 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node39642 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node39645 = (inp[15]) ? node39653 : node39646;
														assign node39646 = (inp[5]) ? node39650 : node39647;
															assign node39647 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node39650 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node39653 = (inp[5]) ? node39657 : node39654;
															assign node39654 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node39657 = (inp[8]) ? 4'b0100 : 4'b0100;
											assign node39660 = (inp[1]) ? node39692 : node39661;
												assign node39661 = (inp[8]) ? node39677 : node39662;
													assign node39662 = (inp[7]) ? node39670 : node39663;
														assign node39663 = (inp[14]) ? node39667 : node39664;
															assign node39664 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node39667 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node39670 = (inp[14]) ? node39674 : node39671;
															assign node39671 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node39674 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node39677 = (inp[7]) ? node39685 : node39678;
														assign node39678 = (inp[14]) ? node39682 : node39679;
															assign node39679 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node39682 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node39685 = (inp[14]) ? node39689 : node39686;
															assign node39686 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node39689 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node39692 = (inp[15]) ? node39706 : node39693;
													assign node39693 = (inp[5]) ? node39699 : node39694;
														assign node39694 = (inp[7]) ? node39696 : 4'b1101;
															assign node39696 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node39699 = (inp[7]) ? node39703 : node39700;
															assign node39700 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node39703 = (inp[8]) ? 4'b1110 : 4'b1110;
													assign node39706 = (inp[5]) ? node39712 : node39707;
														assign node39707 = (inp[7]) ? node39709 : 4'b1110;
															assign node39709 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node39712 = (inp[14]) ? node39716 : node39713;
															assign node39713 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node39716 = (inp[8]) ? 4'b1100 : 4'b1100;
								assign node39719 = (inp[0]) ? node39969 : node39720;
									assign node39720 = (inp[15]) ? node39846 : node39721;
										assign node39721 = (inp[5]) ? node39783 : node39722;
											assign node39722 = (inp[14]) ? node39754 : node39723;
												assign node39723 = (inp[6]) ? node39739 : node39724;
													assign node39724 = (inp[1]) ? node39732 : node39725;
														assign node39725 = (inp[7]) ? node39729 : node39726;
															assign node39726 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node39729 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node39732 = (inp[13]) ? node39736 : node39733;
															assign node39733 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node39736 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node39739 = (inp[1]) ? node39747 : node39740;
														assign node39740 = (inp[7]) ? node39744 : node39741;
															assign node39741 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node39744 = (inp[8]) ? 4'b0111 : 4'b1110;
														assign node39747 = (inp[13]) ? node39751 : node39748;
															assign node39748 = (inp[7]) ? 4'b0110 : 4'b1110;
															assign node39751 = (inp[8]) ? 4'b0110 : 4'b0110;
												assign node39754 = (inp[6]) ? node39770 : node39755;
													assign node39755 = (inp[1]) ? node39763 : node39756;
														assign node39756 = (inp[13]) ? node39760 : node39757;
															assign node39757 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node39760 = (inp[8]) ? 4'b1110 : 4'b0110;
														assign node39763 = (inp[7]) ? node39767 : node39764;
															assign node39764 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node39767 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node39770 = (inp[1]) ? node39776 : node39771;
														assign node39771 = (inp[13]) ? node39773 : 4'b1111;
															assign node39773 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node39776 = (inp[8]) ? node39780 : node39777;
															assign node39777 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node39780 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node39783 = (inp[14]) ? node39815 : node39784;
												assign node39784 = (inp[6]) ? node39800 : node39785;
													assign node39785 = (inp[13]) ? node39793 : node39786;
														assign node39786 = (inp[8]) ? node39790 : node39787;
															assign node39787 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node39790 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node39793 = (inp[1]) ? node39797 : node39794;
															assign node39794 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node39797 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node39800 = (inp[1]) ? node39808 : node39801;
														assign node39801 = (inp[8]) ? node39805 : node39802;
															assign node39802 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node39805 = (inp[7]) ? 4'b0101 : 4'b1100;
														assign node39808 = (inp[13]) ? node39812 : node39809;
															assign node39809 = (inp[7]) ? 4'b0100 : 4'b1100;
															assign node39812 = (inp[8]) ? 4'b0101 : 4'b0100;
												assign node39815 = (inp[6]) ? node39831 : node39816;
													assign node39816 = (inp[13]) ? node39824 : node39817;
														assign node39817 = (inp[1]) ? node39821 : node39818;
															assign node39818 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node39821 = (inp[8]) ? 4'b1100 : 4'b0100;
														assign node39824 = (inp[8]) ? node39828 : node39825;
															assign node39825 = (inp[7]) ? 4'b1101 : 4'b0100;
															assign node39828 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node39831 = (inp[1]) ? node39839 : node39832;
														assign node39832 = (inp[13]) ? node39836 : node39833;
															assign node39833 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node39836 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node39839 = (inp[8]) ? node39843 : node39840;
															assign node39840 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node39843 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node39846 = (inp[5]) ? node39906 : node39847;
											assign node39847 = (inp[1]) ? node39879 : node39848;
												assign node39848 = (inp[6]) ? node39864 : node39849;
													assign node39849 = (inp[13]) ? node39857 : node39850;
														assign node39850 = (inp[8]) ? node39854 : node39851;
															assign node39851 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node39854 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node39857 = (inp[8]) ? node39861 : node39858;
															assign node39858 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node39861 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node39864 = (inp[13]) ? node39872 : node39865;
														assign node39865 = (inp[8]) ? node39869 : node39866;
															assign node39866 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node39869 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node39872 = (inp[7]) ? node39876 : node39873;
															assign node39873 = (inp[8]) ? 4'b0100 : 4'b1100;
															assign node39876 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node39879 = (inp[6]) ? node39895 : node39880;
													assign node39880 = (inp[13]) ? node39888 : node39881;
														assign node39881 = (inp[14]) ? node39885 : node39882;
															assign node39882 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node39885 = (inp[7]) ? 4'b1100 : 4'b0100;
														assign node39888 = (inp[7]) ? node39892 : node39889;
															assign node39889 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node39892 = (inp[8]) ? 4'b1100 : 4'b1100;
													assign node39895 = (inp[13]) ? node39901 : node39896;
														assign node39896 = (inp[7]) ? node39898 : 4'b1100;
															assign node39898 = (inp[8]) ? 4'b0100 : 4'b1100;
														assign node39901 = (inp[14]) ? node39903 : 4'b0100;
															assign node39903 = (inp[7]) ? 4'b0100 : 4'b0100;
											assign node39906 = (inp[1]) ? node39938 : node39907;
												assign node39907 = (inp[6]) ? node39923 : node39908;
													assign node39908 = (inp[13]) ? node39916 : node39909;
														assign node39909 = (inp[7]) ? node39913 : node39910;
															assign node39910 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node39913 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node39916 = (inp[7]) ? node39920 : node39917;
															assign node39917 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node39920 = (inp[8]) ? 4'b1110 : 4'b0110;
													assign node39923 = (inp[13]) ? node39931 : node39924;
														assign node39924 = (inp[8]) ? node39928 : node39925;
															assign node39925 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node39928 = (inp[14]) ? 4'b1110 : 4'b1110;
														assign node39931 = (inp[14]) ? node39935 : node39932;
															assign node39932 = (inp[7]) ? 4'b0110 : 4'b1110;
															assign node39935 = (inp[8]) ? 4'b0110 : 4'b0110;
												assign node39938 = (inp[6]) ? node39954 : node39939;
													assign node39939 = (inp[13]) ? node39947 : node39940;
														assign node39940 = (inp[14]) ? node39944 : node39941;
															assign node39941 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node39944 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node39947 = (inp[8]) ? node39951 : node39948;
															assign node39948 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node39951 = (inp[14]) ? 4'b1110 : 4'b1110;
													assign node39954 = (inp[13]) ? node39962 : node39955;
														assign node39955 = (inp[14]) ? node39959 : node39956;
															assign node39956 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node39959 = (inp[8]) ? 4'b0110 : 4'b1110;
														assign node39962 = (inp[8]) ? node39966 : node39963;
															assign node39963 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node39966 = (inp[14]) ? 4'b0110 : 4'b0110;
									assign node39969 = (inp[6]) ? node40097 : node39970;
										assign node39970 = (inp[1]) ? node40034 : node39971;
											assign node39971 = (inp[13]) ? node40003 : node39972;
												assign node39972 = (inp[14]) ? node39988 : node39973;
													assign node39973 = (inp[7]) ? node39981 : node39974;
														assign node39974 = (inp[8]) ? node39978 : node39975;
															assign node39975 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node39978 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node39981 = (inp[8]) ? node39985 : node39982;
															assign node39982 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node39985 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node39988 = (inp[8]) ? node39996 : node39989;
														assign node39989 = (inp[7]) ? node39993 : node39990;
															assign node39990 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node39993 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node39996 = (inp[7]) ? node40000 : node39997;
															assign node39997 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node40000 = (inp[5]) ? 4'b0100 : 4'b0100;
												assign node40003 = (inp[7]) ? node40019 : node40004;
													assign node40004 = (inp[15]) ? node40012 : node40005;
														assign node40005 = (inp[5]) ? node40009 : node40006;
															assign node40006 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node40009 = (inp[8]) ? 4'b1111 : 4'b0110;
														assign node40012 = (inp[5]) ? node40016 : node40013;
															assign node40013 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node40016 = (inp[8]) ? 4'b0100 : 4'b0100;
													assign node40019 = (inp[14]) ? node40027 : node40020;
														assign node40020 = (inp[8]) ? node40024 : node40021;
															assign node40021 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node40024 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node40027 = (inp[8]) ? node40031 : node40028;
															assign node40028 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node40031 = (inp[5]) ? 4'b1100 : 4'b1100;
											assign node40034 = (inp[13]) ? node40066 : node40035;
												assign node40035 = (inp[8]) ? node40051 : node40036;
													assign node40036 = (inp[7]) ? node40044 : node40037;
														assign node40037 = (inp[14]) ? node40041 : node40038;
															assign node40038 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node40041 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node40044 = (inp[14]) ? node40048 : node40045;
															assign node40045 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node40048 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node40051 = (inp[7]) ? node40059 : node40052;
														assign node40052 = (inp[14]) ? node40056 : node40053;
															assign node40053 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node40056 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node40059 = (inp[14]) ? node40063 : node40060;
															assign node40060 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node40063 = (inp[15]) ? 4'b1100 : 4'b1100;
												assign node40066 = (inp[8]) ? node40082 : node40067;
													assign node40067 = (inp[14]) ? node40075 : node40068;
														assign node40068 = (inp[7]) ? node40072 : node40069;
															assign node40069 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node40072 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node40075 = (inp[7]) ? node40079 : node40076;
															assign node40076 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node40079 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node40082 = (inp[14]) ? node40090 : node40083;
														assign node40083 = (inp[7]) ? node40087 : node40084;
															assign node40084 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node40087 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node40090 = (inp[7]) ? node40094 : node40091;
															assign node40091 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node40094 = (inp[5]) ? 4'b1100 : 4'b1100;
										assign node40097 = (inp[13]) ? node40159 : node40098;
											assign node40098 = (inp[1]) ? node40128 : node40099;
												assign node40099 = (inp[5]) ? node40115 : node40100;
													assign node40100 = (inp[15]) ? node40108 : node40101;
														assign node40101 = (inp[7]) ? node40105 : node40102;
															assign node40102 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node40105 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node40108 = (inp[7]) ? node40112 : node40109;
															assign node40109 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node40112 = (inp[8]) ? 4'b1110 : 4'b1110;
													assign node40115 = (inp[15]) ? node40121 : node40116;
														assign node40116 = (inp[8]) ? node40118 : 4'b1111;
															assign node40118 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node40121 = (inp[8]) ? node40125 : node40122;
															assign node40122 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node40125 = (inp[14]) ? 4'b1100 : 4'b1100;
												assign node40128 = (inp[7]) ? node40144 : node40129;
													assign node40129 = (inp[8]) ? node40137 : node40130;
														assign node40130 = (inp[14]) ? node40134 : node40131;
															assign node40131 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node40134 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node40137 = (inp[14]) ? node40141 : node40138;
															assign node40138 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node40141 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node40144 = (inp[14]) ? node40152 : node40145;
														assign node40145 = (inp[8]) ? node40149 : node40146;
															assign node40146 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node40149 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node40152 = (inp[8]) ? node40156 : node40153;
															assign node40153 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node40156 = (inp[5]) ? 4'b0110 : 4'b0100;
											assign node40159 = (inp[1]) ? node40191 : node40160;
												assign node40160 = (inp[7]) ? node40176 : node40161;
													assign node40161 = (inp[14]) ? node40169 : node40162;
														assign node40162 = (inp[8]) ? node40166 : node40163;
															assign node40163 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node40166 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node40169 = (inp[8]) ? node40173 : node40170;
															assign node40170 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node40173 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node40176 = (inp[14]) ? node40184 : node40177;
														assign node40177 = (inp[8]) ? node40181 : node40178;
															assign node40178 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node40181 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node40184 = (inp[8]) ? node40188 : node40185;
															assign node40185 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node40188 = (inp[15]) ? 4'b0100 : 4'b0100;
												assign node40191 = (inp[14]) ? node40203 : node40192;
													assign node40192 = (inp[8]) ? node40200 : node40193;
														assign node40193 = (inp[7]) ? node40197 : node40194;
															assign node40194 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node40197 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node40200 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node40203 = (inp[15]) ? node40211 : node40204;
														assign node40204 = (inp[5]) ? node40208 : node40205;
															assign node40205 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node40208 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node40211 = (inp[5]) ? node40215 : node40212;
															assign node40212 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node40215 = (inp[8]) ? 4'b0100 : 4'b0100;
							assign node40218 = (inp[5]) ? node40706 : node40219;
								assign node40219 = (inp[15]) ? node40471 : node40220;
									assign node40220 = (inp[0]) ? node40346 : node40221;
										assign node40221 = (inp[1]) ? node40283 : node40222;
											assign node40222 = (inp[11]) ? node40254 : node40223;
												assign node40223 = (inp[6]) ? node40239 : node40224;
													assign node40224 = (inp[13]) ? node40232 : node40225;
														assign node40225 = (inp[7]) ? node40229 : node40226;
															assign node40226 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node40229 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node40232 = (inp[7]) ? node40236 : node40233;
															assign node40233 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node40236 = (inp[8]) ? 4'b0100 : 4'b1100;
													assign node40239 = (inp[13]) ? node40247 : node40240;
														assign node40240 = (inp[7]) ? node40244 : node40241;
															assign node40241 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node40244 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node40247 = (inp[7]) ? node40251 : node40248;
															assign node40248 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node40251 = (inp[8]) ? 4'b1100 : 4'b0100;
												assign node40254 = (inp[6]) ? node40270 : node40255;
													assign node40255 = (inp[13]) ? node40263 : node40256;
														assign node40256 = (inp[8]) ? node40260 : node40257;
															assign node40257 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node40260 = (inp[14]) ? 4'b0100 : 4'b0100;
														assign node40263 = (inp[14]) ? node40267 : node40264;
															assign node40264 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node40267 = (inp[8]) ? 4'b1101 : 4'b0100;
													assign node40270 = (inp[13]) ? node40276 : node40271;
														assign node40271 = (inp[8]) ? node40273 : 4'b1101;
															assign node40273 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node40276 = (inp[7]) ? node40280 : node40277;
															assign node40277 = (inp[8]) ? 4'b0100 : 4'b1100;
															assign node40280 = (inp[8]) ? 4'b0100 : 4'b0100;
											assign node40283 = (inp[8]) ? node40315 : node40284;
												assign node40284 = (inp[11]) ? node40300 : node40285;
													assign node40285 = (inp[6]) ? node40293 : node40286;
														assign node40286 = (inp[13]) ? node40290 : node40287;
															assign node40287 = (inp[7]) ? 4'b0100 : 4'b1100;
															assign node40290 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node40293 = (inp[13]) ? node40297 : node40294;
															assign node40294 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node40297 = (inp[7]) ? 4'b1100 : 4'b1100;
													assign node40300 = (inp[6]) ? node40308 : node40301;
														assign node40301 = (inp[13]) ? node40305 : node40302;
															assign node40302 = (inp[14]) ? 4'b1101 : 4'b0100;
															assign node40305 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node40308 = (inp[13]) ? node40312 : node40309;
															assign node40309 = (inp[7]) ? 4'b0100 : 4'b1100;
															assign node40312 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node40315 = (inp[7]) ? node40331 : node40316;
													assign node40316 = (inp[14]) ? node40324 : node40317;
														assign node40317 = (inp[11]) ? node40321 : node40318;
															assign node40318 = (inp[13]) ? 4'b0100 : 4'b0100;
															assign node40321 = (inp[13]) ? 4'b0100 : 4'b0100;
														assign node40324 = (inp[13]) ? node40328 : node40325;
															assign node40325 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node40328 = (inp[11]) ? 4'b0101 : 4'b0101;
													assign node40331 = (inp[14]) ? node40339 : node40332;
														assign node40332 = (inp[13]) ? node40336 : node40333;
															assign node40333 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node40336 = (inp[6]) ? 4'b0101 : 4'b0101;
														assign node40339 = (inp[13]) ? node40343 : node40340;
															assign node40340 = (inp[11]) ? 4'b0100 : 4'b0100;
															assign node40343 = (inp[6]) ? 4'b0100 : 4'b0100;
										assign node40346 = (inp[14]) ? node40410 : node40347;
											assign node40347 = (inp[6]) ? node40379 : node40348;
												assign node40348 = (inp[11]) ? node40364 : node40349;
													assign node40349 = (inp[13]) ? node40357 : node40350;
														assign node40350 = (inp[8]) ? node40354 : node40351;
															assign node40351 = (inp[7]) ? 4'b1110 : 4'b1111;
															assign node40354 = (inp[7]) ? 4'b0111 : 4'b1110;
														assign node40357 = (inp[1]) ? node40361 : node40358;
															assign node40358 = (inp[7]) ? 4'b0110 : 4'b1110;
															assign node40361 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node40364 = (inp[13]) ? node40372 : node40365;
														assign node40365 = (inp[1]) ? node40369 : node40366;
															assign node40366 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node40369 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node40372 = (inp[1]) ? node40376 : node40373;
															assign node40373 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node40376 = (inp[8]) ? 4'b1111 : 4'b1110;
												assign node40379 = (inp[11]) ? node40395 : node40380;
													assign node40380 = (inp[13]) ? node40388 : node40381;
														assign node40381 = (inp[8]) ? node40385 : node40382;
															assign node40382 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node40385 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node40388 = (inp[1]) ? node40392 : node40389;
															assign node40389 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node40392 = (inp[7]) ? 4'b1110 : 4'b1110;
													assign node40395 = (inp[13]) ? node40403 : node40396;
														assign node40396 = (inp[1]) ? node40400 : node40397;
															assign node40397 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node40400 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node40403 = (inp[1]) ? node40407 : node40404;
															assign node40404 = (inp[7]) ? 4'b0110 : 4'b1110;
															assign node40407 = (inp[8]) ? 4'b0110 : 4'b0110;
											assign node40410 = (inp[6]) ? node40442 : node40411;
												assign node40411 = (inp[1]) ? node40427 : node40412;
													assign node40412 = (inp[11]) ? node40420 : node40413;
														assign node40413 = (inp[13]) ? node40417 : node40414;
															assign node40414 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node40417 = (inp[7]) ? 4'b0110 : 4'b1110;
														assign node40420 = (inp[13]) ? node40424 : node40421;
															assign node40421 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node40424 = (inp[8]) ? 4'b1110 : 4'b0110;
													assign node40427 = (inp[11]) ? node40435 : node40428;
														assign node40428 = (inp[8]) ? node40432 : node40429;
															assign node40429 = (inp[7]) ? 4'b0111 : 4'b1110;
															assign node40432 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node40435 = (inp[13]) ? node40439 : node40436;
															assign node40436 = (inp[8]) ? 4'b1111 : 4'b0110;
															assign node40439 = (inp[8]) ? 4'b1110 : 4'b1110;
												assign node40442 = (inp[11]) ? node40458 : node40443;
													assign node40443 = (inp[1]) ? node40451 : node40444;
														assign node40444 = (inp[13]) ? node40448 : node40445;
															assign node40445 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node40448 = (inp[8]) ? 4'b1111 : 4'b0110;
														assign node40451 = (inp[7]) ? node40455 : node40452;
															assign node40452 = (inp[8]) ? 4'b1111 : 4'b0110;
															assign node40455 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node40458 = (inp[1]) ? node40464 : node40459;
														assign node40459 = (inp[13]) ? 4'b0111 : node40460;
															assign node40460 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node40464 = (inp[13]) ? node40468 : node40465;
															assign node40465 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node40468 = (inp[8]) ? 4'b0110 : 4'b0110;
									assign node40471 = (inp[0]) ? node40587 : node40472;
										assign node40472 = (inp[7]) ? node40530 : node40473;
											assign node40473 = (inp[13]) ? node40501 : node40474;
												assign node40474 = (inp[1]) ? node40486 : node40475;
													assign node40475 = (inp[14]) ? node40481 : node40476;
														assign node40476 = (inp[8]) ? 4'b1110 : node40477;
															assign node40477 = (inp[6]) ? 4'b0111 : 4'b0111;
														assign node40481 = (inp[8]) ? node40483 : 4'b1110;
															assign node40483 = (inp[6]) ? 4'b1111 : 4'b0111;
													assign node40486 = (inp[14]) ? node40494 : node40487;
														assign node40487 = (inp[8]) ? node40491 : node40488;
															assign node40488 = (inp[6]) ? 4'b1111 : 4'b0111;
															assign node40491 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node40494 = (inp[8]) ? node40498 : node40495;
															assign node40495 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node40498 = (inp[6]) ? 4'b0111 : 4'b0111;
												assign node40501 = (inp[11]) ? node40515 : node40502;
													assign node40502 = (inp[6]) ? node40508 : node40503;
														assign node40503 = (inp[1]) ? 4'b0110 : node40504;
															assign node40504 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node40508 = (inp[1]) ? node40512 : node40509;
															assign node40509 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node40512 = (inp[8]) ? 4'b1110 : 4'b1110;
													assign node40515 = (inp[14]) ? node40523 : node40516;
														assign node40516 = (inp[8]) ? node40520 : node40517;
															assign node40517 = (inp[1]) ? 4'b1111 : 4'b0111;
															assign node40520 = (inp[1]) ? 4'b0110 : 4'b0110;
														assign node40523 = (inp[8]) ? node40527 : node40524;
															assign node40524 = (inp[6]) ? 4'b1110 : 4'b0110;
															assign node40527 = (inp[6]) ? 4'b0111 : 4'b1111;
											assign node40530 = (inp[6]) ? node40558 : node40531;
												assign node40531 = (inp[11]) ? node40547 : node40532;
													assign node40532 = (inp[1]) ? node40540 : node40533;
														assign node40533 = (inp[14]) ? node40537 : node40534;
															assign node40534 = (inp[8]) ? 4'b0111 : 4'b1110;
															assign node40537 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node40540 = (inp[13]) ? node40544 : node40541;
															assign node40541 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node40544 = (inp[8]) ? 4'b0110 : 4'b0110;
													assign node40547 = (inp[1]) ? node40555 : node40548;
														assign node40548 = (inp[13]) ? node40552 : node40549;
															assign node40549 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node40552 = (inp[14]) ? 4'b1111 : 4'b0110;
														assign node40555 = (inp[13]) ? 4'b1110 : 4'b1111;
												assign node40558 = (inp[11]) ? node40572 : node40559;
													assign node40559 = (inp[13]) ? node40567 : node40560;
														assign node40560 = (inp[1]) ? node40564 : node40561;
															assign node40561 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node40564 = (inp[14]) ? 4'b1110 : 4'b0110;
														assign node40567 = (inp[8]) ? node40569 : 4'b1111;
															assign node40569 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node40572 = (inp[1]) ? node40580 : node40573;
														assign node40573 = (inp[13]) ? node40577 : node40574;
															assign node40574 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node40577 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node40580 = (inp[14]) ? node40584 : node40581;
															assign node40581 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node40584 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node40587 = (inp[1]) ? node40649 : node40588;
											assign node40588 = (inp[7]) ? node40620 : node40589;
												assign node40589 = (inp[13]) ? node40605 : node40590;
													assign node40590 = (inp[8]) ? node40598 : node40591;
														assign node40591 = (inp[14]) ? node40595 : node40592;
															assign node40592 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node40595 = (inp[6]) ? 4'b0100 : 4'b0100;
														assign node40598 = (inp[14]) ? node40602 : node40599;
															assign node40599 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node40602 = (inp[11]) ? 4'b0101 : 4'b0101;
													assign node40605 = (inp[6]) ? node40613 : node40606;
														assign node40606 = (inp[11]) ? node40610 : node40607;
															assign node40607 = (inp[8]) ? 4'b0100 : 4'b1100;
															assign node40610 = (inp[14]) ? 4'b0100 : 4'b0100;
														assign node40613 = (inp[11]) ? node40617 : node40614;
															assign node40614 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node40617 = (inp[14]) ? 4'b1100 : 4'b1100;
												assign node40620 = (inp[13]) ? node40634 : node40621;
													assign node40621 = (inp[8]) ? node40627 : node40622;
														assign node40622 = (inp[14]) ? 4'b1101 : node40623;
															assign node40623 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node40627 = (inp[14]) ? node40631 : node40628;
															assign node40628 = (inp[11]) ? 4'b0101 : 4'b1101;
															assign node40631 = (inp[11]) ? 4'b0100 : 4'b0100;
													assign node40634 = (inp[11]) ? node40642 : node40635;
														assign node40635 = (inp[6]) ? node40639 : node40636;
															assign node40636 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node40639 = (inp[8]) ? 4'b1100 : 4'b0100;
														assign node40642 = (inp[6]) ? node40646 : node40643;
															assign node40643 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node40646 = (inp[14]) ? 4'b0100 : 4'b0100;
											assign node40649 = (inp[6]) ? node40679 : node40650;
												assign node40650 = (inp[11]) ? node40666 : node40651;
													assign node40651 = (inp[13]) ? node40659 : node40652;
														assign node40652 = (inp[7]) ? node40656 : node40653;
															assign node40653 = (inp[8]) ? 4'b0100 : 4'b1100;
															assign node40656 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node40659 = (inp[8]) ? node40663 : node40660;
															assign node40660 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node40663 = (inp[7]) ? 4'b0100 : 4'b0100;
													assign node40666 = (inp[13]) ? node40672 : node40667;
														assign node40667 = (inp[8]) ? node40669 : 4'b0100;
															assign node40669 = (inp[7]) ? 4'b1100 : 4'b0100;
														assign node40672 = (inp[8]) ? node40676 : node40673;
															assign node40673 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node40676 = (inp[14]) ? 4'b1100 : 4'b1100;
												assign node40679 = (inp[11]) ? node40693 : node40680;
													assign node40680 = (inp[13]) ? node40688 : node40681;
														assign node40681 = (inp[8]) ? node40685 : node40682;
															assign node40682 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node40685 = (inp[7]) ? 4'b1100 : 4'b0100;
														assign node40688 = (inp[14]) ? node40690 : 4'b1101;
															assign node40690 = (inp[8]) ? 4'b1100 : 4'b1100;
													assign node40693 = (inp[13]) ? node40699 : node40694;
														assign node40694 = (inp[14]) ? 4'b0101 : node40695;
															assign node40695 = (inp[7]) ? 4'b0100 : 4'b1100;
														assign node40699 = (inp[7]) ? node40703 : node40700;
															assign node40700 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node40703 = (inp[14]) ? 4'b0100 : 4'b0101;
								assign node40706 = (inp[0]) ? node40956 : node40707;
									assign node40707 = (inp[15]) ? node40829 : node40708;
										assign node40708 = (inp[13]) ? node40768 : node40709;
											assign node40709 = (inp[7]) ? node40737 : node40710;
												assign node40710 = (inp[14]) ? node40726 : node40711;
													assign node40711 = (inp[8]) ? node40719 : node40712;
														assign node40712 = (inp[6]) ? node40716 : node40713;
															assign node40713 = (inp[11]) ? 4'b0101 : 4'b1101;
															assign node40716 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node40719 = (inp[6]) ? node40723 : node40720;
															assign node40720 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node40723 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node40726 = (inp[8]) ? node40734 : node40727;
														assign node40727 = (inp[6]) ? node40731 : node40728;
															assign node40728 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node40731 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node40734 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node40737 = (inp[14]) ? node40753 : node40738;
													assign node40738 = (inp[8]) ? node40746 : node40739;
														assign node40739 = (inp[1]) ? node40743 : node40740;
															assign node40740 = (inp[11]) ? 4'b0100 : 4'b0100;
															assign node40743 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node40746 = (inp[6]) ? node40750 : node40747;
															assign node40747 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node40750 = (inp[11]) ? 4'b0101 : 4'b0101;
													assign node40753 = (inp[8]) ? node40761 : node40754;
														assign node40754 = (inp[6]) ? node40758 : node40755;
															assign node40755 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node40758 = (inp[11]) ? 4'b0101 : 4'b0101;
														assign node40761 = (inp[6]) ? node40765 : node40762;
															assign node40762 = (inp[1]) ? 4'b0100 : 4'b1100;
															assign node40765 = (inp[11]) ? 4'b0100 : 4'b0100;
											assign node40768 = (inp[1]) ? node40798 : node40769;
												assign node40769 = (inp[6]) ? node40785 : node40770;
													assign node40770 = (inp[14]) ? node40778 : node40771;
														assign node40771 = (inp[11]) ? node40775 : node40772;
															assign node40772 = (inp[7]) ? 4'b0100 : 4'b1100;
															assign node40775 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node40778 = (inp[11]) ? node40782 : node40779;
															assign node40779 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node40782 = (inp[7]) ? 4'b1100 : 4'b0100;
													assign node40785 = (inp[8]) ? node40793 : node40786;
														assign node40786 = (inp[11]) ? node40790 : node40787;
															assign node40787 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node40790 = (inp[7]) ? 4'b0101 : 4'b1100;
														assign node40793 = (inp[11]) ? node40795 : 4'b1101;
															assign node40795 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node40798 = (inp[7]) ? node40814 : node40799;
													assign node40799 = (inp[8]) ? node40807 : node40800;
														assign node40800 = (inp[14]) ? node40804 : node40801;
															assign node40801 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node40804 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node40807 = (inp[14]) ? node40811 : node40808;
															assign node40808 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node40811 = (inp[6]) ? 4'b0101 : 4'b0101;
													assign node40814 = (inp[6]) ? node40822 : node40815;
														assign node40815 = (inp[11]) ? node40819 : node40816;
															assign node40816 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node40819 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node40822 = (inp[11]) ? node40826 : node40823;
															assign node40823 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node40826 = (inp[14]) ? 4'b0100 : 4'b0100;
										assign node40829 = (inp[7]) ? node40893 : node40830;
											assign node40830 = (inp[1]) ? node40862 : node40831;
												assign node40831 = (inp[8]) ? node40847 : node40832;
													assign node40832 = (inp[14]) ? node40840 : node40833;
														assign node40833 = (inp[6]) ? node40837 : node40834;
															assign node40834 = (inp[11]) ? 4'b0111 : 4'b1111;
															assign node40837 = (inp[11]) ? 4'b1111 : 4'b0111;
														assign node40840 = (inp[13]) ? node40844 : node40841;
															assign node40841 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node40844 = (inp[11]) ? 4'b0110 : 4'b0110;
													assign node40847 = (inp[14]) ? node40855 : node40848;
														assign node40848 = (inp[11]) ? node40852 : node40849;
															assign node40849 = (inp[6]) ? 4'b0110 : 4'b1110;
															assign node40852 = (inp[6]) ? 4'b1110 : 4'b0110;
														assign node40855 = (inp[6]) ? node40859 : node40856;
															assign node40856 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node40859 = (inp[13]) ? 4'b0111 : 4'b0111;
												assign node40862 = (inp[6]) ? node40878 : node40863;
													assign node40863 = (inp[13]) ? node40871 : node40864;
														assign node40864 = (inp[11]) ? node40868 : node40865;
															assign node40865 = (inp[8]) ? 4'b0110 : 4'b1110;
															assign node40868 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node40871 = (inp[11]) ? node40875 : node40872;
															assign node40872 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node40875 = (inp[14]) ? 4'b1110 : 4'b1110;
													assign node40878 = (inp[11]) ? node40886 : node40879;
														assign node40879 = (inp[13]) ? node40883 : node40880;
															assign node40880 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node40883 = (inp[14]) ? 4'b1110 : 4'b1110;
														assign node40886 = (inp[14]) ? node40890 : node40887;
															assign node40887 = (inp[13]) ? 4'b0110 : 4'b1110;
															assign node40890 = (inp[8]) ? 4'b0111 : 4'b0110;
											assign node40893 = (inp[1]) ? node40925 : node40894;
												assign node40894 = (inp[11]) ? node40910 : node40895;
													assign node40895 = (inp[6]) ? node40903 : node40896;
														assign node40896 = (inp[13]) ? node40900 : node40897;
															assign node40897 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node40900 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node40903 = (inp[13]) ? node40907 : node40904;
															assign node40904 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node40907 = (inp[8]) ? 4'b1110 : 4'b0110;
													assign node40910 = (inp[6]) ? node40918 : node40911;
														assign node40911 = (inp[13]) ? node40915 : node40912;
															assign node40912 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node40915 = (inp[8]) ? 4'b1110 : 4'b0110;
														assign node40918 = (inp[13]) ? node40922 : node40919;
															assign node40919 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node40922 = (inp[8]) ? 4'b0110 : 4'b0110;
												assign node40925 = (inp[13]) ? node40941 : node40926;
													assign node40926 = (inp[8]) ? node40934 : node40927;
														assign node40927 = (inp[14]) ? node40931 : node40928;
															assign node40928 = (inp[11]) ? 4'b0110 : 4'b1110;
															assign node40931 = (inp[6]) ? 4'b0111 : 4'b0111;
														assign node40934 = (inp[14]) ? node40938 : node40935;
															assign node40935 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node40938 = (inp[6]) ? 4'b0110 : 4'b0110;
													assign node40941 = (inp[14]) ? node40949 : node40942;
														assign node40942 = (inp[8]) ? node40946 : node40943;
															assign node40943 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node40946 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node40949 = (inp[8]) ? node40953 : node40950;
															assign node40950 = (inp[6]) ? 4'b0111 : 4'b1111;
															assign node40953 = (inp[11]) ? 4'b0110 : 4'b1110;
									assign node40956 = (inp[15]) ? node41078 : node40957;
										assign node40957 = (inp[11]) ? node41017 : node40958;
											assign node40958 = (inp[7]) ? node40986 : node40959;
												assign node40959 = (inp[6]) ? node40975 : node40960;
													assign node40960 = (inp[13]) ? node40968 : node40961;
														assign node40961 = (inp[14]) ? node40965 : node40962;
															assign node40962 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node40965 = (inp[8]) ? 4'b0111 : 4'b1110;
														assign node40968 = (inp[1]) ? node40972 : node40969;
															assign node40969 = (inp[8]) ? 4'b0111 : 4'b1110;
															assign node40972 = (inp[14]) ? 4'b0110 : 4'b0110;
													assign node40975 = (inp[8]) ? node40979 : node40976;
														assign node40976 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node40979 = (inp[14]) ? node40983 : node40980;
															assign node40980 = (inp[13]) ? 4'b0110 : 4'b0110;
															assign node40983 = (inp[13]) ? 4'b1111 : 4'b0111;
												assign node40986 = (inp[6]) ? node41002 : node40987;
													assign node40987 = (inp[1]) ? node40995 : node40988;
														assign node40988 = (inp[13]) ? node40992 : node40989;
															assign node40989 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node40992 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node40995 = (inp[8]) ? node40999 : node40996;
															assign node40996 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node40999 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node41002 = (inp[1]) ? node41010 : node41003;
														assign node41003 = (inp[13]) ? node41007 : node41004;
															assign node41004 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node41007 = (inp[14]) ? 4'b1110 : 4'b0110;
														assign node41010 = (inp[14]) ? node41014 : node41011;
															assign node41011 = (inp[8]) ? 4'b1111 : 4'b0110;
															assign node41014 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node41017 = (inp[6]) ? node41049 : node41018;
												assign node41018 = (inp[1]) ? node41034 : node41019;
													assign node41019 = (inp[13]) ? node41027 : node41020;
														assign node41020 = (inp[14]) ? node41024 : node41021;
															assign node41021 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node41024 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node41027 = (inp[14]) ? node41031 : node41028;
															assign node41028 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node41031 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node41034 = (inp[13]) ? node41042 : node41035;
														assign node41035 = (inp[8]) ? node41039 : node41036;
															assign node41036 = (inp[14]) ? 4'b1111 : 4'b0110;
															assign node41039 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node41042 = (inp[7]) ? node41046 : node41043;
															assign node41043 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node41046 = (inp[14]) ? 4'b1110 : 4'b1110;
												assign node41049 = (inp[13]) ? node41063 : node41050;
													assign node41050 = (inp[1]) ? node41058 : node41051;
														assign node41051 = (inp[14]) ? node41055 : node41052;
															assign node41052 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node41055 = (inp[7]) ? 4'b1110 : 4'b1110;
														assign node41058 = (inp[14]) ? 4'b0110 : node41059;
															assign node41059 = (inp[7]) ? 4'b0110 : 4'b1110;
													assign node41063 = (inp[1]) ? node41071 : node41064;
														assign node41064 = (inp[7]) ? node41068 : node41065;
															assign node41065 = (inp[8]) ? 4'b0110 : 4'b1110;
															assign node41068 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node41071 = (inp[8]) ? node41075 : node41072;
															assign node41072 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node41075 = (inp[7]) ? 4'b0110 : 4'b0110;
										assign node41078 = (inp[1]) ? node41142 : node41079;
											assign node41079 = (inp[7]) ? node41111 : node41080;
												assign node41080 = (inp[14]) ? node41096 : node41081;
													assign node41081 = (inp[8]) ? node41089 : node41082;
														assign node41082 = (inp[13]) ? node41086 : node41083;
															assign node41083 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node41086 = (inp[6]) ? 4'b0101 : 4'b0101;
														assign node41089 = (inp[6]) ? node41093 : node41090;
															assign node41090 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node41093 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node41096 = (inp[8]) ? node41104 : node41097;
														assign node41097 = (inp[11]) ? node41101 : node41098;
															assign node41098 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node41101 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node41104 = (inp[13]) ? node41108 : node41105;
															assign node41105 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node41108 = (inp[6]) ? 4'b0101 : 4'b0101;
												assign node41111 = (inp[13]) ? node41127 : node41112;
													assign node41112 = (inp[6]) ? node41120 : node41113;
														assign node41113 = (inp[11]) ? node41117 : node41114;
															assign node41114 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node41117 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node41120 = (inp[11]) ? node41124 : node41121;
															assign node41121 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node41124 = (inp[8]) ? 4'b1100 : 4'b1100;
													assign node41127 = (inp[8]) ? node41135 : node41128;
														assign node41128 = (inp[14]) ? node41132 : node41129;
															assign node41129 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node41132 = (inp[6]) ? 4'b0101 : 4'b0101;
														assign node41135 = (inp[14]) ? node41139 : node41136;
															assign node41136 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node41139 = (inp[11]) ? 4'b0100 : 4'b0100;
											assign node41142 = (inp[6]) ? node41174 : node41143;
												assign node41143 = (inp[11]) ? node41159 : node41144;
													assign node41144 = (inp[13]) ? node41152 : node41145;
														assign node41145 = (inp[7]) ? node41149 : node41146;
															assign node41146 = (inp[14]) ? 4'b0101 : 4'b1100;
															assign node41149 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node41152 = (inp[14]) ? node41156 : node41153;
															assign node41153 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node41156 = (inp[7]) ? 4'b0100 : 4'b0100;
													assign node41159 = (inp[13]) ? node41167 : node41160;
														assign node41160 = (inp[8]) ? node41164 : node41161;
															assign node41161 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node41164 = (inp[14]) ? 4'b1101 : 4'b0100;
														assign node41167 = (inp[14]) ? node41171 : node41168;
															assign node41168 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node41171 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node41174 = (inp[11]) ? node41188 : node41175;
													assign node41175 = (inp[7]) ? node41183 : node41176;
														assign node41176 = (inp[13]) ? node41180 : node41177;
															assign node41177 = (inp[14]) ? 4'b1101 : 4'b0100;
															assign node41180 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node41183 = (inp[14]) ? node41185 : 4'b1101;
															assign node41185 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node41188 = (inp[13]) ? node41194 : node41189;
														assign node41189 = (inp[14]) ? 4'b0101 : node41190;
															assign node41190 = (inp[7]) ? 4'b0101 : 4'b1100;
														assign node41194 = (inp[8]) ? node41198 : node41195;
															assign node41195 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node41198 = (inp[14]) ? 4'b0100 : 4'b0101;
						assign node41201 = (inp[14]) ? node42129 : node41202;
							assign node41202 = (inp[8]) ? node41660 : node41203;
								assign node41203 = (inp[7]) ? node41431 : node41204;
									assign node41204 = (inp[3]) ? node41328 : node41205;
										assign node41205 = (inp[15]) ? node41269 : node41206;
											assign node41206 = (inp[6]) ? node41238 : node41207;
												assign node41207 = (inp[11]) ? node41223 : node41208;
													assign node41208 = (inp[13]) ? node41216 : node41209;
														assign node41209 = (inp[0]) ? node41213 : node41210;
															assign node41210 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node41213 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node41216 = (inp[1]) ? node41220 : node41217;
															assign node41217 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node41220 = (inp[5]) ? 4'b0100 : 4'b0100;
													assign node41223 = (inp[1]) ? node41231 : node41224;
														assign node41224 = (inp[5]) ? node41228 : node41225;
															assign node41225 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node41228 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node41231 = (inp[13]) ? node41235 : node41232;
															assign node41232 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node41235 = (inp[0]) ? 4'b1100 : 4'b1100;
												assign node41238 = (inp[11]) ? node41254 : node41239;
													assign node41239 = (inp[13]) ? node41247 : node41240;
														assign node41240 = (inp[0]) ? node41244 : node41241;
															assign node41241 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node41244 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node41247 = (inp[1]) ? node41251 : node41248;
															assign node41248 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node41251 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node41254 = (inp[1]) ? node41262 : node41255;
														assign node41255 = (inp[0]) ? node41259 : node41256;
															assign node41256 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node41259 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node41262 = (inp[13]) ? node41266 : node41263;
															assign node41263 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node41266 = (inp[5]) ? 4'b0100 : 4'b0100;
											assign node41269 = (inp[5]) ? node41299 : node41270;
												assign node41270 = (inp[0]) ? node41284 : node41271;
													assign node41271 = (inp[1]) ? node41279 : node41272;
														assign node41272 = (inp[6]) ? node41276 : node41273;
															assign node41273 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node41276 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node41279 = (inp[6]) ? node41281 : 4'b0100;
															assign node41281 = (inp[13]) ? 4'b0100 : 4'b0100;
													assign node41284 = (inp[13]) ? node41292 : node41285;
														assign node41285 = (inp[1]) ? node41289 : node41286;
															assign node41286 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node41289 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node41292 = (inp[6]) ? node41296 : node41293;
															assign node41293 = (inp[11]) ? 4'b0110 : 4'b1110;
															assign node41296 = (inp[1]) ? 4'b0110 : 4'b0110;
												assign node41299 = (inp[0]) ? node41315 : node41300;
													assign node41300 = (inp[11]) ? node41308 : node41301;
														assign node41301 = (inp[6]) ? node41305 : node41302;
															assign node41302 = (inp[1]) ? 4'b0110 : 4'b1110;
															assign node41305 = (inp[1]) ? 4'b1110 : 4'b0110;
														assign node41308 = (inp[6]) ? node41312 : node41309;
															assign node41309 = (inp[13]) ? 4'b0110 : 4'b0110;
															assign node41312 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node41315 = (inp[6]) ? node41323 : node41316;
														assign node41316 = (inp[11]) ? node41320 : node41317;
															assign node41317 = (inp[1]) ? 4'b0100 : 4'b1100;
															assign node41320 = (inp[1]) ? 4'b0100 : 4'b0100;
														assign node41323 = (inp[1]) ? node41325 : 4'b0100;
															assign node41325 = (inp[13]) ? 4'b0100 : 4'b1100;
										assign node41328 = (inp[15]) ? node41376 : node41329;
											assign node41329 = (inp[0]) ? node41353 : node41330;
												assign node41330 = (inp[1]) ? node41338 : node41331;
													assign node41331 = (inp[11]) ? node41335 : node41332;
														assign node41332 = (inp[6]) ? 4'b0100 : 4'b1100;
														assign node41335 = (inp[6]) ? 4'b1100 : 4'b0100;
													assign node41338 = (inp[11]) ? node41346 : node41339;
														assign node41339 = (inp[5]) ? node41343 : node41340;
															assign node41340 = (inp[13]) ? 4'b0100 : 4'b0100;
															assign node41343 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node41346 = (inp[13]) ? node41350 : node41347;
															assign node41347 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node41350 = (inp[6]) ? 4'b0100 : 4'b1100;
												assign node41353 = (inp[6]) ? node41365 : node41354;
													assign node41354 = (inp[11]) ? node41360 : node41355;
														assign node41355 = (inp[1]) ? node41357 : 4'b1110;
															assign node41357 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node41360 = (inp[13]) ? node41362 : 4'b0110;
															assign node41362 = (inp[1]) ? 4'b1110 : 4'b0110;
													assign node41365 = (inp[11]) ? node41371 : node41366;
														assign node41366 = (inp[1]) ? node41368 : 4'b0110;
															assign node41368 = (inp[13]) ? 4'b1110 : 4'b0110;
														assign node41371 = (inp[13]) ? node41373 : 4'b1110;
															assign node41373 = (inp[1]) ? 4'b0110 : 4'b1110;
											assign node41376 = (inp[0]) ? node41400 : node41377;
												assign node41377 = (inp[13]) ? node41385 : node41378;
													assign node41378 = (inp[6]) ? node41382 : node41379;
														assign node41379 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node41382 = (inp[11]) ? 4'b1110 : 4'b0110;
													assign node41385 = (inp[11]) ? node41393 : node41386;
														assign node41386 = (inp[5]) ? node41390 : node41387;
															assign node41387 = (inp[1]) ? 4'b0110 : 4'b0110;
															assign node41390 = (inp[1]) ? 4'b0110 : 4'b1110;
														assign node41393 = (inp[6]) ? node41397 : node41394;
															assign node41394 = (inp[1]) ? 4'b1110 : 4'b0110;
															assign node41397 = (inp[1]) ? 4'b0110 : 4'b1110;
												assign node41400 = (inp[5]) ? node41416 : node41401;
													assign node41401 = (inp[13]) ? node41409 : node41402;
														assign node41402 = (inp[11]) ? node41406 : node41403;
															assign node41403 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node41406 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node41409 = (inp[11]) ? node41413 : node41410;
															assign node41410 = (inp[1]) ? 4'b0100 : 4'b1100;
															assign node41413 = (inp[6]) ? 4'b0100 : 4'b0100;
													assign node41416 = (inp[11]) ? node41424 : node41417;
														assign node41417 = (inp[6]) ? node41421 : node41418;
															assign node41418 = (inp[1]) ? 4'b0100 : 4'b1100;
															assign node41421 = (inp[13]) ? 4'b0100 : 4'b0100;
														assign node41424 = (inp[6]) ? node41428 : node41425;
															assign node41425 = (inp[1]) ? 4'b0100 : 4'b0100;
															assign node41428 = (inp[1]) ? 4'b0100 : 4'b1100;
									assign node41431 = (inp[5]) ? node41553 : node41432;
										assign node41432 = (inp[1]) ? node41494 : node41433;
											assign node41433 = (inp[3]) ? node41463 : node41434;
												assign node41434 = (inp[13]) ? node41448 : node41435;
													assign node41435 = (inp[0]) ? node41443 : node41436;
														assign node41436 = (inp[15]) ? node41440 : node41437;
															assign node41437 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node41440 = (inp[11]) ? 4'b0101 : 4'b0101;
														assign node41443 = (inp[15]) ? 4'b1111 : node41444;
															assign node41444 = (inp[6]) ? 4'b0101 : 4'b0101;
													assign node41448 = (inp[15]) ? node41456 : node41449;
														assign node41449 = (inp[0]) ? node41453 : node41450;
															assign node41450 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node41453 = (inp[11]) ? 4'b0101 : 4'b0101;
														assign node41456 = (inp[0]) ? node41460 : node41457;
															assign node41457 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node41460 = (inp[11]) ? 4'b0111 : 4'b0111;
												assign node41463 = (inp[11]) ? node41479 : node41464;
													assign node41464 = (inp[0]) ? node41472 : node41465;
														assign node41465 = (inp[15]) ? node41469 : node41466;
															assign node41466 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node41469 = (inp[6]) ? 4'b0111 : 4'b0111;
														assign node41472 = (inp[15]) ? node41476 : node41473;
															assign node41473 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node41476 = (inp[13]) ? 4'b0101 : 4'b0101;
													assign node41479 = (inp[6]) ? node41487 : node41480;
														assign node41480 = (inp[13]) ? node41484 : node41481;
															assign node41481 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node41484 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node41487 = (inp[13]) ? node41491 : node41488;
															assign node41488 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node41491 = (inp[15]) ? 4'b0101 : 4'b0101;
											assign node41494 = (inp[13]) ? node41526 : node41495;
												assign node41495 = (inp[15]) ? node41511 : node41496;
													assign node41496 = (inp[6]) ? node41504 : node41497;
														assign node41497 = (inp[11]) ? node41501 : node41498;
															assign node41498 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node41501 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node41504 = (inp[11]) ? node41508 : node41505;
															assign node41505 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node41508 = (inp[3]) ? 4'b0101 : 4'b0101;
													assign node41511 = (inp[6]) ? node41519 : node41512;
														assign node41512 = (inp[11]) ? node41516 : node41513;
															assign node41513 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node41516 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node41519 = (inp[11]) ? node41523 : node41520;
															assign node41520 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node41523 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node41526 = (inp[11]) ? node41542 : node41527;
													assign node41527 = (inp[6]) ? node41535 : node41528;
														assign node41528 = (inp[3]) ? node41532 : node41529;
															assign node41529 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node41532 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node41535 = (inp[15]) ? node41539 : node41536;
															assign node41536 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node41539 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node41542 = (inp[6]) ? node41548 : node41543;
														assign node41543 = (inp[15]) ? 4'b1101 : node41544;
															assign node41544 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node41548 = (inp[15]) ? node41550 : 4'b0101;
															assign node41550 = (inp[3]) ? 4'b0101 : 4'b0101;
										assign node41553 = (inp[13]) ? node41615 : node41554;
											assign node41554 = (inp[6]) ? node41584 : node41555;
												assign node41555 = (inp[3]) ? node41569 : node41556;
													assign node41556 = (inp[1]) ? node41564 : node41557;
														assign node41557 = (inp[11]) ? node41561 : node41558;
															assign node41558 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node41561 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node41564 = (inp[11]) ? node41566 : 4'b0111;
															assign node41566 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node41569 = (inp[11]) ? node41577 : node41570;
														assign node41570 = (inp[1]) ? node41574 : node41571;
															assign node41571 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node41574 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node41577 = (inp[1]) ? node41581 : node41578;
															assign node41578 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node41581 = (inp[0]) ? 4'b1101 : 4'b1101;
												assign node41584 = (inp[1]) ? node41600 : node41585;
													assign node41585 = (inp[11]) ? node41593 : node41586;
														assign node41586 = (inp[3]) ? node41590 : node41587;
															assign node41587 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node41590 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node41593 = (inp[0]) ? node41597 : node41594;
															assign node41594 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node41597 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node41600 = (inp[11]) ? node41608 : node41601;
														assign node41601 = (inp[0]) ? node41605 : node41602;
															assign node41602 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node41605 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node41608 = (inp[15]) ? node41612 : node41609;
															assign node41609 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node41612 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node41615 = (inp[11]) ? node41637 : node41616;
												assign node41616 = (inp[6]) ? node41624 : node41617;
													assign node41617 = (inp[0]) ? node41621 : node41618;
														assign node41618 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node41621 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node41624 = (inp[3]) ? node41632 : node41625;
														assign node41625 = (inp[0]) ? node41629 : node41626;
															assign node41626 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node41629 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node41632 = (inp[1]) ? 4'b1101 : node41633;
															assign node41633 = (inp[0]) ? 4'b1101 : 4'b1101;
												assign node41637 = (inp[6]) ? node41653 : node41638;
													assign node41638 = (inp[1]) ? node41646 : node41639;
														assign node41639 = (inp[15]) ? node41643 : node41640;
															assign node41640 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node41643 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node41646 = (inp[15]) ? node41650 : node41647;
															assign node41647 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node41650 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node41653 = (inp[0]) ? node41657 : node41654;
														assign node41654 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node41657 = (inp[15]) ? 4'b0101 : 4'b0111;
								assign node41660 = (inp[7]) ? node41896 : node41661;
									assign node41661 = (inp[13]) ? node41785 : node41662;
										assign node41662 = (inp[15]) ? node41724 : node41663;
											assign node41663 = (inp[0]) ? node41695 : node41664;
												assign node41664 = (inp[5]) ? node41680 : node41665;
													assign node41665 = (inp[3]) ? node41673 : node41666;
														assign node41666 = (inp[11]) ? node41670 : node41667;
															assign node41667 = (inp[6]) ? 4'b0111 : 4'b1111;
															assign node41670 = (inp[1]) ? 4'b0111 : 4'b0111;
														assign node41673 = (inp[11]) ? node41677 : node41674;
															assign node41674 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node41677 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node41680 = (inp[11]) ? node41688 : node41681;
														assign node41681 = (inp[6]) ? node41685 : node41682;
															assign node41682 = (inp[1]) ? 4'b0101 : 4'b1101;
															assign node41685 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node41688 = (inp[6]) ? node41692 : node41689;
															assign node41689 = (inp[1]) ? 4'b1101 : 4'b0101;
															assign node41692 = (inp[1]) ? 4'b0101 : 4'b1101;
												assign node41695 = (inp[3]) ? node41709 : node41696;
													assign node41696 = (inp[5]) ? node41704 : node41697;
														assign node41697 = (inp[11]) ? node41701 : node41698;
															assign node41698 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node41701 = (inp[6]) ? 4'b0101 : 4'b0101;
														assign node41704 = (inp[6]) ? 4'b1111 : node41705;
															assign node41705 = (inp[1]) ? 4'b0111 : 4'b0111;
													assign node41709 = (inp[1]) ? node41717 : node41710;
														assign node41710 = (inp[5]) ? node41714 : node41711;
															assign node41711 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node41714 = (inp[6]) ? 4'b0111 : 4'b0111;
														assign node41717 = (inp[6]) ? node41721 : node41718;
															assign node41718 = (inp[11]) ? 4'b1111 : 4'b0111;
															assign node41721 = (inp[11]) ? 4'b0111 : 4'b1111;
											assign node41724 = (inp[0]) ? node41756 : node41725;
												assign node41725 = (inp[5]) ? node41741 : node41726;
													assign node41726 = (inp[3]) ? node41734 : node41727;
														assign node41727 = (inp[6]) ? node41731 : node41728;
															assign node41728 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node41731 = (inp[1]) ? 4'b0101 : 4'b0101;
														assign node41734 = (inp[1]) ? node41738 : node41735;
															assign node41735 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node41738 = (inp[6]) ? 4'b0111 : 4'b0111;
													assign node41741 = (inp[11]) ? node41749 : node41742;
														assign node41742 = (inp[3]) ? node41746 : node41743;
															assign node41743 = (inp[1]) ? 4'b0111 : 4'b0111;
															assign node41746 = (inp[6]) ? 4'b0111 : 4'b0111;
														assign node41749 = (inp[6]) ? node41753 : node41750;
															assign node41750 = (inp[1]) ? 4'b1111 : 4'b0111;
															assign node41753 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node41756 = (inp[3]) ? node41770 : node41757;
													assign node41757 = (inp[5]) ? node41765 : node41758;
														assign node41758 = (inp[1]) ? node41762 : node41759;
															assign node41759 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node41762 = (inp[6]) ? 4'b0111 : 4'b0111;
														assign node41765 = (inp[1]) ? node41767 : 4'b0101;
															assign node41767 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node41770 = (inp[1]) ? node41778 : node41771;
														assign node41771 = (inp[5]) ? node41775 : node41772;
															assign node41772 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node41775 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node41778 = (inp[5]) ? node41782 : node41779;
															assign node41779 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node41782 = (inp[6]) ? 4'b0101 : 4'b0101;
										assign node41785 = (inp[3]) ? node41849 : node41786;
											assign node41786 = (inp[5]) ? node41818 : node41787;
												assign node41787 = (inp[11]) ? node41803 : node41788;
													assign node41788 = (inp[6]) ? node41796 : node41789;
														assign node41789 = (inp[15]) ? node41793 : node41790;
															assign node41790 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node41793 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node41796 = (inp[15]) ? node41800 : node41797;
															assign node41797 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node41800 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node41803 = (inp[6]) ? node41811 : node41804;
														assign node41804 = (inp[0]) ? node41808 : node41805;
															assign node41805 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node41808 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node41811 = (inp[1]) ? node41815 : node41812;
															assign node41812 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node41815 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node41818 = (inp[0]) ? node41834 : node41819;
													assign node41819 = (inp[15]) ? node41827 : node41820;
														assign node41820 = (inp[11]) ? node41824 : node41821;
															assign node41821 = (inp[6]) ? 4'b1101 : 4'b0101;
															assign node41824 = (inp[6]) ? 4'b0101 : 4'b1101;
														assign node41827 = (inp[1]) ? node41831 : node41828;
															assign node41828 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node41831 = (inp[11]) ? 4'b0111 : 4'b0111;
													assign node41834 = (inp[15]) ? node41842 : node41835;
														assign node41835 = (inp[1]) ? node41839 : node41836;
															assign node41836 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node41839 = (inp[11]) ? 4'b0111 : 4'b0111;
														assign node41842 = (inp[6]) ? node41846 : node41843;
															assign node41843 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node41846 = (inp[11]) ? 4'b0101 : 4'b1101;
											assign node41849 = (inp[6]) ? node41865 : node41850;
												assign node41850 = (inp[11]) ? node41858 : node41851;
													assign node41851 = (inp[15]) ? node41855 : node41852;
														assign node41852 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node41855 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node41858 = (inp[0]) ? node41862 : node41859;
														assign node41859 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node41862 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node41865 = (inp[11]) ? node41881 : node41866;
													assign node41866 = (inp[5]) ? node41874 : node41867;
														assign node41867 = (inp[0]) ? node41871 : node41868;
															assign node41868 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node41871 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node41874 = (inp[1]) ? node41878 : node41875;
															assign node41875 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node41878 = (inp[0]) ? 4'b1101 : 4'b1101;
													assign node41881 = (inp[1]) ? node41889 : node41882;
														assign node41882 = (inp[0]) ? node41886 : node41883;
															assign node41883 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node41886 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node41889 = (inp[15]) ? node41893 : node41890;
															assign node41890 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node41893 = (inp[0]) ? 4'b0101 : 4'b0111;
									assign node41896 = (inp[13]) ? node42020 : node41897;
										assign node41897 = (inp[0]) ? node41961 : node41898;
											assign node41898 = (inp[15]) ? node41930 : node41899;
												assign node41899 = (inp[3]) ? node41915 : node41900;
													assign node41900 = (inp[5]) ? node41908 : node41901;
														assign node41901 = (inp[1]) ? node41905 : node41902;
															assign node41902 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node41905 = (inp[6]) ? 4'b0110 : 4'b0110;
														assign node41908 = (inp[11]) ? node41912 : node41909;
															assign node41909 = (inp[1]) ? 4'b0100 : 4'b0100;
															assign node41912 = (inp[6]) ? 4'b0100 : 4'b0100;
													assign node41915 = (inp[6]) ? node41923 : node41916;
														assign node41916 = (inp[5]) ? node41920 : node41917;
															assign node41917 = (inp[1]) ? 4'b0100 : 4'b1100;
															assign node41920 = (inp[1]) ? 4'b1100 : 4'b0100;
														assign node41923 = (inp[5]) ? node41927 : node41924;
															assign node41924 = (inp[11]) ? 4'b0100 : 4'b0100;
															assign node41927 = (inp[11]) ? 4'b0100 : 4'b0100;
												assign node41930 = (inp[3]) ? node41946 : node41931;
													assign node41931 = (inp[5]) ? node41939 : node41932;
														assign node41932 = (inp[1]) ? node41936 : node41933;
															assign node41933 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node41936 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node41939 = (inp[6]) ? node41943 : node41940;
															assign node41940 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node41943 = (inp[1]) ? 4'b0110 : 4'b0110;
													assign node41946 = (inp[1]) ? node41954 : node41947;
														assign node41947 = (inp[5]) ? node41951 : node41948;
															assign node41948 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node41951 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node41954 = (inp[11]) ? node41958 : node41955;
															assign node41955 = (inp[6]) ? 4'b1110 : 4'b0110;
															assign node41958 = (inp[6]) ? 4'b0110 : 4'b1110;
											assign node41961 = (inp[15]) ? node41991 : node41962;
												assign node41962 = (inp[5]) ? node41976 : node41963;
													assign node41963 = (inp[3]) ? node41969 : node41964;
														assign node41964 = (inp[6]) ? node41966 : 4'b0100;
															assign node41966 = (inp[1]) ? 4'b0100 : 4'b0100;
														assign node41969 = (inp[1]) ? node41973 : node41970;
															assign node41970 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node41973 = (inp[6]) ? 4'b1110 : 4'b0110;
													assign node41976 = (inp[1]) ? node41984 : node41977;
														assign node41977 = (inp[6]) ? node41981 : node41978;
															assign node41978 = (inp[11]) ? 4'b0110 : 4'b1110;
															assign node41981 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node41984 = (inp[3]) ? node41988 : node41985;
															assign node41985 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node41988 = (inp[6]) ? 4'b0110 : 4'b0110;
												assign node41991 = (inp[3]) ? node42005 : node41992;
													assign node41992 = (inp[5]) ? node42000 : node41993;
														assign node41993 = (inp[6]) ? node41997 : node41994;
															assign node41994 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node41997 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node42000 = (inp[6]) ? 4'b0100 : node42001;
															assign node42001 = (inp[1]) ? 4'b1100 : 4'b0100;
													assign node42005 = (inp[1]) ? node42013 : node42006;
														assign node42006 = (inp[11]) ? node42010 : node42007;
															assign node42007 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node42010 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node42013 = (inp[11]) ? node42017 : node42014;
															assign node42014 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node42017 = (inp[6]) ? 4'b0100 : 4'b1100;
										assign node42020 = (inp[0]) ? node42076 : node42021;
											assign node42021 = (inp[15]) ? node42053 : node42022;
												assign node42022 = (inp[5]) ? node42038 : node42023;
													assign node42023 = (inp[3]) ? node42031 : node42024;
														assign node42024 = (inp[1]) ? node42028 : node42025;
															assign node42025 = (inp[11]) ? 4'b0110 : 4'b1110;
															assign node42028 = (inp[6]) ? 4'b0110 : 4'b0110;
														assign node42031 = (inp[6]) ? node42035 : node42032;
															assign node42032 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node42035 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node42038 = (inp[3]) ? node42046 : node42039;
														assign node42039 = (inp[6]) ? node42043 : node42040;
															assign node42040 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node42043 = (inp[11]) ? 4'b0100 : 4'b1100;
														assign node42046 = (inp[11]) ? node42050 : node42047;
															assign node42047 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node42050 = (inp[6]) ? 4'b0100 : 4'b1100;
												assign node42053 = (inp[3]) ? node42069 : node42054;
													assign node42054 = (inp[5]) ? node42062 : node42055;
														assign node42055 = (inp[6]) ? node42059 : node42056;
															assign node42056 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node42059 = (inp[11]) ? 4'b0100 : 4'b1100;
														assign node42062 = (inp[1]) ? node42066 : node42063;
															assign node42063 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node42066 = (inp[11]) ? 4'b0110 : 4'b0110;
													assign node42069 = (inp[11]) ? node42073 : node42070;
														assign node42070 = (inp[6]) ? 4'b1110 : 4'b0110;
														assign node42073 = (inp[6]) ? 4'b0110 : 4'b1110;
											assign node42076 = (inp[15]) ? node42106 : node42077;
												assign node42077 = (inp[5]) ? node42091 : node42078;
													assign node42078 = (inp[3]) ? node42086 : node42079;
														assign node42079 = (inp[1]) ? node42083 : node42080;
															assign node42080 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node42083 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node42086 = (inp[1]) ? node42088 : 4'b1110;
															assign node42088 = (inp[11]) ? 4'b0110 : 4'b0110;
													assign node42091 = (inp[3]) ? node42099 : node42092;
														assign node42092 = (inp[11]) ? node42096 : node42093;
															assign node42093 = (inp[6]) ? 4'b1110 : 4'b0110;
															assign node42096 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node42099 = (inp[6]) ? node42103 : node42100;
															assign node42100 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node42103 = (inp[11]) ? 4'b0110 : 4'b1110;
												assign node42106 = (inp[5]) ? node42122 : node42107;
													assign node42107 = (inp[3]) ? node42115 : node42108;
														assign node42108 = (inp[1]) ? node42112 : node42109;
															assign node42109 = (inp[11]) ? 4'b0110 : 4'b1110;
															assign node42112 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node42115 = (inp[11]) ? node42119 : node42116;
															assign node42116 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node42119 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node42122 = (inp[6]) ? node42126 : node42123;
														assign node42123 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node42126 = (inp[11]) ? 4'b0100 : 4'b1100;
							assign node42129 = (inp[0]) ? node42619 : node42130;
								assign node42130 = (inp[15]) ? node42380 : node42131;
									assign node42131 = (inp[3]) ? node42257 : node42132;
										assign node42132 = (inp[5]) ? node42196 : node42133;
											assign node42133 = (inp[11]) ? node42165 : node42134;
												assign node42134 = (inp[6]) ? node42150 : node42135;
													assign node42135 = (inp[1]) ? node42143 : node42136;
														assign node42136 = (inp[13]) ? node42140 : node42137;
															assign node42137 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node42140 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node42143 = (inp[13]) ? node42147 : node42144;
															assign node42144 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node42147 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node42150 = (inp[13]) ? node42158 : node42151;
														assign node42151 = (inp[1]) ? node42155 : node42152;
															assign node42152 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node42155 = (inp[8]) ? 4'b1111 : 4'b0110;
														assign node42158 = (inp[1]) ? node42162 : node42159;
															assign node42159 = (inp[8]) ? 4'b1111 : 4'b0110;
															assign node42162 = (inp[8]) ? 4'b1110 : 4'b1110;
												assign node42165 = (inp[6]) ? node42181 : node42166;
													assign node42166 = (inp[13]) ? node42174 : node42167;
														assign node42167 = (inp[1]) ? node42171 : node42168;
															assign node42168 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node42171 = (inp[7]) ? 4'b1111 : 4'b0110;
														assign node42174 = (inp[1]) ? node42178 : node42175;
															assign node42175 = (inp[8]) ? 4'b1111 : 4'b0110;
															assign node42178 = (inp[7]) ? 4'b1110 : 4'b1110;
													assign node42181 = (inp[1]) ? node42189 : node42182;
														assign node42182 = (inp[13]) ? node42186 : node42183;
															assign node42183 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node42186 = (inp[7]) ? 4'b0110 : 4'b1110;
														assign node42189 = (inp[8]) ? node42193 : node42190;
															assign node42190 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node42193 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node42196 = (inp[11]) ? node42228 : node42197;
												assign node42197 = (inp[6]) ? node42213 : node42198;
													assign node42198 = (inp[1]) ? node42206 : node42199;
														assign node42199 = (inp[13]) ? node42203 : node42200;
															assign node42200 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node42203 = (inp[8]) ? 4'b0100 : 4'b1100;
														assign node42206 = (inp[7]) ? node42210 : node42207;
															assign node42207 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node42210 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node42213 = (inp[13]) ? node42221 : node42214;
														assign node42214 = (inp[1]) ? node42218 : node42215;
															assign node42215 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node42218 = (inp[8]) ? 4'b1100 : 4'b0100;
														assign node42221 = (inp[1]) ? node42225 : node42222;
															assign node42222 = (inp[8]) ? 4'b1100 : 4'b0100;
															assign node42225 = (inp[8]) ? 4'b1100 : 4'b1100;
												assign node42228 = (inp[6]) ? node42242 : node42229;
													assign node42229 = (inp[13]) ? node42235 : node42230;
														assign node42230 = (inp[1]) ? node42232 : 4'b0101;
															assign node42232 = (inp[7]) ? 4'b1100 : 4'b0100;
														assign node42235 = (inp[7]) ? node42239 : node42236;
															assign node42236 = (inp[8]) ? 4'b1101 : 4'b0100;
															assign node42239 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node42242 = (inp[1]) ? node42250 : node42243;
														assign node42243 = (inp[13]) ? node42247 : node42244;
															assign node42244 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node42247 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node42250 = (inp[13]) ? node42254 : node42251;
															assign node42251 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node42254 = (inp[8]) ? 4'b0101 : 4'b0100;
										assign node42257 = (inp[5]) ? node42319 : node42258;
											assign node42258 = (inp[8]) ? node42290 : node42259;
												assign node42259 = (inp[7]) ? node42275 : node42260;
													assign node42260 = (inp[13]) ? node42268 : node42261;
														assign node42261 = (inp[6]) ? node42265 : node42262;
															assign node42262 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node42265 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node42268 = (inp[11]) ? node42272 : node42269;
															assign node42269 = (inp[1]) ? 4'b0100 : 4'b0100;
															assign node42272 = (inp[6]) ? 4'b0100 : 4'b0100;
													assign node42275 = (inp[11]) ? node42283 : node42276;
														assign node42276 = (inp[6]) ? node42280 : node42277;
															assign node42277 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node42280 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node42283 = (inp[6]) ? node42287 : node42284;
															assign node42284 = (inp[13]) ? 4'b1101 : 4'b0101;
															assign node42287 = (inp[13]) ? 4'b0101 : 4'b0101;
												assign node42290 = (inp[7]) ? node42306 : node42291;
													assign node42291 = (inp[1]) ? node42299 : node42292;
														assign node42292 = (inp[6]) ? node42296 : node42293;
															assign node42293 = (inp[13]) ? 4'b0101 : 4'b0101;
															assign node42296 = (inp[11]) ? 4'b0101 : 4'b0101;
														assign node42299 = (inp[6]) ? node42303 : node42300;
															assign node42300 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node42303 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node42306 = (inp[6]) ? node42314 : node42307;
														assign node42307 = (inp[11]) ? node42311 : node42308;
															assign node42308 = (inp[13]) ? 4'b0100 : 4'b0100;
															assign node42311 = (inp[1]) ? 4'b1100 : 4'b0100;
														assign node42314 = (inp[11]) ? node42316 : 4'b1100;
															assign node42316 = (inp[1]) ? 4'b0100 : 4'b1100;
											assign node42319 = (inp[13]) ? node42349 : node42320;
												assign node42320 = (inp[7]) ? node42334 : node42321;
													assign node42321 = (inp[8]) ? node42327 : node42322;
														assign node42322 = (inp[1]) ? node42324 : 4'b1100;
															assign node42324 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node42327 = (inp[6]) ? node42331 : node42328;
															assign node42328 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node42331 = (inp[1]) ? 4'b0101 : 4'b0101;
													assign node42334 = (inp[8]) ? node42342 : node42335;
														assign node42335 = (inp[1]) ? node42339 : node42336;
															assign node42336 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node42339 = (inp[6]) ? 4'b0101 : 4'b0101;
														assign node42342 = (inp[1]) ? node42346 : node42343;
															assign node42343 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node42346 = (inp[11]) ? 4'b0100 : 4'b0100;
												assign node42349 = (inp[1]) ? node42365 : node42350;
													assign node42350 = (inp[11]) ? node42358 : node42351;
														assign node42351 = (inp[6]) ? node42355 : node42352;
															assign node42352 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node42355 = (inp[7]) ? 4'b1101 : 4'b0100;
														assign node42358 = (inp[6]) ? node42362 : node42359;
															assign node42359 = (inp[7]) ? 4'b1100 : 4'b0100;
															assign node42362 = (inp[7]) ? 4'b0100 : 4'b1100;
													assign node42365 = (inp[8]) ? node42373 : node42366;
														assign node42366 = (inp[7]) ? node42370 : node42367;
															assign node42367 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node42370 = (inp[11]) ? 4'b0101 : 4'b0101;
														assign node42373 = (inp[7]) ? node42377 : node42374;
															assign node42374 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node42377 = (inp[6]) ? 4'b1100 : 4'b0100;
									assign node42380 = (inp[5]) ? node42504 : node42381;
										assign node42381 = (inp[3]) ? node42441 : node42382;
											assign node42382 = (inp[1]) ? node42412 : node42383;
												assign node42383 = (inp[7]) ? node42397 : node42384;
													assign node42384 = (inp[8]) ? node42392 : node42385;
														assign node42385 = (inp[13]) ? node42389 : node42386;
															assign node42386 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node42389 = (inp[6]) ? 4'b0100 : 4'b0100;
														assign node42392 = (inp[13]) ? 4'b0101 : node42393;
															assign node42393 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node42397 = (inp[8]) ? node42405 : node42398;
														assign node42398 = (inp[11]) ? node42402 : node42399;
															assign node42399 = (inp[6]) ? 4'b0101 : 4'b0101;
															assign node42402 = (inp[13]) ? 4'b1101 : 4'b0101;
														assign node42405 = (inp[13]) ? node42409 : node42406;
															assign node42406 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node42409 = (inp[6]) ? 4'b0100 : 4'b1100;
												assign node42412 = (inp[6]) ? node42428 : node42413;
													assign node42413 = (inp[11]) ? node42421 : node42414;
														assign node42414 = (inp[13]) ? node42418 : node42415;
															assign node42415 = (inp[7]) ? 4'b0100 : 4'b1100;
															assign node42418 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node42421 = (inp[8]) ? node42425 : node42422;
															assign node42422 = (inp[7]) ? 4'b1101 : 4'b0100;
															assign node42425 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node42428 = (inp[11]) ? node42434 : node42429;
														assign node42429 = (inp[8]) ? 4'b1101 : node42430;
															assign node42430 = (inp[7]) ? 4'b1101 : 4'b0100;
														assign node42434 = (inp[13]) ? node42438 : node42435;
															assign node42435 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node42438 = (inp[8]) ? 4'b0100 : 4'b0100;
											assign node42441 = (inp[11]) ? node42473 : node42442;
												assign node42442 = (inp[6]) ? node42458 : node42443;
													assign node42443 = (inp[1]) ? node42451 : node42444;
														assign node42444 = (inp[13]) ? node42448 : node42445;
															assign node42445 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node42448 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node42451 = (inp[13]) ? node42455 : node42452;
															assign node42452 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node42455 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node42458 = (inp[1]) ? node42466 : node42459;
														assign node42459 = (inp[13]) ? node42463 : node42460;
															assign node42460 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node42463 = (inp[7]) ? 4'b1110 : 4'b0110;
														assign node42466 = (inp[13]) ? node42470 : node42467;
															assign node42467 = (inp[8]) ? 4'b1111 : 4'b0110;
															assign node42470 = (inp[8]) ? 4'b1110 : 4'b1110;
												assign node42473 = (inp[6]) ? node42489 : node42474;
													assign node42474 = (inp[1]) ? node42482 : node42475;
														assign node42475 = (inp[13]) ? node42479 : node42476;
															assign node42476 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node42479 = (inp[7]) ? 4'b1110 : 4'b0110;
														assign node42482 = (inp[8]) ? node42486 : node42483;
															assign node42483 = (inp[7]) ? 4'b1111 : 4'b0110;
															assign node42486 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node42489 = (inp[1]) ? node42497 : node42490;
														assign node42490 = (inp[13]) ? node42494 : node42491;
															assign node42491 = (inp[7]) ? 4'b1110 : 4'b1110;
															assign node42494 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node42497 = (inp[7]) ? node42501 : node42498;
															assign node42498 = (inp[8]) ? 4'b0111 : 4'b1110;
															assign node42501 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node42504 = (inp[1]) ? node42566 : node42505;
											assign node42505 = (inp[3]) ? node42535 : node42506;
												assign node42506 = (inp[8]) ? node42520 : node42507;
													assign node42507 = (inp[7]) ? node42513 : node42508;
														assign node42508 = (inp[11]) ? node42510 : 4'b0110;
															assign node42510 = (inp[6]) ? 4'b1110 : 4'b0110;
														assign node42513 = (inp[13]) ? node42517 : node42514;
															assign node42514 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node42517 = (inp[11]) ? 4'b0111 : 4'b0111;
													assign node42520 = (inp[7]) ? node42528 : node42521;
														assign node42521 = (inp[6]) ? node42525 : node42522;
															assign node42522 = (inp[13]) ? 4'b0111 : 4'b0111;
															assign node42525 = (inp[13]) ? 4'b0111 : 4'b0111;
														assign node42528 = (inp[11]) ? node42532 : node42529;
															assign node42529 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node42532 = (inp[13]) ? 4'b0110 : 4'b0110;
												assign node42535 = (inp[13]) ? node42551 : node42536;
													assign node42536 = (inp[6]) ? node42544 : node42537;
														assign node42537 = (inp[11]) ? node42541 : node42538;
															assign node42538 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node42541 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node42544 = (inp[11]) ? node42548 : node42545;
															assign node42545 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node42548 = (inp[8]) ? 4'b1110 : 4'b1110;
													assign node42551 = (inp[6]) ? node42559 : node42552;
														assign node42552 = (inp[11]) ? node42556 : node42553;
															assign node42553 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node42556 = (inp[7]) ? 4'b1110 : 4'b0110;
														assign node42559 = (inp[11]) ? node42563 : node42560;
															assign node42560 = (inp[7]) ? 4'b1111 : 4'b0110;
															assign node42563 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node42566 = (inp[8]) ? node42588 : node42567;
												assign node42567 = (inp[7]) ? node42581 : node42568;
													assign node42568 = (inp[11]) ? node42574 : node42569;
														assign node42569 = (inp[3]) ? 4'b1110 : node42570;
															assign node42570 = (inp[6]) ? 4'b0110 : 4'b0110;
														assign node42574 = (inp[3]) ? node42578 : node42575;
															assign node42575 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node42578 = (inp[6]) ? 4'b0110 : 4'b0110;
													assign node42581 = (inp[6]) ? node42585 : node42582;
														assign node42582 = (inp[11]) ? 4'b1111 : 4'b0111;
														assign node42585 = (inp[11]) ? 4'b0111 : 4'b1111;
												assign node42588 = (inp[7]) ? node42604 : node42589;
													assign node42589 = (inp[13]) ? node42597 : node42590;
														assign node42590 = (inp[11]) ? node42594 : node42591;
															assign node42591 = (inp[6]) ? 4'b1111 : 4'b0111;
															assign node42594 = (inp[6]) ? 4'b0111 : 4'b1111;
														assign node42597 = (inp[11]) ? node42601 : node42598;
															assign node42598 = (inp[6]) ? 4'b1111 : 4'b0111;
															assign node42601 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node42604 = (inp[13]) ? node42612 : node42605;
														assign node42605 = (inp[6]) ? node42609 : node42606;
															assign node42606 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node42609 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node42612 = (inp[3]) ? node42616 : node42613;
															assign node42613 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node42616 = (inp[11]) ? 4'b0110 : 4'b0110;
								assign node42619 = (inp[15]) ? node42843 : node42620;
									assign node42620 = (inp[5]) ? node42742 : node42621;
										assign node42621 = (inp[3]) ? node42681 : node42622;
											assign node42622 = (inp[13]) ? node42652 : node42623;
												assign node42623 = (inp[8]) ? node42639 : node42624;
													assign node42624 = (inp[7]) ? node42632 : node42625;
														assign node42625 = (inp[1]) ? node42629 : node42626;
															assign node42626 = (inp[6]) ? 4'b0100 : 4'b0100;
															assign node42629 = (inp[11]) ? 4'b0100 : 4'b0100;
														assign node42632 = (inp[6]) ? node42636 : node42633;
															assign node42633 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node42636 = (inp[1]) ? 4'b0101 : 4'b0101;
													assign node42639 = (inp[7]) ? node42647 : node42640;
														assign node42640 = (inp[6]) ? node42644 : node42641;
															assign node42641 = (inp[11]) ? 4'b0101 : 4'b0101;
															assign node42644 = (inp[11]) ? 4'b0101 : 4'b0101;
														assign node42647 = (inp[11]) ? node42649 : 4'b0100;
															assign node42649 = (inp[1]) ? 4'b0100 : 4'b0100;
												assign node42652 = (inp[8]) ? node42666 : node42653;
													assign node42653 = (inp[7]) ? node42659 : node42654;
														assign node42654 = (inp[1]) ? node42656 : 4'b1100;
															assign node42656 = (inp[6]) ? 4'b0100 : 4'b0100;
														assign node42659 = (inp[11]) ? node42663 : node42660;
															assign node42660 = (inp[6]) ? 4'b1101 : 4'b0101;
															assign node42663 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node42666 = (inp[7]) ? node42674 : node42667;
														assign node42667 = (inp[11]) ? node42671 : node42668;
															assign node42668 = (inp[6]) ? 4'b1101 : 4'b0101;
															assign node42671 = (inp[6]) ? 4'b0101 : 4'b1101;
														assign node42674 = (inp[6]) ? node42678 : node42675;
															assign node42675 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node42678 = (inp[11]) ? 4'b0100 : 4'b1100;
											assign node42681 = (inp[1]) ? node42711 : node42682;
												assign node42682 = (inp[13]) ? node42698 : node42683;
													assign node42683 = (inp[7]) ? node42691 : node42684;
														assign node42684 = (inp[8]) ? node42688 : node42685;
															assign node42685 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node42688 = (inp[11]) ? 4'b0111 : 4'b0111;
														assign node42691 = (inp[8]) ? node42695 : node42692;
															assign node42692 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node42695 = (inp[11]) ? 4'b0110 : 4'b0110;
													assign node42698 = (inp[11]) ? node42706 : node42699;
														assign node42699 = (inp[6]) ? node42703 : node42700;
															assign node42700 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node42703 = (inp[8]) ? 4'b1110 : 4'b0110;
														assign node42706 = (inp[6]) ? 4'b0111 : node42707;
															assign node42707 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node42711 = (inp[13]) ? node42727 : node42712;
													assign node42712 = (inp[8]) ? node42720 : node42713;
														assign node42713 = (inp[7]) ? node42717 : node42714;
															assign node42714 = (inp[6]) ? 4'b0110 : 4'b0110;
															assign node42717 = (inp[6]) ? 4'b0111 : 4'b0111;
														assign node42720 = (inp[7]) ? node42724 : node42721;
															assign node42721 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node42724 = (inp[11]) ? 4'b0110 : 4'b0110;
													assign node42727 = (inp[11]) ? node42735 : node42728;
														assign node42728 = (inp[6]) ? node42732 : node42729;
															assign node42729 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node42732 = (inp[7]) ? 4'b1110 : 4'b1110;
														assign node42735 = (inp[6]) ? node42739 : node42736;
															assign node42736 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node42739 = (inp[7]) ? 4'b0110 : 4'b0110;
										assign node42742 = (inp[7]) ? node42796 : node42743;
											assign node42743 = (inp[8]) ? node42767 : node42744;
												assign node42744 = (inp[6]) ? node42756 : node42745;
													assign node42745 = (inp[11]) ? node42751 : node42746;
														assign node42746 = (inp[1]) ? node42748 : 4'b1110;
															assign node42748 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node42751 = (inp[1]) ? node42753 : 4'b0110;
															assign node42753 = (inp[13]) ? 4'b1110 : 4'b0110;
													assign node42756 = (inp[11]) ? node42762 : node42757;
														assign node42757 = (inp[1]) ? node42759 : 4'b0110;
															assign node42759 = (inp[13]) ? 4'b1110 : 4'b0110;
														assign node42762 = (inp[1]) ? node42764 : 4'b1110;
															assign node42764 = (inp[13]) ? 4'b0110 : 4'b1110;
												assign node42767 = (inp[3]) ? node42783 : node42768;
													assign node42768 = (inp[13]) ? node42776 : node42769;
														assign node42769 = (inp[11]) ? node42773 : node42770;
															assign node42770 = (inp[1]) ? 4'b0111 : 4'b0111;
															assign node42773 = (inp[1]) ? 4'b0111 : 4'b0111;
														assign node42776 = (inp[1]) ? node42780 : node42777;
															assign node42777 = (inp[11]) ? 4'b0111 : 4'b0111;
															assign node42780 = (inp[11]) ? 4'b1111 : 4'b0111;
													assign node42783 = (inp[6]) ? node42789 : node42784;
														assign node42784 = (inp[11]) ? 4'b1111 : node42785;
															assign node42785 = (inp[13]) ? 4'b0111 : 4'b0111;
														assign node42789 = (inp[11]) ? node42793 : node42790;
															assign node42790 = (inp[1]) ? 4'b1111 : 4'b0111;
															assign node42793 = (inp[1]) ? 4'b0111 : 4'b0111;
											assign node42796 = (inp[8]) ? node42820 : node42797;
												assign node42797 = (inp[6]) ? node42809 : node42798;
													assign node42798 = (inp[11]) ? node42804 : node42799;
														assign node42799 = (inp[13]) ? 4'b0111 : node42800;
															assign node42800 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node42804 = (inp[1]) ? 4'b1111 : node42805;
															assign node42805 = (inp[13]) ? 4'b1111 : 4'b0111;
													assign node42809 = (inp[11]) ? node42815 : node42810;
														assign node42810 = (inp[13]) ? 4'b1111 : node42811;
															assign node42811 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node42815 = (inp[13]) ? 4'b0111 : node42816;
															assign node42816 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node42820 = (inp[11]) ? node42832 : node42821;
													assign node42821 = (inp[6]) ? node42827 : node42822;
														assign node42822 = (inp[1]) ? 4'b0110 : node42823;
															assign node42823 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node42827 = (inp[13]) ? 4'b1110 : node42828;
															assign node42828 = (inp[1]) ? 4'b1110 : 4'b0110;
													assign node42832 = (inp[6]) ? node42838 : node42833;
														assign node42833 = (inp[13]) ? 4'b1110 : node42834;
															assign node42834 = (inp[1]) ? 4'b1110 : 4'b0110;
														assign node42838 = (inp[13]) ? 4'b0110 : node42839;
															assign node42839 = (inp[1]) ? 4'b0110 : 4'b1110;
									assign node42843 = (inp[5]) ? node42967 : node42844;
										assign node42844 = (inp[3]) ? node42908 : node42845;
											assign node42845 = (inp[1]) ? node42877 : node42846;
												assign node42846 = (inp[6]) ? node42862 : node42847;
													assign node42847 = (inp[11]) ? node42855 : node42848;
														assign node42848 = (inp[13]) ? node42852 : node42849;
															assign node42849 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node42852 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node42855 = (inp[8]) ? node42859 : node42856;
															assign node42856 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node42859 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node42862 = (inp[11]) ? node42870 : node42863;
														assign node42863 = (inp[13]) ? node42867 : node42864;
															assign node42864 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node42867 = (inp[8]) ? 4'b1110 : 4'b0110;
														assign node42870 = (inp[13]) ? node42874 : node42871;
															assign node42871 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node42874 = (inp[7]) ? 4'b0110 : 4'b1110;
												assign node42877 = (inp[8]) ? node42893 : node42878;
													assign node42878 = (inp[7]) ? node42886 : node42879;
														assign node42879 = (inp[6]) ? node42883 : node42880;
															assign node42880 = (inp[13]) ? 4'b0110 : 4'b0110;
															assign node42883 = (inp[13]) ? 4'b1110 : 4'b0110;
														assign node42886 = (inp[13]) ? node42890 : node42887;
															assign node42887 = (inp[6]) ? 4'b0111 : 4'b0111;
															assign node42890 = (inp[6]) ? 4'b0111 : 4'b0111;
													assign node42893 = (inp[7]) ? node42901 : node42894;
														assign node42894 = (inp[6]) ? node42898 : node42895;
															assign node42895 = (inp[11]) ? 4'b1111 : 4'b0111;
															assign node42898 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node42901 = (inp[13]) ? node42905 : node42902;
															assign node42902 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node42905 = (inp[6]) ? 4'b0110 : 4'b0110;
											assign node42908 = (inp[6]) ? node42938 : node42909;
												assign node42909 = (inp[11]) ? node42923 : node42910;
													assign node42910 = (inp[1]) ? node42918 : node42911;
														assign node42911 = (inp[13]) ? node42915 : node42912;
															assign node42912 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node42915 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node42918 = (inp[8]) ? node42920 : 4'b0101;
															assign node42920 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node42923 = (inp[1]) ? node42931 : node42924;
														assign node42924 = (inp[13]) ? node42928 : node42925;
															assign node42925 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node42928 = (inp[8]) ? 4'b1100 : 4'b0100;
														assign node42931 = (inp[13]) ? node42935 : node42932;
															assign node42932 = (inp[7]) ? 4'b1100 : 4'b0100;
															assign node42935 = (inp[7]) ? 4'b1100 : 4'b1100;
												assign node42938 = (inp[11]) ? node42952 : node42939;
													assign node42939 = (inp[13]) ? node42947 : node42940;
														assign node42940 = (inp[7]) ? node42944 : node42941;
															assign node42941 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node42944 = (inp[1]) ? 4'b1100 : 4'b0100;
														assign node42947 = (inp[7]) ? node42949 : 4'b1101;
															assign node42949 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node42952 = (inp[13]) ? node42960 : node42953;
														assign node42953 = (inp[1]) ? node42957 : node42954;
															assign node42954 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node42957 = (inp[7]) ? 4'b0100 : 4'b1100;
														assign node42960 = (inp[8]) ? node42964 : node42961;
															assign node42961 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node42964 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node42967 = (inp[7]) ? node43011 : node42968;
											assign node42968 = (inp[8]) ? node42990 : node42969;
												assign node42969 = (inp[6]) ? node42981 : node42970;
													assign node42970 = (inp[11]) ? node42976 : node42971;
														assign node42971 = (inp[1]) ? node42973 : 4'b1100;
															assign node42973 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node42976 = (inp[13]) ? node42978 : 4'b0100;
															assign node42978 = (inp[1]) ? 4'b1100 : 4'b0100;
													assign node42981 = (inp[11]) ? node42985 : node42982;
														assign node42982 = (inp[1]) ? 4'b1100 : 4'b0100;
														assign node42985 = (inp[13]) ? node42987 : 4'b1100;
															assign node42987 = (inp[1]) ? 4'b0100 : 4'b1100;
												assign node42990 = (inp[6]) ? node43000 : node42991;
													assign node42991 = (inp[11]) ? node42995 : node42992;
														assign node42992 = (inp[13]) ? 4'b0101 : 4'b1101;
														assign node42995 = (inp[13]) ? 4'b1101 : node42996;
															assign node42996 = (inp[1]) ? 4'b1101 : 4'b0101;
													assign node43000 = (inp[11]) ? node43006 : node43001;
														assign node43001 = (inp[13]) ? 4'b1101 : node43002;
															assign node43002 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node43006 = (inp[1]) ? 4'b0101 : node43007;
															assign node43007 = (inp[13]) ? 4'b0101 : 4'b1101;
											assign node43011 = (inp[8]) ? node43043 : node43012;
												assign node43012 = (inp[3]) ? node43028 : node43013;
													assign node43013 = (inp[6]) ? node43021 : node43014;
														assign node43014 = (inp[11]) ? node43018 : node43015;
															assign node43015 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node43018 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node43021 = (inp[11]) ? node43025 : node43022;
															assign node43022 = (inp[1]) ? 4'b1101 : 4'b0101;
															assign node43025 = (inp[13]) ? 4'b0101 : 4'b0101;
													assign node43028 = (inp[11]) ? node43036 : node43029;
														assign node43029 = (inp[6]) ? node43033 : node43030;
															assign node43030 = (inp[1]) ? 4'b0101 : 4'b0101;
															assign node43033 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node43036 = (inp[6]) ? node43040 : node43037;
															assign node43037 = (inp[1]) ? 4'b1101 : 4'b0101;
															assign node43040 = (inp[13]) ? 4'b0101 : 4'b0101;
												assign node43043 = (inp[6]) ? node43055 : node43044;
													assign node43044 = (inp[11]) ? node43050 : node43045;
														assign node43045 = (inp[13]) ? 4'b0100 : node43046;
															assign node43046 = (inp[1]) ? 4'b0100 : 4'b1100;
														assign node43050 = (inp[1]) ? 4'b1100 : node43051;
															assign node43051 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node43055 = (inp[11]) ? node43061 : node43056;
														assign node43056 = (inp[1]) ? 4'b1100 : node43057;
															assign node43057 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node43061 = (inp[1]) ? 4'b0100 : node43062;
															assign node43062 = (inp[13]) ? 4'b0100 : 4'b1100;
			assign node43066 = (inp[10]) ? node50268 : node43067;
				assign node43067 = (inp[12]) ? node46691 : node43068;
					assign node43068 = (inp[6]) ? node44850 : node43069;
						assign node43069 = (inp[11]) ? node43951 : node43070;
							assign node43070 = (inp[1]) ? node43500 : node43071;
								assign node43071 = (inp[13]) ? node43279 : node43072;
									assign node43072 = (inp[15]) ? node43178 : node43073;
										assign node43073 = (inp[0]) ? node43123 : node43074;
											assign node43074 = (inp[3]) ? node43102 : node43075;
												assign node43075 = (inp[5]) ? node43089 : node43076;
													assign node43076 = (inp[2]) ? node43084 : node43077;
														assign node43077 = (inp[8]) ? node43081 : node43078;
															assign node43078 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node43081 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node43084 = (inp[14]) ? node43086 : 4'b1110;
															assign node43086 = (inp[7]) ? 4'b1110 : 4'b1110;
													assign node43089 = (inp[2]) ? node43095 : node43090;
														assign node43090 = (inp[14]) ? 4'b1101 : node43091;
															assign node43091 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node43095 = (inp[8]) ? node43099 : node43096;
															assign node43096 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node43099 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node43102 = (inp[2]) ? node43116 : node43103;
													assign node43103 = (inp[7]) ? node43109 : node43104;
														assign node43104 = (inp[5]) ? 4'b1100 : node43105;
															assign node43105 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node43109 = (inp[14]) ? node43113 : node43110;
															assign node43110 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node43113 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node43116 = (inp[8]) ? node43120 : node43117;
														assign node43117 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node43120 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node43123 = (inp[3]) ? node43155 : node43124;
												assign node43124 = (inp[5]) ? node43140 : node43125;
													assign node43125 = (inp[8]) ? node43133 : node43126;
														assign node43126 = (inp[7]) ? node43130 : node43127;
															assign node43127 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node43130 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node43133 = (inp[7]) ? node43137 : node43134;
															assign node43134 = (inp[14]) ? 4'b1101 : 4'b1100;
															assign node43137 = (inp[14]) ? 4'b1100 : 4'b1100;
													assign node43140 = (inp[8]) ? node43148 : node43141;
														assign node43141 = (inp[7]) ? node43145 : node43142;
															assign node43142 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node43145 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node43148 = (inp[7]) ? node43152 : node43149;
															assign node43149 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node43152 = (inp[2]) ? 4'b1110 : 4'b1110;
												assign node43155 = (inp[8]) ? node43167 : node43156;
													assign node43156 = (inp[7]) ? node43162 : node43157;
														assign node43157 = (inp[14]) ? 4'b1110 : node43158;
															assign node43158 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node43162 = (inp[14]) ? 4'b1111 : node43163;
															assign node43163 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node43167 = (inp[7]) ? node43173 : node43168;
														assign node43168 = (inp[14]) ? 4'b1111 : node43169;
															assign node43169 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node43173 = (inp[2]) ? 4'b1110 : node43174;
															assign node43174 = (inp[14]) ? 4'b1110 : 4'b1111;
										assign node43178 = (inp[0]) ? node43226 : node43179;
											assign node43179 = (inp[3]) ? node43207 : node43180;
												assign node43180 = (inp[5]) ? node43194 : node43181;
													assign node43181 = (inp[14]) ? node43187 : node43182;
														assign node43182 = (inp[7]) ? 4'b1101 : node43183;
															assign node43183 = (inp[2]) ? 4'b1100 : 4'b1100;
														assign node43187 = (inp[7]) ? node43191 : node43188;
															assign node43188 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node43191 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node43194 = (inp[7]) ? node43200 : node43195;
														assign node43195 = (inp[14]) ? node43197 : 4'b1110;
															assign node43197 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node43200 = (inp[8]) ? node43204 : node43201;
															assign node43201 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node43204 = (inp[2]) ? 4'b1110 : 4'b1110;
												assign node43207 = (inp[8]) ? node43215 : node43208;
													assign node43208 = (inp[7]) ? 4'b1111 : node43209;
														assign node43209 = (inp[2]) ? 4'b1110 : node43210;
															assign node43210 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node43215 = (inp[7]) ? node43221 : node43216;
														assign node43216 = (inp[2]) ? 4'b1111 : node43217;
															assign node43217 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node43221 = (inp[14]) ? 4'b1110 : node43222;
															assign node43222 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node43226 = (inp[3]) ? node43256 : node43227;
												assign node43227 = (inp[5]) ? node43241 : node43228;
													assign node43228 = (inp[7]) ? node43234 : node43229;
														assign node43229 = (inp[2]) ? node43231 : 4'b1110;
															assign node43231 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node43234 = (inp[8]) ? node43238 : node43235;
															assign node43235 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node43238 = (inp[2]) ? 4'b1110 : 4'b1110;
													assign node43241 = (inp[2]) ? node43249 : node43242;
														assign node43242 = (inp[7]) ? node43246 : node43243;
															assign node43243 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node43246 = (inp[14]) ? 4'b1100 : 4'b1100;
														assign node43249 = (inp[8]) ? node43253 : node43250;
															assign node43250 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node43253 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node43256 = (inp[14]) ? node43272 : node43257;
													assign node43257 = (inp[8]) ? node43265 : node43258;
														assign node43258 = (inp[2]) ? node43262 : node43259;
															assign node43259 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node43262 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node43265 = (inp[5]) ? node43269 : node43266;
															assign node43266 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node43269 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node43272 = (inp[8]) ? node43276 : node43273;
														assign node43273 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node43276 = (inp[7]) ? 4'b1100 : 4'b1101;
									assign node43279 = (inp[8]) ? node43395 : node43280;
										assign node43280 = (inp[7]) ? node43342 : node43281;
											assign node43281 = (inp[2]) ? node43311 : node43282;
												assign node43282 = (inp[14]) ? node43298 : node43283;
													assign node43283 = (inp[5]) ? node43291 : node43284;
														assign node43284 = (inp[3]) ? node43288 : node43285;
															assign node43285 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node43288 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node43291 = (inp[3]) ? node43295 : node43292;
															assign node43292 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node43295 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node43298 = (inp[15]) ? node43306 : node43299;
														assign node43299 = (inp[0]) ? node43303 : node43300;
															assign node43300 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node43303 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node43306 = (inp[0]) ? node43308 : 4'b1110;
															assign node43308 = (inp[3]) ? 4'b1100 : 4'b1100;
												assign node43311 = (inp[14]) ? node43327 : node43312;
													assign node43312 = (inp[5]) ? node43320 : node43313;
														assign node43313 = (inp[0]) ? node43317 : node43314;
															assign node43314 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node43317 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node43320 = (inp[0]) ? node43324 : node43321;
															assign node43321 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node43324 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node43327 = (inp[3]) ? node43335 : node43328;
														assign node43328 = (inp[0]) ? node43332 : node43329;
															assign node43329 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node43332 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node43335 = (inp[15]) ? node43339 : node43336;
															assign node43336 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node43339 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node43342 = (inp[2]) ? node43372 : node43343;
												assign node43343 = (inp[14]) ? node43359 : node43344;
													assign node43344 = (inp[5]) ? node43352 : node43345;
														assign node43345 = (inp[3]) ? node43349 : node43346;
															assign node43346 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node43349 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node43352 = (inp[0]) ? node43356 : node43353;
															assign node43353 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node43356 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node43359 = (inp[5]) ? node43367 : node43360;
														assign node43360 = (inp[3]) ? node43364 : node43361;
															assign node43361 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node43364 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node43367 = (inp[3]) ? node43369 : 4'b0101;
															assign node43369 = (inp[15]) ? 4'b0101 : 4'b0101;
												assign node43372 = (inp[5]) ? node43388 : node43373;
													assign node43373 = (inp[3]) ? node43381 : node43374;
														assign node43374 = (inp[15]) ? node43378 : node43375;
															assign node43375 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node43378 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node43381 = (inp[15]) ? node43385 : node43382;
															assign node43382 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node43385 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node43388 = (inp[15]) ? node43392 : node43389;
														assign node43389 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node43392 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node43395 = (inp[7]) ? node43449 : node43396;
											assign node43396 = (inp[2]) ? node43426 : node43397;
												assign node43397 = (inp[14]) ? node43411 : node43398;
													assign node43398 = (inp[0]) ? node43404 : node43399;
														assign node43399 = (inp[15]) ? node43401 : 4'b1100;
															assign node43401 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node43404 = (inp[15]) ? node43408 : node43405;
															assign node43405 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node43408 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node43411 = (inp[5]) ? node43419 : node43412;
														assign node43412 = (inp[3]) ? node43416 : node43413;
															assign node43413 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node43416 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node43419 = (inp[15]) ? node43423 : node43420;
															assign node43420 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node43423 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node43426 = (inp[5]) ? node43442 : node43427;
													assign node43427 = (inp[15]) ? node43435 : node43428;
														assign node43428 = (inp[0]) ? node43432 : node43429;
															assign node43429 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node43432 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node43435 = (inp[0]) ? node43439 : node43436;
															assign node43436 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node43439 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node43442 = (inp[15]) ? node43446 : node43443;
														assign node43443 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node43446 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node43449 = (inp[14]) ? node43477 : node43450;
												assign node43450 = (inp[2]) ? node43464 : node43451;
													assign node43451 = (inp[15]) ? node43457 : node43452;
														assign node43452 = (inp[0]) ? 4'b0111 : node43453;
															assign node43453 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node43457 = (inp[0]) ? node43461 : node43458;
															assign node43458 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node43461 = (inp[3]) ? 4'b0101 : 4'b0101;
													assign node43464 = (inp[0]) ? node43470 : node43465;
														assign node43465 = (inp[3]) ? 4'b0110 : node43466;
															assign node43466 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node43470 = (inp[15]) ? node43474 : node43471;
															assign node43471 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node43474 = (inp[3]) ? 4'b0100 : 4'b0100;
												assign node43477 = (inp[3]) ? node43493 : node43478;
													assign node43478 = (inp[15]) ? node43486 : node43479;
														assign node43479 = (inp[5]) ? node43483 : node43480;
															assign node43480 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node43483 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node43486 = (inp[5]) ? node43490 : node43487;
															assign node43487 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node43490 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node43493 = (inp[0]) ? node43497 : node43494;
														assign node43494 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node43497 = (inp[15]) ? 4'b0100 : 4'b0110;
								assign node43500 = (inp[13]) ? node43734 : node43501;
									assign node43501 = (inp[7]) ? node43625 : node43502;
										assign node43502 = (inp[8]) ? node43564 : node43503;
											assign node43503 = (inp[14]) ? node43533 : node43504;
												assign node43504 = (inp[2]) ? node43520 : node43505;
													assign node43505 = (inp[0]) ? node43513 : node43506;
														assign node43506 = (inp[15]) ? node43510 : node43507;
															assign node43507 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node43510 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node43513 = (inp[15]) ? node43517 : node43514;
															assign node43514 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node43517 = (inp[5]) ? 4'b1101 : 4'b1101;
													assign node43520 = (inp[0]) ? node43526 : node43521;
														assign node43521 = (inp[15]) ? 4'b1110 : node43522;
															assign node43522 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node43526 = (inp[15]) ? node43530 : node43527;
															assign node43527 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node43530 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node43533 = (inp[2]) ? node43549 : node43534;
													assign node43534 = (inp[5]) ? node43542 : node43535;
														assign node43535 = (inp[3]) ? node43539 : node43536;
															assign node43536 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node43539 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node43542 = (inp[15]) ? node43546 : node43543;
															assign node43543 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node43546 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node43549 = (inp[5]) ? node43557 : node43550;
														assign node43550 = (inp[3]) ? node43554 : node43551;
															assign node43551 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node43554 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node43557 = (inp[0]) ? node43561 : node43558;
															assign node43558 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node43561 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node43564 = (inp[14]) ? node43594 : node43565;
												assign node43565 = (inp[2]) ? node43581 : node43566;
													assign node43566 = (inp[3]) ? node43574 : node43567;
														assign node43567 = (inp[5]) ? node43571 : node43568;
															assign node43568 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node43571 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node43574 = (inp[0]) ? node43578 : node43575;
															assign node43575 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node43578 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node43581 = (inp[15]) ? node43589 : node43582;
														assign node43582 = (inp[0]) ? node43586 : node43583;
															assign node43583 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node43586 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node43589 = (inp[0]) ? 4'b0101 : node43590;
															assign node43590 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node43594 = (inp[3]) ? node43610 : node43595;
													assign node43595 = (inp[0]) ? node43603 : node43596;
														assign node43596 = (inp[5]) ? node43600 : node43597;
															assign node43597 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node43600 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node43603 = (inp[15]) ? node43607 : node43604;
															assign node43604 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node43607 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node43610 = (inp[5]) ? node43618 : node43611;
														assign node43611 = (inp[15]) ? node43615 : node43612;
															assign node43612 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node43615 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node43618 = (inp[15]) ? node43622 : node43619;
															assign node43619 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node43622 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node43625 = (inp[8]) ? node43683 : node43626;
											assign node43626 = (inp[2]) ? node43652 : node43627;
												assign node43627 = (inp[14]) ? node43639 : node43628;
													assign node43628 = (inp[15]) ? node43634 : node43629;
														assign node43629 = (inp[0]) ? node43631 : 4'b1100;
															assign node43631 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node43634 = (inp[5]) ? node43636 : 4'b1110;
															assign node43636 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node43639 = (inp[0]) ? node43645 : node43640;
														assign node43640 = (inp[15]) ? 4'b0111 : node43641;
															assign node43641 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node43645 = (inp[15]) ? node43649 : node43646;
															assign node43646 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node43649 = (inp[3]) ? 4'b0101 : 4'b0101;
												assign node43652 = (inp[3]) ? node43668 : node43653;
													assign node43653 = (inp[5]) ? node43661 : node43654;
														assign node43654 = (inp[14]) ? node43658 : node43655;
															assign node43655 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node43658 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node43661 = (inp[15]) ? node43665 : node43662;
															assign node43662 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node43665 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node43668 = (inp[14]) ? node43676 : node43669;
														assign node43669 = (inp[15]) ? node43673 : node43670;
															assign node43670 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node43673 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node43676 = (inp[0]) ? node43680 : node43677;
															assign node43677 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node43680 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node43683 = (inp[14]) ? node43711 : node43684;
												assign node43684 = (inp[2]) ? node43698 : node43685;
													assign node43685 = (inp[5]) ? node43693 : node43686;
														assign node43686 = (inp[3]) ? node43690 : node43687;
															assign node43687 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node43690 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node43693 = (inp[3]) ? node43695 : 4'b0101;
															assign node43695 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node43698 = (inp[0]) ? node43704 : node43699;
														assign node43699 = (inp[15]) ? node43701 : 4'b0100;
															assign node43701 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node43704 = (inp[15]) ? node43708 : node43705;
															assign node43705 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node43708 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node43711 = (inp[15]) ? node43723 : node43712;
													assign node43712 = (inp[0]) ? node43718 : node43713;
														assign node43713 = (inp[5]) ? 4'b0100 : node43714;
															assign node43714 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node43718 = (inp[3]) ? 4'b0110 : node43719;
															assign node43719 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node43723 = (inp[0]) ? node43729 : node43724;
														assign node43724 = (inp[5]) ? 4'b0110 : node43725;
															assign node43725 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node43729 = (inp[5]) ? 4'b0100 : node43730;
															assign node43730 = (inp[3]) ? 4'b0100 : 4'b0110;
									assign node43734 = (inp[8]) ? node43846 : node43735;
										assign node43735 = (inp[7]) ? node43793 : node43736;
											assign node43736 = (inp[14]) ? node43762 : node43737;
												assign node43737 = (inp[2]) ? node43749 : node43738;
													assign node43738 = (inp[15]) ? node43744 : node43739;
														assign node43739 = (inp[0]) ? 4'b0111 : node43740;
															assign node43740 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node43744 = (inp[0]) ? 4'b0101 : node43745;
															assign node43745 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node43749 = (inp[3]) ? node43755 : node43750;
														assign node43750 = (inp[5]) ? 4'b0100 : node43751;
															assign node43751 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node43755 = (inp[5]) ? node43759 : node43756;
															assign node43756 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node43759 = (inp[15]) ? 4'b0100 : 4'b0100;
												assign node43762 = (inp[5]) ? node43778 : node43763;
													assign node43763 = (inp[15]) ? node43771 : node43764;
														assign node43764 = (inp[2]) ? node43768 : node43765;
															assign node43765 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node43768 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node43771 = (inp[0]) ? node43775 : node43772;
															assign node43772 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node43775 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node43778 = (inp[3]) ? node43786 : node43779;
														assign node43779 = (inp[2]) ? node43783 : node43780;
															assign node43780 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node43783 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node43786 = (inp[15]) ? node43790 : node43787;
															assign node43787 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node43790 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node43793 = (inp[14]) ? node43823 : node43794;
												assign node43794 = (inp[2]) ? node43810 : node43795;
													assign node43795 = (inp[3]) ? node43803 : node43796;
														assign node43796 = (inp[15]) ? node43800 : node43797;
															assign node43797 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node43800 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node43803 = (inp[5]) ? node43807 : node43804;
															assign node43804 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node43807 = (inp[0]) ? 4'b0100 : 4'b0100;
													assign node43810 = (inp[5]) ? node43816 : node43811;
														assign node43811 = (inp[0]) ? node43813 : 4'b0101;
															assign node43813 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node43816 = (inp[3]) ? node43820 : node43817;
															assign node43817 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node43820 = (inp[0]) ? 4'b0101 : 4'b0101;
												assign node43823 = (inp[0]) ? node43835 : node43824;
													assign node43824 = (inp[15]) ? node43830 : node43825;
														assign node43825 = (inp[5]) ? 4'b0101 : node43826;
															assign node43826 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node43830 = (inp[5]) ? 4'b0111 : node43831;
															assign node43831 = (inp[2]) ? 4'b0101 : 4'b0111;
													assign node43835 = (inp[15]) ? node43841 : node43836;
														assign node43836 = (inp[3]) ? 4'b0111 : node43837;
															assign node43837 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node43841 = (inp[3]) ? 4'b0101 : node43842;
															assign node43842 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node43846 = (inp[7]) ? node43902 : node43847;
											assign node43847 = (inp[2]) ? node43879 : node43848;
												assign node43848 = (inp[14]) ? node43864 : node43849;
													assign node43849 = (inp[0]) ? node43857 : node43850;
														assign node43850 = (inp[15]) ? node43854 : node43851;
															assign node43851 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node43854 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node43857 = (inp[15]) ? node43861 : node43858;
															assign node43858 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node43861 = (inp[3]) ? 4'b0100 : 4'b0100;
													assign node43864 = (inp[5]) ? node43872 : node43865;
														assign node43865 = (inp[3]) ? node43869 : node43866;
															assign node43866 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node43869 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node43872 = (inp[0]) ? node43876 : node43873;
															assign node43873 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node43876 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node43879 = (inp[15]) ? node43891 : node43880;
													assign node43880 = (inp[0]) ? node43886 : node43881;
														assign node43881 = (inp[3]) ? 4'b0101 : node43882;
															assign node43882 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node43886 = (inp[5]) ? 4'b0111 : node43887;
															assign node43887 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node43891 = (inp[0]) ? node43897 : node43892;
														assign node43892 = (inp[5]) ? 4'b0111 : node43893;
															assign node43893 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node43897 = (inp[5]) ? 4'b0101 : node43898;
															assign node43898 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node43902 = (inp[2]) ? node43930 : node43903;
												assign node43903 = (inp[14]) ? node43919 : node43904;
													assign node43904 = (inp[3]) ? node43912 : node43905;
														assign node43905 = (inp[5]) ? node43909 : node43906;
															assign node43906 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node43909 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node43912 = (inp[0]) ? node43916 : node43913;
															assign node43913 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node43916 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node43919 = (inp[5]) ? node43925 : node43920;
														assign node43920 = (inp[0]) ? node43922 : 4'b0110;
															assign node43922 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node43925 = (inp[15]) ? 4'b0100 : node43926;
															assign node43926 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node43930 = (inp[5]) ? node43944 : node43931;
													assign node43931 = (inp[14]) ? node43939 : node43932;
														assign node43932 = (inp[15]) ? node43936 : node43933;
															assign node43933 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node43936 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node43939 = (inp[3]) ? 4'b0110 : node43940;
															assign node43940 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node43944 = (inp[0]) ? node43948 : node43945;
														assign node43945 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node43948 = (inp[15]) ? 4'b0100 : 4'b0110;
							assign node43951 = (inp[1]) ? node44401 : node43952;
								assign node43952 = (inp[13]) ? node44184 : node43953;
									assign node43953 = (inp[5]) ? node44077 : node43954;
										assign node43954 = (inp[7]) ? node44014 : node43955;
											assign node43955 = (inp[8]) ? node43985 : node43956;
												assign node43956 = (inp[14]) ? node43970 : node43957;
													assign node43957 = (inp[2]) ? node43965 : node43958;
														assign node43958 = (inp[15]) ? node43962 : node43959;
															assign node43959 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node43962 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node43965 = (inp[0]) ? 4'b0100 : node43966;
															assign node43966 = (inp[3]) ? 4'b0100 : 4'b0100;
													assign node43970 = (inp[3]) ? node43978 : node43971;
														assign node43971 = (inp[2]) ? node43975 : node43972;
															assign node43972 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node43975 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node43978 = (inp[0]) ? node43982 : node43979;
															assign node43979 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node43982 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node43985 = (inp[14]) ? node43999 : node43986;
													assign node43986 = (inp[2]) ? node43992 : node43987;
														assign node43987 = (inp[3]) ? node43989 : 4'b0110;
															assign node43989 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node43992 = (inp[0]) ? node43996 : node43993;
															assign node43993 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node43996 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node43999 = (inp[2]) ? node44007 : node44000;
														assign node44000 = (inp[15]) ? node44004 : node44001;
															assign node44001 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node44004 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node44007 = (inp[3]) ? node44011 : node44008;
															assign node44008 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node44011 = (inp[15]) ? 4'b0101 : 4'b0101;
											assign node44014 = (inp[8]) ? node44046 : node44015;
												assign node44015 = (inp[2]) ? node44031 : node44016;
													assign node44016 = (inp[14]) ? node44024 : node44017;
														assign node44017 = (inp[0]) ? node44021 : node44018;
															assign node44018 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node44021 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node44024 = (inp[15]) ? node44028 : node44025;
															assign node44025 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node44028 = (inp[3]) ? 4'b0101 : 4'b0101;
													assign node44031 = (inp[15]) ? node44039 : node44032;
														assign node44032 = (inp[14]) ? node44036 : node44033;
															assign node44033 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node44036 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node44039 = (inp[0]) ? node44043 : node44040;
															assign node44040 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node44043 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node44046 = (inp[2]) ? node44062 : node44047;
													assign node44047 = (inp[14]) ? node44055 : node44048;
														assign node44048 = (inp[0]) ? node44052 : node44049;
															assign node44049 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node44052 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node44055 = (inp[0]) ? node44059 : node44056;
															assign node44056 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node44059 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node44062 = (inp[0]) ? node44070 : node44063;
														assign node44063 = (inp[14]) ? node44067 : node44064;
															assign node44064 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node44067 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node44070 = (inp[3]) ? node44074 : node44071;
															assign node44071 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node44074 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node44077 = (inp[0]) ? node44131 : node44078;
											assign node44078 = (inp[15]) ? node44102 : node44079;
												assign node44079 = (inp[7]) ? node44091 : node44080;
													assign node44080 = (inp[8]) ? node44086 : node44081;
														assign node44081 = (inp[2]) ? 4'b0100 : node44082;
															assign node44082 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node44086 = (inp[2]) ? 4'b0101 : node44087;
															assign node44087 = (inp[14]) ? 4'b0101 : 4'b0100;
													assign node44091 = (inp[8]) ? node44097 : node44092;
														assign node44092 = (inp[2]) ? 4'b0101 : node44093;
															assign node44093 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node44097 = (inp[14]) ? 4'b0100 : node44098;
															assign node44098 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node44102 = (inp[2]) ? node44118 : node44103;
													assign node44103 = (inp[8]) ? node44111 : node44104;
														assign node44104 = (inp[3]) ? node44108 : node44105;
															assign node44105 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node44108 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node44111 = (inp[3]) ? node44115 : node44112;
															assign node44112 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node44115 = (inp[14]) ? 4'b0110 : 4'b0110;
													assign node44118 = (inp[14]) ? node44124 : node44119;
														assign node44119 = (inp[7]) ? node44121 : 4'b0111;
															assign node44121 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node44124 = (inp[3]) ? node44128 : node44125;
															assign node44125 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node44128 = (inp[8]) ? 4'b0110 : 4'b0110;
											assign node44131 = (inp[15]) ? node44155 : node44132;
												assign node44132 = (inp[2]) ? node44148 : node44133;
													assign node44133 = (inp[3]) ? node44141 : node44134;
														assign node44134 = (inp[8]) ? node44138 : node44135;
															assign node44135 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node44138 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node44141 = (inp[14]) ? node44145 : node44142;
															assign node44142 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node44145 = (inp[8]) ? 4'b0110 : 4'b0110;
													assign node44148 = (inp[8]) ? node44152 : node44149;
														assign node44149 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node44152 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node44155 = (inp[14]) ? node44171 : node44156;
													assign node44156 = (inp[7]) ? node44164 : node44157;
														assign node44157 = (inp[8]) ? node44161 : node44158;
															assign node44158 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node44161 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node44164 = (inp[2]) ? node44168 : node44165;
															assign node44165 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node44168 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node44171 = (inp[3]) ? node44179 : node44172;
														assign node44172 = (inp[8]) ? node44176 : node44173;
															assign node44173 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node44176 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node44179 = (inp[7]) ? 4'b0100 : node44180;
															assign node44180 = (inp[8]) ? 4'b0101 : 4'b0100;
									assign node44184 = (inp[7]) ? node44294 : node44185;
										assign node44185 = (inp[8]) ? node44241 : node44186;
											assign node44186 = (inp[14]) ? node44218 : node44187;
												assign node44187 = (inp[2]) ? node44203 : node44188;
													assign node44188 = (inp[5]) ? node44196 : node44189;
														assign node44189 = (inp[3]) ? node44193 : node44190;
															assign node44190 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node44193 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node44196 = (inp[0]) ? node44200 : node44197;
															assign node44197 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node44200 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node44203 = (inp[3]) ? node44211 : node44204;
														assign node44204 = (inp[0]) ? node44208 : node44205;
															assign node44205 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node44208 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node44211 = (inp[0]) ? node44215 : node44212;
															assign node44212 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node44215 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node44218 = (inp[3]) ? node44234 : node44219;
													assign node44219 = (inp[5]) ? node44227 : node44220;
														assign node44220 = (inp[0]) ? node44224 : node44221;
															assign node44221 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node44224 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node44227 = (inp[2]) ? node44231 : node44228;
															assign node44228 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node44231 = (inp[0]) ? 4'b0100 : 4'b0100;
													assign node44234 = (inp[0]) ? node44238 : node44235;
														assign node44235 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node44238 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node44241 = (inp[2]) ? node44273 : node44242;
												assign node44242 = (inp[14]) ? node44258 : node44243;
													assign node44243 = (inp[0]) ? node44251 : node44244;
														assign node44244 = (inp[15]) ? node44248 : node44245;
															assign node44245 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node44248 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node44251 = (inp[15]) ? node44255 : node44252;
															assign node44252 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node44255 = (inp[3]) ? 4'b0100 : 4'b0100;
													assign node44258 = (inp[15]) ? node44266 : node44259;
														assign node44259 = (inp[0]) ? node44263 : node44260;
															assign node44260 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node44263 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node44266 = (inp[0]) ? node44270 : node44267;
															assign node44267 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node44270 = (inp[3]) ? 4'b1101 : 4'b1101;
												assign node44273 = (inp[5]) ? node44287 : node44274;
													assign node44274 = (inp[14]) ? node44282 : node44275;
														assign node44275 = (inp[15]) ? node44279 : node44276;
															assign node44276 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node44279 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node44282 = (inp[15]) ? node44284 : 4'b1111;
															assign node44284 = (inp[0]) ? 4'b1101 : 4'b1101;
													assign node44287 = (inp[15]) ? node44291 : node44288;
														assign node44288 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node44291 = (inp[0]) ? 4'b1101 : 4'b1111;
										assign node44294 = (inp[8]) ? node44352 : node44295;
											assign node44295 = (inp[2]) ? node44323 : node44296;
												assign node44296 = (inp[14]) ? node44310 : node44297;
													assign node44297 = (inp[15]) ? node44305 : node44298;
														assign node44298 = (inp[0]) ? node44302 : node44299;
															assign node44299 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node44302 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node44305 = (inp[0]) ? 4'b0100 : node44306;
															assign node44306 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node44310 = (inp[15]) ? node44316 : node44311;
														assign node44311 = (inp[5]) ? 4'b1101 : node44312;
															assign node44312 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node44316 = (inp[3]) ? node44320 : node44317;
															assign node44317 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node44320 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node44323 = (inp[5]) ? node44337 : node44324;
													assign node44324 = (inp[14]) ? node44332 : node44325;
														assign node44325 = (inp[3]) ? node44329 : node44326;
															assign node44326 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node44329 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node44332 = (inp[0]) ? node44334 : 4'b1111;
															assign node44334 = (inp[15]) ? 4'b1101 : 4'b1101;
													assign node44337 = (inp[3]) ? node44345 : node44338;
														assign node44338 = (inp[0]) ? node44342 : node44339;
															assign node44339 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node44342 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node44345 = (inp[0]) ? node44349 : node44346;
															assign node44346 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node44349 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node44352 = (inp[14]) ? node44378 : node44353;
												assign node44353 = (inp[2]) ? node44365 : node44354;
													assign node44354 = (inp[15]) ? node44358 : node44355;
														assign node44355 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node44358 = (inp[0]) ? node44362 : node44359;
															assign node44359 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node44362 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node44365 = (inp[0]) ? node44373 : node44366;
														assign node44366 = (inp[15]) ? node44370 : node44367;
															assign node44367 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node44370 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node44373 = (inp[15]) ? 4'b1100 : node44374;
															assign node44374 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node44378 = (inp[5]) ? node44394 : node44379;
													assign node44379 = (inp[15]) ? node44387 : node44380;
														assign node44380 = (inp[2]) ? node44384 : node44381;
															assign node44381 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node44384 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node44387 = (inp[2]) ? node44391 : node44388;
															assign node44388 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node44391 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node44394 = (inp[0]) ? node44398 : node44395;
														assign node44395 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node44398 = (inp[15]) ? 4'b1100 : 4'b1110;
								assign node44401 = (inp[13]) ? node44621 : node44402;
									assign node44402 = (inp[8]) ? node44512 : node44403;
										assign node44403 = (inp[7]) ? node44459 : node44404;
											assign node44404 = (inp[14]) ? node44436 : node44405;
												assign node44405 = (inp[2]) ? node44421 : node44406;
													assign node44406 = (inp[15]) ? node44414 : node44407;
														assign node44407 = (inp[0]) ? node44411 : node44408;
															assign node44408 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node44411 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node44414 = (inp[0]) ? node44418 : node44415;
															assign node44415 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node44418 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node44421 = (inp[3]) ? node44429 : node44422;
														assign node44422 = (inp[15]) ? node44426 : node44423;
															assign node44423 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node44426 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node44429 = (inp[0]) ? node44433 : node44430;
															assign node44430 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node44433 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node44436 = (inp[3]) ? node44452 : node44437;
													assign node44437 = (inp[5]) ? node44445 : node44438;
														assign node44438 = (inp[15]) ? node44442 : node44439;
															assign node44439 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node44442 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node44445 = (inp[0]) ? node44449 : node44446;
															assign node44446 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node44449 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node44452 = (inp[0]) ? node44456 : node44453;
														assign node44453 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node44456 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node44459 = (inp[2]) ? node44489 : node44460;
												assign node44460 = (inp[14]) ? node44474 : node44461;
													assign node44461 = (inp[5]) ? node44467 : node44462;
														assign node44462 = (inp[0]) ? 4'b0100 : node44463;
															assign node44463 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node44467 = (inp[3]) ? node44471 : node44468;
															assign node44468 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node44471 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node44474 = (inp[3]) ? node44482 : node44475;
														assign node44475 = (inp[0]) ? node44479 : node44476;
															assign node44476 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node44479 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node44482 = (inp[15]) ? node44486 : node44483;
															assign node44483 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node44486 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node44489 = (inp[15]) ? node44501 : node44490;
													assign node44490 = (inp[0]) ? node44496 : node44491;
														assign node44491 = (inp[5]) ? 4'b1101 : node44492;
															assign node44492 = (inp[14]) ? 4'b1111 : 4'b1101;
														assign node44496 = (inp[3]) ? 4'b1111 : node44497;
															assign node44497 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node44501 = (inp[0]) ? node44507 : node44502;
														assign node44502 = (inp[3]) ? 4'b1111 : node44503;
															assign node44503 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node44507 = (inp[3]) ? 4'b1101 : node44508;
															assign node44508 = (inp[5]) ? 4'b1101 : 4'b1111;
										assign node44512 = (inp[7]) ? node44566 : node44513;
											assign node44513 = (inp[14]) ? node44543 : node44514;
												assign node44514 = (inp[2]) ? node44528 : node44515;
													assign node44515 = (inp[3]) ? node44521 : node44516;
														assign node44516 = (inp[15]) ? node44518 : 4'b0100;
															assign node44518 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node44521 = (inp[15]) ? node44525 : node44522;
															assign node44522 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node44525 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node44528 = (inp[0]) ? node44536 : node44529;
														assign node44529 = (inp[15]) ? node44533 : node44530;
															assign node44530 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node44533 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node44536 = (inp[15]) ? node44540 : node44537;
															assign node44537 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node44540 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node44543 = (inp[0]) ? node44555 : node44544;
													assign node44544 = (inp[15]) ? node44550 : node44545;
														assign node44545 = (inp[3]) ? 4'b1101 : node44546;
															assign node44546 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node44550 = (inp[3]) ? 4'b1111 : node44551;
															assign node44551 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node44555 = (inp[15]) ? node44561 : node44556;
														assign node44556 = (inp[3]) ? 4'b1111 : node44557;
															assign node44557 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node44561 = (inp[3]) ? 4'b1101 : node44562;
															assign node44562 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node44566 = (inp[2]) ? node44598 : node44567;
												assign node44567 = (inp[14]) ? node44583 : node44568;
													assign node44568 = (inp[0]) ? node44576 : node44569;
														assign node44569 = (inp[15]) ? node44573 : node44570;
															assign node44570 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node44573 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node44576 = (inp[15]) ? node44580 : node44577;
															assign node44577 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node44580 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node44583 = (inp[3]) ? node44591 : node44584;
														assign node44584 = (inp[5]) ? node44588 : node44585;
															assign node44585 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node44588 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node44591 = (inp[5]) ? node44595 : node44592;
															assign node44592 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node44595 = (inp[15]) ? 4'b1100 : 4'b1100;
												assign node44598 = (inp[5]) ? node44614 : node44599;
													assign node44599 = (inp[0]) ? node44607 : node44600;
														assign node44600 = (inp[15]) ? node44604 : node44601;
															assign node44601 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node44604 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node44607 = (inp[15]) ? node44611 : node44608;
															assign node44608 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node44611 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node44614 = (inp[0]) ? node44618 : node44615;
														assign node44615 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node44618 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node44621 = (inp[8]) ? node44739 : node44622;
										assign node44622 = (inp[7]) ? node44684 : node44623;
											assign node44623 = (inp[14]) ? node44653 : node44624;
												assign node44624 = (inp[2]) ? node44638 : node44625;
													assign node44625 = (inp[0]) ? node44633 : node44626;
														assign node44626 = (inp[15]) ? node44630 : node44627;
															assign node44627 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node44630 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node44633 = (inp[15]) ? 4'b1101 : node44634;
															assign node44634 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node44638 = (inp[15]) ? node44646 : node44639;
														assign node44639 = (inp[0]) ? node44643 : node44640;
															assign node44640 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node44643 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node44646 = (inp[0]) ? node44650 : node44647;
															assign node44647 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node44650 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node44653 = (inp[2]) ? node44669 : node44654;
													assign node44654 = (inp[0]) ? node44662 : node44655;
														assign node44655 = (inp[15]) ? node44659 : node44656;
															assign node44656 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node44659 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node44662 = (inp[15]) ? node44666 : node44663;
															assign node44663 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node44666 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node44669 = (inp[15]) ? node44677 : node44670;
														assign node44670 = (inp[0]) ? node44674 : node44671;
															assign node44671 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node44674 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node44677 = (inp[0]) ? node44681 : node44678;
															assign node44678 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node44681 = (inp[3]) ? 4'b1100 : 4'b1100;
											assign node44684 = (inp[14]) ? node44716 : node44685;
												assign node44685 = (inp[2]) ? node44701 : node44686;
													assign node44686 = (inp[0]) ? node44694 : node44687;
														assign node44687 = (inp[15]) ? node44691 : node44688;
															assign node44688 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node44691 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node44694 = (inp[15]) ? node44698 : node44695;
															assign node44695 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node44698 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node44701 = (inp[3]) ? node44709 : node44702;
														assign node44702 = (inp[15]) ? node44706 : node44703;
															assign node44703 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node44706 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node44709 = (inp[0]) ? node44713 : node44710;
															assign node44710 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node44713 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node44716 = (inp[0]) ? node44728 : node44717;
													assign node44717 = (inp[15]) ? node44723 : node44718;
														assign node44718 = (inp[3]) ? 4'b1101 : node44719;
															assign node44719 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node44723 = (inp[5]) ? 4'b1111 : node44724;
															assign node44724 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node44728 = (inp[15]) ? node44734 : node44729;
														assign node44729 = (inp[5]) ? 4'b1111 : node44730;
															assign node44730 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node44734 = (inp[5]) ? 4'b1101 : node44735;
															assign node44735 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node44739 = (inp[7]) ? node44799 : node44740;
											assign node44740 = (inp[14]) ? node44768 : node44741;
												assign node44741 = (inp[2]) ? node44755 : node44742;
													assign node44742 = (inp[0]) ? node44748 : node44743;
														assign node44743 = (inp[5]) ? 4'b1100 : node44744;
															assign node44744 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node44748 = (inp[15]) ? node44752 : node44749;
															assign node44749 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node44752 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node44755 = (inp[5]) ? node44763 : node44756;
														assign node44756 = (inp[0]) ? node44760 : node44757;
															assign node44757 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node44760 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node44763 = (inp[15]) ? 4'b1111 : node44764;
															assign node44764 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node44768 = (inp[5]) ? node44784 : node44769;
													assign node44769 = (inp[3]) ? node44777 : node44770;
														assign node44770 = (inp[2]) ? node44774 : node44771;
															assign node44771 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node44774 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node44777 = (inp[2]) ? node44781 : node44778;
															assign node44778 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node44781 = (inp[0]) ? 4'b1101 : 4'b1101;
													assign node44784 = (inp[3]) ? node44792 : node44785;
														assign node44785 = (inp[2]) ? node44789 : node44786;
															assign node44786 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node44789 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node44792 = (inp[15]) ? node44796 : node44793;
															assign node44793 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node44796 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node44799 = (inp[2]) ? node44827 : node44800;
												assign node44800 = (inp[14]) ? node44812 : node44801;
													assign node44801 = (inp[15]) ? node44807 : node44802;
														assign node44802 = (inp[0]) ? node44804 : 4'b1101;
															assign node44804 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node44807 = (inp[0]) ? 4'b1101 : node44808;
															assign node44808 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node44812 = (inp[5]) ? node44820 : node44813;
														assign node44813 = (inp[0]) ? node44817 : node44814;
															assign node44814 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node44817 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node44820 = (inp[3]) ? node44824 : node44821;
															assign node44821 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node44824 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node44827 = (inp[3]) ? node44843 : node44828;
													assign node44828 = (inp[14]) ? node44836 : node44829;
														assign node44829 = (inp[5]) ? node44833 : node44830;
															assign node44830 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node44833 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node44836 = (inp[0]) ? node44840 : node44837;
															assign node44837 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node44840 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node44843 = (inp[15]) ? node44847 : node44844;
														assign node44844 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node44847 = (inp[0]) ? 4'b1100 : 4'b1110;
						assign node44850 = (inp[11]) ? node45778 : node44851;
							assign node44851 = (inp[13]) ? node45297 : node44852;
								assign node44852 = (inp[1]) ? node45070 : node44853;
									assign node44853 = (inp[14]) ? node44969 : node44854;
										assign node44854 = (inp[7]) ? node44918 : node44855;
											assign node44855 = (inp[0]) ? node44887 : node44856;
												assign node44856 = (inp[15]) ? node44872 : node44857;
													assign node44857 = (inp[3]) ? node44865 : node44858;
														assign node44858 = (inp[5]) ? node44862 : node44859;
															assign node44859 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node44862 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node44865 = (inp[8]) ? node44869 : node44866;
															assign node44866 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node44869 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node44872 = (inp[3]) ? node44880 : node44873;
														assign node44873 = (inp[5]) ? node44877 : node44874;
															assign node44874 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node44877 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node44880 = (inp[5]) ? node44884 : node44881;
															assign node44881 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node44884 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node44887 = (inp[15]) ? node44903 : node44888;
													assign node44888 = (inp[5]) ? node44896 : node44889;
														assign node44889 = (inp[3]) ? node44893 : node44890;
															assign node44890 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node44893 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node44896 = (inp[2]) ? node44900 : node44897;
															assign node44897 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node44900 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node44903 = (inp[3]) ? node44911 : node44904;
														assign node44904 = (inp[5]) ? node44908 : node44905;
															assign node44905 = (inp[2]) ? 4'b0110 : 4'b0110;
															assign node44908 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node44911 = (inp[2]) ? node44915 : node44912;
															assign node44912 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node44915 = (inp[8]) ? 4'b0101 : 4'b0100;
											assign node44918 = (inp[5]) ? node44944 : node44919;
												assign node44919 = (inp[2]) ? node44933 : node44920;
													assign node44920 = (inp[8]) ? node44928 : node44921;
														assign node44921 = (inp[3]) ? node44925 : node44922;
															assign node44922 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node44925 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node44928 = (inp[15]) ? node44930 : 4'b0111;
															assign node44930 = (inp[0]) ? 4'b0101 : 4'b0101;
													assign node44933 = (inp[8]) ? node44939 : node44934;
														assign node44934 = (inp[0]) ? 4'b0111 : node44935;
															assign node44935 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node44939 = (inp[3]) ? 4'b0110 : node44940;
															assign node44940 = (inp[0]) ? 4'b0100 : 4'b0100;
												assign node44944 = (inp[8]) ? node44954 : node44945;
													assign node44945 = (inp[2]) ? 4'b0111 : node44946;
														assign node44946 = (inp[15]) ? node44950 : node44947;
															assign node44947 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node44950 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node44954 = (inp[2]) ? node44962 : node44955;
														assign node44955 = (inp[3]) ? node44959 : node44956;
															assign node44956 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node44959 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node44962 = (inp[0]) ? node44966 : node44963;
															assign node44963 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node44966 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node44969 = (inp[7]) ? node45017 : node44970;
											assign node44970 = (inp[8]) ? node44994 : node44971;
												assign node44971 = (inp[0]) ? node44983 : node44972;
													assign node44972 = (inp[15]) ? node44978 : node44973;
														assign node44973 = (inp[3]) ? 4'b0100 : node44974;
															assign node44974 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node44978 = (inp[3]) ? 4'b0110 : node44979;
															assign node44979 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node44983 = (inp[15]) ? node44989 : node44984;
														assign node44984 = (inp[3]) ? 4'b0110 : node44985;
															assign node44985 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node44989 = (inp[5]) ? 4'b0100 : node44990;
															assign node44990 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node44994 = (inp[15]) ? node45006 : node44995;
													assign node44995 = (inp[0]) ? node45001 : node44996;
														assign node44996 = (inp[3]) ? 4'b0101 : node44997;
															assign node44997 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node45001 = (inp[3]) ? 4'b0111 : node45002;
															assign node45002 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node45006 = (inp[0]) ? node45012 : node45007;
														assign node45007 = (inp[3]) ? 4'b0111 : node45008;
															assign node45008 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node45012 = (inp[5]) ? 4'b0101 : node45013;
															assign node45013 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node45017 = (inp[8]) ? node45047 : node45018;
												assign node45018 = (inp[2]) ? node45032 : node45019;
													assign node45019 = (inp[3]) ? node45025 : node45020;
														assign node45020 = (inp[0]) ? node45022 : 4'b0101;
															assign node45022 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node45025 = (inp[0]) ? node45029 : node45026;
															assign node45026 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node45029 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node45032 = (inp[0]) ? node45040 : node45033;
														assign node45033 = (inp[15]) ? node45037 : node45034;
															assign node45034 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node45037 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node45040 = (inp[15]) ? node45044 : node45041;
															assign node45041 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node45044 = (inp[3]) ? 4'b0101 : 4'b0101;
												assign node45047 = (inp[5]) ? node45063 : node45048;
													assign node45048 = (inp[2]) ? node45056 : node45049;
														assign node45049 = (inp[3]) ? node45053 : node45050;
															assign node45050 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node45053 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node45056 = (inp[3]) ? node45060 : node45057;
															assign node45057 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node45060 = (inp[0]) ? 4'b0100 : 4'b0100;
													assign node45063 = (inp[0]) ? node45067 : node45064;
														assign node45064 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node45067 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node45070 = (inp[7]) ? node45180 : node45071;
										assign node45071 = (inp[8]) ? node45127 : node45072;
											assign node45072 = (inp[2]) ? node45104 : node45073;
												assign node45073 = (inp[14]) ? node45089 : node45074;
													assign node45074 = (inp[0]) ? node45082 : node45075;
														assign node45075 = (inp[15]) ? node45079 : node45076;
															assign node45076 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node45079 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node45082 = (inp[15]) ? node45086 : node45083;
															assign node45083 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node45086 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node45089 = (inp[15]) ? node45097 : node45090;
														assign node45090 = (inp[0]) ? node45094 : node45091;
															assign node45091 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node45094 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node45097 = (inp[0]) ? node45101 : node45098;
															assign node45098 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node45101 = (inp[5]) ? 4'b0100 : 4'b0100;
												assign node45104 = (inp[0]) ? node45116 : node45105;
													assign node45105 = (inp[15]) ? node45111 : node45106;
														assign node45106 = (inp[5]) ? 4'b0100 : node45107;
															assign node45107 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node45111 = (inp[3]) ? 4'b0110 : node45112;
															assign node45112 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node45116 = (inp[15]) ? node45122 : node45117;
														assign node45117 = (inp[5]) ? 4'b0110 : node45118;
															assign node45118 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node45122 = (inp[3]) ? 4'b0100 : node45123;
															assign node45123 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node45127 = (inp[14]) ? node45157 : node45128;
												assign node45128 = (inp[2]) ? node45144 : node45129;
													assign node45129 = (inp[0]) ? node45137 : node45130;
														assign node45130 = (inp[15]) ? node45134 : node45131;
															assign node45131 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node45134 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node45137 = (inp[15]) ? node45141 : node45138;
															assign node45138 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node45141 = (inp[3]) ? 4'b0100 : 4'b0100;
													assign node45144 = (inp[5]) ? node45150 : node45145;
														assign node45145 = (inp[15]) ? node45147 : 4'b1111;
															assign node45147 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node45150 = (inp[3]) ? node45154 : node45151;
															assign node45151 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node45154 = (inp[15]) ? 4'b1101 : 4'b1101;
												assign node45157 = (inp[15]) ? node45169 : node45158;
													assign node45158 = (inp[0]) ? node45164 : node45159;
														assign node45159 = (inp[5]) ? 4'b1101 : node45160;
															assign node45160 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node45164 = (inp[3]) ? 4'b1111 : node45165;
															assign node45165 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node45169 = (inp[0]) ? node45175 : node45170;
														assign node45170 = (inp[3]) ? 4'b1111 : node45171;
															assign node45171 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node45175 = (inp[3]) ? 4'b1101 : node45176;
															assign node45176 = (inp[5]) ? 4'b1101 : 4'b1111;
										assign node45180 = (inp[8]) ? node45236 : node45181;
											assign node45181 = (inp[14]) ? node45213 : node45182;
												assign node45182 = (inp[2]) ? node45198 : node45183;
													assign node45183 = (inp[5]) ? node45191 : node45184;
														assign node45184 = (inp[0]) ? node45188 : node45185;
															assign node45185 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node45188 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node45191 = (inp[3]) ? node45195 : node45192;
															assign node45192 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node45195 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node45198 = (inp[5]) ? node45206 : node45199;
														assign node45199 = (inp[0]) ? node45203 : node45200;
															assign node45200 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node45203 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node45206 = (inp[3]) ? node45210 : node45207;
															assign node45207 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node45210 = (inp[15]) ? 4'b1101 : 4'b1101;
												assign node45213 = (inp[3]) ? node45229 : node45214;
													assign node45214 = (inp[5]) ? node45222 : node45215;
														assign node45215 = (inp[2]) ? node45219 : node45216;
															assign node45216 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node45219 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node45222 = (inp[2]) ? node45226 : node45223;
															assign node45223 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node45226 = (inp[0]) ? 4'b1101 : 4'b1101;
													assign node45229 = (inp[15]) ? node45233 : node45230;
														assign node45230 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node45233 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node45236 = (inp[14]) ? node45266 : node45237;
												assign node45237 = (inp[2]) ? node45253 : node45238;
													assign node45238 = (inp[0]) ? node45246 : node45239;
														assign node45239 = (inp[15]) ? node45243 : node45240;
															assign node45240 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node45243 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node45246 = (inp[15]) ? node45250 : node45247;
															assign node45247 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node45250 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node45253 = (inp[0]) ? node45259 : node45254;
														assign node45254 = (inp[15]) ? node45256 : 4'b1100;
															assign node45256 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node45259 = (inp[15]) ? node45263 : node45260;
															assign node45260 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node45263 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node45266 = (inp[2]) ? node45282 : node45267;
													assign node45267 = (inp[3]) ? node45275 : node45268;
														assign node45268 = (inp[0]) ? node45272 : node45269;
															assign node45269 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node45272 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node45275 = (inp[0]) ? node45279 : node45276;
															assign node45276 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node45279 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node45282 = (inp[15]) ? node45290 : node45283;
														assign node45283 = (inp[0]) ? node45287 : node45284;
															assign node45284 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node45287 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node45290 = (inp[0]) ? node45294 : node45291;
															assign node45291 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node45294 = (inp[5]) ? 4'b1100 : 4'b1110;
								assign node45297 = (inp[1]) ? node45529 : node45298;
									assign node45298 = (inp[7]) ? node45414 : node45299;
										assign node45299 = (inp[8]) ? node45353 : node45300;
											assign node45300 = (inp[14]) ? node45330 : node45301;
												assign node45301 = (inp[2]) ? node45317 : node45302;
													assign node45302 = (inp[0]) ? node45310 : node45303;
														assign node45303 = (inp[15]) ? node45307 : node45304;
															assign node45304 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node45307 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node45310 = (inp[15]) ? node45314 : node45311;
															assign node45311 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node45314 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node45317 = (inp[0]) ? node45325 : node45318;
														assign node45318 = (inp[15]) ? node45322 : node45319;
															assign node45319 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node45322 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node45325 = (inp[15]) ? node45327 : 4'b0110;
															assign node45327 = (inp[3]) ? 4'b0100 : 4'b0100;
												assign node45330 = (inp[15]) ? node45342 : node45331;
													assign node45331 = (inp[0]) ? node45337 : node45332;
														assign node45332 = (inp[5]) ? 4'b0100 : node45333;
															assign node45333 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node45337 = (inp[5]) ? 4'b0110 : node45338;
															assign node45338 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node45342 = (inp[0]) ? node45348 : node45343;
														assign node45343 = (inp[3]) ? 4'b0110 : node45344;
															assign node45344 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node45348 = (inp[3]) ? 4'b0100 : node45349;
															assign node45349 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node45353 = (inp[14]) ? node45385 : node45354;
												assign node45354 = (inp[2]) ? node45370 : node45355;
													assign node45355 = (inp[3]) ? node45363 : node45356;
														assign node45356 = (inp[5]) ? node45360 : node45357;
															assign node45357 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node45360 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node45363 = (inp[15]) ? node45367 : node45364;
															assign node45364 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node45367 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node45370 = (inp[3]) ? node45378 : node45371;
														assign node45371 = (inp[15]) ? node45375 : node45372;
															assign node45372 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node45375 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node45378 = (inp[0]) ? node45382 : node45379;
															assign node45379 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node45382 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node45385 = (inp[5]) ? node45399 : node45386;
													assign node45386 = (inp[2]) ? node45394 : node45387;
														assign node45387 = (inp[3]) ? node45391 : node45388;
															assign node45388 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node45391 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node45394 = (inp[15]) ? 4'b1101 : node45395;
															assign node45395 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node45399 = (inp[2]) ? node45407 : node45400;
														assign node45400 = (inp[15]) ? node45404 : node45401;
															assign node45401 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node45404 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node45407 = (inp[3]) ? node45411 : node45408;
															assign node45408 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node45411 = (inp[0]) ? 4'b1101 : 4'b1111;
										assign node45414 = (inp[8]) ? node45474 : node45415;
											assign node45415 = (inp[2]) ? node45443 : node45416;
												assign node45416 = (inp[14]) ? node45430 : node45417;
													assign node45417 = (inp[15]) ? node45425 : node45418;
														assign node45418 = (inp[0]) ? node45422 : node45419;
															assign node45419 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node45422 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node45425 = (inp[0]) ? node45427 : 4'b0110;
															assign node45427 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node45430 = (inp[5]) ? node45438 : node45431;
														assign node45431 = (inp[3]) ? node45435 : node45432;
															assign node45432 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node45435 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node45438 = (inp[15]) ? node45440 : 4'b1101;
															assign node45440 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node45443 = (inp[14]) ? node45459 : node45444;
													assign node45444 = (inp[3]) ? node45452 : node45445;
														assign node45445 = (inp[0]) ? node45449 : node45446;
															assign node45446 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node45449 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node45452 = (inp[15]) ? node45456 : node45453;
															assign node45453 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node45456 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node45459 = (inp[5]) ? node45467 : node45460;
														assign node45460 = (inp[0]) ? node45464 : node45461;
															assign node45461 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node45464 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node45467 = (inp[0]) ? node45471 : node45468;
															assign node45468 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node45471 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node45474 = (inp[14]) ? node45506 : node45475;
												assign node45475 = (inp[2]) ? node45491 : node45476;
													assign node45476 = (inp[3]) ? node45484 : node45477;
														assign node45477 = (inp[5]) ? node45481 : node45478;
															assign node45478 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node45481 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node45484 = (inp[15]) ? node45488 : node45485;
															assign node45485 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node45488 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node45491 = (inp[3]) ? node45499 : node45492;
														assign node45492 = (inp[5]) ? node45496 : node45493;
															assign node45493 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node45496 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node45499 = (inp[0]) ? node45503 : node45500;
															assign node45500 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node45503 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node45506 = (inp[0]) ? node45518 : node45507;
													assign node45507 = (inp[15]) ? node45513 : node45508;
														assign node45508 = (inp[5]) ? 4'b1100 : node45509;
															assign node45509 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node45513 = (inp[5]) ? 4'b1110 : node45514;
															assign node45514 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node45518 = (inp[15]) ? node45524 : node45519;
														assign node45519 = (inp[5]) ? 4'b1110 : node45520;
															assign node45520 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node45524 = (inp[3]) ? 4'b1100 : node45525;
															assign node45525 = (inp[5]) ? 4'b1100 : 4'b1110;
									assign node45529 = (inp[3]) ? node45653 : node45530;
										assign node45530 = (inp[2]) ? node45592 : node45531;
											assign node45531 = (inp[15]) ? node45563 : node45532;
												assign node45532 = (inp[0]) ? node45548 : node45533;
													assign node45533 = (inp[5]) ? node45541 : node45534;
														assign node45534 = (inp[7]) ? node45538 : node45535;
															assign node45535 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node45538 = (inp[14]) ? 4'b1110 : 4'b1110;
														assign node45541 = (inp[7]) ? node45545 : node45542;
															assign node45542 = (inp[14]) ? 4'b1100 : 4'b1100;
															assign node45545 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node45548 = (inp[5]) ? node45556 : node45549;
														assign node45549 = (inp[14]) ? node45553 : node45550;
															assign node45550 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node45553 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node45556 = (inp[14]) ? node45560 : node45557;
															assign node45557 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node45560 = (inp[7]) ? 4'b1110 : 4'b1110;
												assign node45563 = (inp[5]) ? node45577 : node45564;
													assign node45564 = (inp[0]) ? node45570 : node45565;
														assign node45565 = (inp[7]) ? node45567 : 4'b1100;
															assign node45567 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node45570 = (inp[7]) ? node45574 : node45571;
															assign node45571 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node45574 = (inp[14]) ? 4'b1110 : 4'b1110;
													assign node45577 = (inp[0]) ? node45585 : node45578;
														assign node45578 = (inp[8]) ? node45582 : node45579;
															assign node45579 = (inp[14]) ? 4'b1110 : 4'b1110;
															assign node45582 = (inp[14]) ? 4'b1110 : 4'b1110;
														assign node45585 = (inp[14]) ? node45589 : node45586;
															assign node45586 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node45589 = (inp[8]) ? 4'b1100 : 4'b1100;
											assign node45592 = (inp[0]) ? node45622 : node45593;
												assign node45593 = (inp[15]) ? node45609 : node45594;
													assign node45594 = (inp[5]) ? node45602 : node45595;
														assign node45595 = (inp[7]) ? node45599 : node45596;
															assign node45596 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node45599 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node45602 = (inp[7]) ? node45606 : node45603;
															assign node45603 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node45606 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node45609 = (inp[5]) ? node45617 : node45610;
														assign node45610 = (inp[14]) ? node45614 : node45611;
															assign node45611 = (inp[7]) ? 4'b1100 : 4'b1100;
															assign node45614 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node45617 = (inp[7]) ? 4'b1111 : node45618;
															assign node45618 = (inp[8]) ? 4'b1111 : 4'b1110;
												assign node45622 = (inp[8]) ? node45638 : node45623;
													assign node45623 = (inp[7]) ? node45631 : node45624;
														assign node45624 = (inp[14]) ? node45628 : node45625;
															assign node45625 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node45628 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node45631 = (inp[15]) ? node45635 : node45632;
															assign node45632 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node45635 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node45638 = (inp[7]) ? node45646 : node45639;
														assign node45639 = (inp[5]) ? node45643 : node45640;
															assign node45640 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node45643 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node45646 = (inp[15]) ? node45650 : node45647;
															assign node45647 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node45650 = (inp[5]) ? 4'b1100 : 4'b1110;
										assign node45653 = (inp[5]) ? node45715 : node45654;
											assign node45654 = (inp[7]) ? node45686 : node45655;
												assign node45655 = (inp[8]) ? node45671 : node45656;
													assign node45656 = (inp[2]) ? node45664 : node45657;
														assign node45657 = (inp[14]) ? node45661 : node45658;
															assign node45658 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node45661 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node45664 = (inp[14]) ? node45668 : node45665;
															assign node45665 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node45668 = (inp[0]) ? 4'b1100 : 4'b1100;
													assign node45671 = (inp[2]) ? node45679 : node45672;
														assign node45672 = (inp[14]) ? node45676 : node45673;
															assign node45673 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node45676 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node45679 = (inp[0]) ? node45683 : node45680;
															assign node45680 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node45683 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node45686 = (inp[8]) ? node45700 : node45687;
													assign node45687 = (inp[2]) ? node45693 : node45688;
														assign node45688 = (inp[14]) ? node45690 : 4'b1100;
															assign node45690 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node45693 = (inp[15]) ? node45697 : node45694;
															assign node45694 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node45697 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node45700 = (inp[2]) ? node45708 : node45701;
														assign node45701 = (inp[14]) ? node45705 : node45702;
															assign node45702 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node45705 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node45708 = (inp[0]) ? node45712 : node45709;
															assign node45709 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node45712 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node45715 = (inp[7]) ? node45747 : node45716;
												assign node45716 = (inp[8]) ? node45732 : node45717;
													assign node45717 = (inp[2]) ? node45725 : node45718;
														assign node45718 = (inp[14]) ? node45722 : node45719;
															assign node45719 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node45722 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node45725 = (inp[14]) ? node45729 : node45726;
															assign node45726 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node45729 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node45732 = (inp[2]) ? node45740 : node45733;
														assign node45733 = (inp[14]) ? node45737 : node45734;
															assign node45734 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node45737 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node45740 = (inp[14]) ? node45744 : node45741;
															assign node45741 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node45744 = (inp[0]) ? 4'b1101 : 4'b1101;
												assign node45747 = (inp[8]) ? node45763 : node45748;
													assign node45748 = (inp[14]) ? node45756 : node45749;
														assign node45749 = (inp[2]) ? node45753 : node45750;
															assign node45750 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node45753 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node45756 = (inp[15]) ? node45760 : node45757;
															assign node45757 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node45760 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node45763 = (inp[2]) ? node45771 : node45764;
														assign node45764 = (inp[14]) ? node45768 : node45765;
															assign node45765 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node45768 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node45771 = (inp[0]) ? node45775 : node45772;
															assign node45772 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node45775 = (inp[15]) ? 4'b1100 : 4'b1110;
							assign node45778 = (inp[1]) ? node46218 : node45779;
								assign node45779 = (inp[13]) ? node45997 : node45780;
									assign node45780 = (inp[7]) ? node45884 : node45781;
										assign node45781 = (inp[8]) ? node45833 : node45782;
											assign node45782 = (inp[2]) ? node45810 : node45783;
												assign node45783 = (inp[14]) ? node45799 : node45784;
													assign node45784 = (inp[0]) ? node45792 : node45785;
														assign node45785 = (inp[15]) ? node45789 : node45786;
															assign node45786 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node45789 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node45792 = (inp[15]) ? node45796 : node45793;
															assign node45793 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node45796 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node45799 = (inp[15]) ? node45803 : node45800;
														assign node45800 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node45803 = (inp[0]) ? node45807 : node45804;
															assign node45804 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node45807 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node45810 = (inp[5]) ? node45826 : node45811;
													assign node45811 = (inp[15]) ? node45819 : node45812;
														assign node45812 = (inp[14]) ? node45816 : node45813;
															assign node45813 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node45816 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node45819 = (inp[0]) ? node45823 : node45820;
															assign node45820 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node45823 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node45826 = (inp[0]) ? node45830 : node45827;
														assign node45827 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node45830 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node45833 = (inp[14]) ? node45861 : node45834;
												assign node45834 = (inp[2]) ? node45846 : node45835;
													assign node45835 = (inp[15]) ? node45841 : node45836;
														assign node45836 = (inp[0]) ? node45838 : 4'b1100;
															assign node45838 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node45841 = (inp[0]) ? node45843 : 4'b1110;
															assign node45843 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node45846 = (inp[5]) ? node45854 : node45847;
														assign node45847 = (inp[15]) ? node45851 : node45848;
															assign node45848 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node45851 = (inp[3]) ? 4'b1101 : 4'b1101;
														assign node45854 = (inp[15]) ? node45858 : node45855;
															assign node45855 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node45858 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node45861 = (inp[15]) ? node45873 : node45862;
													assign node45862 = (inp[0]) ? node45868 : node45863;
														assign node45863 = (inp[5]) ? 4'b1101 : node45864;
															assign node45864 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node45868 = (inp[3]) ? 4'b1111 : node45869;
															assign node45869 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node45873 = (inp[0]) ? node45879 : node45874;
														assign node45874 = (inp[5]) ? 4'b1111 : node45875;
															assign node45875 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node45879 = (inp[3]) ? 4'b1101 : node45880;
															assign node45880 = (inp[5]) ? 4'b1101 : 4'b1111;
										assign node45884 = (inp[8]) ? node45938 : node45885;
											assign node45885 = (inp[2]) ? node45915 : node45886;
												assign node45886 = (inp[14]) ? node45902 : node45887;
													assign node45887 = (inp[15]) ? node45895 : node45888;
														assign node45888 = (inp[0]) ? node45892 : node45889;
															assign node45889 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node45892 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node45895 = (inp[0]) ? node45899 : node45896;
															assign node45896 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node45899 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node45902 = (inp[3]) ? node45910 : node45903;
														assign node45903 = (inp[0]) ? node45907 : node45904;
															assign node45904 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node45907 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node45910 = (inp[5]) ? 4'b1111 : node45911;
															assign node45911 = (inp[15]) ? 4'b1101 : 4'b1101;
												assign node45915 = (inp[15]) ? node45927 : node45916;
													assign node45916 = (inp[0]) ? node45922 : node45917;
														assign node45917 = (inp[3]) ? 4'b1101 : node45918;
															assign node45918 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node45922 = (inp[3]) ? 4'b1111 : node45923;
															assign node45923 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node45927 = (inp[0]) ? node45933 : node45928;
														assign node45928 = (inp[3]) ? 4'b1111 : node45929;
															assign node45929 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node45933 = (inp[3]) ? 4'b1101 : node45934;
															assign node45934 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node45938 = (inp[14]) ? node45968 : node45939;
												assign node45939 = (inp[2]) ? node45953 : node45940;
													assign node45940 = (inp[0]) ? node45948 : node45941;
														assign node45941 = (inp[15]) ? node45945 : node45942;
															assign node45942 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node45945 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node45948 = (inp[5]) ? 4'b1111 : node45949;
															assign node45949 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node45953 = (inp[0]) ? node45961 : node45954;
														assign node45954 = (inp[15]) ? node45958 : node45955;
															assign node45955 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node45958 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node45961 = (inp[15]) ? node45965 : node45962;
															assign node45962 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node45965 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node45968 = (inp[2]) ? node45984 : node45969;
													assign node45969 = (inp[15]) ? node45977 : node45970;
														assign node45970 = (inp[0]) ? node45974 : node45971;
															assign node45971 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node45974 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node45977 = (inp[0]) ? node45981 : node45978;
															assign node45978 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node45981 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node45984 = (inp[15]) ? node45990 : node45985;
														assign node45985 = (inp[0]) ? node45987 : 4'b1100;
															assign node45987 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node45990 = (inp[0]) ? node45994 : node45991;
															assign node45991 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node45994 = (inp[5]) ? 4'b1100 : 4'b1100;
									assign node45997 = (inp[8]) ? node46111 : node45998;
										assign node45998 = (inp[7]) ? node46058 : node45999;
											assign node45999 = (inp[2]) ? node46027 : node46000;
												assign node46000 = (inp[14]) ? node46014 : node46001;
													assign node46001 = (inp[3]) ? node46007 : node46002;
														assign node46002 = (inp[5]) ? 4'b1111 : node46003;
															assign node46003 = (inp[0]) ? 4'b1101 : 4'b1101;
														assign node46007 = (inp[0]) ? node46011 : node46008;
															assign node46008 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node46011 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node46014 = (inp[15]) ? node46020 : node46015;
														assign node46015 = (inp[0]) ? node46017 : 4'b1100;
															assign node46017 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node46020 = (inp[0]) ? node46024 : node46021;
															assign node46021 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node46024 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node46027 = (inp[5]) ? node46043 : node46028;
													assign node46028 = (inp[15]) ? node46036 : node46029;
														assign node46029 = (inp[14]) ? node46033 : node46030;
															assign node46030 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node46033 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node46036 = (inp[3]) ? node46040 : node46037;
															assign node46037 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node46040 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node46043 = (inp[14]) ? node46051 : node46044;
														assign node46044 = (inp[0]) ? node46048 : node46045;
															assign node46045 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node46048 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node46051 = (inp[0]) ? node46055 : node46052;
															assign node46052 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node46055 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node46058 = (inp[2]) ? node46088 : node46059;
												assign node46059 = (inp[14]) ? node46073 : node46060;
													assign node46060 = (inp[5]) ? node46066 : node46061;
														assign node46061 = (inp[3]) ? node46063 : 4'b1110;
															assign node46063 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node46066 = (inp[0]) ? node46070 : node46067;
															assign node46067 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node46070 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node46073 = (inp[5]) ? node46081 : node46074;
														assign node46074 = (inp[3]) ? node46078 : node46075;
															assign node46075 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node46078 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node46081 = (inp[15]) ? node46085 : node46082;
															assign node46082 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node46085 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node46088 = (inp[0]) ? node46100 : node46089;
													assign node46089 = (inp[15]) ? node46095 : node46090;
														assign node46090 = (inp[5]) ? 4'b0101 : node46091;
															assign node46091 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node46095 = (inp[5]) ? 4'b0111 : node46096;
															assign node46096 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node46100 = (inp[15]) ? node46106 : node46101;
														assign node46101 = (inp[3]) ? 4'b0111 : node46102;
															assign node46102 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node46106 = (inp[3]) ? 4'b0101 : node46107;
															assign node46107 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node46111 = (inp[7]) ? node46163 : node46112;
											assign node46112 = (inp[14]) ? node46140 : node46113;
												assign node46113 = (inp[2]) ? node46127 : node46114;
													assign node46114 = (inp[15]) ? node46122 : node46115;
														assign node46115 = (inp[0]) ? node46119 : node46116;
															assign node46116 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node46119 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node46122 = (inp[0]) ? node46124 : 4'b1110;
															assign node46124 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node46127 = (inp[0]) ? node46133 : node46128;
														assign node46128 = (inp[15]) ? node46130 : 4'b0101;
															assign node46130 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node46133 = (inp[15]) ? node46137 : node46134;
															assign node46134 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node46137 = (inp[3]) ? 4'b0101 : 4'b0101;
												assign node46140 = (inp[3]) ? node46156 : node46141;
													assign node46141 = (inp[2]) ? node46149 : node46142;
														assign node46142 = (inp[5]) ? node46146 : node46143;
															assign node46143 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node46146 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node46149 = (inp[5]) ? node46153 : node46150;
															assign node46150 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node46153 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node46156 = (inp[0]) ? node46160 : node46157;
														assign node46157 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node46160 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node46163 = (inp[14]) ? node46195 : node46164;
												assign node46164 = (inp[2]) ? node46180 : node46165;
													assign node46165 = (inp[5]) ? node46173 : node46166;
														assign node46166 = (inp[15]) ? node46170 : node46167;
															assign node46167 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node46170 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node46173 = (inp[15]) ? node46177 : node46174;
															assign node46174 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node46177 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node46180 = (inp[3]) ? node46188 : node46181;
														assign node46181 = (inp[0]) ? node46185 : node46182;
															assign node46182 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node46185 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node46188 = (inp[5]) ? node46192 : node46189;
															assign node46189 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node46192 = (inp[15]) ? 4'b0100 : 4'b0100;
												assign node46195 = (inp[5]) ? node46211 : node46196;
													assign node46196 = (inp[15]) ? node46204 : node46197;
														assign node46197 = (inp[0]) ? node46201 : node46198;
															assign node46198 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node46201 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node46204 = (inp[3]) ? node46208 : node46205;
															assign node46205 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node46208 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node46211 = (inp[15]) ? node46215 : node46212;
														assign node46212 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node46215 = (inp[0]) ? 4'b0100 : 4'b0110;
								assign node46218 = (inp[13]) ? node46444 : node46219;
									assign node46219 = (inp[8]) ? node46331 : node46220;
										assign node46220 = (inp[7]) ? node46276 : node46221;
											assign node46221 = (inp[14]) ? node46249 : node46222;
												assign node46222 = (inp[2]) ? node46234 : node46223;
													assign node46223 = (inp[0]) ? node46229 : node46224;
														assign node46224 = (inp[15]) ? 4'b1111 : node46225;
															assign node46225 = (inp[5]) ? 4'b1101 : 4'b1101;
														assign node46229 = (inp[15]) ? 4'b1101 : node46230;
															assign node46230 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node46234 = (inp[5]) ? node46242 : node46235;
														assign node46235 = (inp[15]) ? node46239 : node46236;
															assign node46236 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node46239 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node46242 = (inp[3]) ? node46246 : node46243;
															assign node46243 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node46246 = (inp[15]) ? 4'b1100 : 4'b1100;
												assign node46249 = (inp[2]) ? node46265 : node46250;
													assign node46250 = (inp[5]) ? node46258 : node46251;
														assign node46251 = (inp[15]) ? node46255 : node46252;
															assign node46252 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node46255 = (inp[3]) ? 4'b1100 : 4'b1100;
														assign node46258 = (inp[3]) ? node46262 : node46259;
															assign node46259 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node46262 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node46265 = (inp[15]) ? node46271 : node46266;
														assign node46266 = (inp[5]) ? 4'b1110 : node46267;
															assign node46267 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node46271 = (inp[0]) ? 4'b1100 : node46272;
															assign node46272 = (inp[5]) ? 4'b1110 : 4'b1100;
											assign node46276 = (inp[2]) ? node46308 : node46277;
												assign node46277 = (inp[14]) ? node46293 : node46278;
													assign node46278 = (inp[5]) ? node46286 : node46279;
														assign node46279 = (inp[0]) ? node46283 : node46280;
															assign node46280 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node46283 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node46286 = (inp[0]) ? node46290 : node46287;
															assign node46287 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node46290 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node46293 = (inp[5]) ? node46301 : node46294;
														assign node46294 = (inp[15]) ? node46298 : node46295;
															assign node46295 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node46298 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node46301 = (inp[0]) ? node46305 : node46302;
															assign node46302 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node46305 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node46308 = (inp[0]) ? node46320 : node46309;
													assign node46309 = (inp[15]) ? node46315 : node46310;
														assign node46310 = (inp[5]) ? 4'b0101 : node46311;
															assign node46311 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node46315 = (inp[5]) ? 4'b0111 : node46316;
															assign node46316 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node46320 = (inp[15]) ? node46326 : node46321;
														assign node46321 = (inp[3]) ? 4'b0111 : node46322;
															assign node46322 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node46326 = (inp[3]) ? 4'b0101 : node46327;
															assign node46327 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node46331 = (inp[7]) ? node46389 : node46332;
											assign node46332 = (inp[14]) ? node46360 : node46333;
												assign node46333 = (inp[2]) ? node46345 : node46334;
													assign node46334 = (inp[0]) ? node46340 : node46335;
														assign node46335 = (inp[15]) ? node46337 : 4'b1100;
															assign node46337 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node46340 = (inp[15]) ? node46342 : 4'b1110;
															assign node46342 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node46345 = (inp[0]) ? node46353 : node46346;
														assign node46346 = (inp[15]) ? node46350 : node46347;
															assign node46347 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node46350 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node46353 = (inp[15]) ? node46357 : node46354;
															assign node46354 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node46357 = (inp[3]) ? 4'b0101 : 4'b0101;
												assign node46360 = (inp[2]) ? node46376 : node46361;
													assign node46361 = (inp[3]) ? node46369 : node46362;
														assign node46362 = (inp[15]) ? node46366 : node46363;
															assign node46363 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node46366 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node46369 = (inp[0]) ? node46373 : node46370;
															assign node46370 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node46373 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node46376 = (inp[5]) ? node46384 : node46377;
														assign node46377 = (inp[0]) ? node46381 : node46378;
															assign node46378 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node46381 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node46384 = (inp[3]) ? 4'b0111 : node46385;
															assign node46385 = (inp[0]) ? 4'b0101 : 4'b0101;
											assign node46389 = (inp[14]) ? node46421 : node46390;
												assign node46390 = (inp[2]) ? node46406 : node46391;
													assign node46391 = (inp[0]) ? node46399 : node46392;
														assign node46392 = (inp[15]) ? node46396 : node46393;
															assign node46393 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node46396 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node46399 = (inp[15]) ? node46403 : node46400;
															assign node46400 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node46403 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node46406 = (inp[15]) ? node46414 : node46407;
														assign node46407 = (inp[0]) ? node46411 : node46408;
															assign node46408 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node46411 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node46414 = (inp[0]) ? node46418 : node46415;
															assign node46415 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node46418 = (inp[3]) ? 4'b0100 : 4'b0100;
												assign node46421 = (inp[5]) ? node46437 : node46422;
													assign node46422 = (inp[15]) ? node46430 : node46423;
														assign node46423 = (inp[3]) ? node46427 : node46424;
															assign node46424 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node46427 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node46430 = (inp[0]) ? node46434 : node46431;
															assign node46431 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node46434 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node46437 = (inp[0]) ? node46441 : node46438;
														assign node46438 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node46441 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node46444 = (inp[5]) ? node46564 : node46445;
										assign node46445 = (inp[7]) ? node46505 : node46446;
											assign node46446 = (inp[8]) ? node46478 : node46447;
												assign node46447 = (inp[14]) ? node46463 : node46448;
													assign node46448 = (inp[2]) ? node46456 : node46449;
														assign node46449 = (inp[0]) ? node46453 : node46450;
															assign node46450 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node46453 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node46456 = (inp[15]) ? node46460 : node46457;
															assign node46457 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node46460 = (inp[3]) ? 4'b0100 : 4'b0100;
													assign node46463 = (inp[15]) ? node46471 : node46464;
														assign node46464 = (inp[0]) ? node46468 : node46465;
															assign node46465 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node46468 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node46471 = (inp[0]) ? node46475 : node46472;
															assign node46472 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node46475 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node46478 = (inp[14]) ? node46492 : node46479;
													assign node46479 = (inp[2]) ? node46487 : node46480;
														assign node46480 = (inp[0]) ? node46484 : node46481;
															assign node46481 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node46484 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node46487 = (inp[3]) ? node46489 : 4'b0111;
															assign node46489 = (inp[0]) ? 4'b0101 : 4'b0101;
													assign node46492 = (inp[0]) ? node46498 : node46493;
														assign node46493 = (inp[2]) ? node46495 : 4'b0111;
															assign node46495 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node46498 = (inp[15]) ? node46502 : node46499;
															assign node46499 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node46502 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node46505 = (inp[8]) ? node46535 : node46506;
												assign node46506 = (inp[14]) ? node46520 : node46507;
													assign node46507 = (inp[2]) ? node46515 : node46508;
														assign node46508 = (inp[0]) ? node46512 : node46509;
															assign node46509 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node46512 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node46515 = (inp[15]) ? node46517 : 4'b0101;
															assign node46517 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node46520 = (inp[15]) ? node46528 : node46521;
														assign node46521 = (inp[3]) ? node46525 : node46522;
															assign node46522 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node46525 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node46528 = (inp[2]) ? node46532 : node46529;
															assign node46529 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node46532 = (inp[3]) ? 4'b0101 : 4'b0101;
												assign node46535 = (inp[2]) ? node46549 : node46536;
													assign node46536 = (inp[14]) ? node46544 : node46537;
														assign node46537 = (inp[15]) ? node46541 : node46538;
															assign node46538 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node46541 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node46544 = (inp[3]) ? node46546 : 4'b0110;
															assign node46546 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node46549 = (inp[15]) ? node46557 : node46550;
														assign node46550 = (inp[3]) ? node46554 : node46551;
															assign node46551 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node46554 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node46557 = (inp[0]) ? node46561 : node46558;
															assign node46558 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node46561 = (inp[3]) ? 4'b0100 : 4'b0110;
										assign node46564 = (inp[2]) ? node46628 : node46565;
											assign node46565 = (inp[8]) ? node46597 : node46566;
												assign node46566 = (inp[14]) ? node46582 : node46567;
													assign node46567 = (inp[7]) ? node46575 : node46568;
														assign node46568 = (inp[15]) ? node46572 : node46569;
															assign node46569 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node46572 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node46575 = (inp[3]) ? node46579 : node46576;
															assign node46576 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node46579 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node46582 = (inp[7]) ? node46590 : node46583;
														assign node46583 = (inp[3]) ? node46587 : node46584;
															assign node46584 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node46587 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node46590 = (inp[15]) ? node46594 : node46591;
															assign node46591 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node46594 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node46597 = (inp[15]) ? node46613 : node46598;
													assign node46598 = (inp[0]) ? node46606 : node46599;
														assign node46599 = (inp[7]) ? node46603 : node46600;
															assign node46600 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node46603 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node46606 = (inp[14]) ? node46610 : node46607;
															assign node46607 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node46610 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node46613 = (inp[0]) ? node46621 : node46614;
														assign node46614 = (inp[7]) ? node46618 : node46615;
															assign node46615 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node46618 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node46621 = (inp[3]) ? node46625 : node46622;
															assign node46622 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node46625 = (inp[7]) ? 4'b0100 : 4'b0100;
											assign node46628 = (inp[3]) ? node46660 : node46629;
												assign node46629 = (inp[0]) ? node46645 : node46630;
													assign node46630 = (inp[15]) ? node46638 : node46631;
														assign node46631 = (inp[14]) ? node46635 : node46632;
															assign node46632 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node46635 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node46638 = (inp[14]) ? node46642 : node46639;
															assign node46639 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node46642 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node46645 = (inp[15]) ? node46653 : node46646;
														assign node46646 = (inp[8]) ? node46650 : node46647;
															assign node46647 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node46650 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node46653 = (inp[7]) ? node46657 : node46654;
															assign node46654 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node46657 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node46660 = (inp[15]) ? node46676 : node46661;
													assign node46661 = (inp[0]) ? node46669 : node46662;
														assign node46662 = (inp[8]) ? node46666 : node46663;
															assign node46663 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node46666 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node46669 = (inp[8]) ? node46673 : node46670;
															assign node46670 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node46673 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node46676 = (inp[0]) ? node46684 : node46677;
														assign node46677 = (inp[14]) ? node46681 : node46678;
															assign node46678 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node46681 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node46684 = (inp[8]) ? node46688 : node46685;
															assign node46685 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node46688 = (inp[7]) ? 4'b0100 : 4'b0101;
					assign node46691 = (inp[6]) ? node48475 : node46692;
						assign node46692 = (inp[11]) ? node47574 : node46693;
							assign node46693 = (inp[1]) ? node47127 : node46694;
								assign node46694 = (inp[13]) ? node46908 : node46695;
									assign node46695 = (inp[7]) ? node46803 : node46696;
										assign node46696 = (inp[8]) ? node46752 : node46697;
											assign node46697 = (inp[14]) ? node46723 : node46698;
												assign node46698 = (inp[2]) ? node46710 : node46699;
													assign node46699 = (inp[15]) ? node46705 : node46700;
														assign node46700 = (inp[0]) ? node46702 : 4'b1101;
															assign node46702 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node46705 = (inp[0]) ? node46707 : 4'b1111;
															assign node46707 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node46710 = (inp[3]) ? node46718 : node46711;
														assign node46711 = (inp[0]) ? node46715 : node46712;
															assign node46712 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node46715 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node46718 = (inp[5]) ? 4'b1100 : node46719;
															assign node46719 = (inp[0]) ? 4'b1100 : 4'b1100;
												assign node46723 = (inp[3]) ? node46739 : node46724;
													assign node46724 = (inp[5]) ? node46732 : node46725;
														assign node46725 = (inp[2]) ? node46729 : node46726;
															assign node46726 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node46729 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node46732 = (inp[0]) ? node46736 : node46733;
															assign node46733 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node46736 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node46739 = (inp[5]) ? node46745 : node46740;
														assign node46740 = (inp[15]) ? node46742 : 4'b1100;
															assign node46742 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node46745 = (inp[15]) ? node46749 : node46746;
															assign node46746 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node46749 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node46752 = (inp[14]) ? node46780 : node46753;
												assign node46753 = (inp[2]) ? node46765 : node46754;
													assign node46754 = (inp[5]) ? node46760 : node46755;
														assign node46755 = (inp[15]) ? node46757 : 4'b1110;
															assign node46757 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node46760 = (inp[3]) ? node46762 : 4'b1100;
															assign node46762 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node46765 = (inp[5]) ? node46773 : node46766;
														assign node46766 = (inp[0]) ? node46770 : node46767;
															assign node46767 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node46770 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node46773 = (inp[0]) ? node46777 : node46774;
															assign node46774 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node46777 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node46780 = (inp[0]) ? node46792 : node46781;
													assign node46781 = (inp[15]) ? node46787 : node46782;
														assign node46782 = (inp[5]) ? 4'b1101 : node46783;
															assign node46783 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node46787 = (inp[3]) ? 4'b1111 : node46788;
															assign node46788 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node46792 = (inp[15]) ? node46798 : node46793;
														assign node46793 = (inp[5]) ? 4'b1111 : node46794;
															assign node46794 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node46798 = (inp[3]) ? 4'b1101 : node46799;
															assign node46799 = (inp[5]) ? 4'b1101 : 4'b1111;
										assign node46803 = (inp[8]) ? node46855 : node46804;
											assign node46804 = (inp[14]) ? node46834 : node46805;
												assign node46805 = (inp[2]) ? node46821 : node46806;
													assign node46806 = (inp[15]) ? node46814 : node46807;
														assign node46807 = (inp[0]) ? node46811 : node46808;
															assign node46808 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node46811 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node46814 = (inp[0]) ? node46818 : node46815;
															assign node46815 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node46818 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node46821 = (inp[15]) ? node46829 : node46822;
														assign node46822 = (inp[0]) ? node46826 : node46823;
															assign node46823 = (inp[3]) ? 4'b1101 : 4'b1101;
															assign node46826 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node46829 = (inp[0]) ? 4'b1101 : node46830;
															assign node46830 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node46834 = (inp[15]) ? node46846 : node46835;
													assign node46835 = (inp[0]) ? node46841 : node46836;
														assign node46836 = (inp[3]) ? 4'b1101 : node46837;
															assign node46837 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node46841 = (inp[5]) ? 4'b1111 : node46842;
															assign node46842 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node46846 = (inp[0]) ? node46852 : node46847;
														assign node46847 = (inp[3]) ? 4'b1111 : node46848;
															assign node46848 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node46852 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node46855 = (inp[14]) ? node46885 : node46856;
												assign node46856 = (inp[2]) ? node46872 : node46857;
													assign node46857 = (inp[3]) ? node46865 : node46858;
														assign node46858 = (inp[5]) ? node46862 : node46859;
															assign node46859 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node46862 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node46865 = (inp[5]) ? node46869 : node46866;
															assign node46866 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node46869 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node46872 = (inp[15]) ? node46878 : node46873;
														assign node46873 = (inp[0]) ? node46875 : 4'b1100;
															assign node46875 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node46878 = (inp[0]) ? node46882 : node46879;
															assign node46879 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node46882 = (inp[5]) ? 4'b1100 : 4'b1100;
												assign node46885 = (inp[5]) ? node46901 : node46886;
													assign node46886 = (inp[0]) ? node46894 : node46887;
														assign node46887 = (inp[2]) ? node46891 : node46888;
															assign node46888 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node46891 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node46894 = (inp[2]) ? node46898 : node46895;
															assign node46895 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node46898 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node46901 = (inp[0]) ? node46905 : node46902;
														assign node46902 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node46905 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node46908 = (inp[8]) ? node47024 : node46909;
										assign node46909 = (inp[7]) ? node46963 : node46910;
											assign node46910 = (inp[14]) ? node46940 : node46911;
												assign node46911 = (inp[2]) ? node46927 : node46912;
													assign node46912 = (inp[3]) ? node46920 : node46913;
														assign node46913 = (inp[5]) ? node46917 : node46914;
															assign node46914 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node46917 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node46920 = (inp[5]) ? node46924 : node46921;
															assign node46921 = (inp[15]) ? 4'b1101 : 4'b1101;
															assign node46924 = (inp[0]) ? 4'b1101 : 4'b1101;
													assign node46927 = (inp[3]) ? node46933 : node46928;
														assign node46928 = (inp[0]) ? node46930 : 4'b1110;
															assign node46930 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node46933 = (inp[15]) ? node46937 : node46934;
															assign node46934 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node46937 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node46940 = (inp[5]) ? node46956 : node46941;
													assign node46941 = (inp[15]) ? node46949 : node46942;
														assign node46942 = (inp[2]) ? node46946 : node46943;
															assign node46943 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node46946 = (inp[0]) ? 4'b1100 : 4'b1100;
														assign node46949 = (inp[2]) ? node46953 : node46950;
															assign node46950 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node46953 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node46956 = (inp[15]) ? node46960 : node46957;
														assign node46957 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node46960 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node46963 = (inp[2]) ? node46993 : node46964;
												assign node46964 = (inp[14]) ? node46980 : node46965;
													assign node46965 = (inp[15]) ? node46973 : node46966;
														assign node46966 = (inp[0]) ? node46970 : node46967;
															assign node46967 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node46970 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node46973 = (inp[0]) ? node46977 : node46974;
															assign node46974 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node46977 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node46980 = (inp[15]) ? node46986 : node46981;
														assign node46981 = (inp[5]) ? 4'b0111 : node46982;
															assign node46982 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node46986 = (inp[0]) ? node46990 : node46987;
															assign node46987 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node46990 = (inp[5]) ? 4'b0101 : 4'b0101;
												assign node46993 = (inp[14]) ? node47009 : node46994;
													assign node46994 = (inp[0]) ? node47002 : node46995;
														assign node46995 = (inp[15]) ? node46999 : node46996;
															assign node46996 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node46999 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node47002 = (inp[15]) ? node47006 : node47003;
															assign node47003 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node47006 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node47009 = (inp[3]) ? node47017 : node47010;
														assign node47010 = (inp[5]) ? node47014 : node47011;
															assign node47011 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node47014 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node47017 = (inp[15]) ? node47021 : node47018;
															assign node47018 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node47021 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node47024 = (inp[7]) ? node47076 : node47025;
											assign node47025 = (inp[14]) ? node47053 : node47026;
												assign node47026 = (inp[2]) ? node47040 : node47027;
													assign node47027 = (inp[15]) ? node47033 : node47028;
														assign node47028 = (inp[0]) ? node47030 : 4'b1100;
															assign node47030 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node47033 = (inp[0]) ? node47037 : node47034;
															assign node47034 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node47037 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node47040 = (inp[5]) ? node47048 : node47041;
														assign node47041 = (inp[0]) ? node47045 : node47042;
															assign node47042 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node47045 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node47048 = (inp[3]) ? 4'b0111 : node47049;
															assign node47049 = (inp[15]) ? 4'b0101 : 4'b0101;
												assign node47053 = (inp[0]) ? node47065 : node47054;
													assign node47054 = (inp[15]) ? node47060 : node47055;
														assign node47055 = (inp[5]) ? 4'b0101 : node47056;
															assign node47056 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node47060 = (inp[3]) ? 4'b0111 : node47061;
															assign node47061 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node47065 = (inp[15]) ? node47071 : node47066;
														assign node47066 = (inp[3]) ? 4'b0111 : node47067;
															assign node47067 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node47071 = (inp[5]) ? 4'b0101 : node47072;
															assign node47072 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node47076 = (inp[2]) ? node47104 : node47077;
												assign node47077 = (inp[14]) ? node47093 : node47078;
													assign node47078 = (inp[5]) ? node47086 : node47079;
														assign node47079 = (inp[15]) ? node47083 : node47080;
															assign node47080 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node47083 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node47086 = (inp[15]) ? node47090 : node47087;
															assign node47087 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node47090 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node47093 = (inp[0]) ? node47101 : node47094;
														assign node47094 = (inp[15]) ? node47098 : node47095;
															assign node47095 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node47098 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node47101 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node47104 = (inp[3]) ? node47120 : node47105;
													assign node47105 = (inp[0]) ? node47113 : node47106;
														assign node47106 = (inp[15]) ? node47110 : node47107;
															assign node47107 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node47110 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node47113 = (inp[15]) ? node47117 : node47114;
															assign node47114 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node47117 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node47120 = (inp[15]) ? node47124 : node47121;
														assign node47121 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node47124 = (inp[0]) ? 4'b0100 : 4'b0110;
								assign node47127 = (inp[13]) ? node47349 : node47128;
									assign node47128 = (inp[8]) ? node47246 : node47129;
										assign node47129 = (inp[7]) ? node47183 : node47130;
											assign node47130 = (inp[14]) ? node47160 : node47131;
												assign node47131 = (inp[2]) ? node47147 : node47132;
													assign node47132 = (inp[3]) ? node47140 : node47133;
														assign node47133 = (inp[5]) ? node47137 : node47134;
															assign node47134 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node47137 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node47140 = (inp[5]) ? node47144 : node47141;
															assign node47141 = (inp[0]) ? 4'b1101 : 4'b1101;
															assign node47144 = (inp[0]) ? 4'b1101 : 4'b1101;
													assign node47147 = (inp[0]) ? node47155 : node47148;
														assign node47148 = (inp[15]) ? node47152 : node47149;
															assign node47149 = (inp[3]) ? 4'b1100 : 4'b1100;
															assign node47152 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node47155 = (inp[15]) ? node47157 : 4'b1110;
															assign node47157 = (inp[3]) ? 4'b1100 : 4'b1100;
												assign node47160 = (inp[15]) ? node47172 : node47161;
													assign node47161 = (inp[0]) ? node47167 : node47162;
														assign node47162 = (inp[3]) ? 4'b1100 : node47163;
															assign node47163 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node47167 = (inp[5]) ? 4'b1110 : node47168;
															assign node47168 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node47172 = (inp[0]) ? node47178 : node47173;
														assign node47173 = (inp[5]) ? 4'b1110 : node47174;
															assign node47174 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node47178 = (inp[3]) ? 4'b1100 : node47179;
															assign node47179 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node47183 = (inp[14]) ? node47215 : node47184;
												assign node47184 = (inp[2]) ? node47200 : node47185;
													assign node47185 = (inp[3]) ? node47193 : node47186;
														assign node47186 = (inp[15]) ? node47190 : node47187;
															assign node47187 = (inp[0]) ? 4'b1100 : 4'b1100;
															assign node47190 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node47193 = (inp[5]) ? node47197 : node47194;
															assign node47194 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node47197 = (inp[15]) ? 4'b1100 : 4'b1100;
													assign node47200 = (inp[15]) ? node47208 : node47201;
														assign node47201 = (inp[0]) ? node47205 : node47202;
															assign node47202 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node47205 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node47208 = (inp[0]) ? node47212 : node47209;
															assign node47209 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node47212 = (inp[3]) ? 4'b0101 : 4'b0101;
												assign node47215 = (inp[3]) ? node47231 : node47216;
													assign node47216 = (inp[2]) ? node47224 : node47217;
														assign node47217 = (inp[0]) ? node47221 : node47218;
															assign node47218 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node47221 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node47224 = (inp[15]) ? node47228 : node47225;
															assign node47225 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node47228 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node47231 = (inp[5]) ? node47239 : node47232;
														assign node47232 = (inp[15]) ? node47236 : node47233;
															assign node47233 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node47236 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node47239 = (inp[0]) ? node47243 : node47240;
															assign node47240 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node47243 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node47246 = (inp[7]) ? node47300 : node47247;
											assign node47247 = (inp[2]) ? node47277 : node47248;
												assign node47248 = (inp[14]) ? node47262 : node47249;
													assign node47249 = (inp[0]) ? node47255 : node47250;
														assign node47250 = (inp[3]) ? 4'b1100 : node47251;
															assign node47251 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node47255 = (inp[15]) ? node47259 : node47256;
															assign node47256 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node47259 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node47262 = (inp[3]) ? node47270 : node47263;
														assign node47263 = (inp[0]) ? node47267 : node47264;
															assign node47264 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node47267 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node47270 = (inp[0]) ? node47274 : node47271;
															assign node47271 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node47274 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node47277 = (inp[15]) ? node47289 : node47278;
													assign node47278 = (inp[0]) ? node47284 : node47279;
														assign node47279 = (inp[3]) ? 4'b0101 : node47280;
															assign node47280 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node47284 = (inp[3]) ? 4'b0111 : node47285;
															assign node47285 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node47289 = (inp[0]) ? node47295 : node47290;
														assign node47290 = (inp[3]) ? 4'b0111 : node47291;
															assign node47291 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node47295 = (inp[5]) ? 4'b0101 : node47296;
															assign node47296 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node47300 = (inp[2]) ? node47330 : node47301;
												assign node47301 = (inp[14]) ? node47315 : node47302;
													assign node47302 = (inp[15]) ? node47308 : node47303;
														assign node47303 = (inp[0]) ? 4'b0111 : node47304;
															assign node47304 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node47308 = (inp[0]) ? node47312 : node47309;
															assign node47309 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node47312 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node47315 = (inp[3]) ? node47323 : node47316;
														assign node47316 = (inp[0]) ? node47320 : node47317;
															assign node47317 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node47320 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node47323 = (inp[0]) ? node47327 : node47324;
															assign node47324 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node47327 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node47330 = (inp[0]) ? node47342 : node47331;
													assign node47331 = (inp[15]) ? node47337 : node47332;
														assign node47332 = (inp[5]) ? 4'b0100 : node47333;
															assign node47333 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node47337 = (inp[3]) ? 4'b0110 : node47338;
															assign node47338 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node47342 = (inp[15]) ? node47344 : 4'b0110;
														assign node47344 = (inp[3]) ? 4'b0100 : node47345;
															assign node47345 = (inp[5]) ? 4'b0100 : 4'b0110;
									assign node47349 = (inp[0]) ? node47463 : node47350;
										assign node47350 = (inp[15]) ? node47402 : node47351;
											assign node47351 = (inp[3]) ? node47379 : node47352;
												assign node47352 = (inp[5]) ? node47368 : node47353;
													assign node47353 = (inp[2]) ? node47361 : node47354;
														assign node47354 = (inp[8]) ? node47358 : node47355;
															assign node47355 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node47358 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node47361 = (inp[8]) ? node47365 : node47362;
															assign node47362 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node47365 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node47368 = (inp[8]) ? node47374 : node47369;
														assign node47369 = (inp[7]) ? node47371 : 4'b0100;
															assign node47371 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node47374 = (inp[7]) ? node47376 : 4'b0101;
															assign node47376 = (inp[2]) ? 4'b0100 : 4'b0100;
												assign node47379 = (inp[8]) ? node47391 : node47380;
													assign node47380 = (inp[7]) ? node47386 : node47381;
														assign node47381 = (inp[14]) ? 4'b0100 : node47382;
															assign node47382 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node47386 = (inp[14]) ? 4'b0101 : node47387;
															assign node47387 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node47391 = (inp[7]) ? node47397 : node47392;
														assign node47392 = (inp[2]) ? 4'b0101 : node47393;
															assign node47393 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node47397 = (inp[2]) ? 4'b0100 : node47398;
															assign node47398 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node47402 = (inp[5]) ? node47434 : node47403;
												assign node47403 = (inp[3]) ? node47419 : node47404;
													assign node47404 = (inp[7]) ? node47412 : node47405;
														assign node47405 = (inp[8]) ? node47409 : node47406;
															assign node47406 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node47409 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node47412 = (inp[8]) ? node47416 : node47413;
															assign node47413 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node47416 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node47419 = (inp[2]) ? node47427 : node47420;
														assign node47420 = (inp[7]) ? node47424 : node47421;
															assign node47421 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node47424 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node47427 = (inp[8]) ? node47431 : node47428;
															assign node47428 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node47431 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node47434 = (inp[14]) ? node47448 : node47435;
													assign node47435 = (inp[8]) ? node47441 : node47436;
														assign node47436 = (inp[3]) ? 4'b0110 : node47437;
															assign node47437 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node47441 = (inp[7]) ? node47445 : node47442;
															assign node47442 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node47445 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node47448 = (inp[2]) ? node47456 : node47449;
														assign node47449 = (inp[3]) ? node47453 : node47450;
															assign node47450 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node47453 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node47456 = (inp[8]) ? node47460 : node47457;
															assign node47457 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node47460 = (inp[7]) ? 4'b0110 : 4'b0111;
										assign node47463 = (inp[15]) ? node47519 : node47464;
											assign node47464 = (inp[5]) ? node47496 : node47465;
												assign node47465 = (inp[3]) ? node47481 : node47466;
													assign node47466 = (inp[8]) ? node47474 : node47467;
														assign node47467 = (inp[7]) ? node47471 : node47468;
															assign node47468 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node47471 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node47474 = (inp[7]) ? node47478 : node47475;
															assign node47475 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node47478 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node47481 = (inp[2]) ? node47489 : node47482;
														assign node47482 = (inp[8]) ? node47486 : node47483;
															assign node47483 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node47486 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node47489 = (inp[7]) ? node47493 : node47490;
															assign node47490 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node47493 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node47496 = (inp[2]) ? node47512 : node47497;
													assign node47497 = (inp[3]) ? node47505 : node47498;
														assign node47498 = (inp[14]) ? node47502 : node47499;
															assign node47499 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node47502 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node47505 = (inp[14]) ? node47509 : node47506;
															assign node47506 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node47509 = (inp[7]) ? 4'b0110 : 4'b0110;
													assign node47512 = (inp[8]) ? node47516 : node47513;
														assign node47513 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node47516 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node47519 = (inp[5]) ? node47551 : node47520;
												assign node47520 = (inp[3]) ? node47536 : node47521;
													assign node47521 = (inp[2]) ? node47529 : node47522;
														assign node47522 = (inp[7]) ? node47526 : node47523;
															assign node47523 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node47526 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node47529 = (inp[7]) ? node47533 : node47530;
															assign node47530 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node47533 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node47536 = (inp[2]) ? node47544 : node47537;
														assign node47537 = (inp[7]) ? node47541 : node47538;
															assign node47538 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node47541 = (inp[14]) ? 4'b0100 : 4'b0100;
														assign node47544 = (inp[8]) ? node47548 : node47545;
															assign node47545 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node47548 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node47551 = (inp[2]) ? node47567 : node47552;
													assign node47552 = (inp[7]) ? node47560 : node47553;
														assign node47553 = (inp[8]) ? node47557 : node47554;
															assign node47554 = (inp[14]) ? 4'b0100 : 4'b0101;
															assign node47557 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node47560 = (inp[3]) ? node47564 : node47561;
															assign node47561 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node47564 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node47567 = (inp[7]) ? node47571 : node47568;
														assign node47568 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node47571 = (inp[8]) ? 4'b0100 : 4'b0101;
							assign node47574 = (inp[13]) ? node48028 : node47575;
								assign node47575 = (inp[1]) ? node47799 : node47576;
									assign node47576 = (inp[8]) ? node47690 : node47577;
										assign node47577 = (inp[7]) ? node47629 : node47578;
											assign node47578 = (inp[14]) ? node47606 : node47579;
												assign node47579 = (inp[2]) ? node47593 : node47580;
													assign node47580 = (inp[3]) ? node47586 : node47581;
														assign node47581 = (inp[15]) ? 4'b0101 : node47582;
															assign node47582 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node47586 = (inp[15]) ? node47590 : node47587;
															assign node47587 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node47590 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node47593 = (inp[5]) ? node47601 : node47594;
														assign node47594 = (inp[0]) ? node47598 : node47595;
															assign node47595 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node47598 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node47601 = (inp[0]) ? node47603 : 4'b0100;
															assign node47603 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node47606 = (inp[0]) ? node47618 : node47607;
													assign node47607 = (inp[15]) ? node47613 : node47608;
														assign node47608 = (inp[5]) ? 4'b0100 : node47609;
															assign node47609 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node47613 = (inp[3]) ? 4'b0110 : node47614;
															assign node47614 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node47618 = (inp[15]) ? node47624 : node47619;
														assign node47619 = (inp[3]) ? 4'b0110 : node47620;
															assign node47620 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node47624 = (inp[5]) ? 4'b0100 : node47625;
															assign node47625 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node47629 = (inp[2]) ? node47659 : node47630;
												assign node47630 = (inp[14]) ? node47646 : node47631;
													assign node47631 = (inp[3]) ? node47639 : node47632;
														assign node47632 = (inp[15]) ? node47636 : node47633;
															assign node47633 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node47636 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node47639 = (inp[15]) ? node47643 : node47640;
															assign node47640 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node47643 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node47646 = (inp[0]) ? node47654 : node47647;
														assign node47647 = (inp[15]) ? node47651 : node47648;
															assign node47648 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node47651 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node47654 = (inp[15]) ? 4'b0101 : node47655;
															assign node47655 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node47659 = (inp[3]) ? node47675 : node47660;
													assign node47660 = (inp[15]) ? node47668 : node47661;
														assign node47661 = (inp[14]) ? node47665 : node47662;
															assign node47662 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node47665 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node47668 = (inp[0]) ? node47672 : node47669;
															assign node47669 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node47672 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node47675 = (inp[14]) ? node47683 : node47676;
														assign node47676 = (inp[15]) ? node47680 : node47677;
															assign node47677 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node47680 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node47683 = (inp[0]) ? node47687 : node47684;
															assign node47684 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node47687 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node47690 = (inp[7]) ? node47746 : node47691;
											assign node47691 = (inp[14]) ? node47723 : node47692;
												assign node47692 = (inp[2]) ? node47708 : node47693;
													assign node47693 = (inp[3]) ? node47701 : node47694;
														assign node47694 = (inp[5]) ? node47698 : node47695;
															assign node47695 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node47698 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node47701 = (inp[0]) ? node47705 : node47702;
															assign node47702 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node47705 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node47708 = (inp[5]) ? node47716 : node47709;
														assign node47709 = (inp[15]) ? node47713 : node47710;
															assign node47710 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node47713 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node47716 = (inp[0]) ? node47720 : node47717;
															assign node47717 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node47720 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node47723 = (inp[15]) ? node47735 : node47724;
													assign node47724 = (inp[0]) ? node47730 : node47725;
														assign node47725 = (inp[3]) ? 4'b0101 : node47726;
															assign node47726 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node47730 = (inp[3]) ? 4'b0111 : node47731;
															assign node47731 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node47735 = (inp[0]) ? node47741 : node47736;
														assign node47736 = (inp[3]) ? 4'b0111 : node47737;
															assign node47737 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node47741 = (inp[5]) ? 4'b0101 : node47742;
															assign node47742 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node47746 = (inp[14]) ? node47776 : node47747;
												assign node47747 = (inp[2]) ? node47761 : node47748;
													assign node47748 = (inp[0]) ? node47756 : node47749;
														assign node47749 = (inp[15]) ? node47753 : node47750;
															assign node47750 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node47753 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node47756 = (inp[15]) ? 4'b0101 : node47757;
															assign node47757 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node47761 = (inp[15]) ? node47769 : node47762;
														assign node47762 = (inp[0]) ? node47766 : node47763;
															assign node47763 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node47766 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node47769 = (inp[0]) ? node47773 : node47770;
															assign node47770 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node47773 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node47776 = (inp[5]) ? node47792 : node47777;
													assign node47777 = (inp[2]) ? node47785 : node47778;
														assign node47778 = (inp[0]) ? node47782 : node47779;
															assign node47779 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node47782 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node47785 = (inp[0]) ? node47789 : node47786;
															assign node47786 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node47789 = (inp[3]) ? 4'b0100 : 4'b0100;
													assign node47792 = (inp[0]) ? node47796 : node47793;
														assign node47793 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node47796 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node47799 = (inp[8]) ? node47919 : node47800;
										assign node47800 = (inp[7]) ? node47860 : node47801;
											assign node47801 = (inp[2]) ? node47829 : node47802;
												assign node47802 = (inp[14]) ? node47814 : node47803;
													assign node47803 = (inp[0]) ? node47807 : node47804;
														assign node47804 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node47807 = (inp[15]) ? node47811 : node47808;
															assign node47808 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node47811 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node47814 = (inp[3]) ? node47822 : node47815;
														assign node47815 = (inp[0]) ? node47819 : node47816;
															assign node47816 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node47819 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node47822 = (inp[15]) ? node47826 : node47823;
															assign node47823 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node47826 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node47829 = (inp[14]) ? node47845 : node47830;
													assign node47830 = (inp[15]) ? node47838 : node47831;
														assign node47831 = (inp[0]) ? node47835 : node47832;
															assign node47832 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node47835 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node47838 = (inp[0]) ? node47842 : node47839;
															assign node47839 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node47842 = (inp[5]) ? 4'b0100 : 4'b0100;
													assign node47845 = (inp[5]) ? node47853 : node47846;
														assign node47846 = (inp[3]) ? node47850 : node47847;
															assign node47847 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node47850 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node47853 = (inp[3]) ? node47857 : node47854;
															assign node47854 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node47857 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node47860 = (inp[14]) ? node47890 : node47861;
												assign node47861 = (inp[2]) ? node47877 : node47862;
													assign node47862 = (inp[15]) ? node47870 : node47863;
														assign node47863 = (inp[0]) ? node47867 : node47864;
															assign node47864 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node47867 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node47870 = (inp[0]) ? node47874 : node47871;
															assign node47871 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node47874 = (inp[5]) ? 4'b0100 : 4'b0100;
													assign node47877 = (inp[5]) ? node47883 : node47878;
														assign node47878 = (inp[3]) ? 4'b1011 : node47879;
															assign node47879 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node47883 = (inp[0]) ? node47887 : node47884;
															assign node47884 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node47887 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node47890 = (inp[2]) ? node47906 : node47891;
													assign node47891 = (inp[3]) ? node47899 : node47892;
														assign node47892 = (inp[5]) ? node47896 : node47893;
															assign node47893 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node47896 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node47899 = (inp[15]) ? node47903 : node47900;
															assign node47900 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node47903 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node47906 = (inp[5]) ? node47912 : node47907;
														assign node47907 = (inp[0]) ? node47909 : 4'b1001;
															assign node47909 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node47912 = (inp[3]) ? node47916 : node47913;
															assign node47913 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node47916 = (inp[15]) ? 4'b1001 : 4'b1001;
										assign node47919 = (inp[7]) ? node47973 : node47920;
											assign node47920 = (inp[2]) ? node47950 : node47921;
												assign node47921 = (inp[14]) ? node47937 : node47922;
													assign node47922 = (inp[5]) ? node47930 : node47923;
														assign node47923 = (inp[0]) ? node47927 : node47924;
															assign node47924 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node47927 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node47930 = (inp[15]) ? node47934 : node47931;
															assign node47931 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node47934 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node47937 = (inp[5]) ? node47943 : node47938;
														assign node47938 = (inp[3]) ? 4'b1001 : node47939;
															assign node47939 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node47943 = (inp[0]) ? node47947 : node47944;
															assign node47944 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node47947 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node47950 = (inp[0]) ? node47962 : node47951;
													assign node47951 = (inp[15]) ? node47957 : node47952;
														assign node47952 = (inp[5]) ? 4'b1001 : node47953;
															assign node47953 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node47957 = (inp[3]) ? 4'b1011 : node47958;
															assign node47958 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node47962 = (inp[15]) ? node47968 : node47963;
														assign node47963 = (inp[3]) ? 4'b1011 : node47964;
															assign node47964 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node47968 = (inp[5]) ? 4'b1001 : node47969;
															assign node47969 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node47973 = (inp[14]) ? node48005 : node47974;
												assign node47974 = (inp[2]) ? node47990 : node47975;
													assign node47975 = (inp[0]) ? node47983 : node47976;
														assign node47976 = (inp[15]) ? node47980 : node47977;
															assign node47977 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node47980 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node47983 = (inp[15]) ? node47987 : node47984;
															assign node47984 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node47987 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node47990 = (inp[5]) ? node47998 : node47991;
														assign node47991 = (inp[15]) ? node47995 : node47992;
															assign node47992 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node47995 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node47998 = (inp[0]) ? node48002 : node47999;
															assign node47999 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node48002 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node48005 = (inp[3]) ? node48021 : node48006;
													assign node48006 = (inp[5]) ? node48014 : node48007;
														assign node48007 = (inp[0]) ? node48011 : node48008;
															assign node48008 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node48011 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node48014 = (inp[15]) ? node48018 : node48015;
															assign node48015 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node48018 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node48021 = (inp[0]) ? node48025 : node48022;
														assign node48022 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node48025 = (inp[15]) ? 4'b1000 : 4'b1010;
								assign node48028 = (inp[1]) ? node48254 : node48029;
									assign node48029 = (inp[8]) ? node48149 : node48030;
										assign node48030 = (inp[7]) ? node48092 : node48031;
											assign node48031 = (inp[14]) ? node48063 : node48032;
												assign node48032 = (inp[2]) ? node48048 : node48033;
													assign node48033 = (inp[3]) ? node48041 : node48034;
														assign node48034 = (inp[15]) ? node48038 : node48035;
															assign node48035 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node48038 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node48041 = (inp[0]) ? node48045 : node48042;
															assign node48042 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node48045 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node48048 = (inp[5]) ? node48056 : node48049;
														assign node48049 = (inp[3]) ? node48053 : node48050;
															assign node48050 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node48053 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node48056 = (inp[15]) ? node48060 : node48057;
															assign node48057 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node48060 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node48063 = (inp[3]) ? node48079 : node48064;
													assign node48064 = (inp[15]) ? node48072 : node48065;
														assign node48065 = (inp[0]) ? node48069 : node48066;
															assign node48066 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node48069 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node48072 = (inp[5]) ? node48076 : node48073;
															assign node48073 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node48076 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node48079 = (inp[5]) ? node48087 : node48080;
														assign node48080 = (inp[0]) ? node48084 : node48081;
															assign node48081 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node48084 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node48087 = (inp[2]) ? 4'b0100 : node48088;
															assign node48088 = (inp[15]) ? 4'b0100 : 4'b0100;
											assign node48092 = (inp[2]) ? node48120 : node48093;
												assign node48093 = (inp[14]) ? node48109 : node48094;
													assign node48094 = (inp[5]) ? node48102 : node48095;
														assign node48095 = (inp[15]) ? node48099 : node48096;
															assign node48096 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node48099 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node48102 = (inp[0]) ? node48106 : node48103;
															assign node48103 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node48106 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node48109 = (inp[0]) ? node48115 : node48110;
														assign node48110 = (inp[15]) ? node48112 : 4'b1001;
															assign node48112 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node48115 = (inp[15]) ? node48117 : 4'b1011;
															assign node48117 = (inp[3]) ? 4'b1001 : 4'b1001;
												assign node48120 = (inp[3]) ? node48136 : node48121;
													assign node48121 = (inp[5]) ? node48129 : node48122;
														assign node48122 = (inp[15]) ? node48126 : node48123;
															assign node48123 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node48126 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node48129 = (inp[15]) ? node48133 : node48130;
															assign node48130 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node48133 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node48136 = (inp[14]) ? node48144 : node48137;
														assign node48137 = (inp[5]) ? node48141 : node48138;
															assign node48138 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node48141 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node48144 = (inp[5]) ? 4'b1001 : node48145;
															assign node48145 = (inp[0]) ? 4'b1001 : 4'b1001;
										assign node48149 = (inp[7]) ? node48205 : node48150;
											assign node48150 = (inp[14]) ? node48176 : node48151;
												assign node48151 = (inp[2]) ? node48163 : node48152;
													assign node48152 = (inp[0]) ? node48158 : node48153;
														assign node48153 = (inp[15]) ? node48155 : 4'b0100;
															assign node48155 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node48158 = (inp[3]) ? node48160 : 4'b0110;
															assign node48160 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node48163 = (inp[15]) ? node48171 : node48164;
														assign node48164 = (inp[0]) ? node48168 : node48165;
															assign node48165 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node48168 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node48171 = (inp[3]) ? 4'b1011 : node48172;
															assign node48172 = (inp[5]) ? 4'b1001 : 4'b1001;
												assign node48176 = (inp[5]) ? node48192 : node48177;
													assign node48177 = (inp[2]) ? node48185 : node48178;
														assign node48178 = (inp[15]) ? node48182 : node48179;
															assign node48179 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node48182 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node48185 = (inp[0]) ? node48189 : node48186;
															assign node48186 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node48189 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node48192 = (inp[2]) ? node48200 : node48193;
														assign node48193 = (inp[3]) ? node48197 : node48194;
															assign node48194 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node48197 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node48200 = (inp[3]) ? 4'b1011 : node48201;
															assign node48201 = (inp[0]) ? 4'b1001 : 4'b1001;
											assign node48205 = (inp[14]) ? node48231 : node48206;
												assign node48206 = (inp[2]) ? node48220 : node48207;
													assign node48207 = (inp[5]) ? node48215 : node48208;
														assign node48208 = (inp[0]) ? node48212 : node48209;
															assign node48209 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node48212 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node48215 = (inp[15]) ? node48217 : 4'b1011;
															assign node48217 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node48220 = (inp[15]) ? node48226 : node48221;
														assign node48221 = (inp[0]) ? node48223 : 4'b1000;
															assign node48223 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node48226 = (inp[0]) ? node48228 : 4'b1010;
															assign node48228 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node48231 = (inp[0]) ? node48243 : node48232;
													assign node48232 = (inp[15]) ? node48238 : node48233;
														assign node48233 = (inp[3]) ? 4'b1000 : node48234;
															assign node48234 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node48238 = (inp[5]) ? 4'b1010 : node48239;
															assign node48239 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node48243 = (inp[15]) ? node48249 : node48244;
														assign node48244 = (inp[5]) ? 4'b1010 : node48245;
															assign node48245 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node48249 = (inp[5]) ? 4'b1000 : node48250;
															assign node48250 = (inp[3]) ? 4'b1000 : 4'b1010;
									assign node48254 = (inp[0]) ? node48366 : node48255;
										assign node48255 = (inp[15]) ? node48309 : node48256;
											assign node48256 = (inp[3]) ? node48286 : node48257;
												assign node48257 = (inp[5]) ? node48273 : node48258;
													assign node48258 = (inp[7]) ? node48266 : node48259;
														assign node48259 = (inp[8]) ? node48263 : node48260;
															assign node48260 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node48263 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node48266 = (inp[8]) ? node48270 : node48267;
															assign node48267 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node48270 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node48273 = (inp[8]) ? node48279 : node48274;
														assign node48274 = (inp[14]) ? 4'b1001 : node48275;
															assign node48275 = (inp[2]) ? 4'b1000 : 4'b1000;
														assign node48279 = (inp[7]) ? node48283 : node48280;
															assign node48280 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node48283 = (inp[14]) ? 4'b1000 : 4'b1000;
												assign node48286 = (inp[8]) ? node48298 : node48287;
													assign node48287 = (inp[7]) ? node48293 : node48288;
														assign node48288 = (inp[2]) ? 4'b1000 : node48289;
															assign node48289 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node48293 = (inp[2]) ? 4'b1001 : node48294;
															assign node48294 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node48298 = (inp[7]) ? node48304 : node48299;
														assign node48299 = (inp[14]) ? 4'b1001 : node48300;
															assign node48300 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node48304 = (inp[2]) ? 4'b1000 : node48305;
															assign node48305 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node48309 = (inp[3]) ? node48337 : node48310;
												assign node48310 = (inp[5]) ? node48324 : node48311;
													assign node48311 = (inp[2]) ? node48319 : node48312;
														assign node48312 = (inp[14]) ? node48316 : node48313;
															assign node48313 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node48316 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node48319 = (inp[7]) ? 4'b1001 : node48320;
															assign node48320 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node48324 = (inp[2]) ? node48332 : node48325;
														assign node48325 = (inp[7]) ? node48329 : node48326;
															assign node48326 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node48329 = (inp[14]) ? 4'b1010 : 4'b1010;
														assign node48332 = (inp[7]) ? node48334 : 4'b1011;
															assign node48334 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node48337 = (inp[2]) ? node48353 : node48338;
													assign node48338 = (inp[7]) ? node48346 : node48339;
														assign node48339 = (inp[5]) ? node48343 : node48340;
															assign node48340 = (inp[8]) ? 4'b1010 : 4'b1010;
															assign node48343 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node48346 = (inp[5]) ? node48350 : node48347;
															assign node48347 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node48350 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node48353 = (inp[14]) ? node48361 : node48354;
														assign node48354 = (inp[5]) ? node48358 : node48355;
															assign node48355 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node48358 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node48361 = (inp[8]) ? node48363 : 4'b1011;
															assign node48363 = (inp[7]) ? 4'b1010 : 4'b1011;
										assign node48366 = (inp[15]) ? node48420 : node48367;
											assign node48367 = (inp[3]) ? node48397 : node48368;
												assign node48368 = (inp[5]) ? node48382 : node48369;
													assign node48369 = (inp[8]) ? node48377 : node48370;
														assign node48370 = (inp[7]) ? node48374 : node48371;
															assign node48371 = (inp[2]) ? 4'b1000 : 4'b1000;
															assign node48374 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node48377 = (inp[7]) ? node48379 : 4'b1001;
															assign node48379 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node48382 = (inp[14]) ? node48390 : node48383;
														assign node48383 = (inp[8]) ? node48387 : node48384;
															assign node48384 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node48387 = (inp[2]) ? 4'b1010 : 4'b1010;
														assign node48390 = (inp[2]) ? node48394 : node48391;
															assign node48391 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node48394 = (inp[7]) ? 4'b1010 : 4'b1010;
												assign node48397 = (inp[7]) ? node48409 : node48398;
													assign node48398 = (inp[8]) ? node48404 : node48399;
														assign node48399 = (inp[14]) ? 4'b1010 : node48400;
															assign node48400 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node48404 = (inp[2]) ? 4'b1011 : node48405;
															assign node48405 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node48409 = (inp[8]) ? node48415 : node48410;
														assign node48410 = (inp[14]) ? 4'b1011 : node48411;
															assign node48411 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node48415 = (inp[2]) ? 4'b1010 : node48416;
															assign node48416 = (inp[14]) ? 4'b1010 : 4'b1011;
											assign node48420 = (inp[3]) ? node48452 : node48421;
												assign node48421 = (inp[5]) ? node48437 : node48422;
													assign node48422 = (inp[2]) ? node48430 : node48423;
														assign node48423 = (inp[14]) ? node48427 : node48424;
															assign node48424 = (inp[8]) ? 4'b1010 : 4'b1010;
															assign node48427 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node48430 = (inp[14]) ? node48434 : node48431;
															assign node48431 = (inp[8]) ? 4'b1010 : 4'b1010;
															assign node48434 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node48437 = (inp[14]) ? node48445 : node48438;
														assign node48438 = (inp[8]) ? node48442 : node48439;
															assign node48439 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node48442 = (inp[2]) ? 4'b1000 : 4'b1000;
														assign node48445 = (inp[7]) ? node48449 : node48446;
															assign node48446 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node48449 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node48452 = (inp[7]) ? node48464 : node48453;
													assign node48453 = (inp[8]) ? node48459 : node48454;
														assign node48454 = (inp[2]) ? 4'b1000 : node48455;
															assign node48455 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node48459 = (inp[2]) ? 4'b1001 : node48460;
															assign node48460 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node48464 = (inp[8]) ? node48470 : node48465;
														assign node48465 = (inp[2]) ? 4'b1001 : node48466;
															assign node48466 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node48470 = (inp[2]) ? 4'b1000 : node48471;
															assign node48471 = (inp[14]) ? 4'b1000 : 4'b1001;
						assign node48475 = (inp[11]) ? node49393 : node48476;
							assign node48476 = (inp[13]) ? node48930 : node48477;
								assign node48477 = (inp[1]) ? node48709 : node48478;
									assign node48478 = (inp[5]) ? node48596 : node48479;
										assign node48479 = (inp[15]) ? node48535 : node48480;
											assign node48480 = (inp[2]) ? node48506 : node48481;
												assign node48481 = (inp[3]) ? node48497 : node48482;
													assign node48482 = (inp[0]) ? node48490 : node48483;
														assign node48483 = (inp[8]) ? node48487 : node48484;
															assign node48484 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node48487 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node48490 = (inp[7]) ? node48494 : node48491;
															assign node48491 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node48494 = (inp[14]) ? 4'b0100 : 4'b0100;
													assign node48497 = (inp[0]) ? node48499 : 4'b0100;
														assign node48499 = (inp[7]) ? node48503 : node48500;
															assign node48500 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node48503 = (inp[14]) ? 4'b0110 : 4'b0110;
												assign node48506 = (inp[3]) ? node48520 : node48507;
													assign node48507 = (inp[0]) ? node48515 : node48508;
														assign node48508 = (inp[14]) ? node48512 : node48509;
															assign node48509 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node48512 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node48515 = (inp[14]) ? 4'b0100 : node48516;
															assign node48516 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node48520 = (inp[0]) ? node48528 : node48521;
														assign node48521 = (inp[7]) ? node48525 : node48522;
															assign node48522 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node48525 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node48528 = (inp[14]) ? node48532 : node48529;
															assign node48529 = (inp[8]) ? 4'b0110 : 4'b0110;
															assign node48532 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node48535 = (inp[3]) ? node48567 : node48536;
												assign node48536 = (inp[0]) ? node48552 : node48537;
													assign node48537 = (inp[7]) ? node48545 : node48538;
														assign node48538 = (inp[8]) ? node48542 : node48539;
															assign node48539 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node48542 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node48545 = (inp[8]) ? node48549 : node48546;
															assign node48546 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node48549 = (inp[2]) ? 4'b0100 : 4'b0100;
													assign node48552 = (inp[2]) ? node48560 : node48553;
														assign node48553 = (inp[7]) ? node48557 : node48554;
															assign node48554 = (inp[14]) ? 4'b0110 : 4'b0110;
															assign node48557 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node48560 = (inp[14]) ? node48564 : node48561;
															assign node48561 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node48564 = (inp[8]) ? 4'b0110 : 4'b0110;
												assign node48567 = (inp[0]) ? node48581 : node48568;
													assign node48568 = (inp[14]) ? node48574 : node48569;
														assign node48569 = (inp[7]) ? node48571 : 4'b0110;
															assign node48571 = (inp[8]) ? 4'b0110 : 4'b0110;
														assign node48574 = (inp[8]) ? node48578 : node48575;
															assign node48575 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node48578 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node48581 = (inp[2]) ? node48589 : node48582;
														assign node48582 = (inp[7]) ? node48586 : node48583;
															assign node48583 = (inp[8]) ? 4'b0100 : 4'b0100;
															assign node48586 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node48589 = (inp[14]) ? node48593 : node48590;
															assign node48590 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node48593 = (inp[7]) ? 4'b0100 : 4'b0100;
										assign node48596 = (inp[8]) ? node48650 : node48597;
											assign node48597 = (inp[7]) ? node48629 : node48598;
												assign node48598 = (inp[14]) ? node48614 : node48599;
													assign node48599 = (inp[2]) ? node48607 : node48600;
														assign node48600 = (inp[3]) ? node48604 : node48601;
															assign node48601 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node48604 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node48607 = (inp[15]) ? node48611 : node48608;
															assign node48608 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node48611 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node48614 = (inp[3]) ? node48622 : node48615;
														assign node48615 = (inp[2]) ? node48619 : node48616;
															assign node48616 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node48619 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node48622 = (inp[15]) ? node48626 : node48623;
															assign node48623 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node48626 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node48629 = (inp[14]) ? node48643 : node48630;
													assign node48630 = (inp[2]) ? node48638 : node48631;
														assign node48631 = (inp[0]) ? node48635 : node48632;
															assign node48632 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node48635 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node48638 = (inp[3]) ? node48640 : 4'b0101;
															assign node48640 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node48643 = (inp[0]) ? node48647 : node48644;
														assign node48644 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node48647 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node48650 = (inp[7]) ? node48680 : node48651;
												assign node48651 = (inp[2]) ? node48665 : node48652;
													assign node48652 = (inp[14]) ? node48658 : node48653;
														assign node48653 = (inp[15]) ? 4'b0100 : node48654;
															assign node48654 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node48658 = (inp[3]) ? node48662 : node48659;
															assign node48659 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node48662 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node48665 = (inp[14]) ? node48673 : node48666;
														assign node48666 = (inp[15]) ? node48670 : node48667;
															assign node48667 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node48670 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node48673 = (inp[3]) ? node48677 : node48674;
															assign node48674 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node48677 = (inp[0]) ? 4'b0101 : 4'b0101;
												assign node48680 = (inp[14]) ? node48694 : node48681;
													assign node48681 = (inp[2]) ? node48689 : node48682;
														assign node48682 = (inp[15]) ? node48686 : node48683;
															assign node48683 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node48686 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node48689 = (inp[3]) ? node48691 : 4'b0100;
															assign node48691 = (inp[0]) ? 4'b0100 : 4'b0100;
													assign node48694 = (inp[2]) ? node48702 : node48695;
														assign node48695 = (inp[15]) ? node48699 : node48696;
															assign node48696 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node48699 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node48702 = (inp[3]) ? node48706 : node48703;
															assign node48703 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node48706 = (inp[0]) ? 4'b0100 : 4'b0100;
									assign node48709 = (inp[7]) ? node48829 : node48710;
										assign node48710 = (inp[8]) ? node48770 : node48711;
											assign node48711 = (inp[14]) ? node48739 : node48712;
												assign node48712 = (inp[2]) ? node48726 : node48713;
													assign node48713 = (inp[3]) ? node48721 : node48714;
														assign node48714 = (inp[0]) ? node48718 : node48715;
															assign node48715 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node48718 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node48721 = (inp[5]) ? node48723 : 4'b0111;
															assign node48723 = (inp[0]) ? 4'b0101 : 4'b0101;
													assign node48726 = (inp[5]) ? node48734 : node48727;
														assign node48727 = (inp[15]) ? node48731 : node48728;
															assign node48728 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node48731 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node48734 = (inp[3]) ? node48736 : 4'b0110;
															assign node48736 = (inp[15]) ? 4'b0100 : 4'b0100;
												assign node48739 = (inp[2]) ? node48755 : node48740;
													assign node48740 = (inp[15]) ? node48748 : node48741;
														assign node48741 = (inp[0]) ? node48745 : node48742;
															assign node48742 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node48745 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node48748 = (inp[0]) ? node48752 : node48749;
															assign node48749 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node48752 = (inp[3]) ? 4'b0100 : 4'b0100;
													assign node48755 = (inp[5]) ? node48763 : node48756;
														assign node48756 = (inp[3]) ? node48760 : node48757;
															assign node48757 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node48760 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node48763 = (inp[15]) ? node48767 : node48764;
															assign node48764 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node48767 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node48770 = (inp[2]) ? node48800 : node48771;
												assign node48771 = (inp[14]) ? node48787 : node48772;
													assign node48772 = (inp[5]) ? node48780 : node48773;
														assign node48773 = (inp[15]) ? node48777 : node48774;
															assign node48774 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node48777 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node48780 = (inp[0]) ? node48784 : node48781;
															assign node48781 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node48784 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node48787 = (inp[0]) ? node48795 : node48788;
														assign node48788 = (inp[15]) ? node48792 : node48789;
															assign node48789 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node48792 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node48795 = (inp[15]) ? node48797 : 4'b1011;
															assign node48797 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node48800 = (inp[3]) ? node48814 : node48801;
													assign node48801 = (inp[15]) ? node48809 : node48802;
														assign node48802 = (inp[0]) ? node48806 : node48803;
															assign node48803 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node48806 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node48809 = (inp[5]) ? node48811 : 4'b1011;
															assign node48811 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node48814 = (inp[14]) ? node48822 : node48815;
														assign node48815 = (inp[5]) ? node48819 : node48816;
															assign node48816 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node48819 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node48822 = (inp[5]) ? node48826 : node48823;
															assign node48823 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node48826 = (inp[15]) ? 4'b1001 : 4'b1001;
										assign node48829 = (inp[8]) ? node48879 : node48830;
											assign node48830 = (inp[2]) ? node48856 : node48831;
												assign node48831 = (inp[14]) ? node48843 : node48832;
													assign node48832 = (inp[15]) ? node48838 : node48833;
														assign node48833 = (inp[0]) ? node48835 : 4'b0100;
															assign node48835 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node48838 = (inp[3]) ? node48840 : 4'b0110;
															assign node48840 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node48843 = (inp[0]) ? node48851 : node48844;
														assign node48844 = (inp[15]) ? node48848 : node48845;
															assign node48845 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node48848 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node48851 = (inp[15]) ? 4'b1001 : node48852;
															assign node48852 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node48856 = (inp[15]) ? node48868 : node48857;
													assign node48857 = (inp[0]) ? node48863 : node48858;
														assign node48858 = (inp[3]) ? 4'b1001 : node48859;
															assign node48859 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node48863 = (inp[5]) ? 4'b1011 : node48864;
															assign node48864 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node48868 = (inp[0]) ? node48874 : node48869;
														assign node48869 = (inp[5]) ? 4'b1011 : node48870;
															assign node48870 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node48874 = (inp[5]) ? 4'b1001 : node48875;
															assign node48875 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node48879 = (inp[14]) ? node48907 : node48880;
												assign node48880 = (inp[2]) ? node48894 : node48881;
													assign node48881 = (inp[15]) ? node48887 : node48882;
														assign node48882 = (inp[0]) ? node48884 : 4'b1001;
															assign node48884 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node48887 = (inp[0]) ? node48891 : node48888;
															assign node48888 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node48891 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node48894 = (inp[0]) ? node48902 : node48895;
														assign node48895 = (inp[15]) ? node48899 : node48896;
															assign node48896 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node48899 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node48902 = (inp[15]) ? 4'b1000 : node48903;
															assign node48903 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node48907 = (inp[15]) ? node48919 : node48908;
													assign node48908 = (inp[0]) ? node48914 : node48909;
														assign node48909 = (inp[5]) ? 4'b1000 : node48910;
															assign node48910 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node48914 = (inp[5]) ? 4'b1010 : node48915;
															assign node48915 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node48919 = (inp[0]) ? node48925 : node48920;
														assign node48920 = (inp[3]) ? 4'b1010 : node48921;
															assign node48921 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node48925 = (inp[5]) ? 4'b1000 : node48926;
															assign node48926 = (inp[3]) ? 4'b1000 : 4'b1010;
								assign node48930 = (inp[1]) ? node49144 : node48931;
									assign node48931 = (inp[8]) ? node49041 : node48932;
										assign node48932 = (inp[7]) ? node48988 : node48933;
											assign node48933 = (inp[2]) ? node48965 : node48934;
												assign node48934 = (inp[14]) ? node48950 : node48935;
													assign node48935 = (inp[0]) ? node48943 : node48936;
														assign node48936 = (inp[15]) ? node48940 : node48937;
															assign node48937 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node48940 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node48943 = (inp[15]) ? node48947 : node48944;
															assign node48944 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node48947 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node48950 = (inp[5]) ? node48958 : node48951;
														assign node48951 = (inp[3]) ? node48955 : node48952;
															assign node48952 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node48955 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node48958 = (inp[3]) ? node48962 : node48959;
															assign node48959 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node48962 = (inp[0]) ? 4'b0100 : 4'b0100;
												assign node48965 = (inp[15]) ? node48977 : node48966;
													assign node48966 = (inp[0]) ? node48972 : node48967;
														assign node48967 = (inp[3]) ? 4'b0100 : node48968;
															assign node48968 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node48972 = (inp[3]) ? 4'b0110 : node48973;
															assign node48973 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node48977 = (inp[0]) ? node48983 : node48978;
														assign node48978 = (inp[5]) ? 4'b0110 : node48979;
															assign node48979 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node48983 = (inp[5]) ? 4'b0100 : node48984;
															assign node48984 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node48988 = (inp[2]) ? node49018 : node48989;
												assign node48989 = (inp[14]) ? node49005 : node48990;
													assign node48990 = (inp[3]) ? node48998 : node48991;
														assign node48991 = (inp[15]) ? node48995 : node48992;
															assign node48992 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node48995 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node48998 = (inp[5]) ? node49002 : node48999;
															assign node48999 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node49002 = (inp[0]) ? 4'b0100 : 4'b0100;
													assign node49005 = (inp[0]) ? node49011 : node49006;
														assign node49006 = (inp[15]) ? node49008 : 4'b1001;
															assign node49008 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node49011 = (inp[15]) ? node49015 : node49012;
															assign node49012 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node49015 = (inp[5]) ? 4'b1001 : 4'b1001;
												assign node49018 = (inp[0]) ? node49030 : node49019;
													assign node49019 = (inp[15]) ? node49025 : node49020;
														assign node49020 = (inp[3]) ? 4'b1001 : node49021;
															assign node49021 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node49025 = (inp[5]) ? 4'b1011 : node49026;
															assign node49026 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node49030 = (inp[15]) ? node49036 : node49031;
														assign node49031 = (inp[5]) ? 4'b1011 : node49032;
															assign node49032 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node49036 = (inp[5]) ? 4'b1001 : node49037;
															assign node49037 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node49041 = (inp[7]) ? node49095 : node49042;
											assign node49042 = (inp[2]) ? node49072 : node49043;
												assign node49043 = (inp[14]) ? node49059 : node49044;
													assign node49044 = (inp[3]) ? node49052 : node49045;
														assign node49045 = (inp[15]) ? node49049 : node49046;
															assign node49046 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node49049 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node49052 = (inp[15]) ? node49056 : node49053;
															assign node49053 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node49056 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node49059 = (inp[0]) ? node49067 : node49060;
														assign node49060 = (inp[15]) ? node49064 : node49061;
															assign node49061 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node49064 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node49067 = (inp[15]) ? node49069 : 4'b1011;
															assign node49069 = (inp[3]) ? 4'b1001 : 4'b1001;
												assign node49072 = (inp[0]) ? node49084 : node49073;
													assign node49073 = (inp[15]) ? node49079 : node49074;
														assign node49074 = (inp[5]) ? 4'b1001 : node49075;
															assign node49075 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node49079 = (inp[5]) ? 4'b1011 : node49080;
															assign node49080 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node49084 = (inp[15]) ? node49090 : node49085;
														assign node49085 = (inp[5]) ? 4'b1011 : node49086;
															assign node49086 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node49090 = (inp[3]) ? 4'b1001 : node49091;
															assign node49091 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node49095 = (inp[14]) ? node49121 : node49096;
												assign node49096 = (inp[2]) ? node49110 : node49097;
													assign node49097 = (inp[15]) ? node49105 : node49098;
														assign node49098 = (inp[0]) ? node49102 : node49099;
															assign node49099 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node49102 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node49105 = (inp[3]) ? 4'b1001 : node49106;
															assign node49106 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node49110 = (inp[15]) ? node49116 : node49111;
														assign node49111 = (inp[0]) ? 4'b1010 : node49112;
															assign node49112 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node49116 = (inp[0]) ? 4'b1000 : node49117;
															assign node49117 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node49121 = (inp[0]) ? node49133 : node49122;
													assign node49122 = (inp[15]) ? node49128 : node49123;
														assign node49123 = (inp[5]) ? 4'b1000 : node49124;
															assign node49124 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node49128 = (inp[3]) ? 4'b1010 : node49129;
															assign node49129 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node49133 = (inp[15]) ? node49139 : node49134;
														assign node49134 = (inp[5]) ? 4'b1010 : node49135;
															assign node49135 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node49139 = (inp[3]) ? 4'b1000 : node49140;
															assign node49140 = (inp[5]) ? 4'b1000 : 4'b1010;
									assign node49144 = (inp[5]) ? node49272 : node49145;
										assign node49145 = (inp[15]) ? node49209 : node49146;
											assign node49146 = (inp[8]) ? node49178 : node49147;
												assign node49147 = (inp[7]) ? node49163 : node49148;
													assign node49148 = (inp[2]) ? node49156 : node49149;
														assign node49149 = (inp[14]) ? node49153 : node49150;
															assign node49150 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node49153 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node49156 = (inp[14]) ? node49160 : node49157;
															assign node49157 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node49160 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node49163 = (inp[2]) ? node49171 : node49164;
														assign node49164 = (inp[14]) ? node49168 : node49165;
															assign node49165 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node49168 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node49171 = (inp[3]) ? node49175 : node49172;
															assign node49172 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node49175 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node49178 = (inp[7]) ? node49194 : node49179;
													assign node49179 = (inp[14]) ? node49187 : node49180;
														assign node49180 = (inp[2]) ? node49184 : node49181;
															assign node49181 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node49184 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node49187 = (inp[2]) ? node49191 : node49188;
															assign node49188 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node49191 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node49194 = (inp[2]) ? node49202 : node49195;
														assign node49195 = (inp[14]) ? node49199 : node49196;
															assign node49196 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node49199 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node49202 = (inp[0]) ? node49206 : node49203;
															assign node49203 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node49206 = (inp[3]) ? 4'b1010 : 4'b1000;
											assign node49209 = (inp[2]) ? node49241 : node49210;
												assign node49210 = (inp[14]) ? node49226 : node49211;
													assign node49211 = (inp[8]) ? node49219 : node49212;
														assign node49212 = (inp[7]) ? node49216 : node49213;
															assign node49213 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node49216 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node49219 = (inp[7]) ? node49223 : node49220;
															assign node49220 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node49223 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node49226 = (inp[3]) ? node49234 : node49227;
														assign node49227 = (inp[0]) ? node49231 : node49228;
															assign node49228 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node49231 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node49234 = (inp[0]) ? node49238 : node49235;
															assign node49235 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node49238 = (inp[8]) ? 4'b1000 : 4'b1000;
												assign node49241 = (inp[7]) ? node49257 : node49242;
													assign node49242 = (inp[8]) ? node49250 : node49243;
														assign node49243 = (inp[3]) ? node49247 : node49244;
															assign node49244 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node49247 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node49250 = (inp[14]) ? node49254 : node49251;
															assign node49251 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node49254 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node49257 = (inp[8]) ? node49265 : node49258;
														assign node49258 = (inp[14]) ? node49262 : node49259;
															assign node49259 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node49262 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node49265 = (inp[0]) ? node49269 : node49266;
															assign node49266 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node49269 = (inp[3]) ? 4'b1000 : 4'b1010;
										assign node49272 = (inp[2]) ? node49332 : node49273;
											assign node49273 = (inp[7]) ? node49303 : node49274;
												assign node49274 = (inp[3]) ? node49290 : node49275;
													assign node49275 = (inp[0]) ? node49283 : node49276;
														assign node49276 = (inp[15]) ? node49280 : node49277;
															assign node49277 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node49280 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node49283 = (inp[15]) ? node49287 : node49284;
															assign node49284 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node49287 = (inp[14]) ? 4'b1000 : 4'b1000;
													assign node49290 = (inp[8]) ? node49298 : node49291;
														assign node49291 = (inp[14]) ? node49295 : node49292;
															assign node49292 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node49295 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node49298 = (inp[14]) ? 4'b1011 : node49299;
															assign node49299 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node49303 = (inp[8]) ? node49319 : node49304;
													assign node49304 = (inp[14]) ? node49312 : node49305;
														assign node49305 = (inp[3]) ? node49309 : node49306;
															assign node49306 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node49309 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node49312 = (inp[0]) ? node49316 : node49313;
															assign node49313 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node49316 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node49319 = (inp[14]) ? node49327 : node49320;
														assign node49320 = (inp[15]) ? node49324 : node49321;
															assign node49321 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node49324 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node49327 = (inp[3]) ? node49329 : 4'b1000;
															assign node49329 = (inp[15]) ? 4'b1000 : 4'b1000;
											assign node49332 = (inp[3]) ? node49362 : node49333;
												assign node49333 = (inp[14]) ? node49347 : node49334;
													assign node49334 = (inp[15]) ? node49342 : node49335;
														assign node49335 = (inp[0]) ? node49339 : node49336;
															assign node49336 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node49339 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node49342 = (inp[0]) ? 4'b1000 : node49343;
															assign node49343 = (inp[8]) ? 4'b1010 : 4'b1010;
													assign node49347 = (inp[8]) ? node49355 : node49348;
														assign node49348 = (inp[7]) ? node49352 : node49349;
															assign node49349 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node49352 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node49355 = (inp[7]) ? node49359 : node49356;
															assign node49356 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node49359 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node49362 = (inp[8]) ? node49378 : node49363;
													assign node49363 = (inp[7]) ? node49371 : node49364;
														assign node49364 = (inp[0]) ? node49368 : node49365;
															assign node49365 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node49368 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node49371 = (inp[15]) ? node49375 : node49372;
															assign node49372 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node49375 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node49378 = (inp[7]) ? node49386 : node49379;
														assign node49379 = (inp[14]) ? node49383 : node49380;
															assign node49380 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node49383 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node49386 = (inp[0]) ? node49390 : node49387;
															assign node49387 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node49390 = (inp[15]) ? 4'b1000 : 4'b1010;
							assign node49393 = (inp[13]) ? node49829 : node49394;
								assign node49394 = (inp[1]) ? node49614 : node49395;
									assign node49395 = (inp[0]) ? node49511 : node49396;
										assign node49396 = (inp[15]) ? node49456 : node49397;
											assign node49397 = (inp[5]) ? node49429 : node49398;
												assign node49398 = (inp[3]) ? node49414 : node49399;
													assign node49399 = (inp[2]) ? node49407 : node49400;
														assign node49400 = (inp[8]) ? node49404 : node49401;
															assign node49401 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node49404 = (inp[14]) ? 4'b1010 : 4'b1010;
														assign node49407 = (inp[8]) ? node49411 : node49408;
															assign node49408 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node49411 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node49414 = (inp[7]) ? node49422 : node49415;
														assign node49415 = (inp[8]) ? node49419 : node49416;
															assign node49416 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node49419 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node49422 = (inp[8]) ? node49426 : node49423;
															assign node49423 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node49426 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node49429 = (inp[3]) ? node49443 : node49430;
													assign node49430 = (inp[7]) ? node49438 : node49431;
														assign node49431 = (inp[8]) ? node49435 : node49432;
															assign node49432 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node49435 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node49438 = (inp[8]) ? 4'b1000 : node49439;
															assign node49439 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node49443 = (inp[8]) ? node49449 : node49444;
														assign node49444 = (inp[2]) ? node49446 : 4'b1001;
															assign node49446 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node49449 = (inp[7]) ? node49453 : node49450;
															assign node49450 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node49453 = (inp[14]) ? 4'b1000 : 4'b1000;
											assign node49456 = (inp[5]) ? node49488 : node49457;
												assign node49457 = (inp[3]) ? node49473 : node49458;
													assign node49458 = (inp[14]) ? node49466 : node49459;
														assign node49459 = (inp[7]) ? node49463 : node49460;
															assign node49460 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node49463 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node49466 = (inp[8]) ? node49470 : node49467;
															assign node49467 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node49470 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node49473 = (inp[2]) ? node49481 : node49474;
														assign node49474 = (inp[14]) ? node49478 : node49475;
															assign node49475 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node49478 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node49481 = (inp[8]) ? node49485 : node49482;
															assign node49482 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node49485 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node49488 = (inp[8]) ? node49500 : node49489;
													assign node49489 = (inp[7]) ? node49495 : node49490;
														assign node49490 = (inp[14]) ? 4'b1010 : node49491;
															assign node49491 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node49495 = (inp[2]) ? 4'b1011 : node49496;
															assign node49496 = (inp[3]) ? 4'b1010 : 4'b1011;
													assign node49500 = (inp[7]) ? node49506 : node49501;
														assign node49501 = (inp[2]) ? 4'b1011 : node49502;
															assign node49502 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node49506 = (inp[2]) ? 4'b1010 : node49507;
															assign node49507 = (inp[14]) ? 4'b1010 : 4'b1011;
										assign node49511 = (inp[15]) ? node49561 : node49512;
											assign node49512 = (inp[3]) ? node49540 : node49513;
												assign node49513 = (inp[5]) ? node49525 : node49514;
													assign node49514 = (inp[2]) ? node49520 : node49515;
														assign node49515 = (inp[7]) ? 4'b1001 : node49516;
															assign node49516 = (inp[14]) ? 4'b1000 : 4'b1000;
														assign node49520 = (inp[14]) ? 4'b1000 : node49521;
															assign node49521 = (inp[8]) ? 4'b1000 : 4'b1000;
													assign node49525 = (inp[14]) ? node49533 : node49526;
														assign node49526 = (inp[7]) ? node49530 : node49527;
															assign node49527 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node49530 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node49533 = (inp[7]) ? node49537 : node49534;
															assign node49534 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node49537 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node49540 = (inp[8]) ? node49552 : node49541;
													assign node49541 = (inp[7]) ? node49547 : node49542;
														assign node49542 = (inp[14]) ? 4'b1010 : node49543;
															assign node49543 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node49547 = (inp[2]) ? 4'b1011 : node49548;
															assign node49548 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node49552 = (inp[7]) ? node49556 : node49553;
														assign node49553 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node49556 = (inp[2]) ? 4'b1010 : node49557;
															assign node49557 = (inp[14]) ? 4'b1010 : 4'b1011;
											assign node49561 = (inp[5]) ? node49591 : node49562;
												assign node49562 = (inp[3]) ? node49576 : node49563;
													assign node49563 = (inp[7]) ? node49571 : node49564;
														assign node49564 = (inp[8]) ? node49568 : node49565;
															assign node49565 = (inp[14]) ? 4'b1010 : 4'b1011;
															assign node49568 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node49571 = (inp[8]) ? node49573 : 4'b1011;
															assign node49573 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node49576 = (inp[14]) ? node49584 : node49577;
														assign node49577 = (inp[8]) ? node49581 : node49578;
															assign node49578 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node49581 = (inp[2]) ? 4'b1000 : 4'b1000;
														assign node49584 = (inp[7]) ? node49588 : node49585;
															assign node49585 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node49588 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node49591 = (inp[14]) ? node49607 : node49592;
													assign node49592 = (inp[3]) ? node49600 : node49593;
														assign node49593 = (inp[7]) ? node49597 : node49594;
															assign node49594 = (inp[2]) ? 4'b1000 : 4'b1000;
															assign node49597 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node49600 = (inp[2]) ? node49604 : node49601;
															assign node49601 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node49604 = (inp[8]) ? 4'b1000 : 4'b1000;
													assign node49607 = (inp[8]) ? node49611 : node49608;
														assign node49608 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node49611 = (inp[7]) ? 4'b1000 : 4'b1001;
									assign node49614 = (inp[7]) ? node49720 : node49615;
										assign node49615 = (inp[8]) ? node49671 : node49616;
											assign node49616 = (inp[2]) ? node49648 : node49617;
												assign node49617 = (inp[14]) ? node49633 : node49618;
													assign node49618 = (inp[15]) ? node49626 : node49619;
														assign node49619 = (inp[0]) ? node49623 : node49620;
															assign node49620 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node49623 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node49626 = (inp[0]) ? node49630 : node49627;
															assign node49627 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node49630 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node49633 = (inp[5]) ? node49641 : node49634;
														assign node49634 = (inp[3]) ? node49638 : node49635;
															assign node49635 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node49638 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node49641 = (inp[15]) ? node49645 : node49642;
															assign node49642 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node49645 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node49648 = (inp[0]) ? node49660 : node49649;
													assign node49649 = (inp[15]) ? node49655 : node49650;
														assign node49650 = (inp[3]) ? 4'b1000 : node49651;
															assign node49651 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node49655 = (inp[5]) ? 4'b1010 : node49656;
															assign node49656 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node49660 = (inp[15]) ? node49666 : node49661;
														assign node49661 = (inp[3]) ? 4'b1010 : node49662;
															assign node49662 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node49666 = (inp[5]) ? 4'b1000 : node49667;
															assign node49667 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node49671 = (inp[14]) ? node49699 : node49672;
												assign node49672 = (inp[2]) ? node49686 : node49673;
													assign node49673 = (inp[3]) ? node49681 : node49674;
														assign node49674 = (inp[15]) ? node49678 : node49675;
															assign node49675 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node49678 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node49681 = (inp[5]) ? node49683 : 4'b1010;
															assign node49683 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node49686 = (inp[15]) ? node49692 : node49687;
														assign node49687 = (inp[0]) ? 4'b0011 : node49688;
															assign node49688 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node49692 = (inp[0]) ? node49696 : node49693;
															assign node49693 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node49696 = (inp[3]) ? 4'b0001 : 4'b0001;
												assign node49699 = (inp[0]) ? node49709 : node49700;
													assign node49700 = (inp[15]) ? node49704 : node49701;
														assign node49701 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node49704 = (inp[5]) ? 4'b0011 : node49705;
															assign node49705 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node49709 = (inp[15]) ? node49715 : node49710;
														assign node49710 = (inp[5]) ? 4'b0011 : node49711;
															assign node49711 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node49715 = (inp[3]) ? 4'b0001 : node49716;
															assign node49716 = (inp[5]) ? 4'b0001 : 4'b0011;
										assign node49720 = (inp[8]) ? node49776 : node49721;
											assign node49721 = (inp[14]) ? node49749 : node49722;
												assign node49722 = (inp[2]) ? node49738 : node49723;
													assign node49723 = (inp[0]) ? node49731 : node49724;
														assign node49724 = (inp[15]) ? node49728 : node49725;
															assign node49725 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node49728 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node49731 = (inp[15]) ? node49735 : node49732;
															assign node49732 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node49735 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node49738 = (inp[0]) ? node49744 : node49739;
														assign node49739 = (inp[15]) ? 4'b0011 : node49740;
															assign node49740 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node49744 = (inp[15]) ? 4'b0001 : node49745;
															assign node49745 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node49749 = (inp[2]) ? node49765 : node49750;
													assign node49750 = (inp[0]) ? node49758 : node49751;
														assign node49751 = (inp[15]) ? node49755 : node49752;
															assign node49752 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node49755 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node49758 = (inp[15]) ? node49762 : node49759;
															assign node49759 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node49762 = (inp[5]) ? 4'b0001 : 4'b0001;
													assign node49765 = (inp[15]) ? node49773 : node49766;
														assign node49766 = (inp[0]) ? node49770 : node49767;
															assign node49767 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node49770 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node49773 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node49776 = (inp[2]) ? node49808 : node49777;
												assign node49777 = (inp[14]) ? node49793 : node49778;
													assign node49778 = (inp[15]) ? node49786 : node49779;
														assign node49779 = (inp[0]) ? node49783 : node49780;
															assign node49780 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node49783 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node49786 = (inp[0]) ? node49790 : node49787;
															assign node49787 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node49790 = (inp[5]) ? 4'b0001 : 4'b0001;
													assign node49793 = (inp[3]) ? node49801 : node49794;
														assign node49794 = (inp[0]) ? node49798 : node49795;
															assign node49795 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node49798 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node49801 = (inp[15]) ? node49805 : node49802;
															assign node49802 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node49805 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node49808 = (inp[3]) ? node49822 : node49809;
													assign node49809 = (inp[14]) ? node49817 : node49810;
														assign node49810 = (inp[5]) ? node49814 : node49811;
															assign node49811 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node49814 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node49817 = (inp[15]) ? node49819 : 4'b0010;
															assign node49819 = (inp[5]) ? 4'b0000 : 4'b0000;
													assign node49822 = (inp[0]) ? node49826 : node49823;
														assign node49823 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node49826 = (inp[15]) ? 4'b0000 : 4'b0010;
								assign node49829 = (inp[1]) ? node50057 : node49830;
									assign node49830 = (inp[7]) ? node49944 : node49831;
										assign node49831 = (inp[8]) ? node49885 : node49832;
											assign node49832 = (inp[2]) ? node49862 : node49833;
												assign node49833 = (inp[14]) ? node49847 : node49834;
													assign node49834 = (inp[5]) ? node49842 : node49835;
														assign node49835 = (inp[15]) ? node49839 : node49836;
															assign node49836 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node49839 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node49842 = (inp[3]) ? 4'b1011 : node49843;
															assign node49843 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node49847 = (inp[5]) ? node49855 : node49848;
														assign node49848 = (inp[3]) ? node49852 : node49849;
															assign node49849 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node49852 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node49855 = (inp[15]) ? node49859 : node49856;
															assign node49856 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node49859 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node49862 = (inp[0]) ? node49874 : node49863;
													assign node49863 = (inp[15]) ? node49869 : node49864;
														assign node49864 = (inp[3]) ? 4'b1000 : node49865;
															assign node49865 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node49869 = (inp[3]) ? 4'b1010 : node49870;
															assign node49870 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node49874 = (inp[15]) ? node49880 : node49875;
														assign node49875 = (inp[3]) ? 4'b1010 : node49876;
															assign node49876 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node49880 = (inp[5]) ? 4'b1000 : node49881;
															assign node49881 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node49885 = (inp[2]) ? node49917 : node49886;
												assign node49886 = (inp[14]) ? node49902 : node49887;
													assign node49887 = (inp[5]) ? node49895 : node49888;
														assign node49888 = (inp[0]) ? node49892 : node49889;
															assign node49889 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node49892 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node49895 = (inp[3]) ? node49899 : node49896;
															assign node49896 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node49899 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node49902 = (inp[3]) ? node49910 : node49903;
														assign node49903 = (inp[15]) ? node49907 : node49904;
															assign node49904 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node49907 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node49910 = (inp[5]) ? node49914 : node49911;
															assign node49911 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node49914 = (inp[0]) ? 4'b0001 : 4'b0001;
												assign node49917 = (inp[5]) ? node49931 : node49918;
													assign node49918 = (inp[0]) ? node49924 : node49919;
														assign node49919 = (inp[14]) ? 4'b0001 : node49920;
															assign node49920 = (inp[3]) ? 4'b0001 : 4'b0001;
														assign node49924 = (inp[3]) ? node49928 : node49925;
															assign node49925 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node49928 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node49931 = (inp[3]) ? node49937 : node49932;
														assign node49932 = (inp[14]) ? 4'b0011 : node49933;
															assign node49933 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node49937 = (inp[15]) ? node49941 : node49938;
															assign node49938 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node49941 = (inp[0]) ? 4'b0001 : 4'b0011;
										assign node49944 = (inp[8]) ? node49996 : node49945;
											assign node49945 = (inp[2]) ? node49975 : node49946;
												assign node49946 = (inp[14]) ? node49960 : node49947;
													assign node49947 = (inp[15]) ? node49953 : node49948;
														assign node49948 = (inp[3]) ? 4'b1000 : node49949;
															assign node49949 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node49953 = (inp[0]) ? node49957 : node49954;
															assign node49954 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node49957 = (inp[3]) ? 4'b1000 : 4'b1000;
													assign node49960 = (inp[3]) ? node49968 : node49961;
														assign node49961 = (inp[15]) ? node49965 : node49962;
															assign node49962 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node49965 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node49968 = (inp[15]) ? node49972 : node49969;
															assign node49969 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node49972 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node49975 = (inp[15]) ? node49985 : node49976;
													assign node49976 = (inp[0]) ? node49980 : node49977;
														assign node49977 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node49980 = (inp[3]) ? 4'b0011 : node49981;
															assign node49981 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node49985 = (inp[0]) ? node49991 : node49986;
														assign node49986 = (inp[3]) ? 4'b0011 : node49987;
															assign node49987 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node49991 = (inp[3]) ? 4'b0001 : node49992;
															assign node49992 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node49996 = (inp[14]) ? node50026 : node49997;
												assign node49997 = (inp[2]) ? node50013 : node49998;
													assign node49998 = (inp[3]) ? node50006 : node49999;
														assign node49999 = (inp[5]) ? node50003 : node50000;
															assign node50000 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node50003 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node50006 = (inp[15]) ? node50010 : node50007;
															assign node50007 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node50010 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node50013 = (inp[15]) ? node50019 : node50014;
														assign node50014 = (inp[0]) ? 4'b0010 : node50015;
															assign node50015 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node50019 = (inp[0]) ? node50023 : node50020;
															assign node50020 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node50023 = (inp[3]) ? 4'b0000 : 4'b0000;
												assign node50026 = (inp[2]) ? node50042 : node50027;
													assign node50027 = (inp[15]) ? node50035 : node50028;
														assign node50028 = (inp[0]) ? node50032 : node50029;
															assign node50029 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node50032 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node50035 = (inp[0]) ? node50039 : node50036;
															assign node50036 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node50039 = (inp[3]) ? 4'b0000 : 4'b0000;
													assign node50042 = (inp[5]) ? node50050 : node50043;
														assign node50043 = (inp[15]) ? node50047 : node50044;
															assign node50044 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node50047 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node50050 = (inp[3]) ? node50054 : node50051;
															assign node50051 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node50054 = (inp[15]) ? 4'b0000 : 4'b0000;
									assign node50057 = (inp[7]) ? node50159 : node50058;
										assign node50058 = (inp[8]) ? node50114 : node50059;
											assign node50059 = (inp[2]) ? node50091 : node50060;
												assign node50060 = (inp[14]) ? node50076 : node50061;
													assign node50061 = (inp[15]) ? node50069 : node50062;
														assign node50062 = (inp[0]) ? node50066 : node50063;
															assign node50063 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node50066 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node50069 = (inp[0]) ? node50073 : node50070;
															assign node50070 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node50073 = (inp[5]) ? 4'b0001 : 4'b0001;
													assign node50076 = (inp[0]) ? node50084 : node50077;
														assign node50077 = (inp[15]) ? node50081 : node50078;
															assign node50078 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node50081 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node50084 = (inp[15]) ? node50088 : node50085;
															assign node50085 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node50088 = (inp[3]) ? 4'b0000 : 4'b0000;
												assign node50091 = (inp[0]) ? node50103 : node50092;
													assign node50092 = (inp[15]) ? node50098 : node50093;
														assign node50093 = (inp[5]) ? 4'b0000 : node50094;
															assign node50094 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node50098 = (inp[3]) ? 4'b0010 : node50099;
															assign node50099 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node50103 = (inp[15]) ? node50109 : node50104;
														assign node50104 = (inp[3]) ? 4'b0010 : node50105;
															assign node50105 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node50109 = (inp[3]) ? 4'b0000 : node50110;
															assign node50110 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node50114 = (inp[2]) ? node50138 : node50115;
												assign node50115 = (inp[14]) ? node50129 : node50116;
													assign node50116 = (inp[3]) ? node50122 : node50117;
														assign node50117 = (inp[15]) ? node50119 : 4'b0010;
															assign node50119 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node50122 = (inp[15]) ? node50126 : node50123;
															assign node50123 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node50126 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node50129 = (inp[0]) ? node50135 : node50130;
														assign node50130 = (inp[15]) ? node50132 : 4'b0001;
															assign node50132 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node50135 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node50138 = (inp[3]) ? node50152 : node50139;
													assign node50139 = (inp[14]) ? node50145 : node50140;
														assign node50140 = (inp[15]) ? 4'b0011 : node50141;
															assign node50141 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node50145 = (inp[5]) ? node50149 : node50146;
															assign node50146 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node50149 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node50152 = (inp[0]) ? node50156 : node50153;
														assign node50153 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node50156 = (inp[15]) ? 4'b0001 : 4'b0011;
										assign node50159 = (inp[8]) ? node50217 : node50160;
											assign node50160 = (inp[14]) ? node50188 : node50161;
												assign node50161 = (inp[2]) ? node50175 : node50162;
													assign node50162 = (inp[5]) ? node50168 : node50163;
														assign node50163 = (inp[0]) ? node50165 : 4'b0000;
															assign node50165 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node50168 = (inp[0]) ? node50172 : node50169;
															assign node50169 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node50172 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node50175 = (inp[15]) ? node50181 : node50176;
														assign node50176 = (inp[0]) ? node50178 : 4'b0001;
															assign node50178 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node50181 = (inp[0]) ? node50185 : node50182;
															assign node50182 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node50185 = (inp[3]) ? 4'b0001 : 4'b0001;
												assign node50188 = (inp[2]) ? node50202 : node50189;
													assign node50189 = (inp[15]) ? node50197 : node50190;
														assign node50190 = (inp[0]) ? node50194 : node50191;
															assign node50191 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node50194 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node50197 = (inp[0]) ? 4'b0001 : node50198;
															assign node50198 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node50202 = (inp[3]) ? node50210 : node50203;
														assign node50203 = (inp[0]) ? node50207 : node50204;
															assign node50204 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node50207 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node50210 = (inp[15]) ? node50214 : node50211;
															assign node50211 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node50214 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node50217 = (inp[2]) ? node50245 : node50218;
												assign node50218 = (inp[14]) ? node50234 : node50219;
													assign node50219 = (inp[3]) ? node50227 : node50220;
														assign node50220 = (inp[0]) ? node50224 : node50221;
															assign node50221 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node50224 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node50227 = (inp[0]) ? node50231 : node50228;
															assign node50228 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node50231 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node50234 = (inp[0]) ? node50240 : node50235;
														assign node50235 = (inp[15]) ? node50237 : 4'b0000;
															assign node50237 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node50240 = (inp[15]) ? node50242 : 4'b0010;
															assign node50242 = (inp[3]) ? 4'b0000 : 4'b0000;
												assign node50245 = (inp[3]) ? node50261 : node50246;
													assign node50246 = (inp[15]) ? node50254 : node50247;
														assign node50247 = (inp[5]) ? node50251 : node50248;
															assign node50248 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node50251 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node50254 = (inp[5]) ? node50258 : node50255;
															assign node50255 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node50258 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node50261 = (inp[15]) ? node50265 : node50262;
														assign node50262 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node50265 = (inp[0]) ? 4'b0000 : 4'b0010;
				assign node50268 = (inp[12]) ? node53934 : node50269;
					assign node50269 = (inp[6]) ? node52145 : node50270;
						assign node50270 = (inp[11]) ? node51184 : node50271;
							assign node50271 = (inp[13]) ? node50723 : node50272;
								assign node50272 = (inp[1]) ? node50492 : node50273;
									assign node50273 = (inp[15]) ? node50387 : node50274;
										assign node50274 = (inp[0]) ? node50332 : node50275;
											assign node50275 = (inp[3]) ? node50305 : node50276;
												assign node50276 = (inp[5]) ? node50292 : node50277;
													assign node50277 = (inp[14]) ? node50285 : node50278;
														assign node50278 = (inp[7]) ? node50282 : node50279;
															assign node50279 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node50282 = (inp[8]) ? 4'b1110 : 4'b1110;
														assign node50285 = (inp[8]) ? node50289 : node50286;
															assign node50286 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node50289 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node50292 = (inp[14]) ? node50298 : node50293;
														assign node50293 = (inp[8]) ? node50295 : 4'b1101;
															assign node50295 = (inp[2]) ? 4'b1100 : 4'b1100;
														assign node50298 = (inp[7]) ? node50302 : node50299;
															assign node50299 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node50302 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node50305 = (inp[5]) ? node50319 : node50306;
													assign node50306 = (inp[14]) ? node50314 : node50307;
														assign node50307 = (inp[7]) ? node50311 : node50308;
															assign node50308 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node50311 = (inp[2]) ? 4'b1100 : 4'b1100;
														assign node50314 = (inp[8]) ? node50316 : 4'b1101;
															assign node50316 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node50319 = (inp[14]) ? node50325 : node50320;
														assign node50320 = (inp[7]) ? 4'b1101 : node50321;
															assign node50321 = (inp[2]) ? 4'b1100 : 4'b1100;
														assign node50325 = (inp[8]) ? node50329 : node50326;
															assign node50326 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node50329 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node50332 = (inp[5]) ? node50364 : node50333;
												assign node50333 = (inp[3]) ? node50349 : node50334;
													assign node50334 = (inp[14]) ? node50342 : node50335;
														assign node50335 = (inp[7]) ? node50339 : node50336;
															assign node50336 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node50339 = (inp[8]) ? 4'b1100 : 4'b1100;
														assign node50342 = (inp[8]) ? node50346 : node50343;
															assign node50343 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node50346 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node50349 = (inp[2]) ? node50357 : node50350;
														assign node50350 = (inp[7]) ? node50354 : node50351;
															assign node50351 = (inp[8]) ? 4'b1110 : 4'b1110;
															assign node50354 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node50357 = (inp[8]) ? node50361 : node50358;
															assign node50358 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node50361 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node50364 = (inp[7]) ? node50376 : node50365;
													assign node50365 = (inp[8]) ? node50371 : node50366;
														assign node50366 = (inp[2]) ? 4'b1110 : node50367;
															assign node50367 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node50371 = (inp[2]) ? 4'b1111 : node50372;
															assign node50372 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node50376 = (inp[8]) ? node50382 : node50377;
														assign node50377 = (inp[2]) ? 4'b1111 : node50378;
															assign node50378 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node50382 = (inp[14]) ? 4'b1110 : node50383;
															assign node50383 = (inp[2]) ? 4'b1110 : 4'b1111;
										assign node50387 = (inp[0]) ? node50441 : node50388;
											assign node50388 = (inp[3]) ? node50418 : node50389;
												assign node50389 = (inp[5]) ? node50405 : node50390;
													assign node50390 = (inp[2]) ? node50398 : node50391;
														assign node50391 = (inp[7]) ? node50395 : node50392;
															assign node50392 = (inp[8]) ? 4'b1100 : 4'b1100;
															assign node50395 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node50398 = (inp[7]) ? node50402 : node50399;
															assign node50399 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node50402 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node50405 = (inp[7]) ? node50413 : node50406;
														assign node50406 = (inp[8]) ? node50410 : node50407;
															assign node50407 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node50410 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node50413 = (inp[8]) ? 4'b1110 : node50414;
															assign node50414 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node50418 = (inp[8]) ? node50430 : node50419;
													assign node50419 = (inp[7]) ? node50425 : node50420;
														assign node50420 = (inp[2]) ? 4'b1110 : node50421;
															assign node50421 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node50425 = (inp[14]) ? 4'b1111 : node50426;
															assign node50426 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node50430 = (inp[7]) ? node50436 : node50431;
														assign node50431 = (inp[2]) ? 4'b1111 : node50432;
															assign node50432 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node50436 = (inp[2]) ? 4'b1110 : node50437;
															assign node50437 = (inp[5]) ? 4'b1110 : 4'b1111;
											assign node50441 = (inp[5]) ? node50469 : node50442;
												assign node50442 = (inp[3]) ? node50456 : node50443;
													assign node50443 = (inp[7]) ? node50451 : node50444;
														assign node50444 = (inp[8]) ? node50448 : node50445;
															assign node50445 = (inp[2]) ? 4'b1110 : 4'b1110;
															assign node50448 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node50451 = (inp[8]) ? 4'b1110 : node50452;
															assign node50452 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node50456 = (inp[8]) ? node50462 : node50457;
														assign node50457 = (inp[14]) ? 4'b1101 : node50458;
															assign node50458 = (inp[7]) ? 4'b1100 : 4'b1100;
														assign node50462 = (inp[7]) ? node50466 : node50463;
															assign node50463 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node50466 = (inp[14]) ? 4'b1100 : 4'b1100;
												assign node50469 = (inp[8]) ? node50481 : node50470;
													assign node50470 = (inp[7]) ? node50476 : node50471;
														assign node50471 = (inp[2]) ? 4'b1100 : node50472;
															assign node50472 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node50476 = (inp[2]) ? 4'b1101 : node50477;
															assign node50477 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node50481 = (inp[7]) ? node50487 : node50482;
														assign node50482 = (inp[2]) ? 4'b1101 : node50483;
															assign node50483 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node50487 = (inp[2]) ? 4'b1100 : node50488;
															assign node50488 = (inp[14]) ? 4'b1100 : 4'b1101;
									assign node50492 = (inp[7]) ? node50608 : node50493;
										assign node50493 = (inp[8]) ? node50545 : node50494;
											assign node50494 = (inp[14]) ? node50522 : node50495;
												assign node50495 = (inp[2]) ? node50511 : node50496;
													assign node50496 = (inp[5]) ? node50504 : node50497;
														assign node50497 = (inp[3]) ? node50501 : node50498;
															assign node50498 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node50501 = (inp[15]) ? 4'b1101 : 4'b1101;
														assign node50504 = (inp[0]) ? node50508 : node50505;
															assign node50505 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node50508 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node50511 = (inp[15]) ? node50515 : node50512;
														assign node50512 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node50515 = (inp[0]) ? node50519 : node50516;
															assign node50516 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node50519 = (inp[3]) ? 4'b1100 : 4'b1100;
												assign node50522 = (inp[15]) ? node50534 : node50523;
													assign node50523 = (inp[0]) ? node50529 : node50524;
														assign node50524 = (inp[5]) ? 4'b1100 : node50525;
															assign node50525 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node50529 = (inp[5]) ? 4'b1110 : node50530;
															assign node50530 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node50534 = (inp[0]) ? node50540 : node50535;
														assign node50535 = (inp[5]) ? 4'b1110 : node50536;
															assign node50536 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node50540 = (inp[3]) ? 4'b1100 : node50541;
															assign node50541 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node50545 = (inp[14]) ? node50577 : node50546;
												assign node50546 = (inp[2]) ? node50562 : node50547;
													assign node50547 = (inp[15]) ? node50555 : node50548;
														assign node50548 = (inp[0]) ? node50552 : node50549;
															assign node50549 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node50552 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node50555 = (inp[0]) ? node50559 : node50556;
															assign node50556 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node50559 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node50562 = (inp[5]) ? node50570 : node50563;
														assign node50563 = (inp[3]) ? node50567 : node50564;
															assign node50564 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node50567 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node50570 = (inp[15]) ? node50574 : node50571;
															assign node50571 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node50574 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node50577 = (inp[2]) ? node50593 : node50578;
													assign node50578 = (inp[5]) ? node50586 : node50579;
														assign node50579 = (inp[3]) ? node50583 : node50580;
															assign node50580 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node50583 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node50586 = (inp[0]) ? node50590 : node50587;
															assign node50587 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node50590 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node50593 = (inp[15]) ? node50601 : node50594;
														assign node50594 = (inp[0]) ? node50598 : node50595;
															assign node50595 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node50598 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node50601 = (inp[0]) ? node50605 : node50602;
															assign node50602 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node50605 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node50608 = (inp[8]) ? node50670 : node50609;
											assign node50609 = (inp[14]) ? node50639 : node50610;
												assign node50610 = (inp[2]) ? node50624 : node50611;
													assign node50611 = (inp[15]) ? node50617 : node50612;
														assign node50612 = (inp[0]) ? node50614 : 4'b1100;
															assign node50614 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node50617 = (inp[0]) ? node50621 : node50618;
															assign node50618 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node50621 = (inp[3]) ? 4'b1100 : 4'b1100;
													assign node50624 = (inp[5]) ? node50632 : node50625;
														assign node50625 = (inp[15]) ? node50629 : node50626;
															assign node50626 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node50629 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node50632 = (inp[15]) ? node50636 : node50633;
															assign node50633 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node50636 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node50639 = (inp[2]) ? node50655 : node50640;
													assign node50640 = (inp[5]) ? node50648 : node50641;
														assign node50641 = (inp[0]) ? node50645 : node50642;
															assign node50642 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node50645 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node50648 = (inp[15]) ? node50652 : node50649;
															assign node50649 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node50652 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node50655 = (inp[15]) ? node50663 : node50656;
														assign node50656 = (inp[0]) ? node50660 : node50657;
															assign node50657 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node50660 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node50663 = (inp[0]) ? node50667 : node50664;
															assign node50664 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node50667 = (inp[3]) ? 4'b0101 : 4'b0101;
											assign node50670 = (inp[2]) ? node50700 : node50671;
												assign node50671 = (inp[14]) ? node50687 : node50672;
													assign node50672 = (inp[3]) ? node50680 : node50673;
														assign node50673 = (inp[0]) ? node50677 : node50674;
															assign node50674 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node50677 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node50680 = (inp[15]) ? node50684 : node50681;
															assign node50681 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node50684 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node50687 = (inp[3]) ? node50693 : node50688;
														assign node50688 = (inp[0]) ? node50690 : 4'b0110;
															assign node50690 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node50693 = (inp[5]) ? node50697 : node50694;
															assign node50694 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node50697 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node50700 = (inp[0]) ? node50712 : node50701;
													assign node50701 = (inp[15]) ? node50707 : node50702;
														assign node50702 = (inp[3]) ? 4'b0100 : node50703;
															assign node50703 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node50707 = (inp[3]) ? 4'b0110 : node50708;
															assign node50708 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node50712 = (inp[15]) ? node50718 : node50713;
														assign node50713 = (inp[3]) ? 4'b0110 : node50714;
															assign node50714 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node50718 = (inp[3]) ? 4'b0100 : node50719;
															assign node50719 = (inp[5]) ? 4'b0100 : 4'b0110;
								assign node50723 = (inp[1]) ? node50945 : node50724;
									assign node50724 = (inp[8]) ? node50838 : node50725;
										assign node50725 = (inp[7]) ? node50785 : node50726;
											assign node50726 = (inp[14]) ? node50754 : node50727;
												assign node50727 = (inp[2]) ? node50743 : node50728;
													assign node50728 = (inp[15]) ? node50736 : node50729;
														assign node50729 = (inp[0]) ? node50733 : node50730;
															assign node50730 = (inp[5]) ? 4'b1101 : 4'b1101;
															assign node50733 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node50736 = (inp[0]) ? node50740 : node50737;
															assign node50737 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node50740 = (inp[3]) ? 4'b1101 : 4'b1101;
													assign node50743 = (inp[15]) ? node50749 : node50744;
														assign node50744 = (inp[0]) ? 4'b1110 : node50745;
															assign node50745 = (inp[5]) ? 4'b1100 : 4'b1100;
														assign node50749 = (inp[0]) ? 4'b1100 : node50750;
															assign node50750 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node50754 = (inp[5]) ? node50770 : node50755;
													assign node50755 = (inp[0]) ? node50763 : node50756;
														assign node50756 = (inp[3]) ? node50760 : node50757;
															assign node50757 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node50760 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node50763 = (inp[15]) ? node50767 : node50764;
															assign node50764 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node50767 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node50770 = (inp[3]) ? node50778 : node50771;
														assign node50771 = (inp[0]) ? node50775 : node50772;
															assign node50772 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node50775 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node50778 = (inp[2]) ? node50782 : node50779;
															assign node50779 = (inp[15]) ? 4'b1100 : 4'b1100;
															assign node50782 = (inp[15]) ? 4'b1100 : 4'b1100;
											assign node50785 = (inp[14]) ? node50815 : node50786;
												assign node50786 = (inp[2]) ? node50802 : node50787;
													assign node50787 = (inp[15]) ? node50795 : node50788;
														assign node50788 = (inp[0]) ? node50792 : node50789;
															assign node50789 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node50792 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node50795 = (inp[0]) ? node50799 : node50796;
															assign node50796 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node50799 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node50802 = (inp[0]) ? node50810 : node50803;
														assign node50803 = (inp[15]) ? node50807 : node50804;
															assign node50804 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node50807 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node50810 = (inp[5]) ? 4'b0101 : node50811;
															assign node50811 = (inp[3]) ? 4'b0101 : 4'b0101;
												assign node50815 = (inp[0]) ? node50827 : node50816;
													assign node50816 = (inp[15]) ? node50822 : node50817;
														assign node50817 = (inp[3]) ? 4'b0101 : node50818;
															assign node50818 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node50822 = (inp[3]) ? 4'b0111 : node50823;
															assign node50823 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node50827 = (inp[15]) ? node50833 : node50828;
														assign node50828 = (inp[3]) ? 4'b0111 : node50829;
															assign node50829 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node50833 = (inp[3]) ? 4'b0101 : node50834;
															assign node50834 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node50838 = (inp[7]) ? node50890 : node50839;
											assign node50839 = (inp[14]) ? node50867 : node50840;
												assign node50840 = (inp[2]) ? node50854 : node50841;
													assign node50841 = (inp[3]) ? node50849 : node50842;
														assign node50842 = (inp[0]) ? node50846 : node50843;
															assign node50843 = (inp[5]) ? 4'b1100 : 4'b1100;
															assign node50846 = (inp[15]) ? 4'b1100 : 4'b1100;
														assign node50849 = (inp[15]) ? 4'b1110 : node50850;
															assign node50850 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node50854 = (inp[15]) ? node50860 : node50855;
														assign node50855 = (inp[0]) ? 4'b0111 : node50856;
															assign node50856 = (inp[3]) ? 4'b0101 : 4'b0101;
														assign node50860 = (inp[0]) ? node50864 : node50861;
															assign node50861 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node50864 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node50867 = (inp[15]) ? node50879 : node50868;
													assign node50868 = (inp[0]) ? node50874 : node50869;
														assign node50869 = (inp[3]) ? 4'b0101 : node50870;
															assign node50870 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node50874 = (inp[5]) ? 4'b0111 : node50875;
															assign node50875 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node50879 = (inp[0]) ? node50885 : node50880;
														assign node50880 = (inp[5]) ? 4'b0111 : node50881;
															assign node50881 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node50885 = (inp[3]) ? 4'b0101 : node50886;
															assign node50886 = (inp[5]) ? 4'b0101 : 4'b0111;
											assign node50890 = (inp[14]) ? node50922 : node50891;
												assign node50891 = (inp[2]) ? node50907 : node50892;
													assign node50892 = (inp[0]) ? node50900 : node50893;
														assign node50893 = (inp[15]) ? node50897 : node50894;
															assign node50894 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node50897 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node50900 = (inp[15]) ? node50904 : node50901;
															assign node50901 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node50904 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node50907 = (inp[0]) ? node50915 : node50908;
														assign node50908 = (inp[15]) ? node50912 : node50909;
															assign node50909 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node50912 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node50915 = (inp[15]) ? node50919 : node50916;
															assign node50916 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node50919 = (inp[5]) ? 4'b0100 : 4'b0100;
												assign node50922 = (inp[15]) ? node50934 : node50923;
													assign node50923 = (inp[0]) ? node50929 : node50924;
														assign node50924 = (inp[3]) ? 4'b0100 : node50925;
															assign node50925 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node50929 = (inp[5]) ? 4'b0110 : node50930;
															assign node50930 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node50934 = (inp[0]) ? node50940 : node50935;
														assign node50935 = (inp[3]) ? 4'b0110 : node50936;
															assign node50936 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node50940 = (inp[3]) ? 4'b0100 : node50941;
															assign node50941 = (inp[5]) ? 4'b0100 : 4'b0110;
									assign node50945 = (inp[3]) ? node51067 : node50946;
										assign node50946 = (inp[8]) ? node51006 : node50947;
											assign node50947 = (inp[7]) ? node50977 : node50948;
												assign node50948 = (inp[2]) ? node50964 : node50949;
													assign node50949 = (inp[14]) ? node50957 : node50950;
														assign node50950 = (inp[0]) ? node50954 : node50951;
															assign node50951 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node50954 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node50957 = (inp[5]) ? node50961 : node50958;
															assign node50958 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node50961 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node50964 = (inp[14]) ? node50972 : node50965;
														assign node50965 = (inp[15]) ? node50969 : node50966;
															assign node50966 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node50969 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node50972 = (inp[0]) ? node50974 : 4'b0100;
															assign node50974 = (inp[15]) ? 4'b0100 : 4'b0100;
												assign node50977 = (inp[2]) ? node50991 : node50978;
													assign node50978 = (inp[14]) ? node50986 : node50979;
														assign node50979 = (inp[15]) ? node50983 : node50980;
															assign node50980 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node50983 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node50986 = (inp[5]) ? node50988 : 4'b0101;
															assign node50988 = (inp[0]) ? 4'b0101 : 4'b0101;
													assign node50991 = (inp[14]) ? node50999 : node50992;
														assign node50992 = (inp[15]) ? node50996 : node50993;
															assign node50993 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node50996 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node50999 = (inp[15]) ? node51003 : node51000;
															assign node51000 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node51003 = (inp[0]) ? 4'b0101 : 4'b0101;
											assign node51006 = (inp[7]) ? node51036 : node51007;
												assign node51007 = (inp[14]) ? node51023 : node51008;
													assign node51008 = (inp[2]) ? node51016 : node51009;
														assign node51009 = (inp[15]) ? node51013 : node51010;
															assign node51010 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node51013 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node51016 = (inp[15]) ? node51020 : node51017;
															assign node51017 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node51020 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node51023 = (inp[5]) ? node51031 : node51024;
														assign node51024 = (inp[0]) ? node51028 : node51025;
															assign node51025 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node51028 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node51031 = (inp[2]) ? 4'b0101 : node51032;
															assign node51032 = (inp[0]) ? 4'b0101 : 4'b0101;
												assign node51036 = (inp[14]) ? node51052 : node51037;
													assign node51037 = (inp[2]) ? node51045 : node51038;
														assign node51038 = (inp[15]) ? node51042 : node51039;
															assign node51039 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node51042 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node51045 = (inp[15]) ? node51049 : node51046;
															assign node51046 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node51049 = (inp[0]) ? 4'b0100 : 4'b0100;
													assign node51052 = (inp[15]) ? node51060 : node51053;
														assign node51053 = (inp[0]) ? node51057 : node51054;
															assign node51054 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node51057 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node51060 = (inp[5]) ? node51064 : node51061;
															assign node51061 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node51064 = (inp[0]) ? 4'b0100 : 4'b0110;
										assign node51067 = (inp[15]) ? node51127 : node51068;
											assign node51068 = (inp[0]) ? node51098 : node51069;
												assign node51069 = (inp[2]) ? node51083 : node51070;
													assign node51070 = (inp[14]) ? node51078 : node51071;
														assign node51071 = (inp[7]) ? node51075 : node51072;
															assign node51072 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node51075 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node51078 = (inp[7]) ? node51080 : 4'b0101;
															assign node51080 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node51083 = (inp[5]) ? node51091 : node51084;
														assign node51084 = (inp[7]) ? node51088 : node51085;
															assign node51085 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node51088 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node51091 = (inp[7]) ? node51095 : node51092;
															assign node51092 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node51095 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node51098 = (inp[5]) ? node51114 : node51099;
													assign node51099 = (inp[2]) ? node51107 : node51100;
														assign node51100 = (inp[8]) ? node51104 : node51101;
															assign node51101 = (inp[7]) ? 4'b0110 : 4'b0110;
															assign node51104 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node51107 = (inp[14]) ? node51111 : node51108;
															assign node51108 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node51111 = (inp[8]) ? 4'b0110 : 4'b0110;
													assign node51114 = (inp[2]) ? node51120 : node51115;
														assign node51115 = (inp[8]) ? node51117 : 4'b0110;
															assign node51117 = (inp[7]) ? 4'b0110 : 4'b0110;
														assign node51120 = (inp[7]) ? node51124 : node51121;
															assign node51121 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node51124 = (inp[8]) ? 4'b0110 : 4'b0111;
											assign node51127 = (inp[0]) ? node51157 : node51128;
												assign node51128 = (inp[14]) ? node51142 : node51129;
													assign node51129 = (inp[8]) ? node51137 : node51130;
														assign node51130 = (inp[7]) ? node51134 : node51131;
															assign node51131 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node51134 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node51137 = (inp[2]) ? node51139 : 4'b0110;
															assign node51139 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node51142 = (inp[5]) ? node51150 : node51143;
														assign node51143 = (inp[8]) ? node51147 : node51144;
															assign node51144 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node51147 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node51150 = (inp[7]) ? node51154 : node51151;
															assign node51151 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node51154 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node51157 = (inp[14]) ? node51169 : node51158;
													assign node51158 = (inp[7]) ? node51164 : node51159;
														assign node51159 = (inp[5]) ? 4'b0101 : node51160;
															assign node51160 = (inp[2]) ? 4'b0100 : 4'b0100;
														assign node51164 = (inp[5]) ? node51166 : 4'b0101;
															assign node51166 = (inp[8]) ? 4'b0100 : 4'b0100;
													assign node51169 = (inp[2]) ? node51177 : node51170;
														assign node51170 = (inp[5]) ? node51174 : node51171;
															assign node51171 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node51174 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node51177 = (inp[8]) ? node51181 : node51178;
															assign node51178 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node51181 = (inp[7]) ? 4'b0100 : 4'b0101;
							assign node51184 = (inp[1]) ? node51668 : node51185;
								assign node51185 = (inp[13]) ? node51433 : node51186;
									assign node51186 = (inp[3]) ? node51306 : node51187;
										assign node51187 = (inp[15]) ? node51245 : node51188;
											assign node51188 = (inp[0]) ? node51216 : node51189;
												assign node51189 = (inp[5]) ? node51201 : node51190;
													assign node51190 = (inp[7]) ? node51196 : node51191;
														assign node51191 = (inp[8]) ? 4'b0111 : node51192;
															assign node51192 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node51196 = (inp[8]) ? 4'b0110 : node51197;
															assign node51197 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node51201 = (inp[2]) ? node51209 : node51202;
														assign node51202 = (inp[14]) ? node51206 : node51203;
															assign node51203 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node51206 = (inp[7]) ? 4'b0100 : 4'b0100;
														assign node51209 = (inp[7]) ? node51213 : node51210;
															assign node51210 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node51213 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node51216 = (inp[5]) ? node51232 : node51217;
													assign node51217 = (inp[14]) ? node51225 : node51218;
														assign node51218 = (inp[2]) ? node51222 : node51219;
															assign node51219 = (inp[7]) ? 4'b0100 : 4'b0100;
															assign node51222 = (inp[8]) ? 4'b0100 : 4'b0100;
														assign node51225 = (inp[8]) ? node51229 : node51226;
															assign node51226 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node51229 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node51232 = (inp[14]) ? node51238 : node51233;
														assign node51233 = (inp[7]) ? 4'b0111 : node51234;
															assign node51234 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node51238 = (inp[8]) ? node51242 : node51239;
															assign node51239 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node51242 = (inp[7]) ? 4'b0110 : 4'b0111;
											assign node51245 = (inp[5]) ? node51275 : node51246;
												assign node51246 = (inp[0]) ? node51262 : node51247;
													assign node51247 = (inp[7]) ? node51255 : node51248;
														assign node51248 = (inp[8]) ? node51252 : node51249;
															assign node51249 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node51252 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node51255 = (inp[8]) ? node51259 : node51256;
															assign node51256 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node51259 = (inp[2]) ? 4'b0100 : 4'b0100;
													assign node51262 = (inp[7]) ? node51268 : node51263;
														assign node51263 = (inp[8]) ? node51265 : 4'b0110;
															assign node51265 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node51268 = (inp[8]) ? node51272 : node51269;
															assign node51269 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node51272 = (inp[14]) ? 4'b0110 : 4'b0110;
												assign node51275 = (inp[0]) ? node51291 : node51276;
													assign node51276 = (inp[2]) ? node51284 : node51277;
														assign node51277 = (inp[8]) ? node51281 : node51278;
															assign node51278 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node51281 = (inp[14]) ? 4'b0110 : 4'b0110;
														assign node51284 = (inp[8]) ? node51288 : node51285;
															assign node51285 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node51288 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node51291 = (inp[7]) ? node51299 : node51292;
														assign node51292 = (inp[8]) ? node51296 : node51293;
															assign node51293 = (inp[14]) ? 4'b0100 : 4'b0100;
															assign node51296 = (inp[14]) ? 4'b0101 : 4'b0100;
														assign node51299 = (inp[8]) ? node51303 : node51300;
															assign node51300 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node51303 = (inp[14]) ? 4'b0100 : 4'b0101;
										assign node51306 = (inp[5]) ? node51370 : node51307;
											assign node51307 = (inp[8]) ? node51339 : node51308;
												assign node51308 = (inp[7]) ? node51324 : node51309;
													assign node51309 = (inp[14]) ? node51317 : node51310;
														assign node51310 = (inp[2]) ? node51314 : node51311;
															assign node51311 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node51314 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node51317 = (inp[15]) ? node51321 : node51318;
															assign node51318 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node51321 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node51324 = (inp[14]) ? node51332 : node51325;
														assign node51325 = (inp[2]) ? node51329 : node51326;
															assign node51326 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node51329 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node51332 = (inp[2]) ? node51336 : node51333;
															assign node51333 = (inp[0]) ? 4'b0101 : 4'b0101;
															assign node51336 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node51339 = (inp[7]) ? node51355 : node51340;
													assign node51340 = (inp[2]) ? node51348 : node51341;
														assign node51341 = (inp[14]) ? node51345 : node51342;
															assign node51342 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node51345 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node51348 = (inp[14]) ? node51352 : node51349;
															assign node51349 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node51352 = (inp[15]) ? 4'b0101 : 4'b0101;
													assign node51355 = (inp[2]) ? node51363 : node51356;
														assign node51356 = (inp[14]) ? node51360 : node51357;
															assign node51357 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node51360 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node51363 = (inp[0]) ? node51367 : node51364;
															assign node51364 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node51367 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node51370 = (inp[8]) ? node51402 : node51371;
												assign node51371 = (inp[7]) ? node51387 : node51372;
													assign node51372 = (inp[14]) ? node51380 : node51373;
														assign node51373 = (inp[2]) ? node51377 : node51374;
															assign node51374 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node51377 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node51380 = (inp[2]) ? node51384 : node51381;
															assign node51381 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node51384 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node51387 = (inp[14]) ? node51395 : node51388;
														assign node51388 = (inp[2]) ? node51392 : node51389;
															assign node51389 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node51392 = (inp[0]) ? 4'b0101 : 4'b0101;
														assign node51395 = (inp[15]) ? node51399 : node51396;
															assign node51396 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node51399 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node51402 = (inp[7]) ? node51418 : node51403;
													assign node51403 = (inp[14]) ? node51411 : node51404;
														assign node51404 = (inp[2]) ? node51408 : node51405;
															assign node51405 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node51408 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node51411 = (inp[2]) ? node51415 : node51412;
															assign node51412 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node51415 = (inp[0]) ? 4'b0101 : 4'b0101;
													assign node51418 = (inp[14]) ? node51426 : node51419;
														assign node51419 = (inp[2]) ? node51423 : node51420;
															assign node51420 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node51423 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node51426 = (inp[2]) ? node51430 : node51427;
															assign node51427 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node51430 = (inp[15]) ? 4'b0110 : 4'b0100;
									assign node51433 = (inp[7]) ? node51543 : node51434;
										assign node51434 = (inp[8]) ? node51490 : node51435;
											assign node51435 = (inp[2]) ? node51467 : node51436;
												assign node51436 = (inp[14]) ? node51452 : node51437;
													assign node51437 = (inp[15]) ? node51445 : node51438;
														assign node51438 = (inp[0]) ? node51442 : node51439;
															assign node51439 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node51442 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node51445 = (inp[0]) ? node51449 : node51446;
															assign node51446 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node51449 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node51452 = (inp[5]) ? node51460 : node51453;
														assign node51453 = (inp[15]) ? node51457 : node51454;
															assign node51454 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node51457 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node51460 = (inp[3]) ? node51464 : node51461;
															assign node51461 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node51464 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node51467 = (inp[3]) ? node51483 : node51468;
													assign node51468 = (inp[0]) ? node51476 : node51469;
														assign node51469 = (inp[14]) ? node51473 : node51470;
															assign node51470 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node51473 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node51476 = (inp[5]) ? node51480 : node51477;
															assign node51477 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node51480 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node51483 = (inp[15]) ? node51487 : node51484;
														assign node51484 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node51487 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node51490 = (inp[14]) ? node51520 : node51491;
												assign node51491 = (inp[2]) ? node51507 : node51492;
													assign node51492 = (inp[3]) ? node51500 : node51493;
														assign node51493 = (inp[5]) ? node51497 : node51494;
															assign node51494 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node51497 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node51500 = (inp[5]) ? node51504 : node51501;
															assign node51501 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node51504 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node51507 = (inp[0]) ? node51513 : node51508;
														assign node51508 = (inp[15]) ? node51510 : 4'b1001;
															assign node51510 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node51513 = (inp[15]) ? node51517 : node51514;
															assign node51514 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node51517 = (inp[5]) ? 4'b1001 : 4'b1001;
												assign node51520 = (inp[15]) ? node51532 : node51521;
													assign node51521 = (inp[0]) ? node51527 : node51522;
														assign node51522 = (inp[3]) ? 4'b1001 : node51523;
															assign node51523 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node51527 = (inp[5]) ? 4'b1011 : node51528;
															assign node51528 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node51532 = (inp[0]) ? node51538 : node51533;
														assign node51533 = (inp[3]) ? 4'b1011 : node51534;
															assign node51534 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node51538 = (inp[5]) ? 4'b1001 : node51539;
															assign node51539 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node51543 = (inp[8]) ? node51607 : node51544;
											assign node51544 = (inp[14]) ? node51576 : node51545;
												assign node51545 = (inp[2]) ? node51561 : node51546;
													assign node51546 = (inp[3]) ? node51554 : node51547;
														assign node51547 = (inp[0]) ? node51551 : node51548;
															assign node51548 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node51551 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node51554 = (inp[5]) ? node51558 : node51555;
															assign node51555 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node51558 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node51561 = (inp[0]) ? node51569 : node51562;
														assign node51562 = (inp[15]) ? node51566 : node51563;
															assign node51563 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node51566 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node51569 = (inp[15]) ? node51573 : node51570;
															assign node51570 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node51573 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node51576 = (inp[2]) ? node51592 : node51577;
													assign node51577 = (inp[0]) ? node51585 : node51578;
														assign node51578 = (inp[15]) ? node51582 : node51579;
															assign node51579 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node51582 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node51585 = (inp[15]) ? node51589 : node51586;
															assign node51586 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node51589 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node51592 = (inp[3]) ? node51600 : node51593;
														assign node51593 = (inp[0]) ? node51597 : node51594;
															assign node51594 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node51597 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node51600 = (inp[0]) ? node51604 : node51601;
															assign node51601 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node51604 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node51607 = (inp[2]) ? node51637 : node51608;
												assign node51608 = (inp[14]) ? node51624 : node51609;
													assign node51609 = (inp[0]) ? node51617 : node51610;
														assign node51610 = (inp[15]) ? node51614 : node51611;
															assign node51611 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node51614 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node51617 = (inp[15]) ? node51621 : node51618;
															assign node51618 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node51621 = (inp[3]) ? 4'b1001 : 4'b1001;
													assign node51624 = (inp[3]) ? node51630 : node51625;
														assign node51625 = (inp[0]) ? node51627 : 4'b1010;
															assign node51627 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node51630 = (inp[5]) ? node51634 : node51631;
															assign node51631 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node51634 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node51637 = (inp[3]) ? node51653 : node51638;
													assign node51638 = (inp[5]) ? node51646 : node51639;
														assign node51639 = (inp[0]) ? node51643 : node51640;
															assign node51640 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node51643 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node51646 = (inp[0]) ? node51650 : node51647;
															assign node51647 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node51650 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node51653 = (inp[5]) ? node51661 : node51654;
														assign node51654 = (inp[14]) ? node51658 : node51655;
															assign node51655 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node51658 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node51661 = (inp[0]) ? node51665 : node51662;
															assign node51662 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node51665 = (inp[15]) ? 4'b1000 : 4'b1010;
								assign node51668 = (inp[13]) ? node51896 : node51669;
									assign node51669 = (inp[8]) ? node51785 : node51670;
										assign node51670 = (inp[7]) ? node51732 : node51671;
											assign node51671 = (inp[2]) ? node51703 : node51672;
												assign node51672 = (inp[14]) ? node51688 : node51673;
													assign node51673 = (inp[0]) ? node51681 : node51674;
														assign node51674 = (inp[15]) ? node51678 : node51675;
															assign node51675 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node51678 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node51681 = (inp[15]) ? node51685 : node51682;
															assign node51682 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node51685 = (inp[5]) ? 4'b0101 : 4'b0101;
													assign node51688 = (inp[5]) ? node51696 : node51689;
														assign node51689 = (inp[15]) ? node51693 : node51690;
															assign node51690 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node51693 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node51696 = (inp[15]) ? node51700 : node51697;
															assign node51697 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node51700 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node51703 = (inp[14]) ? node51719 : node51704;
													assign node51704 = (inp[3]) ? node51712 : node51705;
														assign node51705 = (inp[15]) ? node51709 : node51706;
															assign node51706 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node51709 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node51712 = (inp[0]) ? node51716 : node51713;
															assign node51713 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node51716 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node51719 = (inp[0]) ? node51725 : node51720;
														assign node51720 = (inp[15]) ? node51722 : 4'b0100;
															assign node51722 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node51725 = (inp[15]) ? node51729 : node51726;
															assign node51726 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node51729 = (inp[5]) ? 4'b0100 : 4'b0100;
											assign node51732 = (inp[14]) ? node51762 : node51733;
												assign node51733 = (inp[2]) ? node51749 : node51734;
													assign node51734 = (inp[0]) ? node51742 : node51735;
														assign node51735 = (inp[15]) ? node51739 : node51736;
															assign node51736 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node51739 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node51742 = (inp[15]) ? node51746 : node51743;
															assign node51743 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node51746 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node51749 = (inp[15]) ? node51755 : node51750;
														assign node51750 = (inp[0]) ? 4'b1011 : node51751;
															assign node51751 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node51755 = (inp[0]) ? node51759 : node51756;
															assign node51756 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node51759 = (inp[3]) ? 4'b1001 : 4'b1001;
												assign node51762 = (inp[15]) ? node51774 : node51763;
													assign node51763 = (inp[0]) ? node51769 : node51764;
														assign node51764 = (inp[5]) ? 4'b1001 : node51765;
															assign node51765 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node51769 = (inp[5]) ? 4'b1011 : node51770;
															assign node51770 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node51774 = (inp[0]) ? node51780 : node51775;
														assign node51775 = (inp[3]) ? 4'b1011 : node51776;
															assign node51776 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node51780 = (inp[5]) ? 4'b1001 : node51781;
															assign node51781 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node51785 = (inp[7]) ? node51843 : node51786;
											assign node51786 = (inp[2]) ? node51812 : node51787;
												assign node51787 = (inp[14]) ? node51799 : node51788;
													assign node51788 = (inp[3]) ? node51794 : node51789;
														assign node51789 = (inp[15]) ? node51791 : 4'b0100;
															assign node51791 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node51794 = (inp[0]) ? node51796 : 4'b0110;
															assign node51796 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node51799 = (inp[5]) ? node51805 : node51800;
														assign node51800 = (inp[0]) ? 4'b1011 : node51801;
															assign node51801 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node51805 = (inp[3]) ? node51809 : node51806;
															assign node51806 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node51809 = (inp[15]) ? 4'b1001 : 4'b1001;
												assign node51812 = (inp[3]) ? node51828 : node51813;
													assign node51813 = (inp[14]) ? node51821 : node51814;
														assign node51814 = (inp[15]) ? node51818 : node51815;
															assign node51815 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node51818 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node51821 = (inp[0]) ? node51825 : node51822;
															assign node51822 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node51825 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node51828 = (inp[5]) ? node51836 : node51829;
														assign node51829 = (inp[15]) ? node51833 : node51830;
															assign node51830 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node51833 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node51836 = (inp[0]) ? node51840 : node51837;
															assign node51837 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node51840 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node51843 = (inp[2]) ? node51873 : node51844;
												assign node51844 = (inp[14]) ? node51860 : node51845;
													assign node51845 = (inp[15]) ? node51853 : node51846;
														assign node51846 = (inp[0]) ? node51850 : node51847;
															assign node51847 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node51850 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node51853 = (inp[0]) ? node51857 : node51854;
															assign node51854 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node51857 = (inp[3]) ? 4'b1001 : 4'b1001;
													assign node51860 = (inp[15]) ? node51868 : node51861;
														assign node51861 = (inp[0]) ? node51865 : node51862;
															assign node51862 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node51865 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node51868 = (inp[0]) ? 4'b1000 : node51869;
															assign node51869 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node51873 = (inp[15]) ? node51885 : node51874;
													assign node51874 = (inp[0]) ? node51880 : node51875;
														assign node51875 = (inp[3]) ? 4'b1000 : node51876;
															assign node51876 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node51880 = (inp[5]) ? 4'b1010 : node51881;
															assign node51881 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node51885 = (inp[0]) ? node51891 : node51886;
														assign node51886 = (inp[3]) ? 4'b1010 : node51887;
															assign node51887 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node51891 = (inp[5]) ? 4'b1000 : node51892;
															assign node51892 = (inp[3]) ? 4'b1000 : 4'b1010;
									assign node51896 = (inp[14]) ? node52018 : node51897;
										assign node51897 = (inp[2]) ? node51959 : node51898;
											assign node51898 = (inp[15]) ? node51928 : node51899;
												assign node51899 = (inp[0]) ? node51915 : node51900;
													assign node51900 = (inp[3]) ? node51908 : node51901;
														assign node51901 = (inp[5]) ? node51905 : node51902;
															assign node51902 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node51905 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node51908 = (inp[5]) ? node51912 : node51909;
															assign node51909 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node51912 = (inp[8]) ? 4'b1000 : 4'b1000;
													assign node51915 = (inp[5]) ? node51921 : node51916;
														assign node51916 = (inp[3]) ? node51918 : 4'b1000;
															assign node51918 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node51921 = (inp[3]) ? node51925 : node51922;
															assign node51922 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node51925 = (inp[8]) ? 4'b1010 : 4'b1010;
												assign node51928 = (inp[0]) ? node51944 : node51929;
													assign node51929 = (inp[3]) ? node51937 : node51930;
														assign node51930 = (inp[5]) ? node51934 : node51931;
															assign node51931 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node51934 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node51937 = (inp[8]) ? node51941 : node51938;
															assign node51938 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node51941 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node51944 = (inp[5]) ? node51952 : node51945;
														assign node51945 = (inp[3]) ? node51949 : node51946;
															assign node51946 = (inp[8]) ? 4'b1010 : 4'b1010;
															assign node51949 = (inp[7]) ? 4'b1000 : 4'b1000;
														assign node51952 = (inp[3]) ? node51956 : node51953;
															assign node51953 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node51956 = (inp[8]) ? 4'b1000 : 4'b1000;
											assign node51959 = (inp[8]) ? node51987 : node51960;
												assign node51960 = (inp[7]) ? node51972 : node51961;
													assign node51961 = (inp[15]) ? node51967 : node51962;
														assign node51962 = (inp[0]) ? node51964 : 4'b1000;
															assign node51964 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node51967 = (inp[0]) ? 4'b1000 : node51968;
															assign node51968 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node51972 = (inp[0]) ? node51980 : node51973;
														assign node51973 = (inp[15]) ? node51977 : node51974;
															assign node51974 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node51977 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node51980 = (inp[15]) ? node51984 : node51981;
															assign node51981 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node51984 = (inp[3]) ? 4'b1001 : 4'b1001;
												assign node51987 = (inp[7]) ? node52003 : node51988;
													assign node51988 = (inp[0]) ? node51996 : node51989;
														assign node51989 = (inp[15]) ? node51993 : node51990;
															assign node51990 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node51993 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node51996 = (inp[15]) ? node52000 : node51997;
															assign node51997 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node52000 = (inp[3]) ? 4'b1001 : 4'b1001;
													assign node52003 = (inp[3]) ? node52011 : node52004;
														assign node52004 = (inp[15]) ? node52008 : node52005;
															assign node52005 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node52008 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node52011 = (inp[5]) ? node52015 : node52012;
															assign node52012 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node52015 = (inp[0]) ? 4'b1000 : 4'b1000;
										assign node52018 = (inp[2]) ? node52082 : node52019;
											assign node52019 = (inp[3]) ? node52051 : node52020;
												assign node52020 = (inp[7]) ? node52036 : node52021;
													assign node52021 = (inp[8]) ? node52029 : node52022;
														assign node52022 = (inp[0]) ? node52026 : node52023;
															assign node52023 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node52026 = (inp[5]) ? 4'b1000 : 4'b1000;
														assign node52029 = (inp[0]) ? node52033 : node52030;
															assign node52030 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node52033 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node52036 = (inp[8]) ? node52044 : node52037;
														assign node52037 = (inp[5]) ? node52041 : node52038;
															assign node52038 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node52041 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node52044 = (inp[5]) ? node52048 : node52045;
															assign node52045 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node52048 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node52051 = (inp[15]) ? node52067 : node52052;
													assign node52052 = (inp[0]) ? node52060 : node52053;
														assign node52053 = (inp[5]) ? node52057 : node52054;
															assign node52054 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node52057 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node52060 = (inp[7]) ? node52064 : node52061;
															assign node52061 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node52064 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node52067 = (inp[0]) ? node52075 : node52068;
														assign node52068 = (inp[7]) ? node52072 : node52069;
															assign node52069 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node52072 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node52075 = (inp[8]) ? node52079 : node52076;
															assign node52076 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node52079 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node52082 = (inp[3]) ? node52114 : node52083;
												assign node52083 = (inp[5]) ? node52099 : node52084;
													assign node52084 = (inp[7]) ? node52092 : node52085;
														assign node52085 = (inp[8]) ? node52089 : node52086;
															assign node52086 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node52089 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node52092 = (inp[8]) ? node52096 : node52093;
															assign node52093 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node52096 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node52099 = (inp[15]) ? node52107 : node52100;
														assign node52100 = (inp[0]) ? node52104 : node52101;
															assign node52101 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node52104 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node52107 = (inp[0]) ? node52111 : node52108;
															assign node52108 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node52111 = (inp[8]) ? 4'b1000 : 4'b1000;
												assign node52114 = (inp[8]) ? node52130 : node52115;
													assign node52115 = (inp[7]) ? node52123 : node52116;
														assign node52116 = (inp[5]) ? node52120 : node52117;
															assign node52117 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node52120 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node52123 = (inp[5]) ? node52127 : node52124;
															assign node52124 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node52127 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node52130 = (inp[7]) ? node52138 : node52131;
														assign node52131 = (inp[5]) ? node52135 : node52132;
															assign node52132 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node52135 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node52138 = (inp[15]) ? node52142 : node52139;
															assign node52139 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node52142 = (inp[0]) ? 4'b1000 : 4'b1010;
						assign node52145 = (inp[11]) ? node53031 : node52146;
							assign node52146 = (inp[13]) ? node52572 : node52147;
								assign node52147 = (inp[1]) ? node52357 : node52148;
									assign node52148 = (inp[7]) ? node52254 : node52149;
										assign node52149 = (inp[8]) ? node52203 : node52150;
											assign node52150 = (inp[14]) ? node52180 : node52151;
												assign node52151 = (inp[2]) ? node52167 : node52152;
													assign node52152 = (inp[3]) ? node52160 : node52153;
														assign node52153 = (inp[5]) ? node52157 : node52154;
															assign node52154 = (inp[15]) ? 4'b0101 : 4'b0101;
															assign node52157 = (inp[15]) ? 4'b0101 : 4'b0101;
														assign node52160 = (inp[0]) ? node52164 : node52161;
															assign node52161 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node52164 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node52167 = (inp[0]) ? node52173 : node52168;
														assign node52168 = (inp[5]) ? 4'b0100 : node52169;
															assign node52169 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node52173 = (inp[15]) ? node52177 : node52174;
															assign node52174 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node52177 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node52180 = (inp[5]) ? node52196 : node52181;
													assign node52181 = (inp[15]) ? node52189 : node52182;
														assign node52182 = (inp[0]) ? node52186 : node52183;
															assign node52183 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node52186 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node52189 = (inp[0]) ? node52193 : node52190;
															assign node52190 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node52193 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node52196 = (inp[15]) ? node52200 : node52197;
														assign node52197 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node52200 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node52203 = (inp[14]) ? node52231 : node52204;
												assign node52204 = (inp[2]) ? node52220 : node52205;
													assign node52205 = (inp[3]) ? node52213 : node52206;
														assign node52206 = (inp[15]) ? node52210 : node52207;
															assign node52207 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node52210 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node52213 = (inp[0]) ? node52217 : node52214;
															assign node52214 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node52217 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node52220 = (inp[15]) ? node52226 : node52221;
														assign node52221 = (inp[0]) ? 4'b0111 : node52222;
															assign node52222 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node52226 = (inp[0]) ? node52228 : 4'b0111;
															assign node52228 = (inp[5]) ? 4'b0101 : 4'b0101;
												assign node52231 = (inp[15]) ? node52243 : node52232;
													assign node52232 = (inp[0]) ? node52238 : node52233;
														assign node52233 = (inp[5]) ? 4'b0101 : node52234;
															assign node52234 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node52238 = (inp[5]) ? 4'b0111 : node52239;
															assign node52239 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node52243 = (inp[0]) ? node52249 : node52244;
														assign node52244 = (inp[3]) ? 4'b0111 : node52245;
															assign node52245 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node52249 = (inp[5]) ? 4'b0101 : node52250;
															assign node52250 = (inp[3]) ? 4'b0101 : 4'b0111;
										assign node52254 = (inp[8]) ? node52306 : node52255;
											assign node52255 = (inp[14]) ? node52283 : node52256;
												assign node52256 = (inp[2]) ? node52270 : node52257;
													assign node52257 = (inp[3]) ? node52265 : node52258;
														assign node52258 = (inp[15]) ? node52262 : node52259;
															assign node52259 = (inp[0]) ? 4'b0100 : 4'b0100;
															assign node52262 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node52265 = (inp[0]) ? node52267 : 4'b0110;
															assign node52267 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node52270 = (inp[0]) ? node52276 : node52271;
														assign node52271 = (inp[15]) ? 4'b0111 : node52272;
															assign node52272 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node52276 = (inp[15]) ? node52280 : node52277;
															assign node52277 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node52280 = (inp[3]) ? 4'b0101 : 4'b0101;
												assign node52283 = (inp[15]) ? node52295 : node52284;
													assign node52284 = (inp[0]) ? node52290 : node52285;
														assign node52285 = (inp[3]) ? 4'b0101 : node52286;
															assign node52286 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node52290 = (inp[5]) ? 4'b0111 : node52291;
															assign node52291 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node52295 = (inp[0]) ? node52301 : node52296;
														assign node52296 = (inp[5]) ? 4'b0111 : node52297;
															assign node52297 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node52301 = (inp[3]) ? 4'b0101 : node52302;
															assign node52302 = (inp[5]) ? 4'b0101 : 4'b0111;
											assign node52306 = (inp[2]) ? node52334 : node52307;
												assign node52307 = (inp[14]) ? node52323 : node52308;
													assign node52308 = (inp[3]) ? node52316 : node52309;
														assign node52309 = (inp[0]) ? node52313 : node52310;
															assign node52310 = (inp[5]) ? 4'b0101 : 4'b0101;
															assign node52313 = (inp[5]) ? 4'b0101 : 4'b0101;
														assign node52316 = (inp[0]) ? node52320 : node52317;
															assign node52317 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node52320 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node52323 = (inp[0]) ? node52329 : node52324;
														assign node52324 = (inp[15]) ? node52326 : 4'b0100;
															assign node52326 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node52329 = (inp[15]) ? 4'b0100 : node52330;
															assign node52330 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node52334 = (inp[0]) ? node52346 : node52335;
													assign node52335 = (inp[15]) ? node52341 : node52336;
														assign node52336 = (inp[3]) ? 4'b0100 : node52337;
															assign node52337 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node52341 = (inp[5]) ? 4'b0110 : node52342;
															assign node52342 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node52346 = (inp[15]) ? node52352 : node52347;
														assign node52347 = (inp[5]) ? 4'b0110 : node52348;
															assign node52348 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node52352 = (inp[5]) ? 4'b0100 : node52353;
															assign node52353 = (inp[3]) ? 4'b0100 : 4'b0110;
									assign node52357 = (inp[7]) ? node52465 : node52358;
										assign node52358 = (inp[8]) ? node52416 : node52359;
											assign node52359 = (inp[2]) ? node52385 : node52360;
												assign node52360 = (inp[14]) ? node52372 : node52361;
													assign node52361 = (inp[0]) ? node52367 : node52362;
														assign node52362 = (inp[15]) ? node52364 : 4'b0101;
															assign node52364 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node52367 = (inp[15]) ? node52369 : 4'b0111;
															assign node52369 = (inp[3]) ? 4'b0101 : 4'b0101;
													assign node52372 = (inp[0]) ? node52378 : node52373;
														assign node52373 = (inp[15]) ? 4'b0110 : node52374;
															assign node52374 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node52378 = (inp[15]) ? node52382 : node52379;
															assign node52379 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node52382 = (inp[3]) ? 4'b0100 : 4'b0100;
												assign node52385 = (inp[3]) ? node52401 : node52386;
													assign node52386 = (inp[14]) ? node52394 : node52387;
														assign node52387 = (inp[15]) ? node52391 : node52388;
															assign node52388 = (inp[5]) ? 4'b0100 : 4'b0100;
															assign node52391 = (inp[5]) ? 4'b0100 : 4'b0100;
														assign node52394 = (inp[0]) ? node52398 : node52395;
															assign node52395 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node52398 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node52401 = (inp[14]) ? node52409 : node52402;
														assign node52402 = (inp[5]) ? node52406 : node52403;
															assign node52403 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node52406 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node52409 = (inp[0]) ? node52413 : node52410;
															assign node52410 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node52413 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node52416 = (inp[2]) ? node52444 : node52417;
												assign node52417 = (inp[14]) ? node52431 : node52418;
													assign node52418 = (inp[3]) ? node52424 : node52419;
														assign node52419 = (inp[5]) ? node52421 : 4'b0110;
															assign node52421 = (inp[15]) ? 4'b0100 : 4'b0100;
														assign node52424 = (inp[5]) ? node52428 : node52425;
															assign node52425 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node52428 = (inp[15]) ? 4'b0100 : 4'b0100;
													assign node52431 = (inp[15]) ? node52439 : node52432;
														assign node52432 = (inp[0]) ? node52436 : node52433;
															assign node52433 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node52436 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node52439 = (inp[0]) ? node52441 : 4'b1011;
															assign node52441 = (inp[5]) ? 4'b1001 : 4'b1001;
												assign node52444 = (inp[5]) ? node52458 : node52445;
													assign node52445 = (inp[14]) ? node52453 : node52446;
														assign node52446 = (inp[15]) ? node52450 : node52447;
															assign node52447 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node52450 = (inp[3]) ? 4'b1001 : 4'b1001;
														assign node52453 = (inp[15]) ? 4'b1001 : node52454;
															assign node52454 = (inp[3]) ? 4'b1001 : 4'b1001;
													assign node52458 = (inp[15]) ? node52462 : node52459;
														assign node52459 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node52462 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node52465 = (inp[8]) ? node52519 : node52466;
											assign node52466 = (inp[14]) ? node52496 : node52467;
												assign node52467 = (inp[2]) ? node52483 : node52468;
													assign node52468 = (inp[5]) ? node52476 : node52469;
														assign node52469 = (inp[15]) ? node52473 : node52470;
															assign node52470 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node52473 = (inp[0]) ? 4'b0100 : 4'b0100;
														assign node52476 = (inp[3]) ? node52480 : node52477;
															assign node52477 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node52480 = (inp[0]) ? 4'b0100 : 4'b0100;
													assign node52483 = (inp[3]) ? node52491 : node52484;
														assign node52484 = (inp[0]) ? node52488 : node52485;
															assign node52485 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node52488 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node52491 = (inp[0]) ? 4'b1001 : node52492;
															assign node52492 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node52496 = (inp[0]) ? node52508 : node52497;
													assign node52497 = (inp[15]) ? node52503 : node52498;
														assign node52498 = (inp[5]) ? 4'b1001 : node52499;
															assign node52499 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node52503 = (inp[3]) ? 4'b1011 : node52504;
															assign node52504 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node52508 = (inp[15]) ? node52514 : node52509;
														assign node52509 = (inp[3]) ? 4'b1011 : node52510;
															assign node52510 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node52514 = (inp[3]) ? 4'b1001 : node52515;
															assign node52515 = (inp[2]) ? 4'b1011 : 4'b1001;
											assign node52519 = (inp[14]) ? node52549 : node52520;
												assign node52520 = (inp[2]) ? node52536 : node52521;
													assign node52521 = (inp[15]) ? node52529 : node52522;
														assign node52522 = (inp[0]) ? node52526 : node52523;
															assign node52523 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node52526 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node52529 = (inp[0]) ? node52533 : node52530;
															assign node52530 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node52533 = (inp[3]) ? 4'b1001 : 4'b1001;
													assign node52536 = (inp[15]) ? node52544 : node52537;
														assign node52537 = (inp[0]) ? node52541 : node52538;
															assign node52538 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node52541 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node52544 = (inp[5]) ? 4'b1000 : node52545;
															assign node52545 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node52549 = (inp[15]) ? node52561 : node52550;
													assign node52550 = (inp[0]) ? node52556 : node52551;
														assign node52551 = (inp[5]) ? 4'b1000 : node52552;
															assign node52552 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node52556 = (inp[3]) ? 4'b1010 : node52557;
															assign node52557 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node52561 = (inp[0]) ? node52567 : node52562;
														assign node52562 = (inp[5]) ? 4'b1010 : node52563;
															assign node52563 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node52567 = (inp[5]) ? 4'b1000 : node52568;
															assign node52568 = (inp[3]) ? 4'b1000 : 4'b1010;
								assign node52572 = (inp[1]) ? node52800 : node52573;
									assign node52573 = (inp[7]) ? node52687 : node52574;
										assign node52574 = (inp[8]) ? node52628 : node52575;
											assign node52575 = (inp[2]) ? node52605 : node52576;
												assign node52576 = (inp[14]) ? node52590 : node52577;
													assign node52577 = (inp[0]) ? node52585 : node52578;
														assign node52578 = (inp[15]) ? node52582 : node52579;
															assign node52579 = (inp[3]) ? 4'b0101 : 4'b0101;
															assign node52582 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node52585 = (inp[15]) ? node52587 : 4'b0111;
															assign node52587 = (inp[3]) ? 4'b0101 : 4'b0101;
													assign node52590 = (inp[0]) ? node52598 : node52591;
														assign node52591 = (inp[15]) ? node52595 : node52592;
															assign node52592 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node52595 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node52598 = (inp[15]) ? node52602 : node52599;
															assign node52599 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node52602 = (inp[3]) ? 4'b0100 : 4'b0100;
												assign node52605 = (inp[3]) ? node52621 : node52606;
													assign node52606 = (inp[5]) ? node52614 : node52607;
														assign node52607 = (inp[0]) ? node52611 : node52608;
															assign node52608 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node52611 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node52614 = (inp[15]) ? node52618 : node52615;
															assign node52615 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node52618 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node52621 = (inp[0]) ? node52625 : node52622;
														assign node52622 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node52625 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node52628 = (inp[2]) ? node52658 : node52629;
												assign node52629 = (inp[14]) ? node52645 : node52630;
													assign node52630 = (inp[5]) ? node52638 : node52631;
														assign node52631 = (inp[0]) ? node52635 : node52632;
															assign node52632 = (inp[3]) ? 4'b0100 : 4'b0100;
															assign node52635 = (inp[3]) ? 4'b0100 : 4'b0100;
														assign node52638 = (inp[0]) ? node52642 : node52639;
															assign node52639 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node52642 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node52645 = (inp[15]) ? node52651 : node52646;
														assign node52646 = (inp[0]) ? 4'b1011 : node52647;
															assign node52647 = (inp[5]) ? 4'b1001 : 4'b1001;
														assign node52651 = (inp[0]) ? node52655 : node52652;
															assign node52652 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node52655 = (inp[5]) ? 4'b1001 : 4'b1001;
												assign node52658 = (inp[14]) ? node52674 : node52659;
													assign node52659 = (inp[0]) ? node52667 : node52660;
														assign node52660 = (inp[15]) ? node52664 : node52661;
															assign node52661 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node52664 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node52667 = (inp[15]) ? node52671 : node52668;
															assign node52668 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node52671 = (inp[3]) ? 4'b1001 : 4'b1001;
													assign node52674 = (inp[0]) ? node52680 : node52675;
														assign node52675 = (inp[15]) ? node52677 : 4'b1001;
															assign node52677 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node52680 = (inp[15]) ? node52684 : node52681;
															assign node52681 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node52684 = (inp[3]) ? 4'b1001 : 4'b1001;
										assign node52687 = (inp[8]) ? node52739 : node52688;
											assign node52688 = (inp[14]) ? node52716 : node52689;
												assign node52689 = (inp[2]) ? node52703 : node52690;
													assign node52690 = (inp[5]) ? node52696 : node52691;
														assign node52691 = (inp[15]) ? 4'b0110 : node52692;
															assign node52692 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node52696 = (inp[3]) ? node52700 : node52697;
															assign node52697 = (inp[15]) ? 4'b0100 : 4'b0100;
															assign node52700 = (inp[0]) ? 4'b0100 : 4'b0100;
													assign node52703 = (inp[15]) ? node52711 : node52704;
														assign node52704 = (inp[0]) ? node52708 : node52705;
															assign node52705 = (inp[5]) ? 4'b1001 : 4'b1001;
															assign node52708 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node52711 = (inp[5]) ? 4'b1011 : node52712;
															assign node52712 = (inp[0]) ? 4'b1001 : 4'b1001;
												assign node52716 = (inp[0]) ? node52728 : node52717;
													assign node52717 = (inp[15]) ? node52723 : node52718;
														assign node52718 = (inp[5]) ? 4'b1001 : node52719;
															assign node52719 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node52723 = (inp[3]) ? 4'b1011 : node52724;
															assign node52724 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node52728 = (inp[15]) ? node52734 : node52729;
														assign node52729 = (inp[3]) ? 4'b1011 : node52730;
															assign node52730 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node52734 = (inp[5]) ? 4'b1001 : node52735;
															assign node52735 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node52739 = (inp[2]) ? node52769 : node52740;
												assign node52740 = (inp[14]) ? node52754 : node52741;
													assign node52741 = (inp[0]) ? node52749 : node52742;
														assign node52742 = (inp[15]) ? node52746 : node52743;
															assign node52743 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node52746 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node52749 = (inp[15]) ? 4'b1001 : node52750;
															assign node52750 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node52754 = (inp[5]) ? node52762 : node52755;
														assign node52755 = (inp[0]) ? node52759 : node52756;
															assign node52756 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node52759 = (inp[3]) ? 4'b1000 : 4'b1000;
														assign node52762 = (inp[0]) ? node52766 : node52763;
															assign node52763 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node52766 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node52769 = (inp[3]) ? node52785 : node52770;
													assign node52770 = (inp[0]) ? node52778 : node52771;
														assign node52771 = (inp[5]) ? node52775 : node52772;
															assign node52772 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node52775 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node52778 = (inp[14]) ? node52782 : node52779;
															assign node52779 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node52782 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node52785 = (inp[5]) ? node52793 : node52786;
														assign node52786 = (inp[0]) ? node52790 : node52787;
															assign node52787 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node52790 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node52793 = (inp[15]) ? node52797 : node52794;
															assign node52794 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node52797 = (inp[0]) ? 4'b1000 : 4'b1010;
									assign node52800 = (inp[3]) ? node52924 : node52801;
										assign node52801 = (inp[5]) ? node52861 : node52802;
											assign node52802 = (inp[0]) ? node52830 : node52803;
												assign node52803 = (inp[15]) ? node52817 : node52804;
													assign node52804 = (inp[7]) ? node52812 : node52805;
														assign node52805 = (inp[8]) ? node52809 : node52806;
															assign node52806 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node52809 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node52812 = (inp[8]) ? 4'b1010 : node52813;
															assign node52813 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node52817 = (inp[2]) ? node52823 : node52818;
														assign node52818 = (inp[14]) ? 4'b1000 : node52819;
															assign node52819 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node52823 = (inp[7]) ? node52827 : node52824;
															assign node52824 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node52827 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node52830 = (inp[15]) ? node52846 : node52831;
													assign node52831 = (inp[7]) ? node52839 : node52832;
														assign node52832 = (inp[8]) ? node52836 : node52833;
															assign node52833 = (inp[2]) ? 4'b1000 : 4'b1000;
															assign node52836 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node52839 = (inp[8]) ? node52843 : node52840;
															assign node52840 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node52843 = (inp[2]) ? 4'b1000 : 4'b1000;
													assign node52846 = (inp[14]) ? node52854 : node52847;
														assign node52847 = (inp[7]) ? node52851 : node52848;
															assign node52848 = (inp[8]) ? 4'b1010 : 4'b1010;
															assign node52851 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node52854 = (inp[7]) ? node52858 : node52855;
															assign node52855 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node52858 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node52861 = (inp[15]) ? node52893 : node52862;
												assign node52862 = (inp[0]) ? node52878 : node52863;
													assign node52863 = (inp[2]) ? node52871 : node52864;
														assign node52864 = (inp[14]) ? node52868 : node52865;
															assign node52865 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node52868 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node52871 = (inp[14]) ? node52875 : node52872;
															assign node52872 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node52875 = (inp[7]) ? 4'b1000 : 4'b1000;
													assign node52878 = (inp[2]) ? node52886 : node52879;
														assign node52879 = (inp[14]) ? node52883 : node52880;
															assign node52880 = (inp[8]) ? 4'b1010 : 4'b1010;
															assign node52883 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node52886 = (inp[8]) ? node52890 : node52887;
															assign node52887 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node52890 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node52893 = (inp[0]) ? node52909 : node52894;
													assign node52894 = (inp[14]) ? node52902 : node52895;
														assign node52895 = (inp[8]) ? node52899 : node52896;
															assign node52896 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node52899 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node52902 = (inp[7]) ? node52906 : node52903;
															assign node52903 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node52906 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node52909 = (inp[2]) ? node52917 : node52910;
														assign node52910 = (inp[14]) ? node52914 : node52911;
															assign node52911 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node52914 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node52917 = (inp[14]) ? node52921 : node52918;
															assign node52918 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node52921 = (inp[7]) ? 4'b1000 : 4'b1000;
										assign node52924 = (inp[7]) ? node52970 : node52925;
											assign node52925 = (inp[8]) ? node52949 : node52926;
												assign node52926 = (inp[2]) ? node52942 : node52927;
													assign node52927 = (inp[14]) ? node52935 : node52928;
														assign node52928 = (inp[5]) ? node52932 : node52929;
															assign node52929 = (inp[15]) ? 4'b1001 : 4'b1001;
															assign node52932 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node52935 = (inp[15]) ? node52939 : node52936;
															assign node52936 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node52939 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node52942 = (inp[0]) ? node52946 : node52943;
														assign node52943 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node52946 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node52949 = (inp[2]) ? node52963 : node52950;
													assign node52950 = (inp[14]) ? node52956 : node52951;
														assign node52951 = (inp[0]) ? node52953 : 4'b1010;
															assign node52953 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node52956 = (inp[5]) ? node52960 : node52957;
															assign node52957 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node52960 = (inp[15]) ? 4'b1001 : 4'b1001;
													assign node52963 = (inp[0]) ? node52967 : node52964;
														assign node52964 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node52967 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node52970 = (inp[8]) ? node53000 : node52971;
												assign node52971 = (inp[2]) ? node52985 : node52972;
													assign node52972 = (inp[14]) ? node52980 : node52973;
														assign node52973 = (inp[0]) ? node52977 : node52974;
															assign node52974 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node52977 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node52980 = (inp[0]) ? node52982 : 4'b1011;
															assign node52982 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node52985 = (inp[14]) ? node52993 : node52986;
														assign node52986 = (inp[0]) ? node52990 : node52987;
															assign node52987 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node52990 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node52993 = (inp[0]) ? node52997 : node52994;
															assign node52994 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node52997 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node53000 = (inp[2]) ? node53016 : node53001;
													assign node53001 = (inp[14]) ? node53009 : node53002;
														assign node53002 = (inp[0]) ? node53006 : node53003;
															assign node53003 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node53006 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node53009 = (inp[5]) ? node53013 : node53010;
															assign node53010 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node53013 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node53016 = (inp[5]) ? node53024 : node53017;
														assign node53017 = (inp[15]) ? node53021 : node53018;
															assign node53018 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node53021 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node53024 = (inp[0]) ? node53028 : node53025;
															assign node53025 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node53028 = (inp[15]) ? 4'b1000 : 4'b1010;
							assign node53031 = (inp[13]) ? node53469 : node53032;
								assign node53032 = (inp[1]) ? node53254 : node53033;
									assign node53033 = (inp[15]) ? node53149 : node53034;
										assign node53034 = (inp[0]) ? node53094 : node53035;
											assign node53035 = (inp[5]) ? node53065 : node53036;
												assign node53036 = (inp[3]) ? node53050 : node53037;
													assign node53037 = (inp[14]) ? node53043 : node53038;
														assign node53038 = (inp[2]) ? 4'b1011 : node53039;
															assign node53039 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node53043 = (inp[7]) ? node53047 : node53044;
															assign node53044 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node53047 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node53050 = (inp[7]) ? node53058 : node53051;
														assign node53051 = (inp[8]) ? node53055 : node53052;
															assign node53052 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node53055 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node53058 = (inp[8]) ? node53062 : node53059;
															assign node53059 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node53062 = (inp[14]) ? 4'b1000 : 4'b1000;
												assign node53065 = (inp[3]) ? node53081 : node53066;
													assign node53066 = (inp[7]) ? node53074 : node53067;
														assign node53067 = (inp[8]) ? node53071 : node53068;
															assign node53068 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node53071 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node53074 = (inp[8]) ? node53078 : node53075;
															assign node53075 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node53078 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node53081 = (inp[2]) ? node53087 : node53082;
														assign node53082 = (inp[7]) ? node53084 : 4'b1000;
															assign node53084 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node53087 = (inp[8]) ? node53091 : node53088;
															assign node53088 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node53091 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node53094 = (inp[5]) ? node53120 : node53095;
												assign node53095 = (inp[3]) ? node53111 : node53096;
													assign node53096 = (inp[7]) ? node53104 : node53097;
														assign node53097 = (inp[8]) ? node53101 : node53098;
															assign node53098 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node53101 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node53104 = (inp[8]) ? node53108 : node53105;
															assign node53105 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node53108 = (inp[2]) ? 4'b1000 : 4'b1000;
													assign node53111 = (inp[7]) ? node53117 : node53112;
														assign node53112 = (inp[8]) ? 4'b1011 : node53113;
															assign node53113 = (inp[2]) ? 4'b1010 : 4'b1010;
														assign node53117 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node53120 = (inp[2]) ? node53134 : node53121;
													assign node53121 = (inp[14]) ? node53127 : node53122;
														assign node53122 = (inp[3]) ? node53124 : 4'b1011;
															assign node53124 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node53127 = (inp[8]) ? node53131 : node53128;
															assign node53128 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node53131 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node53134 = (inp[3]) ? node53142 : node53135;
														assign node53135 = (inp[14]) ? node53139 : node53136;
															assign node53136 = (inp[8]) ? 4'b1010 : 4'b1010;
															assign node53139 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node53142 = (inp[7]) ? node53146 : node53143;
															assign node53143 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node53146 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node53149 = (inp[0]) ? node53203 : node53150;
											assign node53150 = (inp[5]) ? node53180 : node53151;
												assign node53151 = (inp[3]) ? node53165 : node53152;
													assign node53152 = (inp[14]) ? node53158 : node53153;
														assign node53153 = (inp[8]) ? 4'b1001 : node53154;
															assign node53154 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node53158 = (inp[8]) ? node53162 : node53159;
															assign node53159 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node53162 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node53165 = (inp[2]) ? node53173 : node53166;
														assign node53166 = (inp[14]) ? node53170 : node53167;
															assign node53167 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node53170 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node53173 = (inp[8]) ? node53177 : node53174;
															assign node53174 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node53177 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node53180 = (inp[8]) ? node53192 : node53181;
													assign node53181 = (inp[7]) ? node53187 : node53182;
														assign node53182 = (inp[2]) ? 4'b1010 : node53183;
															assign node53183 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node53187 = (inp[14]) ? 4'b1011 : node53188;
															assign node53188 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node53192 = (inp[7]) ? node53198 : node53193;
														assign node53193 = (inp[14]) ? 4'b1011 : node53194;
															assign node53194 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node53198 = (inp[14]) ? 4'b1010 : node53199;
															assign node53199 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node53203 = (inp[5]) ? node53231 : node53204;
												assign node53204 = (inp[3]) ? node53218 : node53205;
													assign node53205 = (inp[14]) ? node53211 : node53206;
														assign node53206 = (inp[7]) ? 4'b1011 : node53207;
															assign node53207 = (inp[2]) ? 4'b1010 : 4'b1010;
														assign node53211 = (inp[2]) ? node53215 : node53212;
															assign node53212 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node53215 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node53218 = (inp[2]) ? node53224 : node53219;
														assign node53219 = (inp[8]) ? 4'b1001 : node53220;
															assign node53220 = (inp[7]) ? 4'b1000 : 4'b1000;
														assign node53224 = (inp[8]) ? node53228 : node53225;
															assign node53225 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node53228 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node53231 = (inp[7]) ? node53243 : node53232;
													assign node53232 = (inp[8]) ? node53238 : node53233;
														assign node53233 = (inp[14]) ? 4'b1000 : node53234;
															assign node53234 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node53238 = (inp[2]) ? 4'b1001 : node53239;
															assign node53239 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node53243 = (inp[8]) ? node53249 : node53244;
														assign node53244 = (inp[2]) ? 4'b1001 : node53245;
															assign node53245 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node53249 = (inp[2]) ? 4'b1000 : node53250;
															assign node53250 = (inp[14]) ? 4'b1000 : 4'b1001;
									assign node53254 = (inp[8]) ? node53372 : node53255;
										assign node53255 = (inp[7]) ? node53311 : node53256;
											assign node53256 = (inp[14]) ? node53284 : node53257;
												assign node53257 = (inp[2]) ? node53271 : node53258;
													assign node53258 = (inp[5]) ? node53264 : node53259;
														assign node53259 = (inp[0]) ? node53261 : 4'b1011;
															assign node53261 = (inp[15]) ? 4'b1001 : 4'b1001;
														assign node53264 = (inp[15]) ? node53268 : node53265;
															assign node53265 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node53268 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node53271 = (inp[5]) ? node53279 : node53272;
														assign node53272 = (inp[15]) ? node53276 : node53273;
															assign node53273 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node53276 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node53279 = (inp[3]) ? node53281 : 4'b1000;
															assign node53281 = (inp[0]) ? 4'b1000 : 4'b1000;
												assign node53284 = (inp[2]) ? node53298 : node53285;
													assign node53285 = (inp[15]) ? node53293 : node53286;
														assign node53286 = (inp[0]) ? node53290 : node53287;
															assign node53287 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node53290 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node53293 = (inp[0]) ? 4'b1000 : node53294;
															assign node53294 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node53298 = (inp[0]) ? node53306 : node53299;
														assign node53299 = (inp[15]) ? node53303 : node53300;
															assign node53300 = (inp[3]) ? 4'b1000 : 4'b1000;
															assign node53303 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node53306 = (inp[15]) ? node53308 : 4'b1010;
															assign node53308 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node53311 = (inp[14]) ? node53341 : node53312;
												assign node53312 = (inp[2]) ? node53328 : node53313;
													assign node53313 = (inp[5]) ? node53321 : node53314;
														assign node53314 = (inp[3]) ? node53318 : node53315;
															assign node53315 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node53318 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node53321 = (inp[0]) ? node53325 : node53322;
															assign node53322 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node53325 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node53328 = (inp[15]) ? node53334 : node53329;
														assign node53329 = (inp[0]) ? 4'b0011 : node53330;
															assign node53330 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node53334 = (inp[0]) ? node53338 : node53335;
															assign node53335 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node53338 = (inp[3]) ? 4'b0001 : 4'b0001;
												assign node53341 = (inp[5]) ? node53357 : node53342;
													assign node53342 = (inp[3]) ? node53350 : node53343;
														assign node53343 = (inp[15]) ? node53347 : node53344;
															assign node53344 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node53347 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node53350 = (inp[0]) ? node53354 : node53351;
															assign node53351 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node53354 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node53357 = (inp[2]) ? node53365 : node53358;
														assign node53358 = (inp[3]) ? node53362 : node53359;
															assign node53359 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node53362 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node53365 = (inp[3]) ? node53369 : node53366;
															assign node53366 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node53369 = (inp[0]) ? 4'b0001 : 4'b0001;
										assign node53372 = (inp[7]) ? node53426 : node53373;
											assign node53373 = (inp[2]) ? node53403 : node53374;
												assign node53374 = (inp[14]) ? node53390 : node53375;
													assign node53375 = (inp[3]) ? node53383 : node53376;
														assign node53376 = (inp[5]) ? node53380 : node53377;
															assign node53377 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node53380 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node53383 = (inp[5]) ? node53387 : node53384;
															assign node53384 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node53387 = (inp[15]) ? 4'b1000 : 4'b1000;
													assign node53390 = (inp[3]) ? node53396 : node53391;
														assign node53391 = (inp[15]) ? node53393 : 4'b0001;
															assign node53393 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node53396 = (inp[0]) ? node53400 : node53397;
															assign node53397 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node53400 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node53403 = (inp[15]) ? node53415 : node53404;
													assign node53404 = (inp[0]) ? node53410 : node53405;
														assign node53405 = (inp[3]) ? 4'b0001 : node53406;
															assign node53406 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node53410 = (inp[5]) ? 4'b0011 : node53411;
															assign node53411 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node53415 = (inp[0]) ? node53421 : node53416;
														assign node53416 = (inp[5]) ? 4'b0011 : node53417;
															assign node53417 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node53421 = (inp[5]) ? 4'b0001 : node53422;
															assign node53422 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node53426 = (inp[2]) ? node53450 : node53427;
												assign node53427 = (inp[14]) ? node53437 : node53428;
													assign node53428 = (inp[0]) ? node53432 : node53429;
														assign node53429 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node53432 = (inp[15]) ? 4'b0001 : node53433;
															assign node53433 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node53437 = (inp[15]) ? node53445 : node53438;
														assign node53438 = (inp[0]) ? node53442 : node53439;
															assign node53439 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node53442 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node53445 = (inp[0]) ? node53447 : 4'b0010;
															assign node53447 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node53450 = (inp[15]) ? node53458 : node53451;
													assign node53451 = (inp[0]) ? 4'b0010 : node53452;
														assign node53452 = (inp[5]) ? 4'b0000 : node53453;
															assign node53453 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node53458 = (inp[0]) ? node53464 : node53459;
														assign node53459 = (inp[5]) ? 4'b0010 : node53460;
															assign node53460 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node53464 = (inp[3]) ? 4'b0000 : node53465;
															assign node53465 = (inp[5]) ? 4'b0000 : 4'b0010;
								assign node53469 = (inp[1]) ? node53693 : node53470;
									assign node53470 = (inp[7]) ? node53576 : node53471;
										assign node53471 = (inp[8]) ? node53525 : node53472;
											assign node53472 = (inp[2]) ? node53502 : node53473;
												assign node53473 = (inp[14]) ? node53487 : node53474;
													assign node53474 = (inp[0]) ? node53480 : node53475;
														assign node53475 = (inp[15]) ? node53477 : 4'b1001;
															assign node53477 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node53480 = (inp[15]) ? node53484 : node53481;
															assign node53481 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node53484 = (inp[5]) ? 4'b1001 : 4'b1001;
													assign node53487 = (inp[0]) ? node53495 : node53488;
														assign node53488 = (inp[15]) ? node53492 : node53489;
															assign node53489 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node53492 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node53495 = (inp[15]) ? node53499 : node53496;
															assign node53496 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node53499 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node53502 = (inp[15]) ? node53514 : node53503;
													assign node53503 = (inp[0]) ? node53509 : node53504;
														assign node53504 = (inp[5]) ? 4'b1000 : node53505;
															assign node53505 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node53509 = (inp[3]) ? 4'b1010 : node53510;
															assign node53510 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node53514 = (inp[0]) ? node53520 : node53515;
														assign node53515 = (inp[5]) ? 4'b1010 : node53516;
															assign node53516 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node53520 = (inp[5]) ? 4'b1000 : node53521;
															assign node53521 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node53525 = (inp[2]) ? node53553 : node53526;
												assign node53526 = (inp[14]) ? node53542 : node53527;
													assign node53527 = (inp[0]) ? node53535 : node53528;
														assign node53528 = (inp[15]) ? node53532 : node53529;
															assign node53529 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node53532 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node53535 = (inp[3]) ? node53539 : node53536;
															assign node53536 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node53539 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node53542 = (inp[0]) ? node53548 : node53543;
														assign node53543 = (inp[15]) ? node53545 : 4'b0001;
															assign node53545 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node53548 = (inp[15]) ? node53550 : 4'b0011;
															assign node53550 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node53553 = (inp[15]) ? node53565 : node53554;
													assign node53554 = (inp[0]) ? node53560 : node53555;
														assign node53555 = (inp[5]) ? 4'b0001 : node53556;
															assign node53556 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node53560 = (inp[5]) ? 4'b0011 : node53561;
															assign node53561 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node53565 = (inp[0]) ? node53571 : node53566;
														assign node53566 = (inp[5]) ? 4'b0011 : node53567;
															assign node53567 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node53571 = (inp[3]) ? 4'b0001 : node53572;
															assign node53572 = (inp[5]) ? 4'b0001 : 4'b0011;
										assign node53576 = (inp[8]) ? node53636 : node53577;
											assign node53577 = (inp[14]) ? node53605 : node53578;
												assign node53578 = (inp[2]) ? node53592 : node53579;
													assign node53579 = (inp[15]) ? node53587 : node53580;
														assign node53580 = (inp[0]) ? node53584 : node53581;
															assign node53581 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node53584 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node53587 = (inp[0]) ? node53589 : 4'b1010;
															assign node53589 = (inp[3]) ? 4'b1000 : 4'b1000;
													assign node53592 = (inp[15]) ? node53600 : node53593;
														assign node53593 = (inp[0]) ? node53597 : node53594;
															assign node53594 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node53597 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node53600 = (inp[0]) ? node53602 : 4'b0011;
															assign node53602 = (inp[3]) ? 4'b0001 : 4'b0001;
												assign node53605 = (inp[2]) ? node53621 : node53606;
													assign node53606 = (inp[0]) ? node53614 : node53607;
														assign node53607 = (inp[15]) ? node53611 : node53608;
															assign node53608 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node53611 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node53614 = (inp[15]) ? node53618 : node53615;
															assign node53615 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node53618 = (inp[5]) ? 4'b0001 : 4'b0001;
													assign node53621 = (inp[5]) ? node53629 : node53622;
														assign node53622 = (inp[3]) ? node53626 : node53623;
															assign node53623 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node53626 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node53629 = (inp[3]) ? node53633 : node53630;
															assign node53630 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node53633 = (inp[0]) ? 4'b0001 : 4'b0001;
											assign node53636 = (inp[2]) ? node53664 : node53637;
												assign node53637 = (inp[14]) ? node53651 : node53638;
													assign node53638 = (inp[0]) ? node53644 : node53639;
														assign node53639 = (inp[15]) ? 4'b0011 : node53640;
															assign node53640 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node53644 = (inp[15]) ? node53648 : node53645;
															assign node53645 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node53648 = (inp[5]) ? 4'b0001 : 4'b0001;
													assign node53651 = (inp[0]) ? node53659 : node53652;
														assign node53652 = (inp[15]) ? node53656 : node53653;
															assign node53653 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node53656 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node53659 = (inp[15]) ? 4'b0000 : node53660;
															assign node53660 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node53664 = (inp[5]) ? node53678 : node53665;
													assign node53665 = (inp[14]) ? node53673 : node53666;
														assign node53666 = (inp[0]) ? node53670 : node53667;
															assign node53667 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node53670 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node53673 = (inp[15]) ? node53675 : 4'b0010;
															assign node53675 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node53678 = (inp[14]) ? node53686 : node53679;
														assign node53679 = (inp[15]) ? node53683 : node53680;
															assign node53680 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node53683 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node53686 = (inp[3]) ? node53690 : node53687;
															assign node53687 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node53690 = (inp[15]) ? 4'b0000 : 4'b0000;
									assign node53693 = (inp[3]) ? node53813 : node53694;
										assign node53694 = (inp[15]) ? node53750 : node53695;
											assign node53695 = (inp[7]) ? node53719 : node53696;
												assign node53696 = (inp[8]) ? node53706 : node53697;
													assign node53697 = (inp[5]) ? node53703 : node53698;
														assign node53698 = (inp[0]) ? node53700 : 4'b0010;
															assign node53700 = (inp[2]) ? 4'b0000 : 4'b0000;
														assign node53703 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node53706 = (inp[14]) ? node53714 : node53707;
														assign node53707 = (inp[2]) ? node53711 : node53708;
															assign node53708 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node53711 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node53714 = (inp[2]) ? 4'b0001 : node53715;
															assign node53715 = (inp[0]) ? 4'b0001 : 4'b0001;
												assign node53719 = (inp[8]) ? node53735 : node53720;
													assign node53720 = (inp[14]) ? node53728 : node53721;
														assign node53721 = (inp[2]) ? node53725 : node53722;
															assign node53722 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node53725 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node53728 = (inp[0]) ? node53732 : node53729;
															assign node53729 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node53732 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node53735 = (inp[2]) ? node53743 : node53736;
														assign node53736 = (inp[14]) ? node53740 : node53737;
															assign node53737 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node53740 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node53743 = (inp[5]) ? node53747 : node53744;
															assign node53744 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node53747 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node53750 = (inp[14]) ? node53782 : node53751;
												assign node53751 = (inp[0]) ? node53767 : node53752;
													assign node53752 = (inp[5]) ? node53760 : node53753;
														assign node53753 = (inp[2]) ? node53757 : node53754;
															assign node53754 = (inp[7]) ? 4'b0000 : 4'b0000;
															assign node53757 = (inp[7]) ? 4'b0000 : 4'b0000;
														assign node53760 = (inp[2]) ? node53764 : node53761;
															assign node53761 = (inp[7]) ? 4'b0010 : 4'b0010;
															assign node53764 = (inp[8]) ? 4'b0010 : 4'b0010;
													assign node53767 = (inp[5]) ? node53775 : node53768;
														assign node53768 = (inp[2]) ? node53772 : node53769;
															assign node53769 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node53772 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node53775 = (inp[7]) ? node53779 : node53776;
															assign node53776 = (inp[2]) ? 4'b0000 : 4'b0000;
															assign node53779 = (inp[2]) ? 4'b0000 : 4'b0000;
												assign node53782 = (inp[8]) ? node53798 : node53783;
													assign node53783 = (inp[7]) ? node53791 : node53784;
														assign node53784 = (inp[2]) ? node53788 : node53785;
															assign node53785 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node53788 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node53791 = (inp[5]) ? node53795 : node53792;
															assign node53792 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node53795 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node53798 = (inp[7]) ? node53806 : node53799;
														assign node53799 = (inp[5]) ? node53803 : node53800;
															assign node53800 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node53803 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node53806 = (inp[5]) ? node53810 : node53807;
															assign node53807 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node53810 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node53813 = (inp[0]) ? node53875 : node53814;
											assign node53814 = (inp[15]) ? node53844 : node53815;
												assign node53815 = (inp[5]) ? node53831 : node53816;
													assign node53816 = (inp[2]) ? node53824 : node53817;
														assign node53817 = (inp[7]) ? node53821 : node53818;
															assign node53818 = (inp[14]) ? 4'b0000 : 4'b0000;
															assign node53821 = (inp[14]) ? 4'b0000 : 4'b0000;
														assign node53824 = (inp[7]) ? node53828 : node53825;
															assign node53825 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node53828 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node53831 = (inp[14]) ? node53837 : node53832;
														assign node53832 = (inp[7]) ? node53834 : 4'b0001;
															assign node53834 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node53837 = (inp[8]) ? node53841 : node53838;
															assign node53838 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node53841 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node53844 = (inp[14]) ? node53860 : node53845;
													assign node53845 = (inp[5]) ? node53853 : node53846;
														assign node53846 = (inp[7]) ? node53850 : node53847;
															assign node53847 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node53850 = (inp[2]) ? 4'b0010 : 4'b0010;
														assign node53853 = (inp[8]) ? node53857 : node53854;
															assign node53854 = (inp[2]) ? 4'b0010 : 4'b0010;
															assign node53857 = (inp[7]) ? 4'b0010 : 4'b0010;
													assign node53860 = (inp[2]) ? node53868 : node53861;
														assign node53861 = (inp[7]) ? node53865 : node53862;
															assign node53862 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node53865 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node53868 = (inp[5]) ? node53872 : node53869;
															assign node53869 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node53872 = (inp[7]) ? 4'b0011 : 4'b0010;
											assign node53875 = (inp[15]) ? node53907 : node53876;
												assign node53876 = (inp[5]) ? node53892 : node53877;
													assign node53877 = (inp[8]) ? node53885 : node53878;
														assign node53878 = (inp[7]) ? node53882 : node53879;
															assign node53879 = (inp[14]) ? 4'b0010 : 4'b0010;
															assign node53882 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node53885 = (inp[7]) ? node53889 : node53886;
															assign node53886 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node53889 = (inp[14]) ? 4'b0010 : 4'b0010;
													assign node53892 = (inp[7]) ? node53900 : node53893;
														assign node53893 = (inp[8]) ? node53897 : node53894;
															assign node53894 = (inp[2]) ? 4'b0010 : 4'b0010;
															assign node53897 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node53900 = (inp[8]) ? node53904 : node53901;
															assign node53901 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node53904 = (inp[14]) ? 4'b0010 : 4'b0010;
												assign node53907 = (inp[5]) ? node53921 : node53908;
													assign node53908 = (inp[14]) ? node53914 : node53909;
														assign node53909 = (inp[8]) ? node53911 : 4'b0000;
															assign node53911 = (inp[2]) ? 4'b0000 : 4'b0000;
														assign node53914 = (inp[7]) ? node53918 : node53915;
															assign node53915 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node53918 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node53921 = (inp[2]) ? node53927 : node53922;
														assign node53922 = (inp[8]) ? node53924 : 4'b0000;
															assign node53924 = (inp[7]) ? 4'b0000 : 4'b0000;
														assign node53927 = (inp[14]) ? node53931 : node53928;
															assign node53928 = (inp[8]) ? 4'b0000 : 4'b0000;
															assign node53931 = (inp[8]) ? 4'b0000 : 4'b0000;
					assign node53934 = (inp[13]) ? node55756 : node53935;
						assign node53935 = (inp[1]) ? node54829 : node53936;
							assign node53936 = (inp[6]) ? node54386 : node53937;
								assign node53937 = (inp[11]) ? node54159 : node53938;
									assign node53938 = (inp[0]) ? node54060 : node53939;
										assign node53939 = (inp[15]) ? node54003 : node53940;
											assign node53940 = (inp[5]) ? node53972 : node53941;
												assign node53941 = (inp[3]) ? node53957 : node53942;
													assign node53942 = (inp[2]) ? node53950 : node53943;
														assign node53943 = (inp[7]) ? node53947 : node53944;
															assign node53944 = (inp[14]) ? 4'b1010 : 4'b1011;
															assign node53947 = (inp[8]) ? 4'b1010 : 4'b1010;
														assign node53950 = (inp[14]) ? node53954 : node53951;
															assign node53951 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node53954 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node53957 = (inp[14]) ? node53965 : node53958;
														assign node53958 = (inp[8]) ? node53962 : node53959;
															assign node53959 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node53962 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node53965 = (inp[8]) ? node53969 : node53966;
															assign node53966 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node53969 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node53972 = (inp[2]) ? node53988 : node53973;
													assign node53973 = (inp[14]) ? node53981 : node53974;
														assign node53974 = (inp[3]) ? node53978 : node53975;
															assign node53975 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node53978 = (inp[7]) ? 4'b1000 : 4'b1000;
														assign node53981 = (inp[7]) ? node53985 : node53982;
															assign node53982 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node53985 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node53988 = (inp[3]) ? node53996 : node53989;
														assign node53989 = (inp[7]) ? node53993 : node53990;
															assign node53990 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node53993 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node53996 = (inp[7]) ? node54000 : node53997;
															assign node53997 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node54000 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node54003 = (inp[5]) ? node54031 : node54004;
												assign node54004 = (inp[3]) ? node54018 : node54005;
													assign node54005 = (inp[2]) ? node54011 : node54006;
														assign node54006 = (inp[7]) ? 4'b1000 : node54007;
															assign node54007 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node54011 = (inp[7]) ? node54015 : node54012;
															assign node54012 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node54015 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node54018 = (inp[14]) ? node54024 : node54019;
														assign node54019 = (inp[2]) ? node54021 : 4'b1011;
															assign node54021 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node54024 = (inp[7]) ? node54028 : node54025;
															assign node54025 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node54028 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node54031 = (inp[14]) ? node54045 : node54032;
													assign node54032 = (inp[2]) ? node54040 : node54033;
														assign node54033 = (inp[8]) ? node54037 : node54034;
															assign node54034 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node54037 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node54040 = (inp[7]) ? node54042 : 4'b1010;
															assign node54042 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node54045 = (inp[3]) ? node54053 : node54046;
														assign node54046 = (inp[7]) ? node54050 : node54047;
															assign node54047 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node54050 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node54053 = (inp[7]) ? node54057 : node54054;
															assign node54054 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node54057 = (inp[8]) ? 4'b1010 : 4'b1011;
										assign node54060 = (inp[15]) ? node54108 : node54061;
											assign node54061 = (inp[3]) ? node54085 : node54062;
												assign node54062 = (inp[5]) ? node54072 : node54063;
													assign node54063 = (inp[8]) ? 4'b1000 : node54064;
														assign node54064 = (inp[7]) ? node54068 : node54065;
															assign node54065 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node54068 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node54072 = (inp[2]) ? node54080 : node54073;
														assign node54073 = (inp[8]) ? node54077 : node54074;
															assign node54074 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node54077 = (inp[14]) ? 4'b1010 : 4'b1010;
														assign node54080 = (inp[14]) ? node54082 : 4'b1011;
															assign node54082 = (inp[7]) ? 4'b1010 : 4'b1010;
												assign node54085 = (inp[2]) ? node54101 : node54086;
													assign node54086 = (inp[8]) ? node54094 : node54087;
														assign node54087 = (inp[5]) ? node54091 : node54088;
															assign node54088 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node54091 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node54094 = (inp[5]) ? node54098 : node54095;
															assign node54095 = (inp[7]) ? 4'b1010 : 4'b1010;
															assign node54098 = (inp[7]) ? 4'b1010 : 4'b1010;
													assign node54101 = (inp[7]) ? node54105 : node54102;
														assign node54102 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node54105 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node54108 = (inp[3]) ? node54136 : node54109;
												assign node54109 = (inp[5]) ? node54125 : node54110;
													assign node54110 = (inp[7]) ? node54118 : node54111;
														assign node54111 = (inp[8]) ? node54115 : node54112;
															assign node54112 = (inp[2]) ? 4'b1010 : 4'b1010;
															assign node54115 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node54118 = (inp[8]) ? node54122 : node54119;
															assign node54119 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node54122 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node54125 = (inp[8]) ? node54131 : node54126;
														assign node54126 = (inp[7]) ? node54128 : 4'b1000;
															assign node54128 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node54131 = (inp[14]) ? 4'b1001 : node54132;
															assign node54132 = (inp[2]) ? 4'b1000 : 4'b1000;
												assign node54136 = (inp[14]) ? node54152 : node54137;
													assign node54137 = (inp[5]) ? node54145 : node54138;
														assign node54138 = (inp[2]) ? node54142 : node54139;
															assign node54139 = (inp[7]) ? 4'b1000 : 4'b1000;
															assign node54142 = (inp[8]) ? 4'b1000 : 4'b1000;
														assign node54145 = (inp[7]) ? node54149 : node54146;
															assign node54146 = (inp[2]) ? 4'b1000 : 4'b1000;
															assign node54149 = (inp[8]) ? 4'b1000 : 4'b1000;
													assign node54152 = (inp[7]) ? node54156 : node54153;
														assign node54153 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node54156 = (inp[8]) ? 4'b1000 : 4'b1001;
									assign node54159 = (inp[7]) ? node54265 : node54160;
										assign node54160 = (inp[8]) ? node54210 : node54161;
											assign node54161 = (inp[14]) ? node54189 : node54162;
												assign node54162 = (inp[2]) ? node54176 : node54163;
													assign node54163 = (inp[15]) ? node54169 : node54164;
														assign node54164 = (inp[0]) ? node54166 : 4'b0001;
															assign node54166 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node54169 = (inp[0]) ? node54173 : node54170;
															assign node54170 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node54173 = (inp[3]) ? 4'b0001 : 4'b0001;
													assign node54176 = (inp[15]) ? node54184 : node54177;
														assign node54177 = (inp[0]) ? node54181 : node54178;
															assign node54178 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node54181 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node54184 = (inp[0]) ? node54186 : 4'b0010;
															assign node54186 = (inp[5]) ? 4'b0000 : 4'b0000;
												assign node54189 = (inp[3]) ? node54203 : node54190;
													assign node54190 = (inp[0]) ? node54196 : node54191;
														assign node54191 = (inp[2]) ? 4'b0010 : node54192;
															assign node54192 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node54196 = (inp[15]) ? node54200 : node54197;
															assign node54197 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node54200 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node54203 = (inp[15]) ? node54207 : node54204;
														assign node54204 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node54207 = (inp[0]) ? 4'b0000 : 4'b0010;
											assign node54210 = (inp[2]) ? node54242 : node54211;
												assign node54211 = (inp[14]) ? node54227 : node54212;
													assign node54212 = (inp[5]) ? node54220 : node54213;
														assign node54213 = (inp[15]) ? node54217 : node54214;
															assign node54214 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node54217 = (inp[3]) ? 4'b0000 : 4'b0000;
														assign node54220 = (inp[3]) ? node54224 : node54221;
															assign node54221 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node54224 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node54227 = (inp[0]) ? node54235 : node54228;
														assign node54228 = (inp[15]) ? node54232 : node54229;
															assign node54229 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node54232 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node54235 = (inp[15]) ? node54239 : node54236;
															assign node54236 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node54239 = (inp[3]) ? 4'b0001 : 4'b0001;
												assign node54242 = (inp[15]) ? node54254 : node54243;
													assign node54243 = (inp[0]) ? node54249 : node54244;
														assign node54244 = (inp[5]) ? 4'b0001 : node54245;
															assign node54245 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node54249 = (inp[5]) ? 4'b0011 : node54250;
															assign node54250 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node54254 = (inp[0]) ? node54260 : node54255;
														assign node54255 = (inp[3]) ? 4'b0011 : node54256;
															assign node54256 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node54260 = (inp[5]) ? 4'b0001 : node54261;
															assign node54261 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node54265 = (inp[8]) ? node54327 : node54266;
											assign node54266 = (inp[14]) ? node54296 : node54267;
												assign node54267 = (inp[2]) ? node54283 : node54268;
													assign node54268 = (inp[3]) ? node54276 : node54269;
														assign node54269 = (inp[5]) ? node54273 : node54270;
															assign node54270 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node54273 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node54276 = (inp[5]) ? node54280 : node54277;
															assign node54277 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node54280 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node54283 = (inp[0]) ? node54289 : node54284;
														assign node54284 = (inp[15]) ? node54286 : 4'b0001;
															assign node54286 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node54289 = (inp[15]) ? node54293 : node54290;
															assign node54290 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node54293 = (inp[5]) ? 4'b0001 : 4'b0001;
												assign node54296 = (inp[2]) ? node54312 : node54297;
													assign node54297 = (inp[3]) ? node54305 : node54298;
														assign node54298 = (inp[5]) ? node54302 : node54299;
															assign node54299 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node54302 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node54305 = (inp[15]) ? node54309 : node54306;
															assign node54306 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node54309 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node54312 = (inp[5]) ? node54320 : node54313;
														assign node54313 = (inp[3]) ? node54317 : node54314;
															assign node54314 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node54317 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node54320 = (inp[3]) ? node54324 : node54321;
															assign node54321 = (inp[15]) ? 4'b0001 : 4'b0001;
															assign node54324 = (inp[0]) ? 4'b0001 : 4'b0001;
											assign node54327 = (inp[14]) ? node54355 : node54328;
												assign node54328 = (inp[2]) ? node54344 : node54329;
													assign node54329 = (inp[0]) ? node54337 : node54330;
														assign node54330 = (inp[15]) ? node54334 : node54331;
															assign node54331 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node54334 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node54337 = (inp[15]) ? node54341 : node54338;
															assign node54338 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node54341 = (inp[3]) ? 4'b0001 : 4'b0001;
													assign node54344 = (inp[0]) ? node54350 : node54345;
														assign node54345 = (inp[3]) ? 4'b0000 : node54346;
															assign node54346 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node54350 = (inp[15]) ? node54352 : 4'b0010;
															assign node54352 = (inp[5]) ? 4'b0000 : 4'b0000;
												assign node54355 = (inp[5]) ? node54371 : node54356;
													assign node54356 = (inp[15]) ? node54364 : node54357;
														assign node54357 = (inp[2]) ? node54361 : node54358;
															assign node54358 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node54361 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node54364 = (inp[3]) ? node54368 : node54365;
															assign node54365 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node54368 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node54371 = (inp[2]) ? node54379 : node54372;
														assign node54372 = (inp[0]) ? node54376 : node54373;
															assign node54373 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node54376 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node54379 = (inp[3]) ? node54383 : node54380;
															assign node54380 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node54383 = (inp[15]) ? 4'b0000 : 4'b0000;
								assign node54386 = (inp[11]) ? node54624 : node54387;
									assign node54387 = (inp[8]) ? node54511 : node54388;
										assign node54388 = (inp[7]) ? node54452 : node54389;
											assign node54389 = (inp[14]) ? node54421 : node54390;
												assign node54390 = (inp[2]) ? node54406 : node54391;
													assign node54391 = (inp[0]) ? node54399 : node54392;
														assign node54392 = (inp[15]) ? node54396 : node54393;
															assign node54393 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node54396 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node54399 = (inp[15]) ? node54403 : node54400;
															assign node54400 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node54403 = (inp[5]) ? 4'b0001 : 4'b0001;
													assign node54406 = (inp[3]) ? node54414 : node54407;
														assign node54407 = (inp[5]) ? node54411 : node54408;
															assign node54408 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node54411 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node54414 = (inp[15]) ? node54418 : node54415;
															assign node54415 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node54418 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node54421 = (inp[5]) ? node54437 : node54422;
													assign node54422 = (inp[0]) ? node54430 : node54423;
														assign node54423 = (inp[2]) ? node54427 : node54424;
															assign node54424 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node54427 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node54430 = (inp[15]) ? node54434 : node54431;
															assign node54431 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node54434 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node54437 = (inp[2]) ? node54445 : node54438;
														assign node54438 = (inp[15]) ? node54442 : node54439;
															assign node54439 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node54442 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node54445 = (inp[3]) ? node54449 : node54446;
															assign node54446 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node54449 = (inp[0]) ? 4'b0000 : 4'b0010;
											assign node54452 = (inp[14]) ? node54480 : node54453;
												assign node54453 = (inp[2]) ? node54469 : node54454;
													assign node54454 = (inp[5]) ? node54462 : node54455;
														assign node54455 = (inp[0]) ? node54459 : node54456;
															assign node54456 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node54459 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node54462 = (inp[3]) ? node54466 : node54463;
															assign node54463 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node54466 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node54469 = (inp[0]) ? node54477 : node54470;
														assign node54470 = (inp[15]) ? node54474 : node54471;
															assign node54471 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node54474 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node54477 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node54480 = (inp[3]) ? node54496 : node54481;
													assign node54481 = (inp[2]) ? node54489 : node54482;
														assign node54482 = (inp[15]) ? node54486 : node54483;
															assign node54483 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node54486 = (inp[0]) ? 4'b0001 : 4'b0001;
														assign node54489 = (inp[5]) ? node54493 : node54490;
															assign node54490 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node54493 = (inp[0]) ? 4'b0001 : 4'b0001;
													assign node54496 = (inp[5]) ? node54504 : node54497;
														assign node54497 = (inp[0]) ? node54501 : node54498;
															assign node54498 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node54501 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node54504 = (inp[2]) ? node54508 : node54505;
															assign node54505 = (inp[0]) ? 4'b0001 : 4'b0001;
															assign node54508 = (inp[15]) ? 4'b0001 : 4'b0001;
										assign node54511 = (inp[7]) ? node54567 : node54512;
											assign node54512 = (inp[2]) ? node54544 : node54513;
												assign node54513 = (inp[14]) ? node54529 : node54514;
													assign node54514 = (inp[15]) ? node54522 : node54515;
														assign node54515 = (inp[0]) ? node54519 : node54516;
															assign node54516 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node54519 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node54522 = (inp[0]) ? node54526 : node54523;
															assign node54523 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node54526 = (inp[5]) ? 4'b0000 : 4'b0000;
													assign node54529 = (inp[15]) ? node54537 : node54530;
														assign node54530 = (inp[0]) ? node54534 : node54531;
															assign node54531 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node54534 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node54537 = (inp[0]) ? node54541 : node54538;
															assign node54538 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node54541 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node54544 = (inp[5]) ? node54560 : node54545;
													assign node54545 = (inp[15]) ? node54553 : node54546;
														assign node54546 = (inp[0]) ? node54550 : node54547;
															assign node54547 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node54550 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node54553 = (inp[14]) ? node54557 : node54554;
															assign node54554 = (inp[3]) ? 4'b0001 : 4'b0001;
															assign node54557 = (inp[3]) ? 4'b0001 : 4'b0001;
													assign node54560 = (inp[0]) ? node54564 : node54561;
														assign node54561 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node54564 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node54567 = (inp[14]) ? node54595 : node54568;
												assign node54568 = (inp[2]) ? node54582 : node54569;
													assign node54569 = (inp[3]) ? node54575 : node54570;
														assign node54570 = (inp[0]) ? 4'b0011 : node54571;
															assign node54571 = (inp[15]) ? 4'b0001 : 4'b0001;
														assign node54575 = (inp[0]) ? node54579 : node54576;
															assign node54576 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node54579 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node54582 = (inp[3]) ? node54588 : node54583;
														assign node54583 = (inp[15]) ? node54585 : 4'b0010;
															assign node54585 = (inp[0]) ? 4'b0000 : 4'b0000;
														assign node54588 = (inp[5]) ? node54592 : node54589;
															assign node54589 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node54592 = (inp[0]) ? 4'b0000 : 4'b0000;
												assign node54595 = (inp[2]) ? node54611 : node54596;
													assign node54596 = (inp[0]) ? node54604 : node54597;
														assign node54597 = (inp[15]) ? node54601 : node54598;
															assign node54598 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node54601 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node54604 = (inp[15]) ? node54608 : node54605;
															assign node54605 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node54608 = (inp[3]) ? 4'b0000 : 4'b0000;
													assign node54611 = (inp[3]) ? node54617 : node54612;
														assign node54612 = (inp[5]) ? node54614 : 4'b0000;
															assign node54614 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node54617 = (inp[0]) ? node54621 : node54618;
															assign node54618 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node54621 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node54624 = (inp[15]) ? node54718 : node54625;
										assign node54625 = (inp[0]) ? node54671 : node54626;
											assign node54626 = (inp[3]) ? node54652 : node54627;
												assign node54627 = (inp[5]) ? node54641 : node54628;
													assign node54628 = (inp[2]) ? node54634 : node54629;
														assign node54629 = (inp[14]) ? 4'b1011 : node54630;
															assign node54630 = (inp[7]) ? 4'b1010 : 4'b1010;
														assign node54634 = (inp[8]) ? node54638 : node54635;
															assign node54635 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node54638 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node54641 = (inp[7]) ? node54647 : node54642;
														assign node54642 = (inp[8]) ? node54644 : 4'b1000;
															assign node54644 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node54647 = (inp[8]) ? node54649 : 4'b1001;
															assign node54649 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node54652 = (inp[7]) ? node54660 : node54653;
													assign node54653 = (inp[8]) ? 4'b1001 : node54654;
														assign node54654 = (inp[2]) ? 4'b1000 : node54655;
															assign node54655 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node54660 = (inp[8]) ? node54666 : node54661;
														assign node54661 = (inp[14]) ? 4'b1001 : node54662;
															assign node54662 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node54666 = (inp[14]) ? 4'b1000 : node54667;
															assign node54667 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node54671 = (inp[5]) ? node54695 : node54672;
												assign node54672 = (inp[3]) ? node54684 : node54673;
													assign node54673 = (inp[8]) ? node54679 : node54674;
														assign node54674 = (inp[7]) ? 4'b1001 : node54675;
															assign node54675 = (inp[2]) ? 4'b1000 : 4'b1000;
														assign node54679 = (inp[7]) ? 4'b1000 : node54680;
															assign node54680 = (inp[14]) ? 4'b1001 : 4'b1000;
													assign node54684 = (inp[7]) ? node54690 : node54685;
														assign node54685 = (inp[8]) ? 4'b1011 : node54686;
															assign node54686 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node54690 = (inp[8]) ? 4'b1010 : node54691;
															assign node54691 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node54695 = (inp[7]) ? node54707 : node54696;
													assign node54696 = (inp[8]) ? node54702 : node54697;
														assign node54697 = (inp[14]) ? 4'b1010 : node54698;
															assign node54698 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node54702 = (inp[2]) ? 4'b1011 : node54703;
															assign node54703 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node54707 = (inp[8]) ? node54713 : node54708;
														assign node54708 = (inp[14]) ? 4'b1011 : node54709;
															assign node54709 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node54713 = (inp[2]) ? 4'b1010 : node54714;
															assign node54714 = (inp[14]) ? 4'b1010 : 4'b1011;
										assign node54718 = (inp[0]) ? node54770 : node54719;
											assign node54719 = (inp[5]) ? node54747 : node54720;
												assign node54720 = (inp[3]) ? node54734 : node54721;
													assign node54721 = (inp[2]) ? node54729 : node54722;
														assign node54722 = (inp[7]) ? node54726 : node54723;
															assign node54723 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node54726 = (inp[14]) ? 4'b1000 : 4'b1000;
														assign node54729 = (inp[7]) ? 4'b1001 : node54730;
															assign node54730 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node54734 = (inp[7]) ? node54740 : node54735;
														assign node54735 = (inp[8]) ? node54737 : 4'b1010;
															assign node54737 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node54740 = (inp[8]) ? node54744 : node54741;
															assign node54741 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node54744 = (inp[14]) ? 4'b1010 : 4'b1010;
												assign node54747 = (inp[8]) ? node54759 : node54748;
													assign node54748 = (inp[7]) ? node54754 : node54749;
														assign node54749 = (inp[14]) ? 4'b1010 : node54750;
															assign node54750 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node54754 = (inp[14]) ? 4'b1011 : node54755;
															assign node54755 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node54759 = (inp[7]) ? node54765 : node54760;
														assign node54760 = (inp[14]) ? 4'b1011 : node54761;
															assign node54761 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node54765 = (inp[14]) ? 4'b1010 : node54766;
															assign node54766 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node54770 = (inp[5]) ? node54800 : node54771;
												assign node54771 = (inp[3]) ? node54787 : node54772;
													assign node54772 = (inp[8]) ? node54780 : node54773;
														assign node54773 = (inp[7]) ? node54777 : node54774;
															assign node54774 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node54777 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node54780 = (inp[7]) ? node54784 : node54781;
															assign node54781 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node54784 = (inp[14]) ? 4'b1010 : 4'b1010;
													assign node54787 = (inp[7]) ? node54795 : node54788;
														assign node54788 = (inp[8]) ? node54792 : node54789;
															assign node54789 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node54792 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node54795 = (inp[8]) ? node54797 : 4'b1001;
															assign node54797 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node54800 = (inp[14]) ? node54816 : node54801;
													assign node54801 = (inp[2]) ? node54809 : node54802;
														assign node54802 = (inp[8]) ? node54806 : node54803;
															assign node54803 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node54806 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node54809 = (inp[7]) ? node54813 : node54810;
															assign node54810 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node54813 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node54816 = (inp[2]) ? node54824 : node54817;
														assign node54817 = (inp[3]) ? node54821 : node54818;
															assign node54818 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node54821 = (inp[7]) ? 4'b1000 : 4'b1000;
														assign node54824 = (inp[3]) ? 4'b1001 : node54825;
															assign node54825 = (inp[8]) ? 4'b1000 : 4'b1001;
							assign node54829 = (inp[15]) ? node55273 : node54830;
								assign node54830 = (inp[0]) ? node55048 : node54831;
									assign node54831 = (inp[3]) ? node54953 : node54832;
										assign node54832 = (inp[5]) ? node54896 : node54833;
											assign node54833 = (inp[14]) ? node54865 : node54834;
												assign node54834 = (inp[7]) ? node54850 : node54835;
													assign node54835 = (inp[6]) ? node54843 : node54836;
														assign node54836 = (inp[11]) ? node54840 : node54837;
															assign node54837 = (inp[2]) ? 4'b0011 : 4'b1010;
															assign node54840 = (inp[8]) ? 4'b0010 : 4'b0010;
														assign node54843 = (inp[11]) ? node54847 : node54844;
															assign node54844 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node54847 = (inp[8]) ? 4'b0011 : 4'b1010;
													assign node54850 = (inp[11]) ? node54858 : node54851;
														assign node54851 = (inp[6]) ? node54855 : node54852;
															assign node54852 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node54855 = (inp[8]) ? 4'b1010 : 4'b0010;
														assign node54858 = (inp[6]) ? node54862 : node54859;
															assign node54859 = (inp[8]) ? 4'b1010 : 4'b0010;
															assign node54862 = (inp[2]) ? 4'b0010 : 4'b0010;
												assign node54865 = (inp[6]) ? node54881 : node54866;
													assign node54866 = (inp[11]) ? node54874 : node54867;
														assign node54867 = (inp[7]) ? node54871 : node54868;
															assign node54868 = (inp[8]) ? 4'b0011 : 4'b1010;
															assign node54871 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node54874 = (inp[8]) ? node54878 : node54875;
															assign node54875 = (inp[7]) ? 4'b1011 : 4'b0010;
															assign node54878 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node54881 = (inp[11]) ? node54889 : node54882;
														assign node54882 = (inp[7]) ? node54886 : node54883;
															assign node54883 = (inp[8]) ? 4'b1011 : 4'b0010;
															assign node54886 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node54889 = (inp[8]) ? node54893 : node54890;
															assign node54890 = (inp[7]) ? 4'b0011 : 4'b1010;
															assign node54893 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node54896 = (inp[11]) ? node54924 : node54897;
												assign node54897 = (inp[6]) ? node54911 : node54898;
													assign node54898 = (inp[7]) ? node54906 : node54899;
														assign node54899 = (inp[8]) ? node54903 : node54900;
															assign node54900 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node54903 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node54906 = (inp[8]) ? node54908 : 4'b0001;
															assign node54908 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node54911 = (inp[7]) ? node54919 : node54912;
														assign node54912 = (inp[8]) ? node54916 : node54913;
															assign node54913 = (inp[14]) ? 4'b0000 : 4'b0001;
															assign node54916 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node54919 = (inp[8]) ? node54921 : 4'b1001;
															assign node54921 = (inp[14]) ? 4'b1000 : 4'b1000;
												assign node54924 = (inp[6]) ? node54940 : node54925;
													assign node54925 = (inp[7]) ? node54933 : node54926;
														assign node54926 = (inp[8]) ? node54930 : node54927;
															assign node54927 = (inp[14]) ? 4'b0000 : 4'b0000;
															assign node54930 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node54933 = (inp[8]) ? node54937 : node54934;
															assign node54934 = (inp[2]) ? 4'b1001 : 4'b0000;
															assign node54937 = (inp[14]) ? 4'b1000 : 4'b1000;
													assign node54940 = (inp[8]) ? node54948 : node54941;
														assign node54941 = (inp[7]) ? node54945 : node54942;
															assign node54942 = (inp[2]) ? 4'b1000 : 4'b1000;
															assign node54945 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node54948 = (inp[7]) ? node54950 : 4'b0001;
															assign node54950 = (inp[2]) ? 4'b0000 : 4'b0000;
										assign node54953 = (inp[6]) ? node55001 : node54954;
											assign node54954 = (inp[11]) ? node54978 : node54955;
												assign node54955 = (inp[7]) ? node54967 : node54956;
													assign node54956 = (inp[8]) ? node54962 : node54957;
														assign node54957 = (inp[2]) ? 4'b1000 : node54958;
															assign node54958 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node54962 = (inp[2]) ? 4'b0001 : node54963;
															assign node54963 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node54967 = (inp[8]) ? node54973 : node54968;
														assign node54968 = (inp[2]) ? 4'b0001 : node54969;
															assign node54969 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node54973 = (inp[14]) ? 4'b0000 : node54974;
															assign node54974 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node54978 = (inp[8]) ? node54990 : node54979;
													assign node54979 = (inp[7]) ? node54985 : node54980;
														assign node54980 = (inp[2]) ? 4'b0000 : node54981;
															assign node54981 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node54985 = (inp[2]) ? 4'b1001 : node54986;
															assign node54986 = (inp[14]) ? 4'b1001 : 4'b0000;
													assign node54990 = (inp[7]) ? node54996 : node54991;
														assign node54991 = (inp[14]) ? 4'b1001 : node54992;
															assign node54992 = (inp[2]) ? 4'b1001 : 4'b0000;
														assign node54996 = (inp[14]) ? 4'b1000 : node54997;
															assign node54997 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node55001 = (inp[11]) ? node55025 : node55002;
												assign node55002 = (inp[8]) ? node55014 : node55003;
													assign node55003 = (inp[7]) ? node55009 : node55004;
														assign node55004 = (inp[2]) ? 4'b0000 : node55005;
															assign node55005 = (inp[14]) ? 4'b0000 : 4'b0001;
														assign node55009 = (inp[14]) ? 4'b1001 : node55010;
															assign node55010 = (inp[2]) ? 4'b1001 : 4'b0000;
													assign node55014 = (inp[7]) ? node55020 : node55015;
														assign node55015 = (inp[2]) ? 4'b1001 : node55016;
															assign node55016 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node55020 = (inp[14]) ? 4'b1000 : node55021;
															assign node55021 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node55025 = (inp[8]) ? node55037 : node55026;
													assign node55026 = (inp[7]) ? node55032 : node55027;
														assign node55027 = (inp[14]) ? 4'b1000 : node55028;
															assign node55028 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node55032 = (inp[2]) ? 4'b0001 : node55033;
															assign node55033 = (inp[14]) ? 4'b0001 : 4'b1000;
													assign node55037 = (inp[7]) ? node55043 : node55038;
														assign node55038 = (inp[2]) ? 4'b0001 : node55039;
															assign node55039 = (inp[14]) ? 4'b0001 : 4'b1000;
														assign node55043 = (inp[14]) ? 4'b0000 : node55044;
															assign node55044 = (inp[2]) ? 4'b0000 : 4'b0001;
									assign node55048 = (inp[5]) ? node55164 : node55049;
										assign node55049 = (inp[3]) ? node55113 : node55050;
											assign node55050 = (inp[14]) ? node55082 : node55051;
												assign node55051 = (inp[6]) ? node55067 : node55052;
													assign node55052 = (inp[7]) ? node55060 : node55053;
														assign node55053 = (inp[11]) ? node55057 : node55054;
															assign node55054 = (inp[8]) ? 4'b1000 : 4'b1000;
															assign node55057 = (inp[8]) ? 4'b1001 : 4'b0000;
														assign node55060 = (inp[11]) ? node55064 : node55061;
															assign node55061 = (inp[8]) ? 4'b0000 : 4'b1000;
															assign node55064 = (inp[8]) ? 4'b1000 : 4'b0000;
													assign node55067 = (inp[8]) ? node55075 : node55068;
														assign node55068 = (inp[11]) ? node55072 : node55069;
															assign node55069 = (inp[2]) ? 4'b1001 : 4'b0000;
															assign node55072 = (inp[7]) ? 4'b0000 : 4'b1000;
														assign node55075 = (inp[11]) ? node55079 : node55076;
															assign node55076 = (inp[2]) ? 4'b1000 : 4'b0000;
															assign node55079 = (inp[7]) ? 4'b0000 : 4'b0000;
												assign node55082 = (inp[8]) ? node55098 : node55083;
													assign node55083 = (inp[7]) ? node55091 : node55084;
														assign node55084 = (inp[11]) ? node55088 : node55085;
															assign node55085 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node55088 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node55091 = (inp[6]) ? node55095 : node55092;
															assign node55092 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node55095 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node55098 = (inp[7]) ? node55106 : node55099;
														assign node55099 = (inp[6]) ? node55103 : node55100;
															assign node55100 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node55103 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node55106 = (inp[11]) ? node55110 : node55107;
															assign node55107 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node55110 = (inp[6]) ? 4'b0000 : 4'b1000;
											assign node55113 = (inp[6]) ? node55141 : node55114;
												assign node55114 = (inp[11]) ? node55128 : node55115;
													assign node55115 = (inp[7]) ? node55123 : node55116;
														assign node55116 = (inp[8]) ? node55120 : node55117;
															assign node55117 = (inp[2]) ? 4'b1010 : 4'b1010;
															assign node55120 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node55123 = (inp[2]) ? node55125 : 4'b0011;
															assign node55125 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node55128 = (inp[8]) ? node55134 : node55129;
														assign node55129 = (inp[7]) ? node55131 : 4'b0010;
															assign node55131 = (inp[2]) ? 4'b1011 : 4'b0010;
														assign node55134 = (inp[7]) ? node55138 : node55135;
															assign node55135 = (inp[2]) ? 4'b1011 : 4'b0010;
															assign node55138 = (inp[14]) ? 4'b1010 : 4'b1010;
												assign node55141 = (inp[11]) ? node55153 : node55142;
													assign node55142 = (inp[8]) ? node55148 : node55143;
														assign node55143 = (inp[7]) ? 4'b1011 : node55144;
															assign node55144 = (inp[2]) ? 4'b0010 : 4'b0010;
														assign node55148 = (inp[7]) ? node55150 : 4'b1011;
															assign node55150 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node55153 = (inp[7]) ? node55159 : node55154;
														assign node55154 = (inp[8]) ? 4'b0011 : node55155;
															assign node55155 = (inp[2]) ? 4'b1010 : 4'b1010;
														assign node55159 = (inp[8]) ? node55161 : 4'b0011;
															assign node55161 = (inp[2]) ? 4'b0010 : 4'b0010;
										assign node55164 = (inp[8]) ? node55210 : node55165;
											assign node55165 = (inp[7]) ? node55187 : node55166;
												assign node55166 = (inp[14]) ? node55180 : node55167;
													assign node55167 = (inp[2]) ? node55173 : node55168;
														assign node55168 = (inp[11]) ? node55170 : 4'b1011;
															assign node55170 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node55173 = (inp[3]) ? node55177 : node55174;
															assign node55174 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node55177 = (inp[6]) ? 4'b0010 : 4'b0010;
													assign node55180 = (inp[11]) ? node55184 : node55181;
														assign node55181 = (inp[6]) ? 4'b0010 : 4'b1010;
														assign node55184 = (inp[6]) ? 4'b1010 : 4'b0010;
												assign node55187 = (inp[14]) ? node55203 : node55188;
													assign node55188 = (inp[2]) ? node55196 : node55189;
														assign node55189 = (inp[3]) ? node55193 : node55190;
															assign node55190 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node55193 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node55196 = (inp[6]) ? node55200 : node55197;
															assign node55197 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node55200 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node55203 = (inp[6]) ? node55207 : node55204;
														assign node55204 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node55207 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node55210 = (inp[7]) ? node55242 : node55211;
												assign node55211 = (inp[2]) ? node55227 : node55212;
													assign node55212 = (inp[14]) ? node55220 : node55213;
														assign node55213 = (inp[6]) ? node55217 : node55214;
															assign node55214 = (inp[11]) ? 4'b0010 : 4'b1010;
															assign node55217 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node55220 = (inp[11]) ? node55224 : node55221;
															assign node55221 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node55224 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node55227 = (inp[3]) ? node55235 : node55228;
														assign node55228 = (inp[6]) ? node55232 : node55229;
															assign node55229 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node55232 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node55235 = (inp[6]) ? node55239 : node55236;
															assign node55236 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node55239 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node55242 = (inp[14]) ? node55258 : node55243;
													assign node55243 = (inp[2]) ? node55251 : node55244;
														assign node55244 = (inp[3]) ? node55248 : node55245;
															assign node55245 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node55248 = (inp[11]) ? 4'b0011 : 4'b0011;
														assign node55251 = (inp[3]) ? node55255 : node55252;
															assign node55252 = (inp[11]) ? 4'b0010 : 4'b1010;
															assign node55255 = (inp[11]) ? 4'b0010 : 4'b0010;
													assign node55258 = (inp[3]) ? node55266 : node55259;
														assign node55259 = (inp[6]) ? node55263 : node55260;
															assign node55260 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node55263 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node55266 = (inp[2]) ? node55270 : node55267;
															assign node55267 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node55270 = (inp[6]) ? 4'b0010 : 4'b0010;
								assign node55273 = (inp[0]) ? node55523 : node55274;
									assign node55274 = (inp[5]) ? node55398 : node55275;
										assign node55275 = (inp[3]) ? node55337 : node55276;
											assign node55276 = (inp[6]) ? node55308 : node55277;
												assign node55277 = (inp[11]) ? node55293 : node55278;
													assign node55278 = (inp[7]) ? node55286 : node55279;
														assign node55279 = (inp[8]) ? node55283 : node55280;
															assign node55280 = (inp[2]) ? 4'b1000 : 4'b1000;
															assign node55283 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node55286 = (inp[8]) ? node55290 : node55287;
															assign node55287 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node55290 = (inp[2]) ? 4'b0000 : 4'b0000;
													assign node55293 = (inp[7]) ? node55301 : node55294;
														assign node55294 = (inp[8]) ? node55298 : node55295;
															assign node55295 = (inp[2]) ? 4'b0000 : 4'b0000;
															assign node55298 = (inp[2]) ? 4'b1001 : 4'b0000;
														assign node55301 = (inp[8]) ? node55305 : node55302;
															assign node55302 = (inp[2]) ? 4'b1001 : 4'b0000;
															assign node55305 = (inp[2]) ? 4'b1000 : 4'b1000;
												assign node55308 = (inp[11]) ? node55322 : node55309;
													assign node55309 = (inp[8]) ? node55315 : node55310;
														assign node55310 = (inp[7]) ? node55312 : 4'b0000;
															assign node55312 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node55315 = (inp[7]) ? node55319 : node55316;
															assign node55316 = (inp[2]) ? 4'b1001 : 4'b0000;
															assign node55319 = (inp[14]) ? 4'b1000 : 4'b1000;
													assign node55322 = (inp[8]) ? node55330 : node55323;
														assign node55323 = (inp[7]) ? node55327 : node55324;
															assign node55324 = (inp[2]) ? 4'b1000 : 4'b1000;
															assign node55327 = (inp[14]) ? 4'b0001 : 4'b0000;
														assign node55330 = (inp[7]) ? node55334 : node55331;
															assign node55331 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node55334 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node55337 = (inp[7]) ? node55367 : node55338;
												assign node55338 = (inp[8]) ? node55354 : node55339;
													assign node55339 = (inp[2]) ? node55347 : node55340;
														assign node55340 = (inp[14]) ? node55344 : node55341;
															assign node55341 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node55344 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node55347 = (inp[11]) ? node55351 : node55348;
															assign node55348 = (inp[6]) ? 4'b0010 : 4'b1010;
															assign node55351 = (inp[6]) ? 4'b1010 : 4'b0010;
													assign node55354 = (inp[2]) ? node55362 : node55355;
														assign node55355 = (inp[14]) ? node55359 : node55356;
															assign node55356 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node55359 = (inp[11]) ? 4'b0011 : 4'b0011;
														assign node55362 = (inp[6]) ? 4'b0011 : node55363;
															assign node55363 = (inp[11]) ? 4'b1011 : 4'b0011;
												assign node55367 = (inp[8]) ? node55383 : node55368;
													assign node55368 = (inp[2]) ? node55376 : node55369;
														assign node55369 = (inp[14]) ? node55373 : node55370;
															assign node55370 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node55373 = (inp[11]) ? 4'b0011 : 4'b0011;
														assign node55376 = (inp[11]) ? node55380 : node55377;
															assign node55377 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node55380 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node55383 = (inp[14]) ? node55391 : node55384;
														assign node55384 = (inp[2]) ? node55388 : node55385;
															assign node55385 = (inp[11]) ? 4'b0011 : 4'b1011;
															assign node55388 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node55391 = (inp[11]) ? node55395 : node55392;
															assign node55392 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node55395 = (inp[6]) ? 4'b0010 : 4'b1010;
										assign node55398 = (inp[14]) ? node55460 : node55399;
											assign node55399 = (inp[3]) ? node55429 : node55400;
												assign node55400 = (inp[2]) ? node55416 : node55401;
													assign node55401 = (inp[8]) ? node55409 : node55402;
														assign node55402 = (inp[7]) ? node55406 : node55403;
															assign node55403 = (inp[11]) ? 4'b0011 : 4'b0011;
															assign node55406 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node55409 = (inp[7]) ? node55413 : node55410;
															assign node55410 = (inp[6]) ? 4'b0010 : 4'b1010;
															assign node55413 = (inp[6]) ? 4'b0011 : 4'b0011;
													assign node55416 = (inp[6]) ? node55424 : node55417;
														assign node55417 = (inp[11]) ? node55421 : node55418;
															assign node55418 = (inp[8]) ? 4'b0010 : 4'b1010;
															assign node55421 = (inp[7]) ? 4'b1010 : 4'b0010;
														assign node55424 = (inp[11]) ? 4'b1010 : node55425;
															assign node55425 = (inp[7]) ? 4'b1010 : 4'b0010;
												assign node55429 = (inp[6]) ? node55445 : node55430;
													assign node55430 = (inp[8]) ? node55438 : node55431;
														assign node55431 = (inp[11]) ? node55435 : node55432;
															assign node55432 = (inp[7]) ? 4'b0010 : 4'b1010;
															assign node55435 = (inp[7]) ? 4'b0010 : 4'b0010;
														assign node55438 = (inp[11]) ? node55442 : node55439;
															assign node55439 = (inp[2]) ? 4'b0010 : 4'b1010;
															assign node55442 = (inp[2]) ? 4'b1010 : 4'b0010;
													assign node55445 = (inp[11]) ? node55453 : node55446;
														assign node55446 = (inp[7]) ? node55450 : node55447;
															assign node55447 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node55450 = (inp[8]) ? 4'b1010 : 4'b0010;
														assign node55453 = (inp[2]) ? node55457 : node55454;
															assign node55454 = (inp[7]) ? 4'b0010 : 4'b1010;
															assign node55457 = (inp[8]) ? 4'b0010 : 4'b0010;
											assign node55460 = (inp[3]) ? node55492 : node55461;
												assign node55461 = (inp[8]) ? node55477 : node55462;
													assign node55462 = (inp[7]) ? node55470 : node55463;
														assign node55463 = (inp[11]) ? node55467 : node55464;
															assign node55464 = (inp[6]) ? 4'b0010 : 4'b1010;
															assign node55467 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node55470 = (inp[2]) ? node55474 : node55471;
															assign node55471 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node55474 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node55477 = (inp[7]) ? node55485 : node55478;
														assign node55478 = (inp[6]) ? node55482 : node55479;
															assign node55479 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node55482 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node55485 = (inp[2]) ? node55489 : node55486;
															assign node55486 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node55489 = (inp[6]) ? 4'b0010 : 4'b0010;
												assign node55492 = (inp[2]) ? node55508 : node55493;
													assign node55493 = (inp[7]) ? node55501 : node55494;
														assign node55494 = (inp[8]) ? node55498 : node55495;
															assign node55495 = (inp[6]) ? 4'b0010 : 4'b1010;
															assign node55498 = (inp[6]) ? 4'b0011 : 4'b0011;
														assign node55501 = (inp[8]) ? node55505 : node55502;
															assign node55502 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node55505 = (inp[11]) ? 4'b0010 : 4'b0010;
													assign node55508 = (inp[11]) ? node55516 : node55509;
														assign node55509 = (inp[6]) ? node55513 : node55510;
															assign node55510 = (inp[8]) ? 4'b0010 : 4'b0010;
															assign node55513 = (inp[7]) ? 4'b1010 : 4'b0010;
														assign node55516 = (inp[6]) ? node55520 : node55517;
															assign node55517 = (inp[8]) ? 4'b1010 : 4'b0010;
															assign node55520 = (inp[8]) ? 4'b0010 : 4'b0010;
									assign node55523 = (inp[5]) ? node55647 : node55524;
										assign node55524 = (inp[3]) ? node55586 : node55525;
											assign node55525 = (inp[6]) ? node55557 : node55526;
												assign node55526 = (inp[11]) ? node55542 : node55527;
													assign node55527 = (inp[7]) ? node55535 : node55528;
														assign node55528 = (inp[8]) ? node55532 : node55529;
															assign node55529 = (inp[14]) ? 4'b1010 : 4'b1011;
															assign node55532 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node55535 = (inp[8]) ? node55539 : node55536;
															assign node55536 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node55539 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node55542 = (inp[8]) ? node55550 : node55543;
														assign node55543 = (inp[7]) ? node55547 : node55544;
															assign node55544 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node55547 = (inp[14]) ? 4'b1011 : 4'b0010;
														assign node55550 = (inp[7]) ? node55554 : node55551;
															assign node55551 = (inp[2]) ? 4'b1011 : 4'b0010;
															assign node55554 = (inp[2]) ? 4'b1010 : 4'b1010;
												assign node55557 = (inp[11]) ? node55573 : node55558;
													assign node55558 = (inp[7]) ? node55566 : node55559;
														assign node55559 = (inp[8]) ? node55563 : node55560;
															assign node55560 = (inp[2]) ? 4'b0010 : 4'b0010;
															assign node55563 = (inp[2]) ? 4'b1011 : 4'b0010;
														assign node55566 = (inp[8]) ? node55570 : node55567;
															assign node55567 = (inp[2]) ? 4'b1011 : 4'b0010;
															assign node55570 = (inp[2]) ? 4'b1010 : 4'b1010;
													assign node55573 = (inp[8]) ? node55579 : node55574;
														assign node55574 = (inp[2]) ? 4'b1010 : node55575;
															assign node55575 = (inp[14]) ? 4'b0011 : 4'b1010;
														assign node55579 = (inp[7]) ? node55583 : node55580;
															assign node55580 = (inp[2]) ? 4'b0011 : 4'b1010;
															assign node55583 = (inp[2]) ? 4'b0010 : 4'b0010;
											assign node55586 = (inp[11]) ? node55618 : node55587;
												assign node55587 = (inp[6]) ? node55603 : node55588;
													assign node55588 = (inp[8]) ? node55596 : node55589;
														assign node55589 = (inp[7]) ? node55593 : node55590;
															assign node55590 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node55593 = (inp[2]) ? 4'b0001 : 4'b1000;
														assign node55596 = (inp[7]) ? node55600 : node55597;
															assign node55597 = (inp[2]) ? 4'b0001 : 4'b1000;
															assign node55600 = (inp[2]) ? 4'b0000 : 4'b0000;
													assign node55603 = (inp[7]) ? node55611 : node55604;
														assign node55604 = (inp[8]) ? node55608 : node55605;
															assign node55605 = (inp[2]) ? 4'b0000 : 4'b0000;
															assign node55608 = (inp[14]) ? 4'b1001 : 4'b0000;
														assign node55611 = (inp[8]) ? node55615 : node55612;
															assign node55612 = (inp[2]) ? 4'b1001 : 4'b0000;
															assign node55615 = (inp[2]) ? 4'b1000 : 4'b1000;
												assign node55618 = (inp[8]) ? node55634 : node55619;
													assign node55619 = (inp[7]) ? node55627 : node55620;
														assign node55620 = (inp[6]) ? node55624 : node55621;
															assign node55621 = (inp[14]) ? 4'b0000 : 4'b0000;
															assign node55624 = (inp[2]) ? 4'b1000 : 4'b1000;
														assign node55627 = (inp[14]) ? node55631 : node55628;
															assign node55628 = (inp[2]) ? 4'b1001 : 4'b0000;
															assign node55631 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node55634 = (inp[6]) ? node55640 : node55635;
														assign node55635 = (inp[14]) ? 4'b1001 : node55636;
															assign node55636 = (inp[7]) ? 4'b1000 : 4'b0000;
														assign node55640 = (inp[7]) ? node55644 : node55641;
															assign node55641 = (inp[14]) ? 4'b0001 : 4'b0000;
															assign node55644 = (inp[14]) ? 4'b0000 : 4'b0001;
										assign node55647 = (inp[8]) ? node55709 : node55648;
											assign node55648 = (inp[7]) ? node55680 : node55649;
												assign node55649 = (inp[2]) ? node55665 : node55650;
													assign node55650 = (inp[14]) ? node55658 : node55651;
														assign node55651 = (inp[6]) ? node55655 : node55652;
															assign node55652 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node55655 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node55658 = (inp[3]) ? node55662 : node55659;
															assign node55659 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node55662 = (inp[11]) ? 4'b0000 : 4'b0000;
													assign node55665 = (inp[14]) ? node55673 : node55666;
														assign node55666 = (inp[3]) ? node55670 : node55667;
															assign node55667 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node55670 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node55673 = (inp[3]) ? node55677 : node55674;
															assign node55674 = (inp[11]) ? 4'b1000 : 4'b0000;
															assign node55677 = (inp[6]) ? 4'b0000 : 4'b0000;
												assign node55680 = (inp[2]) ? node55694 : node55681;
													assign node55681 = (inp[14]) ? node55689 : node55682;
														assign node55682 = (inp[11]) ? node55686 : node55683;
															assign node55683 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node55686 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node55689 = (inp[11]) ? 4'b1001 : node55690;
															assign node55690 = (inp[6]) ? 4'b1001 : 4'b0001;
													assign node55694 = (inp[14]) ? node55702 : node55695;
														assign node55695 = (inp[11]) ? node55699 : node55696;
															assign node55696 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node55699 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node55702 = (inp[3]) ? node55706 : node55703;
															assign node55703 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node55706 = (inp[11]) ? 4'b0001 : 4'b0001;
											assign node55709 = (inp[7]) ? node55733 : node55710;
												assign node55710 = (inp[2]) ? node55726 : node55711;
													assign node55711 = (inp[14]) ? node55719 : node55712;
														assign node55712 = (inp[11]) ? node55716 : node55713;
															assign node55713 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node55716 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node55719 = (inp[6]) ? node55723 : node55720;
															assign node55720 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node55723 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node55726 = (inp[6]) ? node55730 : node55727;
														assign node55727 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node55730 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node55733 = (inp[14]) ? node55749 : node55734;
													assign node55734 = (inp[2]) ? node55742 : node55735;
														assign node55735 = (inp[11]) ? node55739 : node55736;
															assign node55736 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node55739 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node55742 = (inp[3]) ? node55746 : node55743;
															assign node55743 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node55746 = (inp[6]) ? 4'b0000 : 4'b0000;
													assign node55749 = (inp[11]) ? node55753 : node55750;
														assign node55750 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node55753 = (inp[6]) ? 4'b0000 : 4'b1000;
						assign node55756 = (inp[8]) ? node56554 : node55757;
							assign node55757 = (inp[7]) ? node56231 : node55758;
								assign node55758 = (inp[14]) ? node56004 : node55759;
									assign node55759 = (inp[2]) ? node55885 : node55760;
										assign node55760 = (inp[15]) ? node55822 : node55761;
											assign node55761 = (inp[0]) ? node55791 : node55762;
												assign node55762 = (inp[5]) ? node55778 : node55763;
													assign node55763 = (inp[3]) ? node55771 : node55764;
														assign node55764 = (inp[6]) ? node55768 : node55765;
															assign node55765 = (inp[1]) ? 4'b1011 : 4'b0011;
															assign node55768 = (inp[1]) ? 4'b0011 : 4'b0011;
														assign node55771 = (inp[11]) ? node55775 : node55772;
															assign node55772 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node55775 = (inp[6]) ? 4'b0001 : 4'b0001;
													assign node55778 = (inp[6]) ? node55786 : node55779;
														assign node55779 = (inp[11]) ? node55783 : node55780;
															assign node55780 = (inp[1]) ? 4'b0001 : 4'b1001;
															assign node55783 = (inp[1]) ? 4'b1001 : 4'b0001;
														assign node55786 = (inp[3]) ? 4'b1001 : node55787;
															assign node55787 = (inp[11]) ? 4'b0001 : 4'b0001;
												assign node55791 = (inp[5]) ? node55807 : node55792;
													assign node55792 = (inp[3]) ? node55800 : node55793;
														assign node55793 = (inp[11]) ? node55797 : node55794;
															assign node55794 = (inp[1]) ? 4'b0001 : 4'b0001;
															assign node55797 = (inp[1]) ? 4'b0001 : 4'b0001;
														assign node55800 = (inp[1]) ? node55804 : node55801;
															assign node55801 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node55804 = (inp[6]) ? 4'b0011 : 4'b0011;
													assign node55807 = (inp[3]) ? node55815 : node55808;
														assign node55808 = (inp[6]) ? node55812 : node55809;
															assign node55809 = (inp[11]) ? 4'b0011 : 4'b0011;
															assign node55812 = (inp[1]) ? 4'b0011 : 4'b0011;
														assign node55815 = (inp[1]) ? node55819 : node55816;
															assign node55816 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node55819 = (inp[6]) ? 4'b0011 : 4'b0011;
											assign node55822 = (inp[0]) ? node55854 : node55823;
												assign node55823 = (inp[5]) ? node55839 : node55824;
													assign node55824 = (inp[3]) ? node55832 : node55825;
														assign node55825 = (inp[1]) ? node55829 : node55826;
															assign node55826 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node55829 = (inp[6]) ? 4'b0001 : 4'b0001;
														assign node55832 = (inp[6]) ? node55836 : node55833;
															assign node55833 = (inp[11]) ? 4'b0011 : 4'b1011;
															assign node55836 = (inp[1]) ? 4'b0011 : 4'b0011;
													assign node55839 = (inp[11]) ? node55847 : node55840;
														assign node55840 = (inp[3]) ? node55844 : node55841;
															assign node55841 = (inp[1]) ? 4'b0011 : 4'b0011;
															assign node55844 = (inp[6]) ? 4'b0011 : 4'b0011;
														assign node55847 = (inp[6]) ? node55851 : node55848;
															assign node55848 = (inp[1]) ? 4'b1011 : 4'b0011;
															assign node55851 = (inp[1]) ? 4'b0011 : 4'b1011;
												assign node55854 = (inp[3]) ? node55870 : node55855;
													assign node55855 = (inp[5]) ? node55863 : node55856;
														assign node55856 = (inp[6]) ? node55860 : node55857;
															assign node55857 = (inp[11]) ? 4'b0011 : 4'b0011;
															assign node55860 = (inp[11]) ? 4'b0011 : 4'b0011;
														assign node55863 = (inp[6]) ? node55867 : node55864;
															assign node55864 = (inp[1]) ? 4'b0001 : 4'b0001;
															assign node55867 = (inp[1]) ? 4'b0001 : 4'b0001;
													assign node55870 = (inp[11]) ? node55878 : node55871;
														assign node55871 = (inp[1]) ? node55875 : node55872;
															assign node55872 = (inp[6]) ? 4'b0001 : 4'b1001;
															assign node55875 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node55878 = (inp[6]) ? node55882 : node55879;
															assign node55879 = (inp[1]) ? 4'b1001 : 4'b0001;
															assign node55882 = (inp[1]) ? 4'b0001 : 4'b1001;
										assign node55885 = (inp[15]) ? node55945 : node55886;
											assign node55886 = (inp[0]) ? node55916 : node55887;
												assign node55887 = (inp[5]) ? node55903 : node55888;
													assign node55888 = (inp[3]) ? node55896 : node55889;
														assign node55889 = (inp[1]) ? node55893 : node55890;
															assign node55890 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node55893 = (inp[11]) ? 4'b0010 : 4'b0010;
														assign node55896 = (inp[6]) ? node55900 : node55897;
															assign node55897 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node55900 = (inp[1]) ? 4'b0000 : 4'b0000;
													assign node55903 = (inp[6]) ? node55909 : node55904;
														assign node55904 = (inp[11]) ? node55906 : 4'b0000;
															assign node55906 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node55909 = (inp[11]) ? node55913 : node55910;
															assign node55910 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node55913 = (inp[1]) ? 4'b0000 : 4'b1000;
												assign node55916 = (inp[3]) ? node55930 : node55917;
													assign node55917 = (inp[5]) ? node55925 : node55918;
														assign node55918 = (inp[11]) ? node55922 : node55919;
															assign node55919 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node55922 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node55925 = (inp[1]) ? 4'b0010 : node55926;
															assign node55926 = (inp[6]) ? 4'b1010 : 4'b0010;
													assign node55930 = (inp[5]) ? node55938 : node55931;
														assign node55931 = (inp[1]) ? node55935 : node55932;
															assign node55932 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node55935 = (inp[11]) ? 4'b0010 : 4'b0010;
														assign node55938 = (inp[11]) ? node55942 : node55939;
															assign node55939 = (inp[1]) ? 4'b1010 : 4'b0010;
															assign node55942 = (inp[6]) ? 4'b0010 : 4'b0010;
											assign node55945 = (inp[0]) ? node55977 : node55946;
												assign node55946 = (inp[5]) ? node55962 : node55947;
													assign node55947 = (inp[3]) ? node55955 : node55948;
														assign node55948 = (inp[11]) ? node55952 : node55949;
															assign node55949 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node55952 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node55955 = (inp[11]) ? node55959 : node55956;
															assign node55956 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node55959 = (inp[1]) ? 4'b0010 : 4'b0010;
													assign node55962 = (inp[11]) ? node55970 : node55963;
														assign node55963 = (inp[1]) ? node55967 : node55964;
															assign node55964 = (inp[6]) ? 4'b0010 : 4'b1010;
															assign node55967 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node55970 = (inp[1]) ? node55974 : node55971;
															assign node55971 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node55974 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node55977 = (inp[3]) ? node55991 : node55978;
													assign node55978 = (inp[5]) ? node55986 : node55979;
														assign node55979 = (inp[11]) ? node55983 : node55980;
															assign node55980 = (inp[1]) ? 4'b0010 : 4'b0010;
															assign node55983 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node55986 = (inp[11]) ? node55988 : 4'b1000;
															assign node55988 = (inp[1]) ? 4'b0000 : 4'b0000;
													assign node55991 = (inp[11]) ? node55997 : node55992;
														assign node55992 = (inp[1]) ? node55994 : 4'b0000;
															assign node55994 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node55997 = (inp[6]) ? node56001 : node55998;
															assign node55998 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node56001 = (inp[1]) ? 4'b0000 : 4'b1000;
									assign node56004 = (inp[6]) ? node56124 : node56005;
										assign node56005 = (inp[0]) ? node56061 : node56006;
											assign node56006 = (inp[15]) ? node56038 : node56007;
												assign node56007 = (inp[5]) ? node56023 : node56008;
													assign node56008 = (inp[3]) ? node56016 : node56009;
														assign node56009 = (inp[11]) ? node56013 : node56010;
															assign node56010 = (inp[1]) ? 4'b0010 : 4'b1010;
															assign node56013 = (inp[1]) ? 4'b1010 : 4'b0010;
														assign node56016 = (inp[11]) ? node56020 : node56017;
															assign node56017 = (inp[1]) ? 4'b0000 : 4'b1000;
															assign node56020 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node56023 = (inp[2]) ? node56031 : node56024;
														assign node56024 = (inp[3]) ? node56028 : node56025;
															assign node56025 = (inp[1]) ? 4'b0000 : 4'b0000;
															assign node56028 = (inp[11]) ? 4'b0000 : 4'b0000;
														assign node56031 = (inp[11]) ? node56035 : node56032;
															assign node56032 = (inp[1]) ? 4'b0000 : 4'b1000;
															assign node56035 = (inp[1]) ? 4'b1000 : 4'b0000;
												assign node56038 = (inp[5]) ? node56054 : node56039;
													assign node56039 = (inp[3]) ? node56047 : node56040;
														assign node56040 = (inp[2]) ? node56044 : node56041;
															assign node56041 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node56044 = (inp[1]) ? 4'b0000 : 4'b1000;
														assign node56047 = (inp[1]) ? node56051 : node56048;
															assign node56048 = (inp[11]) ? 4'b0010 : 4'b1010;
															assign node56051 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node56054 = (inp[1]) ? node56058 : node56055;
														assign node56055 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node56058 = (inp[11]) ? 4'b1010 : 4'b0010;
											assign node56061 = (inp[15]) ? node56093 : node56062;
												assign node56062 = (inp[3]) ? node56078 : node56063;
													assign node56063 = (inp[5]) ? node56071 : node56064;
														assign node56064 = (inp[1]) ? node56068 : node56065;
															assign node56065 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node56068 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node56071 = (inp[11]) ? node56075 : node56072;
															assign node56072 = (inp[1]) ? 4'b0010 : 4'b1010;
															assign node56075 = (inp[1]) ? 4'b1010 : 4'b0010;
													assign node56078 = (inp[2]) ? node56086 : node56079;
														assign node56079 = (inp[1]) ? node56083 : node56080;
															assign node56080 = (inp[11]) ? 4'b0010 : 4'b1010;
															assign node56083 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node56086 = (inp[11]) ? node56090 : node56087;
															assign node56087 = (inp[1]) ? 4'b0010 : 4'b1010;
															assign node56090 = (inp[1]) ? 4'b1010 : 4'b0010;
												assign node56093 = (inp[5]) ? node56109 : node56094;
													assign node56094 = (inp[3]) ? node56102 : node56095;
														assign node56095 = (inp[2]) ? node56099 : node56096;
															assign node56096 = (inp[1]) ? 4'b0010 : 4'b0010;
															assign node56099 = (inp[11]) ? 4'b0010 : 4'b0010;
														assign node56102 = (inp[11]) ? node56106 : node56103;
															assign node56103 = (inp[1]) ? 4'b0000 : 4'b1000;
															assign node56106 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node56109 = (inp[2]) ? node56117 : node56110;
														assign node56110 = (inp[3]) ? node56114 : node56111;
															assign node56111 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node56114 = (inp[1]) ? 4'b0000 : 4'b0000;
														assign node56117 = (inp[3]) ? node56121 : node56118;
															assign node56118 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node56121 = (inp[1]) ? 4'b0000 : 4'b0000;
										assign node56124 = (inp[5]) ? node56184 : node56125;
											assign node56125 = (inp[15]) ? node56155 : node56126;
												assign node56126 = (inp[11]) ? node56142 : node56127;
													assign node56127 = (inp[1]) ? node56135 : node56128;
														assign node56128 = (inp[2]) ? node56132 : node56129;
															assign node56129 = (inp[3]) ? 4'b0000 : 4'b0000;
															assign node56132 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node56135 = (inp[0]) ? node56139 : node56136;
															assign node56136 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node56139 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node56142 = (inp[1]) ? node56150 : node56143;
														assign node56143 = (inp[3]) ? node56147 : node56144;
															assign node56144 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node56147 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node56150 = (inp[2]) ? node56152 : 4'b0000;
															assign node56152 = (inp[3]) ? 4'b0000 : 4'b0000;
												assign node56155 = (inp[3]) ? node56171 : node56156;
													assign node56156 = (inp[0]) ? node56164 : node56157;
														assign node56157 = (inp[2]) ? node56161 : node56158;
															assign node56158 = (inp[1]) ? 4'b0000 : 4'b0000;
															assign node56161 = (inp[11]) ? 4'b0000 : 4'b0000;
														assign node56164 = (inp[1]) ? node56168 : node56165;
															assign node56165 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node56168 = (inp[11]) ? 4'b0010 : 4'b1010;
													assign node56171 = (inp[0]) ? node56179 : node56172;
														assign node56172 = (inp[2]) ? node56176 : node56173;
															assign node56173 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node56176 = (inp[1]) ? 4'b0010 : 4'b0010;
														assign node56179 = (inp[2]) ? 4'b0000 : node56180;
															assign node56180 = (inp[1]) ? 4'b0000 : 4'b0000;
											assign node56184 = (inp[1]) ? node56208 : node56185;
												assign node56185 = (inp[11]) ? node56201 : node56186;
													assign node56186 = (inp[3]) ? node56194 : node56187;
														assign node56187 = (inp[0]) ? node56191 : node56188;
															assign node56188 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node56191 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node56194 = (inp[0]) ? node56198 : node56195;
															assign node56195 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node56198 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node56201 = (inp[15]) ? node56205 : node56202;
														assign node56202 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node56205 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node56208 = (inp[11]) ? node56224 : node56209;
													assign node56209 = (inp[3]) ? node56217 : node56210;
														assign node56210 = (inp[0]) ? node56214 : node56211;
															assign node56211 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node56214 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node56217 = (inp[2]) ? node56221 : node56218;
															assign node56218 = (inp[15]) ? 4'b1000 : 4'b1000;
															assign node56221 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node56224 = (inp[15]) ? node56228 : node56225;
														assign node56225 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node56228 = (inp[0]) ? 4'b0000 : 4'b0010;
								assign node56231 = (inp[14]) ? node56451 : node56232;
									assign node56232 = (inp[2]) ? node56352 : node56233;
										assign node56233 = (inp[1]) ? node56293 : node56234;
											assign node56234 = (inp[0]) ? node56262 : node56235;
												assign node56235 = (inp[15]) ? node56247 : node56236;
													assign node56236 = (inp[5]) ? node56242 : node56237;
														assign node56237 = (inp[3]) ? 4'b1000 : node56238;
															assign node56238 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node56242 = (inp[6]) ? node56244 : 4'b1000;
															assign node56244 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node56247 = (inp[5]) ? node56255 : node56248;
														assign node56248 = (inp[3]) ? node56252 : node56249;
															assign node56249 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node56252 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node56255 = (inp[3]) ? node56259 : node56256;
															assign node56256 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node56259 = (inp[11]) ? 4'b0010 : 4'b0010;
												assign node56262 = (inp[15]) ? node56278 : node56263;
													assign node56263 = (inp[3]) ? node56271 : node56264;
														assign node56264 = (inp[5]) ? node56268 : node56265;
															assign node56265 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node56268 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node56271 = (inp[5]) ? node56275 : node56272;
															assign node56272 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node56275 = (inp[6]) ? 4'b0010 : 4'b0010;
													assign node56278 = (inp[5]) ? node56286 : node56279;
														assign node56279 = (inp[3]) ? node56283 : node56280;
															assign node56280 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node56283 = (inp[11]) ? 4'b0000 : 4'b0000;
														assign node56286 = (inp[3]) ? node56290 : node56287;
															assign node56287 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node56290 = (inp[6]) ? 4'b1000 : 4'b0000;
											assign node56293 = (inp[6]) ? node56323 : node56294;
												assign node56294 = (inp[11]) ? node56310 : node56295;
													assign node56295 = (inp[5]) ? node56303 : node56296;
														assign node56296 = (inp[0]) ? node56300 : node56297;
															assign node56297 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node56300 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node56303 = (inp[3]) ? node56307 : node56304;
															assign node56304 = (inp[0]) ? 4'b0000 : 4'b0000;
															assign node56307 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node56310 = (inp[5]) ? node56316 : node56311;
														assign node56311 = (inp[3]) ? 4'b1000 : node56312;
															assign node56312 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node56316 = (inp[3]) ? node56320 : node56317;
															assign node56317 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node56320 = (inp[15]) ? 4'b1000 : 4'b1000;
												assign node56323 = (inp[11]) ? node56337 : node56324;
													assign node56324 = (inp[5]) ? node56330 : node56325;
														assign node56325 = (inp[3]) ? 4'b1010 : node56326;
															assign node56326 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node56330 = (inp[15]) ? node56334 : node56331;
															assign node56331 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node56334 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node56337 = (inp[3]) ? node56345 : node56338;
														assign node56338 = (inp[5]) ? node56342 : node56339;
															assign node56339 = (inp[15]) ? 4'b0000 : 4'b0000;
															assign node56342 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node56345 = (inp[5]) ? node56349 : node56346;
															assign node56346 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node56349 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node56352 = (inp[6]) ? node56400 : node56353;
											assign node56353 = (inp[11]) ? node56377 : node56354;
												assign node56354 = (inp[15]) ? node56366 : node56355;
													assign node56355 = (inp[0]) ? node56361 : node56356;
														assign node56356 = (inp[3]) ? 4'b0001 : node56357;
															assign node56357 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node56361 = (inp[3]) ? 4'b0011 : node56362;
															assign node56362 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node56366 = (inp[0]) ? node56372 : node56367;
														assign node56367 = (inp[5]) ? 4'b0011 : node56368;
															assign node56368 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node56372 = (inp[5]) ? 4'b0001 : node56373;
															assign node56373 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node56377 = (inp[0]) ? node56389 : node56378;
													assign node56378 = (inp[15]) ? node56384 : node56379;
														assign node56379 = (inp[5]) ? 4'b1001 : node56380;
															assign node56380 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node56384 = (inp[3]) ? 4'b1011 : node56385;
															assign node56385 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node56389 = (inp[15]) ? node56395 : node56390;
														assign node56390 = (inp[3]) ? 4'b1011 : node56391;
															assign node56391 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node56395 = (inp[5]) ? 4'b1001 : node56396;
															assign node56396 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node56400 = (inp[11]) ? node56430 : node56401;
												assign node56401 = (inp[5]) ? node56417 : node56402;
													assign node56402 = (inp[15]) ? node56410 : node56403;
														assign node56403 = (inp[1]) ? node56407 : node56404;
															assign node56404 = (inp[0]) ? 4'b1001 : 4'b1001;
															assign node56407 = (inp[0]) ? 4'b1001 : 4'b1001;
														assign node56410 = (inp[1]) ? node56414 : node56411;
															assign node56411 = (inp[3]) ? 4'b1001 : 4'b1001;
															assign node56414 = (inp[0]) ? 4'b1001 : 4'b1001;
													assign node56417 = (inp[1]) ? node56425 : node56418;
														assign node56418 = (inp[0]) ? node56422 : node56419;
															assign node56419 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node56422 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node56425 = (inp[3]) ? 4'b1011 : node56426;
															assign node56426 = (inp[0]) ? 4'b1001 : 4'b1001;
												assign node56430 = (inp[3]) ? node56444 : node56431;
													assign node56431 = (inp[15]) ? node56437 : node56432;
														assign node56432 = (inp[5]) ? node56434 : 4'b0011;
															assign node56434 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node56437 = (inp[5]) ? node56441 : node56438;
															assign node56438 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node56441 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node56444 = (inp[0]) ? node56448 : node56445;
														assign node56445 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node56448 = (inp[15]) ? 4'b0001 : 4'b0011;
									assign node56451 = (inp[6]) ? node56507 : node56452;
										assign node56452 = (inp[11]) ? node56484 : node56453;
											assign node56453 = (inp[3]) ? node56477 : node56454;
												assign node56454 = (inp[15]) ? node56462 : node56455;
													assign node56455 = (inp[0]) ? node56459 : node56456;
														assign node56456 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node56459 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node56462 = (inp[1]) ? node56470 : node56463;
														assign node56463 = (inp[0]) ? node56467 : node56464;
															assign node56464 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node56467 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node56470 = (inp[5]) ? node56474 : node56471;
															assign node56471 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node56474 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node56477 = (inp[15]) ? node56481 : node56478;
													assign node56478 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node56481 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node56484 = (inp[15]) ? node56496 : node56485;
												assign node56485 = (inp[0]) ? node56491 : node56486;
													assign node56486 = (inp[3]) ? 4'b1001 : node56487;
														assign node56487 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node56491 = (inp[3]) ? 4'b1011 : node56492;
														assign node56492 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node56496 = (inp[0]) ? node56502 : node56497;
													assign node56497 = (inp[5]) ? 4'b1011 : node56498;
														assign node56498 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node56502 = (inp[5]) ? 4'b1001 : node56503;
														assign node56503 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node56507 = (inp[11]) ? node56531 : node56508;
											assign node56508 = (inp[15]) ? node56520 : node56509;
												assign node56509 = (inp[0]) ? node56515 : node56510;
													assign node56510 = (inp[5]) ? 4'b1001 : node56511;
														assign node56511 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node56515 = (inp[3]) ? 4'b1011 : node56516;
														assign node56516 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node56520 = (inp[0]) ? node56526 : node56521;
													assign node56521 = (inp[5]) ? 4'b1011 : node56522;
														assign node56522 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node56526 = (inp[3]) ? 4'b1001 : node56527;
														assign node56527 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node56531 = (inp[0]) ? node56543 : node56532;
												assign node56532 = (inp[15]) ? node56538 : node56533;
													assign node56533 = (inp[5]) ? 4'b0001 : node56534;
														assign node56534 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node56538 = (inp[3]) ? 4'b0011 : node56539;
														assign node56539 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node56543 = (inp[15]) ? node56549 : node56544;
													assign node56544 = (inp[5]) ? 4'b0011 : node56545;
														assign node56545 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node56549 = (inp[5]) ? 4'b0001 : node56550;
														assign node56550 = (inp[3]) ? 4'b0001 : 4'b0011;
							assign node56554 = (inp[7]) ? node56934 : node56555;
								assign node56555 = (inp[2]) ? node56777 : node56556;
									assign node56556 = (inp[14]) ? node56684 : node56557;
										assign node56557 = (inp[11]) ? node56621 : node56558;
											assign node56558 = (inp[0]) ? node56590 : node56559;
												assign node56559 = (inp[15]) ? node56575 : node56560;
													assign node56560 = (inp[3]) ? node56568 : node56561;
														assign node56561 = (inp[5]) ? node56565 : node56562;
															assign node56562 = (inp[1]) ? 4'b0010 : 4'b0010;
															assign node56565 = (inp[1]) ? 4'b0000 : 4'b0000;
														assign node56568 = (inp[1]) ? node56572 : node56569;
															assign node56569 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node56572 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node56575 = (inp[3]) ? node56583 : node56576;
														assign node56576 = (inp[5]) ? node56580 : node56577;
															assign node56577 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node56580 = (inp[1]) ? 4'b0010 : 4'b0010;
														assign node56583 = (inp[6]) ? node56587 : node56584;
															assign node56584 = (inp[1]) ? 4'b0010 : 4'b1010;
															assign node56587 = (inp[1]) ? 4'b1010 : 4'b0010;
												assign node56590 = (inp[15]) ? node56606 : node56591;
													assign node56591 = (inp[3]) ? node56599 : node56592;
														assign node56592 = (inp[5]) ? node56596 : node56593;
															assign node56593 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node56596 = (inp[6]) ? 4'b0010 : 4'b1010;
														assign node56599 = (inp[6]) ? node56603 : node56600;
															assign node56600 = (inp[1]) ? 4'b0010 : 4'b1010;
															assign node56603 = (inp[1]) ? 4'b1010 : 4'b0010;
													assign node56606 = (inp[5]) ? node56614 : node56607;
														assign node56607 = (inp[3]) ? node56611 : node56608;
															assign node56608 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node56611 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node56614 = (inp[6]) ? node56618 : node56615;
															assign node56615 = (inp[1]) ? 4'b0000 : 4'b1000;
															assign node56618 = (inp[1]) ? 4'b1000 : 4'b0000;
											assign node56621 = (inp[0]) ? node56653 : node56622;
												assign node56622 = (inp[15]) ? node56638 : node56623;
													assign node56623 = (inp[3]) ? node56631 : node56624;
														assign node56624 = (inp[5]) ? node56628 : node56625;
															assign node56625 = (inp[1]) ? 4'b0010 : 4'b0010;
															assign node56628 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node56631 = (inp[5]) ? node56635 : node56632;
															assign node56632 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node56635 = (inp[1]) ? 4'b1000 : 4'b0000;
													assign node56638 = (inp[3]) ? node56646 : node56639;
														assign node56639 = (inp[5]) ? node56643 : node56640;
															assign node56640 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node56643 = (inp[1]) ? 4'b0010 : 4'b0010;
														assign node56646 = (inp[5]) ? node56650 : node56647;
															assign node56647 = (inp[1]) ? 4'b0010 : 4'b0010;
															assign node56650 = (inp[6]) ? 4'b0010 : 4'b0010;
												assign node56653 = (inp[15]) ? node56669 : node56654;
													assign node56654 = (inp[3]) ? node56662 : node56655;
														assign node56655 = (inp[5]) ? node56659 : node56656;
															assign node56656 = (inp[1]) ? 4'b0000 : 4'b0000;
															assign node56659 = (inp[6]) ? 4'b0010 : 4'b0010;
														assign node56662 = (inp[6]) ? node56666 : node56663;
															assign node56663 = (inp[1]) ? 4'b1010 : 4'b0010;
															assign node56666 = (inp[1]) ? 4'b0010 : 4'b1010;
													assign node56669 = (inp[5]) ? node56677 : node56670;
														assign node56670 = (inp[3]) ? node56674 : node56671;
															assign node56671 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node56674 = (inp[1]) ? 4'b0000 : 4'b0000;
														assign node56677 = (inp[1]) ? node56681 : node56678;
															assign node56678 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node56681 = (inp[6]) ? 4'b0000 : 4'b1000;
										assign node56684 = (inp[6]) ? node56732 : node56685;
											assign node56685 = (inp[11]) ? node56709 : node56686;
												assign node56686 = (inp[3]) ? node56702 : node56687;
													assign node56687 = (inp[0]) ? node56695 : node56688;
														assign node56688 = (inp[1]) ? node56692 : node56689;
															assign node56689 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node56692 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node56695 = (inp[1]) ? node56699 : node56696;
															assign node56696 = (inp[5]) ? 4'b0001 : 4'b0001;
															assign node56699 = (inp[15]) ? 4'b0001 : 4'b0001;
													assign node56702 = (inp[15]) ? node56706 : node56703;
														assign node56703 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node56706 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node56709 = (inp[0]) ? node56721 : node56710;
													assign node56710 = (inp[15]) ? node56716 : node56711;
														assign node56711 = (inp[5]) ? 4'b1001 : node56712;
															assign node56712 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node56716 = (inp[3]) ? 4'b1011 : node56717;
															assign node56717 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node56721 = (inp[15]) ? node56727 : node56722;
														assign node56722 = (inp[3]) ? 4'b1011 : node56723;
															assign node56723 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node56727 = (inp[5]) ? 4'b1001 : node56728;
															assign node56728 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node56732 = (inp[11]) ? node56756 : node56733;
												assign node56733 = (inp[15]) ? node56745 : node56734;
													assign node56734 = (inp[0]) ? node56740 : node56735;
														assign node56735 = (inp[5]) ? 4'b1001 : node56736;
															assign node56736 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node56740 = (inp[3]) ? 4'b1011 : node56741;
															assign node56741 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node56745 = (inp[0]) ? node56751 : node56746;
														assign node56746 = (inp[5]) ? 4'b1011 : node56747;
															assign node56747 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node56751 = (inp[5]) ? 4'b1001 : node56752;
															assign node56752 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node56756 = (inp[15]) ? node56766 : node56757;
													assign node56757 = (inp[0]) ? node56763 : node56758;
														assign node56758 = (inp[3]) ? 4'b0001 : node56759;
															assign node56759 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node56763 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node56766 = (inp[0]) ? node56772 : node56767;
														assign node56767 = (inp[5]) ? 4'b0011 : node56768;
															assign node56768 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node56772 = (inp[3]) ? 4'b0001 : node56773;
															assign node56773 = (inp[5]) ? 4'b0001 : 4'b0011;
									assign node56777 = (inp[0]) ? node56849 : node56778;
										assign node56778 = (inp[15]) ? node56818 : node56779;
											assign node56779 = (inp[5]) ? node56795 : node56780;
												assign node56780 = (inp[3]) ? node56788 : node56781;
													assign node56781 = (inp[6]) ? node56785 : node56782;
														assign node56782 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node56785 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node56788 = (inp[11]) ? node56792 : node56789;
														assign node56789 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node56792 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node56795 = (inp[14]) ? node56811 : node56796;
													assign node56796 = (inp[3]) ? node56804 : node56797;
														assign node56797 = (inp[11]) ? node56801 : node56798;
															assign node56798 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node56801 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node56804 = (inp[6]) ? node56808 : node56805;
															assign node56805 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node56808 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node56811 = (inp[6]) ? node56815 : node56812;
														assign node56812 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node56815 = (inp[11]) ? 4'b0001 : 4'b1001;
											assign node56818 = (inp[5]) ? node56842 : node56819;
												assign node56819 = (inp[3]) ? node56835 : node56820;
													assign node56820 = (inp[1]) ? node56828 : node56821;
														assign node56821 = (inp[14]) ? node56825 : node56822;
															assign node56822 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node56825 = (inp[6]) ? 4'b0001 : 4'b0001;
														assign node56828 = (inp[6]) ? node56832 : node56829;
															assign node56829 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node56832 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node56835 = (inp[11]) ? node56839 : node56836;
														assign node56836 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node56839 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node56842 = (inp[11]) ? node56846 : node56843;
													assign node56843 = (inp[6]) ? 4'b1011 : 4'b0011;
													assign node56846 = (inp[6]) ? 4'b0011 : 4'b1011;
										assign node56849 = (inp[15]) ? node56895 : node56850;
											assign node56850 = (inp[5]) ? node56866 : node56851;
												assign node56851 = (inp[3]) ? node56859 : node56852;
													assign node56852 = (inp[11]) ? node56856 : node56853;
														assign node56853 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node56856 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node56859 = (inp[6]) ? node56863 : node56860;
														assign node56860 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node56863 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node56866 = (inp[1]) ? node56880 : node56867;
													assign node56867 = (inp[3]) ? node56875 : node56868;
														assign node56868 = (inp[11]) ? node56872 : node56869;
															assign node56869 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node56872 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node56875 = (inp[11]) ? node56877 : 4'b0011;
															assign node56877 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node56880 = (inp[14]) ? node56888 : node56881;
														assign node56881 = (inp[3]) ? node56885 : node56882;
															assign node56882 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node56885 = (inp[6]) ? 4'b0011 : 4'b0011;
														assign node56888 = (inp[3]) ? node56892 : node56889;
															assign node56889 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node56892 = (inp[11]) ? 4'b0011 : 4'b0011;
											assign node56895 = (inp[3]) ? node56919 : node56896;
												assign node56896 = (inp[5]) ? node56912 : node56897;
													assign node56897 = (inp[14]) ? node56905 : node56898;
														assign node56898 = (inp[11]) ? node56902 : node56899;
															assign node56899 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node56902 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node56905 = (inp[6]) ? node56909 : node56906;
															assign node56906 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node56909 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node56912 = (inp[6]) ? node56916 : node56913;
														assign node56913 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node56916 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node56919 = (inp[1]) ? node56927 : node56920;
													assign node56920 = (inp[11]) ? node56924 : node56921;
														assign node56921 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node56924 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node56927 = (inp[6]) ? node56931 : node56928;
														assign node56928 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node56931 = (inp[11]) ? 4'b0001 : 4'b1001;
								assign node56934 = (inp[14]) ? node57134 : node56935;
									assign node56935 = (inp[2]) ? node57037 : node56936;
										assign node56936 = (inp[0]) ? node56982 : node56937;
											assign node56937 = (inp[15]) ? node56959 : node56938;
												assign node56938 = (inp[3]) ? node56952 : node56939;
													assign node56939 = (inp[5]) ? node56947 : node56940;
														assign node56940 = (inp[1]) ? node56944 : node56941;
															assign node56941 = (inp[11]) ? 4'b0011 : 4'b0011;
															assign node56944 = (inp[6]) ? 4'b0011 : 4'b0011;
														assign node56947 = (inp[11]) ? node56949 : 4'b1001;
															assign node56949 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node56952 = (inp[11]) ? node56956 : node56953;
														assign node56953 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node56956 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node56959 = (inp[5]) ? node56975 : node56960;
													assign node56960 = (inp[3]) ? node56968 : node56961;
														assign node56961 = (inp[6]) ? node56965 : node56962;
															assign node56962 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node56965 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node56968 = (inp[1]) ? node56972 : node56969;
															assign node56969 = (inp[6]) ? 4'b0011 : 4'b0011;
															assign node56972 = (inp[6]) ? 4'b0011 : 4'b0011;
													assign node56975 = (inp[6]) ? node56979 : node56976;
														assign node56976 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node56979 = (inp[11]) ? 4'b0011 : 4'b1011;
											assign node56982 = (inp[15]) ? node57006 : node56983;
												assign node56983 = (inp[5]) ? node56999 : node56984;
													assign node56984 = (inp[3]) ? node56992 : node56985;
														assign node56985 = (inp[1]) ? node56989 : node56986;
															assign node56986 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node56989 = (inp[11]) ? 4'b0001 : 4'b0001;
														assign node56992 = (inp[11]) ? node56996 : node56993;
															assign node56993 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node56996 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node56999 = (inp[6]) ? node57003 : node57000;
														assign node57000 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node57003 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node57006 = (inp[5]) ? node57022 : node57007;
													assign node57007 = (inp[3]) ? node57015 : node57008;
														assign node57008 = (inp[1]) ? node57012 : node57009;
															assign node57009 = (inp[11]) ? 4'b0011 : 4'b0011;
															assign node57012 = (inp[6]) ? 4'b0011 : 4'b0011;
														assign node57015 = (inp[1]) ? node57019 : node57016;
															assign node57016 = (inp[6]) ? 4'b0001 : 4'b0001;
															assign node57019 = (inp[6]) ? 4'b0001 : 4'b0001;
													assign node57022 = (inp[3]) ? node57030 : node57023;
														assign node57023 = (inp[11]) ? node57027 : node57024;
															assign node57024 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node57027 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node57030 = (inp[11]) ? node57034 : node57031;
															assign node57031 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node57034 = (inp[6]) ? 4'b0001 : 4'b1001;
										assign node57037 = (inp[3]) ? node57097 : node57038;
											assign node57038 = (inp[0]) ? node57068 : node57039;
												assign node57039 = (inp[15]) ? node57053 : node57040;
													assign node57040 = (inp[5]) ? node57048 : node57041;
														assign node57041 = (inp[11]) ? node57045 : node57042;
															assign node57042 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node57045 = (inp[6]) ? 4'b0010 : 4'b1010;
														assign node57048 = (inp[11]) ? 4'b0000 : node57049;
															assign node57049 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node57053 = (inp[5]) ? node57061 : node57054;
														assign node57054 = (inp[11]) ? node57058 : node57055;
															assign node57055 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node57058 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node57061 = (inp[1]) ? node57065 : node57062;
															assign node57062 = (inp[6]) ? 4'b0010 : 4'b0010;
															assign node57065 = (inp[11]) ? 4'b0010 : 4'b0010;
												assign node57068 = (inp[1]) ? node57084 : node57069;
													assign node57069 = (inp[11]) ? node57077 : node57070;
														assign node57070 = (inp[6]) ? node57074 : node57071;
															assign node57071 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node57074 = (inp[15]) ? 4'b1000 : 4'b1000;
														assign node57077 = (inp[6]) ? node57081 : node57078;
															assign node57078 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node57081 = (inp[15]) ? 4'b0000 : 4'b0000;
													assign node57084 = (inp[15]) ? node57090 : node57085;
														assign node57085 = (inp[5]) ? 4'b0010 : node57086;
															assign node57086 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node57090 = (inp[5]) ? node57094 : node57091;
															assign node57091 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node57094 = (inp[6]) ? 4'b0000 : 4'b0000;
											assign node57097 = (inp[6]) ? node57119 : node57098;
												assign node57098 = (inp[11]) ? node57112 : node57099;
													assign node57099 = (inp[1]) ? node57105 : node57100;
														assign node57100 = (inp[5]) ? 4'b0000 : node57101;
															assign node57101 = (inp[15]) ? 4'b0000 : 4'b0000;
														assign node57105 = (inp[15]) ? node57109 : node57106;
															assign node57106 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node57109 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node57112 = (inp[15]) ? node57116 : node57113;
														assign node57113 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node57116 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node57119 = (inp[11]) ? node57127 : node57120;
													assign node57120 = (inp[15]) ? node57124 : node57121;
														assign node57121 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node57124 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node57127 = (inp[15]) ? node57131 : node57128;
														assign node57128 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node57131 = (inp[0]) ? 4'b0000 : 4'b0010;
									assign node57134 = (inp[0]) ? node57230 : node57135;
										assign node57135 = (inp[15]) ? node57191 : node57136;
											assign node57136 = (inp[5]) ? node57168 : node57137;
												assign node57137 = (inp[3]) ? node57153 : node57138;
													assign node57138 = (inp[1]) ? node57146 : node57139;
														assign node57139 = (inp[11]) ? node57143 : node57140;
															assign node57140 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node57143 = (inp[6]) ? 4'b0010 : 4'b1010;
														assign node57146 = (inp[11]) ? node57150 : node57147;
															assign node57147 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node57150 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node57153 = (inp[2]) ? node57161 : node57154;
														assign node57154 = (inp[1]) ? node57158 : node57155;
															assign node57155 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node57158 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node57161 = (inp[1]) ? node57165 : node57162;
															assign node57162 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node57165 = (inp[6]) ? 4'b0000 : 4'b0000;
												assign node57168 = (inp[3]) ? node57184 : node57169;
													assign node57169 = (inp[2]) ? node57177 : node57170;
														assign node57170 = (inp[1]) ? node57174 : node57171;
															assign node57171 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node57174 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node57177 = (inp[1]) ? node57181 : node57178;
															assign node57178 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node57181 = (inp[11]) ? 4'b0000 : 4'b0000;
													assign node57184 = (inp[11]) ? node57188 : node57185;
														assign node57185 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node57188 = (inp[6]) ? 4'b0000 : 4'b1000;
											assign node57191 = (inp[3]) ? node57223 : node57192;
												assign node57192 = (inp[5]) ? node57208 : node57193;
													assign node57193 = (inp[2]) ? node57201 : node57194;
														assign node57194 = (inp[1]) ? node57198 : node57195;
															assign node57195 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node57198 = (inp[11]) ? 4'b0000 : 4'b0000;
														assign node57201 = (inp[6]) ? node57205 : node57202;
															assign node57202 = (inp[11]) ? 4'b1000 : 4'b0000;
															assign node57205 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node57208 = (inp[1]) ? node57216 : node57209;
														assign node57209 = (inp[6]) ? node57213 : node57210;
															assign node57210 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node57213 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node57216 = (inp[2]) ? node57220 : node57217;
															assign node57217 = (inp[11]) ? 4'b0010 : 4'b0010;
															assign node57220 = (inp[6]) ? 4'b0010 : 4'b0010;
												assign node57223 = (inp[11]) ? node57227 : node57224;
													assign node57224 = (inp[6]) ? 4'b1010 : 4'b0010;
													assign node57227 = (inp[6]) ? 4'b0010 : 4'b1010;
										assign node57230 = (inp[15]) ? node57284 : node57231;
											assign node57231 = (inp[5]) ? node57253 : node57232;
												assign node57232 = (inp[3]) ? node57246 : node57233;
													assign node57233 = (inp[1]) ? node57241 : node57234;
														assign node57234 = (inp[2]) ? node57238 : node57235;
															assign node57235 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node57238 = (inp[6]) ? 4'b0000 : 4'b0000;
														assign node57241 = (inp[2]) ? node57243 : 4'b1000;
															assign node57243 = (inp[11]) ? 4'b0000 : 4'b0000;
													assign node57246 = (inp[6]) ? node57250 : node57247;
														assign node57247 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node57250 = (inp[11]) ? 4'b0010 : 4'b1010;
												assign node57253 = (inp[3]) ? node57269 : node57254;
													assign node57254 = (inp[2]) ? node57262 : node57255;
														assign node57255 = (inp[6]) ? node57259 : node57256;
															assign node57256 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node57259 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node57262 = (inp[11]) ? node57266 : node57263;
															assign node57263 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node57266 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node57269 = (inp[2]) ? node57277 : node57270;
														assign node57270 = (inp[6]) ? node57274 : node57271;
															assign node57271 = (inp[11]) ? 4'b1010 : 4'b0010;
															assign node57274 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node57277 = (inp[11]) ? node57281 : node57278;
															assign node57278 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node57281 = (inp[6]) ? 4'b0010 : 4'b1010;
											assign node57284 = (inp[5]) ? node57306 : node57285;
												assign node57285 = (inp[3]) ? node57293 : node57286;
													assign node57286 = (inp[11]) ? node57290 : node57287;
														assign node57287 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node57290 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node57293 = (inp[2]) ? node57301 : node57294;
														assign node57294 = (inp[1]) ? node57298 : node57295;
															assign node57295 = (inp[6]) ? 4'b0000 : 4'b0000;
															assign node57298 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node57301 = (inp[1]) ? node57303 : 4'b0000;
															assign node57303 = (inp[11]) ? 4'b0000 : 4'b0000;
												assign node57306 = (inp[11]) ? node57310 : node57307;
													assign node57307 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node57310 = (inp[6]) ? 4'b0000 : 4'b1000;

endmodule