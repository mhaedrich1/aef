module dtc_split75_bm91 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node41;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node123;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node234;
	wire [3-1:0] node236;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node285;
	wire [3-1:0] node287;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node299;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node315;
	wire [3-1:0] node317;
	wire [3-1:0] node320;
	wire [3-1:0] node322;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node354;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node377;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node383;
	wire [3-1:0] node386;
	wire [3-1:0] node389;
	wire [3-1:0] node391;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node401;
	wire [3-1:0] node403;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node419;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node429;
	wire [3-1:0] node431;
	wire [3-1:0] node433;
	wire [3-1:0] node436;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node444;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node455;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node463;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node473;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node480;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node488;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node499;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node517;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node526;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node536;
	wire [3-1:0] node539;
	wire [3-1:0] node541;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node561;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node574;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node582;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node589;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node595;
	wire [3-1:0] node598;
	wire [3-1:0] node600;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node612;
	wire [3-1:0] node614;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node621;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node630;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node650;
	wire [3-1:0] node652;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node667;
	wire [3-1:0] node669;
	wire [3-1:0] node671;
	wire [3-1:0] node673;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node681;
	wire [3-1:0] node684;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node693;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node716;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node728;
	wire [3-1:0] node731;
	wire [3-1:0] node734;
	wire [3-1:0] node735;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node742;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node756;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node761;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node768;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node789;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node815;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node822;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node835;
	wire [3-1:0] node837;
	wire [3-1:0] node840;
	wire [3-1:0] node841;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node851;
	wire [3-1:0] node854;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node865;
	wire [3-1:0] node869;
	wire [3-1:0] node870;
	wire [3-1:0] node872;
	wire [3-1:0] node875;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node882;
	wire [3-1:0] node884;
	wire [3-1:0] node886;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node903;
	wire [3-1:0] node905;
	wire [3-1:0] node907;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node918;
	wire [3-1:0] node920;
	wire [3-1:0] node922;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node931;
	wire [3-1:0] node933;
	wire [3-1:0] node936;
	wire [3-1:0] node938;
	wire [3-1:0] node941;
	wire [3-1:0] node942;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node964;
	wire [3-1:0] node967;
	wire [3-1:0] node970;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node977;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node986;
	wire [3-1:0] node988;
	wire [3-1:0] node991;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node1000;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1007;
	wire [3-1:0] node1009;
	wire [3-1:0] node1011;
	wire [3-1:0] node1014;
	wire [3-1:0] node1016;
	wire [3-1:0] node1018;
	wire [3-1:0] node1020;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1027;
	wire [3-1:0] node1031;
	wire [3-1:0] node1033;
	wire [3-1:0] node1034;
	wire [3-1:0] node1037;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1042;
	wire [3-1:0] node1045;
	wire [3-1:0] node1048;
	wire [3-1:0] node1049;
	wire [3-1:0] node1052;
	wire [3-1:0] node1055;
	wire [3-1:0] node1056;
	wire [3-1:0] node1058;
	wire [3-1:0] node1059;
	wire [3-1:0] node1060;
	wire [3-1:0] node1065;
	wire [3-1:0] node1066;
	wire [3-1:0] node1067;
	wire [3-1:0] node1071;
	wire [3-1:0] node1072;
	wire [3-1:0] node1076;
	wire [3-1:0] node1077;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1081;
	wire [3-1:0] node1083;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1089;
	wire [3-1:0] node1091;
	wire [3-1:0] node1094;
	wire [3-1:0] node1095;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1105;
	wire [3-1:0] node1108;
	wire [3-1:0] node1110;
	wire [3-1:0] node1114;
	wire [3-1:0] node1115;
	wire [3-1:0] node1116;
	wire [3-1:0] node1118;
	wire [3-1:0] node1121;
	wire [3-1:0] node1123;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1128;
	wire [3-1:0] node1129;
	wire [3-1:0] node1131;
	wire [3-1:0] node1136;
	wire [3-1:0] node1137;
	wire [3-1:0] node1138;
	wire [3-1:0] node1142;
	wire [3-1:0] node1143;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1152;
	wire [3-1:0] node1155;
	wire [3-1:0] node1156;
	wire [3-1:0] node1160;
	wire [3-1:0] node1161;
	wire [3-1:0] node1162;
	wire [3-1:0] node1166;

	assign outp = (inp[3]) ? node878 : node1;
		assign node1 = (inp[9]) ? node447 : node2;
			assign node2 = (inp[1]) ? node216 : node3;
				assign node3 = (inp[10]) ? node91 : node4;
					assign node4 = (inp[6]) ? node38 : node5;
						assign node5 = (inp[4]) ? node27 : node6;
							assign node6 = (inp[7]) ? node22 : node7;
								assign node7 = (inp[5]) ? node15 : node8;
									assign node8 = (inp[0]) ? node10 : 3'b001;
										assign node10 = (inp[2]) ? 3'b000 : node11;
											assign node11 = (inp[8]) ? 3'b000 : 3'b001;
									assign node15 = (inp[0]) ? node17 : 3'b000;
										assign node17 = (inp[2]) ? 3'b001 : node18;
											assign node18 = (inp[8]) ? 3'b000 : 3'b001;
								assign node22 = (inp[0]) ? node24 : 3'b001;
									assign node24 = (inp[5]) ? 3'b001 : 3'b000;
							assign node27 = (inp[0]) ? node29 : 3'b000;
								assign node29 = (inp[5]) ? 3'b000 : node30;
									assign node30 = (inp[2]) ? 3'b001 : node31;
										assign node31 = (inp[8]) ? 3'b001 : node32;
											assign node32 = (inp[7]) ? 3'b001 : 3'b000;
						assign node38 = (inp[5]) ? node48 : node39;
							assign node39 = (inp[8]) ? node41 : 3'b000;
								assign node41 = (inp[4]) ? node43 : 3'b000;
									assign node43 = (inp[7]) ? 3'b000 : node44;
										assign node44 = (inp[0]) ? 3'b000 : 3'b001;
							assign node48 = (inp[7]) ? node78 : node49;
								assign node49 = (inp[8]) ? node67 : node50;
									assign node50 = (inp[11]) ? node58 : node51;
										assign node51 = (inp[4]) ? node55 : node52;
											assign node52 = (inp[0]) ? 3'b000 : 3'b001;
											assign node55 = (inp[0]) ? 3'b001 : 3'b000;
										assign node58 = (inp[2]) ? node64 : node59;
											assign node59 = (inp[4]) ? 3'b000 : node60;
												assign node60 = (inp[0]) ? 3'b000 : 3'b001;
											assign node64 = (inp[0]) ? 3'b001 : 3'b000;
									assign node67 = (inp[11]) ? node73 : node68;
										assign node68 = (inp[4]) ? 3'b001 : node69;
											assign node69 = (inp[0]) ? 3'b000 : 3'b001;
										assign node73 = (inp[4]) ? node75 : 3'b001;
											assign node75 = (inp[0]) ? 3'b001 : 3'b000;
								assign node78 = (inp[8]) ? node86 : node79;
									assign node79 = (inp[0]) ? node83 : node80;
										assign node80 = (inp[4]) ? 3'b000 : 3'b001;
										assign node83 = (inp[4]) ? 3'b001 : 3'b000;
									assign node86 = (inp[4]) ? node88 : 3'b000;
										assign node88 = (inp[0]) ? 3'b001 : 3'b000;
					assign node91 = (inp[7]) ? node181 : node92;
						assign node92 = (inp[8]) ? node140 : node93;
							assign node93 = (inp[4]) ? node123 : node94;
								assign node94 = (inp[2]) ? node106 : node95;
									assign node95 = (inp[6]) ? node101 : node96;
										assign node96 = (inp[5]) ? node98 : 3'b001;
											assign node98 = (inp[0]) ? 3'b001 : 3'b000;
										assign node101 = (inp[0]) ? 3'b000 : node102;
											assign node102 = (inp[5]) ? 3'b001 : 3'b000;
									assign node106 = (inp[11]) ? node116 : node107;
										assign node107 = (inp[6]) ? 3'b000 : node108;
											assign node108 = (inp[0]) ? node112 : node109;
												assign node109 = (inp[5]) ? 3'b000 : 3'b001;
												assign node112 = (inp[5]) ? 3'b001 : 3'b000;
										assign node116 = (inp[0]) ? 3'b000 : node117;
											assign node117 = (inp[5]) ? node119 : 3'b000;
												assign node119 = (inp[6]) ? 3'b001 : 3'b000;
								assign node123 = (inp[0]) ? node125 : 3'b000;
									assign node125 = (inp[2]) ? node133 : node126;
										assign node126 = (inp[11]) ? node128 : 3'b000;
											assign node128 = (inp[5]) ? node130 : 3'b000;
												assign node130 = (inp[6]) ? 3'b001 : 3'b000;
										assign node133 = (inp[5]) ? node137 : node134;
											assign node134 = (inp[6]) ? 3'b000 : 3'b001;
											assign node137 = (inp[6]) ? 3'b001 : 3'b000;
							assign node140 = (inp[5]) ? node162 : node141;
								assign node141 = (inp[6]) ? node157 : node142;
									assign node142 = (inp[2]) ? node150 : node143;
										assign node143 = (inp[4]) ? node147 : node144;
											assign node144 = (inp[0]) ? 3'b000 : 3'b001;
											assign node147 = (inp[0]) ? 3'b001 : 3'b000;
										assign node150 = (inp[0]) ? node154 : node151;
											assign node151 = (inp[4]) ? 3'b000 : 3'b001;
											assign node154 = (inp[4]) ? 3'b001 : 3'b000;
									assign node157 = (inp[0]) ? 3'b000 : node158;
										assign node158 = (inp[4]) ? 3'b001 : 3'b000;
								assign node162 = (inp[6]) ? node176 : node163;
									assign node163 = (inp[0]) ? node165 : 3'b000;
										assign node165 = (inp[4]) ? node171 : node166;
											assign node166 = (inp[2]) ? 3'b001 : node167;
												assign node167 = (inp[11]) ? 3'b001 : 3'b000;
											assign node171 = (inp[11]) ? 3'b000 : node172;
												assign node172 = (inp[2]) ? 3'b000 : 3'b001;
									assign node176 = (inp[0]) ? node178 : 3'b001;
										assign node178 = (inp[4]) ? 3'b001 : 3'b000;
						assign node181 = (inp[4]) ? node199 : node182;
							assign node182 = (inp[6]) ? node188 : node183;
								assign node183 = (inp[0]) ? node185 : 3'b001;
									assign node185 = (inp[5]) ? 3'b001 : 3'b000;
								assign node188 = (inp[0]) ? node194 : node189;
									assign node189 = (inp[8]) ? 3'b000 : node190;
										assign node190 = (inp[5]) ? 3'b001 : 3'b000;
									assign node194 = (inp[2]) ? 3'b001 : node195;
										assign node195 = (inp[5]) ? 3'b000 : 3'b001;
							assign node199 = (inp[6]) ? node205 : node200;
								assign node200 = (inp[0]) ? node202 : 3'b000;
									assign node202 = (inp[5]) ? 3'b000 : 3'b001;
								assign node205 = (inp[5]) ? node209 : node206;
									assign node206 = (inp[0]) ? 3'b000 : 3'b001;
									assign node209 = (inp[8]) ? 3'b001 : node210;
										assign node210 = (inp[0]) ? 3'b001 : node211;
											assign node211 = (inp[2]) ? 3'b001 : 3'b000;
				assign node216 = (inp[8]) ? node340 : node217;
					assign node217 = (inp[4]) ? node269 : node218;
						assign node218 = (inp[0]) ? node260 : node219;
							assign node219 = (inp[6]) ? node241 : node220;
								assign node220 = (inp[7]) ? node228 : node221;
									assign node221 = (inp[10]) ? 3'b001 : node222;
										assign node222 = (inp[5]) ? 3'b001 : node223;
											assign node223 = (inp[2]) ? 3'b001 : 3'b000;
									assign node228 = (inp[10]) ? node234 : node229;
										assign node229 = (inp[11]) ? 3'b000 : node230;
											assign node230 = (inp[2]) ? 3'b001 : 3'b000;
										assign node234 = (inp[2]) ? node236 : 3'b001;
											assign node236 = (inp[5]) ? node238 : 3'b000;
												assign node238 = (inp[11]) ? 3'b001 : 3'b000;
								assign node241 = (inp[7]) ? node249 : node242;
									assign node242 = (inp[5]) ? 3'b000 : node243;
										assign node243 = (inp[11]) ? node245 : 3'b000;
											assign node245 = (inp[2]) ? 3'b000 : 3'b001;
									assign node249 = (inp[10]) ? node255 : node250;
										assign node250 = (inp[11]) ? node252 : 3'b001;
											assign node252 = (inp[2]) ? 3'b001 : 3'b000;
										assign node255 = (inp[5]) ? 3'b000 : node256;
											assign node256 = (inp[2]) ? 3'b000 : 3'b001;
							assign node260 = (inp[5]) ? node264 : node261;
								assign node261 = (inp[6]) ? 3'b001 : 3'b000;
								assign node264 = (inp[7]) ? 3'b000 : node265;
									assign node265 = (inp[6]) ? 3'b000 : 3'b001;
						assign node269 = (inp[10]) ? node311 : node270;
							assign node270 = (inp[2]) ? node290 : node271;
								assign node271 = (inp[6]) ? node279 : node272;
									assign node272 = (inp[5]) ? node274 : 3'b001;
										assign node274 = (inp[7]) ? 3'b001 : node275;
											assign node275 = (inp[0]) ? 3'b001 : 3'b000;
									assign node279 = (inp[0]) ? node285 : node280;
										assign node280 = (inp[5]) ? node282 : 3'b001;
											assign node282 = (inp[7]) ? 3'b001 : 3'b000;
										assign node285 = (inp[11]) ? node287 : 3'b000;
											assign node287 = (inp[7]) ? 3'b000 : 3'b001;
								assign node290 = (inp[0]) ? node304 : node291;
									assign node291 = (inp[6]) ? node297 : node292;
										assign node292 = (inp[5]) ? node294 : 3'b000;
											assign node294 = (inp[7]) ? 3'b001 : 3'b000;
										assign node297 = (inp[5]) ? node299 : 3'b001;
											assign node299 = (inp[7]) ? node301 : 3'b000;
												assign node301 = (inp[11]) ? 3'b000 : 3'b001;
									assign node304 = (inp[6]) ? node306 : 3'b001;
										assign node306 = (inp[7]) ? 3'b000 : node307;
											assign node307 = (inp[5]) ? 3'b001 : 3'b000;
							assign node311 = (inp[0]) ? node325 : node312;
								assign node312 = (inp[6]) ? node320 : node313;
									assign node313 = (inp[7]) ? node315 : 3'b000;
										assign node315 = (inp[2]) ? node317 : 3'b000;
											assign node317 = (inp[5]) ? 3'b000 : 3'b001;
									assign node320 = (inp[5]) ? node322 : 3'b001;
										assign node322 = (inp[7]) ? 3'b001 : 3'b000;
								assign node325 = (inp[6]) ? node335 : node326;
									assign node326 = (inp[11]) ? node328 : 3'b001;
										assign node328 = (inp[2]) ? 3'b001 : node329;
											assign node329 = (inp[7]) ? 3'b001 : node330;
												assign node330 = (inp[5]) ? 3'b000 : 3'b001;
									assign node335 = (inp[7]) ? 3'b000 : node336;
										assign node336 = (inp[5]) ? 3'b001 : 3'b000;
					assign node340 = (inp[5]) ? node394 : node341;
						assign node341 = (inp[7]) ? node369 : node342;
							assign node342 = (inp[0]) ? node364 : node343;
								assign node343 = (inp[10]) ? node349 : node344;
									assign node344 = (inp[6]) ? 3'b001 : node345;
										assign node345 = (inp[4]) ? 3'b001 : 3'b000;
									assign node349 = (inp[11]) ? node357 : node350;
										assign node350 = (inp[6]) ? node354 : node351;
											assign node351 = (inp[4]) ? 3'b000 : 3'b001;
											assign node354 = (inp[4]) ? 3'b001 : 3'b000;
										assign node357 = (inp[6]) ? node361 : node358;
											assign node358 = (inp[4]) ? 3'b000 : 3'b001;
											assign node361 = (inp[4]) ? 3'b001 : 3'b000;
								assign node364 = (inp[4]) ? 3'b000 : node365;
									assign node365 = (inp[6]) ? 3'b001 : 3'b000;
							assign node369 = (inp[0]) ? node389 : node370;
								assign node370 = (inp[4]) ? node380 : node371;
									assign node371 = (inp[6]) ? node377 : node372;
										assign node372 = (inp[2]) ? 3'b000 : node373;
											assign node373 = (inp[10]) ? 3'b000 : 3'b001;
										assign node377 = (inp[10]) ? 3'b001 : 3'b000;
									assign node380 = (inp[6]) ? node386 : node381;
										assign node381 = (inp[11]) ? node383 : 3'b001;
											assign node383 = (inp[2]) ? 3'b001 : 3'b000;
										assign node386 = (inp[2]) ? 3'b000 : 3'b001;
								assign node389 = (inp[6]) ? node391 : 3'b001;
									assign node391 = (inp[4]) ? 3'b000 : 3'b001;
						assign node394 = (inp[0]) ? node436 : node395;
							assign node395 = (inp[7]) ? node413 : node396;
								assign node396 = (inp[4]) ? node406 : node397;
									assign node397 = (inp[6]) ? node401 : node398;
										assign node398 = (inp[11]) ? 3'b001 : 3'b000;
										assign node401 = (inp[2]) ? node403 : 3'b000;
											assign node403 = (inp[11]) ? 3'b000 : 3'b001;
									assign node406 = (inp[6]) ? 3'b000 : node407;
										assign node407 = (inp[10]) ? 3'b000 : node408;
											assign node408 = (inp[2]) ? 3'b001 : 3'b000;
								assign node413 = (inp[11]) ? node429 : node414;
									assign node414 = (inp[6]) ? node422 : node415;
										assign node415 = (inp[10]) ? node419 : node416;
											assign node416 = (inp[4]) ? 3'b000 : 3'b001;
											assign node419 = (inp[4]) ? 3'b001 : 3'b000;
										assign node422 = (inp[4]) ? 3'b001 : node423;
											assign node423 = (inp[10]) ? 3'b001 : node424;
												assign node424 = (inp[2]) ? 3'b000 : 3'b001;
									assign node429 = (inp[10]) ? node431 : 3'b001;
										assign node431 = (inp[2]) ? node433 : 3'b001;
											assign node433 = (inp[4]) ? 3'b001 : 3'b000;
							assign node436 = (inp[7]) ? node438 : 3'b001;
								assign node438 = (inp[6]) ? node444 : node439;
									assign node439 = (inp[4]) ? 3'b001 : node440;
										assign node440 = (inp[11]) ? 3'b000 : 3'b001;
									assign node444 = (inp[4]) ? 3'b000 : 3'b001;
			assign node447 = (inp[4]) ? node697 : node448;
				assign node448 = (inp[6]) ? node564 : node449;
					assign node449 = (inp[0]) ? node503 : node450;
						assign node450 = (inp[1]) ? node458 : node451;
							assign node451 = (inp[7]) ? node455 : node452;
								assign node452 = (inp[5]) ? 3'b100 : 3'b010;
								assign node455 = (inp[5]) ? 3'b010 : 3'b110;
							assign node458 = (inp[5]) ? node488 : node459;
								assign node459 = (inp[7]) ? node467 : node460;
									assign node460 = (inp[10]) ? 3'b110 : node461;
										assign node461 = (inp[2]) ? node463 : 3'b101;
											assign node463 = (inp[8]) ? 3'b101 : 3'b110;
									assign node467 = (inp[8]) ? node483 : node468;
										assign node468 = (inp[11]) ? node476 : node469;
											assign node469 = (inp[10]) ? node473 : node470;
												assign node470 = (inp[2]) ? 3'b010 : 3'b001;
												assign node473 = (inp[2]) ? 3'b001 : 3'b010;
											assign node476 = (inp[2]) ? node480 : node477;
												assign node477 = (inp[10]) ? 3'b110 : 3'b101;
												assign node480 = (inp[10]) ? 3'b001 : 3'b010;
										assign node483 = (inp[2]) ? 3'b001 : node484;
											assign node484 = (inp[10]) ? 3'b001 : 3'b010;
								assign node488 = (inp[7]) ? node490 : 3'b010;
									assign node490 = (inp[8]) ? 3'b110 : node491;
										assign node491 = (inp[2]) ? node495 : node492;
											assign node492 = (inp[10]) ? 3'b010 : 3'b001;
											assign node495 = (inp[10]) ? node499 : node496;
												assign node496 = (inp[11]) ? 3'b101 : 3'b110;
												assign node499 = (inp[11]) ? 3'b110 : 3'b101;
						assign node503 = (inp[5]) ? node529 : node504;
							assign node504 = (inp[7]) ? node520 : node505;
								assign node505 = (inp[1]) ? node513 : node506;
									assign node506 = (inp[8]) ? 3'b001 : node507;
										assign node507 = (inp[2]) ? 3'b001 : node508;
											assign node508 = (inp[11]) ? 3'b110 : 3'b010;
									assign node513 = (inp[8]) ? node517 : node514;
										assign node514 = (inp[11]) ? 3'b001 : 3'b101;
										assign node517 = (inp[11]) ? 3'b000 : 3'b100;
								assign node520 = (inp[8]) ? node526 : node521;
									assign node521 = (inp[2]) ? 3'b101 : node522;
										assign node522 = (inp[1]) ? 3'b101 : 3'b001;
									assign node526 = (inp[1]) ? 3'b011 : 3'b001;
							assign node529 = (inp[1]) ? node551 : node530;
								assign node530 = (inp[11]) ? node544 : node531;
									assign node531 = (inp[2]) ? node539 : node532;
										assign node532 = (inp[8]) ? node536 : node533;
											assign node533 = (inp[7]) ? 3'b110 : 3'b010;
											assign node536 = (inp[7]) ? 3'b110 : 3'b101;
										assign node539 = (inp[7]) ? node541 : 3'b110;
											assign node541 = (inp[8]) ? 3'b010 : 3'b110;
									assign node544 = (inp[2]) ? 3'b110 : node545;
										assign node545 = (inp[8]) ? 3'b110 : node546;
											assign node546 = (inp[7]) ? 3'b110 : 3'b010;
								assign node551 = (inp[7]) ? node557 : node552;
									assign node552 = (inp[8]) ? 3'b111 : node553;
										assign node553 = (inp[11]) ? 3'b110 : 3'b111;
									assign node557 = (inp[8]) ? node561 : node558;
										assign node558 = (inp[11]) ? 3'b001 : 3'b101;
										assign node561 = (inp[11]) ? 3'b101 : 3'b111;
					assign node564 = (inp[1]) ? node624 : node565;
						assign node565 = (inp[7]) ? node579 : node566;
							assign node566 = (inp[0]) ? 3'b101 : node567;
								assign node567 = (inp[5]) ? node571 : node568;
									assign node568 = (inp[10]) ? 3'b001 : 3'b101;
									assign node571 = (inp[2]) ? 3'b110 : node572;
										assign node572 = (inp[10]) ? node574 : 3'b110;
											assign node574 = (inp[8]) ? 3'b110 : 3'b010;
							assign node579 = (inp[8]) ? node603 : node580;
								assign node580 = (inp[5]) ? node592 : node581;
									assign node581 = (inp[0]) ? node589 : node582;
										assign node582 = (inp[10]) ? node584 : 3'b001;
											assign node584 = (inp[2]) ? 3'b101 : node585;
												assign node585 = (inp[11]) ? 3'b001 : 3'b101;
										assign node589 = (inp[10]) ? 3'b011 : 3'b001;
									assign node592 = (inp[0]) ? node598 : node593;
										assign node593 = (inp[10]) ? node595 : 3'b010;
											assign node595 = (inp[2]) ? 3'b010 : 3'b110;
										assign node598 = (inp[2]) ? node600 : 3'b101;
											assign node600 = (inp[10]) ? 3'b011 : 3'b001;
								assign node603 = (inp[0]) ? node609 : node604;
									assign node604 = (inp[5]) ? 3'b001 : node605;
										assign node605 = (inp[10]) ? 3'b101 : 3'b001;
									assign node609 = (inp[10]) ? node617 : node610;
										assign node610 = (inp[11]) ? node612 : 3'b101;
											assign node612 = (inp[2]) ? node614 : 3'b001;
												assign node614 = (inp[5]) ? 3'b001 : 3'b101;
										assign node617 = (inp[5]) ? node621 : node618;
											assign node618 = (inp[2]) ? 3'b111 : 3'b011;
											assign node621 = (inp[2]) ? 3'b011 : 3'b101;
						assign node624 = (inp[5]) ? node656 : node625;
							assign node625 = (inp[0]) ? node647 : node626;
								assign node626 = (inp[10]) ? node636 : node627;
									assign node627 = (inp[8]) ? node633 : node628;
										assign node628 = (inp[2]) ? node630 : 3'b011;
											assign node630 = (inp[7]) ? 3'b011 : 3'b001;
										assign node633 = (inp[7]) ? 3'b001 : 3'b011;
									assign node636 = (inp[7]) ? node642 : node637;
										assign node637 = (inp[2]) ? 3'b101 : node638;
											assign node638 = (inp[8]) ? 3'b101 : 3'b001;
										assign node642 = (inp[8]) ? 3'b011 : node643;
											assign node643 = (inp[2]) ? 3'b001 : 3'b011;
								assign node647 = (inp[7]) ? 3'b111 : node648;
									assign node648 = (inp[8]) ? node650 : 3'b011;
										assign node650 = (inp[10]) ? node652 : 3'b011;
											assign node652 = (inp[2]) ? 3'b111 : 3'b011;
							assign node656 = (inp[8]) ? node676 : node657;
								assign node657 = (inp[10]) ? node667 : node658;
									assign node658 = (inp[0]) ? 3'b001 : node659;
										assign node659 = (inp[7]) ? node661 : 3'b001;
											assign node661 = (inp[2]) ? 3'b011 : node662;
												assign node662 = (inp[11]) ? 3'b001 : 3'b011;
									assign node667 = (inp[2]) ? node669 : 3'b001;
										assign node669 = (inp[0]) ? node671 : 3'b101;
											assign node671 = (inp[11]) ? node673 : 3'b001;
												assign node673 = (inp[7]) ? 3'b001 : 3'b101;
								assign node676 = (inp[0]) ? 3'b011 : node677;
									assign node677 = (inp[10]) ? node687 : node678;
										assign node678 = (inp[7]) ? node684 : node679;
											assign node679 = (inp[2]) ? node681 : 3'b001;
												assign node681 = (inp[11]) ? 3'b001 : 3'b011;
											assign node684 = (inp[2]) ? 3'b001 : 3'b011;
										assign node687 = (inp[7]) ? node693 : node688;
											assign node688 = (inp[2]) ? 3'b001 : node689;
												assign node689 = (inp[11]) ? 3'b001 : 3'b101;
											assign node693 = (inp[2]) ? 3'b101 : 3'b001;
				assign node697 = (inp[6]) ? node807 : node698;
					assign node698 = (inp[0]) ? node776 : node699;
						assign node699 = (inp[5]) ? node739 : node700;
							assign node700 = (inp[1]) ? node712 : node701;
								assign node701 = (inp[10]) ? node703 : 3'b100;
									assign node703 = (inp[7]) ? 3'b100 : node704;
										assign node704 = (inp[2]) ? node706 : 3'b000;
											assign node706 = (inp[8]) ? 3'b100 : node707;
												assign node707 = (inp[11]) ? 3'b000 : 3'b100;
								assign node712 = (inp[7]) ? node724 : node713;
									assign node713 = (inp[10]) ? node719 : node714;
										assign node714 = (inp[2]) ? node716 : 3'b010;
											assign node716 = (inp[8]) ? 3'b110 : 3'b100;
										assign node719 = (inp[8]) ? 3'b100 : node720;
											assign node720 = (inp[11]) ? 3'b000 : 3'b100;
									assign node724 = (inp[8]) ? node734 : node725;
										assign node725 = (inp[2]) ? node731 : node726;
											assign node726 = (inp[11]) ? node728 : 3'b010;
												assign node728 = (inp[10]) ? 3'b100 : 3'b110;
											assign node731 = (inp[10]) ? 3'b010 : 3'b000;
										assign node734 = (inp[11]) ? 3'b010 : node735;
											assign node735 = (inp[2]) ? 3'b010 : 3'b000;
							assign node739 = (inp[1]) ? node749 : node740;
								assign node740 = (inp[10]) ? node742 : 3'b000;
									assign node742 = (inp[2]) ? node744 : 3'b000;
										assign node744 = (inp[8]) ? 3'b000 : node745;
											assign node745 = (inp[11]) ? 3'b000 : 3'b100;
								assign node749 = (inp[7]) ? node759 : node750;
									assign node750 = (inp[8]) ? node752 : 3'b000;
										assign node752 = (inp[2]) ? node756 : node753;
											assign node753 = (inp[11]) ? 3'b000 : 3'b100;
											assign node756 = (inp[11]) ? 3'b000 : 3'b010;
									assign node759 = (inp[2]) ? node771 : node760;
										assign node760 = (inp[8]) ? node764 : node761;
											assign node761 = (inp[10]) ? 3'b000 : 3'b010;
											assign node764 = (inp[10]) ? node768 : node765;
												assign node765 = (inp[11]) ? 3'b110 : 3'b100;
												assign node768 = (inp[11]) ? 3'b100 : 3'b110;
										assign node771 = (inp[11]) ? 3'b100 : node772;
											assign node772 = (inp[10]) ? 3'b110 : 3'b100;
						assign node776 = (inp[1]) ? node794 : node777;
							assign node777 = (inp[5]) ? node787 : node778;
								assign node778 = (inp[2]) ? 3'b010 : node779;
									assign node779 = (inp[7]) ? 3'b010 : node780;
										assign node780 = (inp[8]) ? 3'b010 : node781;
											assign node781 = (inp[11]) ? 3'b100 : 3'b000;
								assign node787 = (inp[7]) ? 3'b100 : node788;
									assign node788 = (inp[8]) ? 3'b100 : node789;
										assign node789 = (inp[2]) ? 3'b100 : 3'b000;
							assign node794 = (inp[5]) ? node800 : node795;
								assign node795 = (inp[7]) ? 3'b110 : node796;
									assign node796 = (inp[8]) ? 3'b100 : 3'b010;
								assign node800 = (inp[8]) ? 3'b010 : node801;
									assign node801 = (inp[7]) ? 3'b010 : node802;
										assign node802 = (inp[11]) ? 3'b100 : 3'b010;
					assign node807 = (inp[0]) ? node859 : node808;
						assign node808 = (inp[1]) ? node840 : node809;
							assign node809 = (inp[8]) ? node825 : node810;
								assign node810 = (inp[7]) ? node812 : 3'b100;
									assign node812 = (inp[10]) ? node818 : node813;
										assign node813 = (inp[11]) ? node815 : 3'b000;
											assign node815 = (inp[5]) ? 3'b100 : 3'b000;
										assign node818 = (inp[2]) ? node822 : node819;
											assign node819 = (inp[11]) ? 3'b100 : 3'b000;
											assign node822 = (inp[5]) ? 3'b110 : 3'b010;
								assign node825 = (inp[5]) ? node829 : node826;
									assign node826 = (inp[7]) ? 3'b110 : 3'b010;
									assign node829 = (inp[11]) ? node835 : node830;
										assign node830 = (inp[10]) ? 3'b010 : node831;
											assign node831 = (inp[7]) ? 3'b000 : 3'b010;
										assign node835 = (inp[7]) ? node837 : 3'b100;
											assign node837 = (inp[10]) ? 3'b010 : 3'b000;
							assign node840 = (inp[7]) ? node844 : node841;
								assign node841 = (inp[5]) ? 3'b100 : 3'b110;
								assign node844 = (inp[2]) ? node848 : node845;
									assign node845 = (inp[5]) ? 3'b010 : 3'b110;
									assign node848 = (inp[8]) ? node854 : node849;
										assign node849 = (inp[11]) ? node851 : 3'b110;
											assign node851 = (inp[5]) ? 3'b101 : 3'b110;
										assign node854 = (inp[5]) ? node856 : 3'b001;
											assign node856 = (inp[10]) ? 3'b010 : 3'b110;
						assign node859 = (inp[5]) ? node869 : node860;
							assign node860 = (inp[7]) ? node862 : 3'b001;
								assign node862 = (inp[1]) ? 3'b101 : node863;
									assign node863 = (inp[2]) ? node865 : 3'b001;
										assign node865 = (inp[10]) ? 3'b101 : 3'b001;
							assign node869 = (inp[1]) ? node875 : node870;
								assign node870 = (inp[10]) ? node872 : 3'b010;
									assign node872 = (inp[7]) ? 3'b110 : 3'b010;
								assign node875 = (inp[7]) ? 3'b001 : 3'b110;
		assign node878 = (inp[6]) ? node900 : node879;
			assign node879 = (inp[4]) ? 3'b000 : node880;
				assign node880 = (inp[0]) ? node882 : 3'b000;
					assign node882 = (inp[9]) ? node884 : 3'b000;
						assign node884 = (inp[1]) ? node886 : 3'b000;
							assign node886 = (inp[5]) ? node892 : node887;
								assign node887 = (inp[7]) ? 3'b100 : node888;
									assign node888 = (inp[8]) ? 3'b100 : 3'b000;
								assign node892 = (inp[11]) ? 3'b000 : node893;
									assign node893 = (inp[7]) ? 3'b000 : node894;
										assign node894 = (inp[8]) ? 3'b100 : 3'b000;
			assign node900 = (inp[9]) ? node1076 : node901;
				assign node901 = (inp[4]) ? node925 : node902;
					assign node902 = (inp[0]) ? node918 : node903;
						assign node903 = (inp[2]) ? node905 : 3'b010;
							assign node905 = (inp[1]) ? node907 : 3'b010;
								assign node907 = (inp[7]) ? node909 : 3'b010;
									assign node909 = (inp[5]) ? node913 : node910;
										assign node910 = (inp[8]) ? 3'b011 : 3'b010;
										assign node913 = (inp[8]) ? 3'b010 : node914;
											assign node914 = (inp[11]) ? 3'b011 : 3'b010;
						assign node918 = (inp[5]) ? node920 : 3'b011;
							assign node920 = (inp[7]) ? node922 : 3'b010;
								assign node922 = (inp[1]) ? 3'b011 : 3'b010;
					assign node925 = (inp[0]) ? node991 : node926;
						assign node926 = (inp[10]) ? node970 : node927;
							assign node927 = (inp[7]) ? node941 : node928;
								assign node928 = (inp[1]) ? node936 : node929;
									assign node929 = (inp[8]) ? node931 : 3'b000;
										assign node931 = (inp[5]) ? node933 : 3'b010;
											assign node933 = (inp[11]) ? 3'b000 : 3'b010;
									assign node936 = (inp[5]) ? node938 : 3'b000;
										assign node938 = (inp[11]) ? 3'b100 : 3'b000;
								assign node941 = (inp[1]) ? node953 : node942;
									assign node942 = (inp[5]) ? node948 : node943;
										assign node943 = (inp[8]) ? 3'b010 : node944;
											assign node944 = (inp[2]) ? 3'b100 : 3'b110;
										assign node948 = (inp[11]) ? 3'b100 : node949;
											assign node949 = (inp[8]) ? 3'b000 : 3'b100;
									assign node953 = (inp[11]) ? node961 : node954;
										assign node954 = (inp[2]) ? node956 : 3'b010;
											assign node956 = (inp[5]) ? 3'b010 : node957;
												assign node957 = (inp[8]) ? 3'b100 : 3'b010;
										assign node961 = (inp[5]) ? node967 : node962;
											assign node962 = (inp[8]) ? node964 : 3'b010;
												assign node964 = (inp[2]) ? 3'b100 : 3'b010;
											assign node967 = (inp[2]) ? 3'b010 : 3'b100;
							assign node970 = (inp[1]) ? node972 : 3'b000;
								assign node972 = (inp[5]) ? node982 : node973;
									assign node973 = (inp[8]) ? 3'b000 : node974;
										assign node974 = (inp[2]) ? 3'b000 : node975;
											assign node975 = (inp[7]) ? node977 : 3'b000;
												assign node977 = (inp[11]) ? 3'b100 : 3'b000;
									assign node982 = (inp[11]) ? node986 : node983;
										assign node983 = (inp[7]) ? 3'b100 : 3'b000;
										assign node986 = (inp[7]) ? node988 : 3'b100;
											assign node988 = (inp[8]) ? 3'b100 : 3'b000;
						assign node991 = (inp[7]) ? node1023 : node992;
							assign node992 = (inp[10]) ? node1014 : node993;
								assign node993 = (inp[1]) ? node1007 : node994;
									assign node994 = (inp[5]) ? node1000 : node995;
										assign node995 = (inp[8]) ? 3'b010 : node996;
											assign node996 = (inp[2]) ? 3'b100 : 3'b010;
										assign node1000 = (inp[2]) ? node1002 : 3'b100;
											assign node1002 = (inp[11]) ? 3'b100 : node1003;
												assign node1003 = (inp[8]) ? 3'b010 : 3'b100;
									assign node1007 = (inp[2]) ? node1009 : 3'b010;
										assign node1009 = (inp[11]) ? node1011 : 3'b110;
											assign node1011 = (inp[5]) ? 3'b010 : 3'b110;
								assign node1014 = (inp[8]) ? node1016 : 3'b100;
									assign node1016 = (inp[1]) ? node1018 : 3'b100;
										assign node1018 = (inp[5]) ? node1020 : 3'b010;
											assign node1020 = (inp[11]) ? 3'b100 : 3'b010;
							assign node1023 = (inp[10]) ? node1055 : node1024;
								assign node1024 = (inp[1]) ? node1040 : node1025;
									assign node1025 = (inp[11]) ? node1031 : node1026;
										assign node1026 = (inp[2]) ? 3'b110 : node1027;
											assign node1027 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1031 = (inp[2]) ? node1033 : 3'b010;
											assign node1033 = (inp[8]) ? node1037 : node1034;
												assign node1034 = (inp[5]) ? 3'b010 : 3'b110;
												assign node1037 = (inp[5]) ? 3'b110 : 3'b010;
									assign node1040 = (inp[5]) ? node1048 : node1041;
										assign node1041 = (inp[8]) ? node1045 : node1042;
											assign node1042 = (inp[2]) ? 3'b110 : 3'b101;
											assign node1045 = (inp[2]) ? 3'b101 : 3'b001;
										assign node1048 = (inp[11]) ? node1052 : node1049;
											assign node1049 = (inp[2]) ? 3'b001 : 3'b110;
											assign node1052 = (inp[2]) ? 3'b110 : 3'b010;
								assign node1055 = (inp[1]) ? node1065 : node1056;
									assign node1056 = (inp[11]) ? node1058 : 3'b010;
										assign node1058 = (inp[5]) ? 3'b100 : node1059;
											assign node1059 = (inp[8]) ? 3'b010 : node1060;
												assign node1060 = (inp[2]) ? 3'b010 : 3'b100;
									assign node1065 = (inp[5]) ? node1071 : node1066;
										assign node1066 = (inp[8]) ? 3'b110 : node1067;
											assign node1067 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1071 = (inp[11]) ? 3'b010 : node1072;
											assign node1072 = (inp[2]) ? 3'b110 : 3'b010;
				assign node1076 = (inp[0]) ? node1114 : node1077;
					assign node1077 = (inp[4]) ? 3'b000 : node1078;
						assign node1078 = (inp[10]) ? node1094 : node1079;
							assign node1079 = (inp[1]) ? node1081 : 3'b000;
								assign node1081 = (inp[7]) ? node1083 : 3'b000;
									assign node1083 = (inp[2]) ? node1085 : 3'b000;
										assign node1085 = (inp[5]) ? node1089 : node1086;
											assign node1086 = (inp[8]) ? 3'b010 : 3'b000;
											assign node1089 = (inp[11]) ? node1091 : 3'b000;
												assign node1091 = (inp[8]) ? 3'b000 : 3'b010;
							assign node1094 = (inp[1]) ? node1102 : node1095;
								assign node1095 = (inp[8]) ? node1097 : 3'b000;
									assign node1097 = (inp[5]) ? 3'b000 : node1098;
										assign node1098 = (inp[7]) ? 3'b100 : 3'b000;
								assign node1102 = (inp[2]) ? node1108 : node1103;
									assign node1103 = (inp[7]) ? node1105 : 3'b000;
										assign node1105 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1108 = (inp[7]) ? node1110 : 3'b100;
										assign node1110 = (inp[8]) ? 3'b010 : 3'b100;
					assign node1114 = (inp[4]) ? node1126 : node1115;
						assign node1115 = (inp[5]) ? node1121 : node1116;
							assign node1116 = (inp[1]) ? node1118 : 3'b010;
								assign node1118 = (inp[7]) ? 3'b110 : 3'b010;
							assign node1121 = (inp[1]) ? node1123 : 3'b100;
								assign node1123 = (inp[7]) ? 3'b010 : 3'b100;
						assign node1126 = (inp[1]) ? node1136 : node1127;
							assign node1127 = (inp[10]) ? 3'b000 : node1128;
								assign node1128 = (inp[11]) ? 3'b000 : node1129;
									assign node1129 = (inp[7]) ? node1131 : 3'b000;
										assign node1131 = (inp[8]) ? 3'b100 : 3'b000;
							assign node1136 = (inp[7]) ? node1142 : node1137;
								assign node1137 = (inp[10]) ? 3'b000 : node1138;
									assign node1138 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1142 = (inp[10]) ? node1160 : node1143;
									assign node1143 = (inp[5]) ? node1149 : node1144;
										assign node1144 = (inp[8]) ? 3'b010 : node1145;
											assign node1145 = (inp[2]) ? 3'b100 : 3'b110;
										assign node1149 = (inp[11]) ? node1155 : node1150;
											assign node1150 = (inp[8]) ? node1152 : 3'b100;
												assign node1152 = (inp[2]) ? 3'b010 : 3'b100;
											assign node1155 = (inp[2]) ? 3'b100 : node1156;
												assign node1156 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1160 = (inp[5]) ? node1166 : node1161;
										assign node1161 = (inp[8]) ? 3'b100 : node1162;
											assign node1162 = (inp[11]) ? 3'b100 : 3'b000;
										assign node1166 = (inp[2]) ? 3'b100 : 3'b000;

endmodule