module dtc_split05_bm47 (
	input  wire [16-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node6;
	wire [1-1:0] node7;
	wire [1-1:0] node8;
	wire [1-1:0] node9;
	wire [1-1:0] node13;
	wire [1-1:0] node15;
	wire [1-1:0] node17;
	wire [1-1:0] node21;
	wire [1-1:0] node22;
	wire [1-1:0] node23;
	wire [1-1:0] node24;
	wire [1-1:0] node25;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node32;
	wire [1-1:0] node33;
	wire [1-1:0] node37;
	wire [1-1:0] node39;
	wire [1-1:0] node40;
	wire [1-1:0] node42;
	wire [1-1:0] node46;
	wire [1-1:0] node47;
	wire [1-1:0] node48;
	wire [1-1:0] node52;
	wire [1-1:0] node54;
	wire [1-1:0] node56;
	wire [1-1:0] node59;
	wire [1-1:0] node61;
	wire [1-1:0] node62;
	wire [1-1:0] node63;
	wire [1-1:0] node64;
	wire [1-1:0] node65;
	wire [1-1:0] node68;
	wire [1-1:0] node69;
	wire [1-1:0] node73;
	wire [1-1:0] node78;
	wire [1-1:0] node79;
	wire [1-1:0] node80;
	wire [1-1:0] node81;
	wire [1-1:0] node82;
	wire [1-1:0] node84;
	wire [1-1:0] node85;
	wire [1-1:0] node87;
	wire [1-1:0] node90;
	wire [1-1:0] node91;
	wire [1-1:0] node95;
	wire [1-1:0] node96;
	wire [1-1:0] node98;
	wire [1-1:0] node101;
	wire [1-1:0] node102;
	wire [1-1:0] node103;
	wire [1-1:0] node104;
	wire [1-1:0] node106;
	wire [1-1:0] node109;
	wire [1-1:0] node110;
	wire [1-1:0] node115;
	wire [1-1:0] node117;
	wire [1-1:0] node120;
	wire [1-1:0] node121;
	wire [1-1:0] node122;
	wire [1-1:0] node123;
	wire [1-1:0] node125;
	wire [1-1:0] node126;
	wire [1-1:0] node127;
	wire [1-1:0] node132;
	wire [1-1:0] node133;
	wire [1-1:0] node135;
	wire [1-1:0] node138;
	wire [1-1:0] node140;
	wire [1-1:0] node143;
	wire [1-1:0] node145;
	wire [1-1:0] node148;
	wire [1-1:0] node149;
	wire [1-1:0] node150;
	wire [1-1:0] node152;
	wire [1-1:0] node154;
	wire [1-1:0] node156;
	wire [1-1:0] node159;
	wire [1-1:0] node161;
	wire [1-1:0] node163;
	wire [1-1:0] node166;
	wire [1-1:0] node167;
	wire [1-1:0] node168;
	wire [1-1:0] node172;
	wire [1-1:0] node174;
	wire [1-1:0] node177;
	wire [1-1:0] node178;
	wire [1-1:0] node179;
	wire [1-1:0] node180;
	wire [1-1:0] node182;
	wire [1-1:0] node186;
	wire [1-1:0] node187;
	wire [1-1:0] node188;
	wire [1-1:0] node189;
	wire [1-1:0] node191;
	wire [1-1:0] node193;
	wire [1-1:0] node199;
	wire [1-1:0] node200;
	wire [1-1:0] node201;
	wire [1-1:0] node202;
	wire [1-1:0] node206;
	wire [1-1:0] node207;
	wire [1-1:0] node209;
	wire [1-1:0] node212;
	wire [1-1:0] node214;
	wire [1-1:0] node216;
	wire [1-1:0] node219;
	wire [1-1:0] node221;
	wire [1-1:0] node224;
	wire [1-1:0] node225;
	wire [1-1:0] node227;
	wire [1-1:0] node228;
	wire [1-1:0] node229;
	wire [1-1:0] node230;
	wire [1-1:0] node232;
	wire [1-1:0] node233;
	wire [1-1:0] node237;
	wire [1-1:0] node239;
	wire [1-1:0] node242;
	wire [1-1:0] node243;
	wire [1-1:0] node245;
	wire [1-1:0] node250;
	wire [1-1:0] node251;
	wire [1-1:0] node252;
	wire [1-1:0] node253;
	wire [1-1:0] node254;
	wire [1-1:0] node256;
	wire [1-1:0] node257;
	wire [1-1:0] node263;
	wire [1-1:0] node264;
	wire [1-1:0] node265;
	wire [1-1:0] node269;
	wire [1-1:0] node270;
	wire [1-1:0] node272;
	wire [1-1:0] node275;
	wire [1-1:0] node276;
	wire [1-1:0] node280;
	wire [1-1:0] node281;
	wire [1-1:0] node283;
	wire [1-1:0] node285;
	wire [1-1:0] node286;
	wire [1-1:0] node288;
	wire [1-1:0] node290;
	wire [1-1:0] node295;
	wire [1-1:0] node296;
	wire [1-1:0] node297;
	wire [1-1:0] node298;
	wire [1-1:0] node299;
	wire [1-1:0] node300;
	wire [1-1:0] node301;
	wire [1-1:0] node303;
	wire [1-1:0] node304;
	wire [1-1:0] node308;
	wire [1-1:0] node309;
	wire [1-1:0] node310;
	wire [1-1:0] node314;
	wire [1-1:0] node316;
	wire [1-1:0] node319;
	wire [1-1:0] node321;
	wire [1-1:0] node322;
	wire [1-1:0] node326;
	wire [1-1:0] node327;
	wire [1-1:0] node329;
	wire [1-1:0] node330;
	wire [1-1:0] node331;
	wire [1-1:0] node333;
	wire [1-1:0] node337;
	wire [1-1:0] node338;
	wire [1-1:0] node340;
	wire [1-1:0] node341;
	wire [1-1:0] node346;
	wire [1-1:0] node347;
	wire [1-1:0] node348;
	wire [1-1:0] node350;
	wire [1-1:0] node351;
	wire [1-1:0] node355;
	wire [1-1:0] node356;
	wire [1-1:0] node360;
	wire [1-1:0] node362;
	wire [1-1:0] node365;
	wire [1-1:0] node366;
	wire [1-1:0] node367;
	wire [1-1:0] node368;
	wire [1-1:0] node370;
	wire [1-1:0] node371;
	wire [1-1:0] node375;
	wire [1-1:0] node376;
	wire [1-1:0] node377;
	wire [1-1:0] node381;
	wire [1-1:0] node382;
	wire [1-1:0] node386;
	wire [1-1:0] node387;
	wire [1-1:0] node389;
	wire [1-1:0] node390;
	wire [1-1:0] node395;
	wire [1-1:0] node396;
	wire [1-1:0] node397;
	wire [1-1:0] node398;
	wire [1-1:0] node400;
	wire [1-1:0] node401;
	wire [1-1:0] node406;
	wire [1-1:0] node407;
	wire [1-1:0] node408;
	wire [1-1:0] node409;
	wire [1-1:0] node412;
	wire [1-1:0] node417;
	wire [1-1:0] node418;
	wire [1-1:0] node420;
	wire [1-1:0] node424;
	wire [1-1:0] node425;
	wire [1-1:0] node426;
	wire [1-1:0] node427;
	wire [1-1:0] node428;
	wire [1-1:0] node430;
	wire [1-1:0] node431;
	wire [1-1:0] node432;
	wire [1-1:0] node437;
	wire [1-1:0] node439;
	wire [1-1:0] node440;
	wire [1-1:0] node444;
	wire [1-1:0] node445;
	wire [1-1:0] node446;
	wire [1-1:0] node448;
	wire [1-1:0] node452;
	wire [1-1:0] node453;
	wire [1-1:0] node454;
	wire [1-1:0] node458;
	wire [1-1:0] node460;
	wire [1-1:0] node463;
	wire [1-1:0] node464;
	wire [1-1:0] node465;
	wire [1-1:0] node467;
	wire [1-1:0] node468;
	wire [1-1:0] node469;
	wire [1-1:0] node472;
	wire [1-1:0] node476;
	wire [1-1:0] node477;
	wire [1-1:0] node479;
	wire [1-1:0] node481;
	wire [1-1:0] node483;
	wire [1-1:0] node487;
	wire [1-1:0] node489;
	wire [1-1:0] node490;
	wire [1-1:0] node491;
	wire [1-1:0] node495;
	wire [1-1:0] node498;
	wire [1-1:0] node499;
	wire [1-1:0] node500;
	wire [1-1:0] node502;
	wire [1-1:0] node503;
	wire [1-1:0] node507;
	wire [1-1:0] node508;
	wire [1-1:0] node510;
	wire [1-1:0] node512;
	wire [1-1:0] node514;
	wire [1-1:0] node517;
	wire [1-1:0] node519;
	wire [1-1:0] node522;
	wire [1-1:0] node524;
	wire [1-1:0] node526;
	wire [1-1:0] node527;
	wire [1-1:0] node528;
	wire [1-1:0] node529;
	wire [1-1:0] node531;
	wire [1-1:0] node535;
	wire [1-1:0] node537;
	wire [1-1:0] node541;
	wire [1-1:0] node542;
	wire [1-1:0] node543;
	wire [1-1:0] node544;
	wire [1-1:0] node545;
	wire [1-1:0] node546;
	wire [1-1:0] node547;
	wire [1-1:0] node548;
	wire [1-1:0] node552;
	wire [1-1:0] node553;
	wire [1-1:0] node554;
	wire [1-1:0] node555;
	wire [1-1:0] node561;
	wire [1-1:0] node562;
	wire [1-1:0] node563;
	wire [1-1:0] node566;
	wire [1-1:0] node567;
	wire [1-1:0] node570;
	wire [1-1:0] node574;
	wire [1-1:0] node575;
	wire [1-1:0] node577;
	wire [1-1:0] node579;
	wire [1-1:0] node581;
	wire [1-1:0] node584;
	wire [1-1:0] node585;
	wire [1-1:0] node586;
	wire [1-1:0] node591;
	wire [1-1:0] node592;
	wire [1-1:0] node593;
	wire [1-1:0] node594;
	wire [1-1:0] node596;
	wire [1-1:0] node600;
	wire [1-1:0] node603;
	wire [1-1:0] node604;
	wire [1-1:0] node606;
	wire [1-1:0] node610;
	wire [1-1:0] node611;
	wire [1-1:0] node613;
	wire [1-1:0] node614;
	wire [1-1:0] node615;
	wire [1-1:0] node616;
	wire [1-1:0] node618;
	wire [1-1:0] node624;
	wire [1-1:0] node625;
	wire [1-1:0] node626;
	wire [1-1:0] node627;
	wire [1-1:0] node628;
	wire [1-1:0] node633;
	wire [1-1:0] node635;
	wire [1-1:0] node638;
	wire [1-1:0] node639;
	wire [1-1:0] node641;
	wire [1-1:0] node642;
	wire [1-1:0] node643;
	wire [1-1:0] node644;
	wire [1-1:0] node645;
	wire [1-1:0] node653;
	wire [1-1:0] node654;
	wire [1-1:0] node655;
	wire [1-1:0] node656;
	wire [1-1:0] node657;
	wire [1-1:0] node659;
	wire [1-1:0] node660;
	wire [1-1:0] node661;
	wire [1-1:0] node666;
	wire [1-1:0] node667;
	wire [1-1:0] node669;
	wire [1-1:0] node673;
	wire [1-1:0] node675;
	wire [1-1:0] node677;
	wire [1-1:0] node680;
	wire [1-1:0] node681;
	wire [1-1:0] node682;
	wire [1-1:0] node683;
	wire [1-1:0] node687;
	wire [1-1:0] node688;
	wire [1-1:0] node691;
	wire [1-1:0] node693;
	wire [1-1:0] node696;
	wire [1-1:0] node698;
	wire [1-1:0] node699;
	wire [1-1:0] node700;
	wire [1-1:0] node705;
	wire [1-1:0] node706;
	wire [1-1:0] node707;
	wire [1-1:0] node709;
	wire [1-1:0] node710;
	wire [1-1:0] node712;
	wire [1-1:0] node716;
	wire [1-1:0] node717;
	wire [1-1:0] node719;
	wire [1-1:0] node723;
	wire [1-1:0] node725;
	wire [1-1:0] node726;
	wire [1-1:0] node727;
	wire [1-1:0] node728;
	wire [1-1:0] node734;
	wire [1-1:0] node735;
	wire [1-1:0] node736;
	wire [1-1:0] node737;
	wire [1-1:0] node739;
	wire [1-1:0] node740;
	wire [1-1:0] node741;
	wire [1-1:0] node742;
	wire [1-1:0] node746;
	wire [1-1:0] node747;
	wire [1-1:0] node748;
	wire [1-1:0] node752;
	wire [1-1:0] node753;
	wire [1-1:0] node758;
	wire [1-1:0] node759;
	wire [1-1:0] node760;
	wire [1-1:0] node761;
	wire [1-1:0] node762;
	wire [1-1:0] node764;
	wire [1-1:0] node765;
	wire [1-1:0] node767;
	wire [1-1:0] node772;
	wire [1-1:0] node774;
	wire [1-1:0] node777;
	wire [1-1:0] node778;
	wire [1-1:0] node779;
	wire [1-1:0] node780;
	wire [1-1:0] node782;
	wire [1-1:0] node783;
	wire [1-1:0] node789;
	wire [1-1:0] node790;
	wire [1-1:0] node791;
	wire [1-1:0] node795;
	wire [1-1:0] node797;
	wire [1-1:0] node800;
	wire [1-1:0] node801;
	wire [1-1:0] node803;
	wire [1-1:0] node804;
	wire [1-1:0] node805;
	wire [1-1:0] node806;
	wire [1-1:0] node808;
	wire [1-1:0] node811;
	wire [1-1:0] node812;
	wire [1-1:0] node816;
	wire [1-1:0] node819;
	wire [1-1:0] node820;
	wire [1-1:0] node821;
	wire [1-1:0] node827;
	wire [1-1:0] node828;
	wire [1-1:0] node829;
	wire [1-1:0] node830;
	wire [1-1:0] node831;
	wire [1-1:0] node832;
	wire [1-1:0] node833;
	wire [1-1:0] node837;
	wire [1-1:0] node839;
	wire [1-1:0] node841;
	wire [1-1:0] node843;
	wire [1-1:0] node846;
	wire [1-1:0] node848;
	wire [1-1:0] node849;
	wire [1-1:0] node850;
	wire [1-1:0] node854;
	wire [1-1:0] node857;
	wire [1-1:0] node858;
	wire [1-1:0] node859;
	wire [1-1:0] node860;
	wire [1-1:0] node861;
	wire [1-1:0] node862;
	wire [1-1:0] node863;
	wire [1-1:0] node870;
	wire [1-1:0] node871;
	wire [1-1:0] node873;
	wire [1-1:0] node877;
	wire [1-1:0] node878;
	wire [1-1:0] node879;
	wire [1-1:0] node880;
	wire [1-1:0] node884;
	wire [1-1:0] node885;
	wire [1-1:0] node890;
	wire [1-1:0] node891;
	wire [1-1:0] node892;
	wire [1-1:0] node893;
	wire [1-1:0] node894;
	wire [1-1:0] node896;
	wire [1-1:0] node898;
	wire [1-1:0] node901;
	wire [1-1:0] node904;
	wire [1-1:0] node906;
	wire [1-1:0] node909;
	wire [1-1:0] node910;
	wire [1-1:0] node911;
	wire [1-1:0] node912;
	wire [1-1:0] node914;
	wire [1-1:0] node920;
	wire [1-1:0] node921;
	wire [1-1:0] node923;
	wire [1-1:0] node924;
	wire [1-1:0] node925;
	wire [1-1:0] node930;
	wire [1-1:0] node931;
	wire [1-1:0] node932;
	wire [1-1:0] node934;
	wire [1-1:0] node935;
	wire [1-1:0] node939;
	wire [1-1:0] node941;
	wire [1-1:0] node944;
	wire [1-1:0] node946;
	wire [1-1:0] node949;
	wire [1-1:0] node950;
	wire [1-1:0] node951;
	wire [1-1:0] node953;
	wire [1-1:0] node954;
	wire [1-1:0] node956;
	wire [1-1:0] node958;
	wire [1-1:0] node960;
	wire [1-1:0] node964;
	wire [1-1:0] node965;
	wire [1-1:0] node966;
	wire [1-1:0] node968;
	wire [1-1:0] node971;
	wire [1-1:0] node973;
	wire [1-1:0] node975;
	wire [1-1:0] node978;
	wire [1-1:0] node979;
	wire [1-1:0] node980;
	wire [1-1:0] node981;
	wire [1-1:0] node986;
	wire [1-1:0] node988;
	wire [1-1:0] node989;
	wire [1-1:0] node991;
	wire [1-1:0] node992;
	wire [1-1:0] node997;
	wire [1-1:0] node998;
	wire [1-1:0] node999;
	wire [1-1:0] node1000;
	wire [1-1:0] node1002;
	wire [1-1:0] node1003;
	wire [1-1:0] node1008;
	wire [1-1:0] node1009;
	wire [1-1:0] node1011;
	wire [1-1:0] node1014;
	wire [1-1:0] node1016;
	wire [1-1:0] node1018;
	wire [1-1:0] node1021;
	wire [1-1:0] node1022;
	wire [1-1:0] node1024;
	wire [1-1:0] node1026;
	wire [1-1:0] node1027;
	wire [1-1:0] node1031;
	wire [1-1:0] node1032;
	wire [1-1:0] node1033;
	wire [1-1:0] node1035;
	wire [1-1:0] node1039;
	wire [1-1:0] node1040;
	wire [1-1:0] node1044;
	wire [1-1:0] node1045;
	wire [1-1:0] node1046;
	wire [1-1:0] node1048;
	wire [1-1:0] node1049;
	wire [1-1:0] node1050;
	wire [1-1:0] node1052;
	wire [1-1:0] node1055;
	wire [1-1:0] node1056;
	wire [1-1:0] node1060;
	wire [1-1:0] node1062;
	wire [1-1:0] node1066;
	wire [1-1:0] node1067;
	wire [1-1:0] node1068;
	wire [1-1:0] node1069;
	wire [1-1:0] node1070;
	wire [1-1:0] node1072;
	wire [1-1:0] node1075;
	wire [1-1:0] node1076;
	wire [1-1:0] node1077;
	wire [1-1:0] node1081;
	wire [1-1:0] node1083;
	wire [1-1:0] node1087;
	wire [1-1:0] node1088;
	wire [1-1:0] node1089;
	wire [1-1:0] node1091;
	wire [1-1:0] node1094;
	wire [1-1:0] node1096;
	wire [1-1:0] node1099;
	wire [1-1:0] node1100;
	wire [1-1:0] node1104;
	wire [1-1:0] node1105;
	wire [1-1:0] node1107;
	wire [1-1:0] node1108;
	wire [1-1:0] node1109;
	wire [1-1:0] node1111;
	wire [1-1:0] node1114;
	wire [1-1:0] node1115;
	wire [1-1:0] node1119;
	wire [1-1:0] node1120;

	assign outp = (inp[8]) ? node734 : node1;
		assign node1 = (inp[1]) ? node295 : node2;
			assign node2 = (inp[0]) ? node78 : node3;
				assign node3 = (inp[6]) ? node21 : node4;
					assign node4 = (inp[12]) ? node6 : 1'b1;
						assign node6 = (inp[15]) ? 1'b1 : node7;
							assign node7 = (inp[9]) ? node13 : node8;
								assign node8 = (inp[7]) ? 1'b0 : node9;
									assign node9 = (inp[3]) ? 1'b1 : 1'b0;
								assign node13 = (inp[10]) ? node15 : 1'b1;
									assign node15 = (inp[3]) ? node17 : 1'b0;
										assign node17 = (inp[14]) ? 1'b1 : 1'b0;
					assign node21 = (inp[5]) ? node59 : node22;
						assign node22 = (inp[7]) ? node46 : node23;
							assign node23 = (inp[3]) ? node37 : node24;
								assign node24 = (inp[15]) ? node32 : node25;
									assign node25 = (inp[12]) ? 1'b1 : node26;
										assign node26 = (inp[10]) ? 1'b0 : node27;
											assign node27 = (inp[9]) ? 1'b1 : 1'b0;
									assign node32 = (inp[10]) ? 1'b0 : node33;
										assign node33 = (inp[9]) ? 1'b1 : 1'b0;
								assign node37 = (inp[9]) ? node39 : 1'b1;
									assign node39 = (inp[10]) ? 1'b1 : node40;
										assign node40 = (inp[14]) ? node42 : 1'b0;
											assign node42 = (inp[4]) ? 1'b1 : 1'b0;
							assign node46 = (inp[9]) ? node52 : node47;
								assign node47 = (inp[15]) ? 1'b0 : node48;
									assign node48 = (inp[12]) ? 1'b1 : 1'b0;
								assign node52 = (inp[10]) ? node54 : 1'b1;
									assign node54 = (inp[12]) ? node56 : 1'b0;
										assign node56 = (inp[15]) ? 1'b0 : 1'b1;
						assign node59 = (inp[12]) ? node61 : 1'b1;
							assign node61 = (inp[15]) ? 1'b1 : node62;
								assign node62 = (inp[13]) ? 1'b0 : node63;
									assign node63 = (inp[2]) ? node73 : node64;
										assign node64 = (inp[7]) ? node68 : node65;
											assign node65 = (inp[9]) ? 1'b0 : 1'b1;
											assign node68 = (inp[4]) ? 1'b0 : node69;
												assign node69 = (inp[10]) ? 1'b0 : 1'b1;
										assign node73 = (inp[9]) ? 1'b1 : 1'b0;
				assign node78 = (inp[4]) ? node224 : node79;
					assign node79 = (inp[5]) ? node177 : node80;
						assign node80 = (inp[14]) ? node120 : node81;
							assign node81 = (inp[6]) ? node95 : node82;
								assign node82 = (inp[13]) ? node84 : 1'b0;
									assign node84 = (inp[3]) ? node90 : node85;
										assign node85 = (inp[7]) ? node87 : 1'b0;
											assign node87 = (inp[12]) ? 1'b0 : 1'b1;
										assign node90 = (inp[2]) ? 1'b1 : node91;
											assign node91 = (inp[12]) ? 1'b1 : 1'b0;
								assign node95 = (inp[7]) ? node101 : node96;
									assign node96 = (inp[10]) ? node98 : 1'b1;
										assign node98 = (inp[15]) ? 1'b0 : 1'b1;
									assign node101 = (inp[3]) ? node115 : node102;
										assign node102 = (inp[12]) ? 1'b1 : node103;
											assign node103 = (inp[2]) ? node109 : node104;
												assign node104 = (inp[9]) ? node106 : 1'b1;
													assign node106 = (inp[15]) ? 1'b1 : 1'b0;
												assign node109 = (inp[15]) ? 1'b0 : node110;
													assign node110 = (inp[11]) ? 1'b0 : 1'b1;
										assign node115 = (inp[15]) ? node117 : 1'b0;
											assign node117 = (inp[10]) ? 1'b0 : 1'b1;
							assign node120 = (inp[6]) ? node148 : node121;
								assign node121 = (inp[11]) ? node143 : node122;
									assign node122 = (inp[9]) ? node132 : node123;
										assign node123 = (inp[3]) ? node125 : 1'b1;
											assign node125 = (inp[12]) ? 1'b0 : node126;
												assign node126 = (inp[13]) ? 1'b1 : node127;
													assign node127 = (inp[2]) ? 1'b0 : 1'b1;
										assign node132 = (inp[7]) ? node138 : node133;
											assign node133 = (inp[13]) ? node135 : 1'b1;
												assign node135 = (inp[12]) ? 1'b0 : 1'b1;
											assign node138 = (inp[2]) ? node140 : 1'b0;
												assign node140 = (inp[10]) ? 1'b1 : 1'b0;
									assign node143 = (inp[2]) ? node145 : 1'b1;
										assign node145 = (inp[12]) ? 1'b1 : 1'b0;
								assign node148 = (inp[10]) ? node166 : node149;
									assign node149 = (inp[13]) ? node159 : node150;
										assign node150 = (inp[2]) ? node152 : 1'b1;
											assign node152 = (inp[3]) ? node154 : 1'b0;
												assign node154 = (inp[15]) ? node156 : 1'b1;
													assign node156 = (inp[12]) ? 1'b1 : 1'b0;
										assign node159 = (inp[2]) ? node161 : 1'b0;
											assign node161 = (inp[3]) ? node163 : 1'b0;
												assign node163 = (inp[11]) ? 1'b1 : 1'b0;
									assign node166 = (inp[7]) ? node172 : node167;
										assign node167 = (inp[2]) ? 1'b0 : node168;
											assign node168 = (inp[12]) ? 1'b1 : 1'b0;
										assign node172 = (inp[12]) ? node174 : 1'b1;
											assign node174 = (inp[15]) ? 1'b1 : 1'b0;
						assign node177 = (inp[2]) ? node199 : node178;
							assign node178 = (inp[14]) ? node186 : node179;
								assign node179 = (inp[11]) ? 1'b0 : node180;
									assign node180 = (inp[7]) ? node182 : 1'b1;
										assign node182 = (inp[3]) ? 1'b0 : 1'b1;
								assign node186 = (inp[11]) ? 1'b1 : node187;
									assign node187 = (inp[13]) ? 1'b0 : node188;
										assign node188 = (inp[9]) ? 1'b1 : node189;
											assign node189 = (inp[10]) ? node191 : 1'b0;
												assign node191 = (inp[7]) ? node193 : 1'b1;
													assign node193 = (inp[12]) ? 1'b0 : 1'b1;
							assign node199 = (inp[15]) ? node219 : node200;
								assign node200 = (inp[12]) ? node206 : node201;
									assign node201 = (inp[11]) ? 1'b0 : node202;
										assign node202 = (inp[13]) ? 1'b1 : 1'b0;
									assign node206 = (inp[11]) ? node212 : node207;
										assign node207 = (inp[7]) ? node209 : 1'b0;
											assign node209 = (inp[9]) ? 1'b0 : 1'b1;
										assign node212 = (inp[3]) ? node214 : 1'b1;
											assign node214 = (inp[7]) ? node216 : 1'b0;
												assign node216 = (inp[10]) ? 1'b1 : 1'b0;
								assign node219 = (inp[13]) ? node221 : 1'b0;
									assign node221 = (inp[11]) ? 1'b0 : 1'b1;
					assign node224 = (inp[6]) ? node250 : node225;
						assign node225 = (inp[12]) ? node227 : 1'b1;
							assign node227 = (inp[15]) ? 1'b1 : node228;
								assign node228 = (inp[10]) ? node242 : node229;
									assign node229 = (inp[2]) ? node237 : node230;
										assign node230 = (inp[14]) ? node232 : 1'b1;
											assign node232 = (inp[9]) ? 1'b1 : node233;
												assign node233 = (inp[13]) ? 1'b1 : 1'b0;
										assign node237 = (inp[9]) ? node239 : 1'b0;
											assign node239 = (inp[3]) ? 1'b0 : 1'b1;
									assign node242 = (inp[9]) ? 1'b0 : node243;
										assign node243 = (inp[5]) ? node245 : 1'b0;
											assign node245 = (inp[7]) ? 1'b0 : 1'b1;
						assign node250 = (inp[5]) ? node280 : node251;
							assign node251 = (inp[15]) ? node263 : node252;
								assign node252 = (inp[12]) ? 1'b1 : node253;
									assign node253 = (inp[10]) ? 1'b0 : node254;
										assign node254 = (inp[9]) ? node256 : 1'b0;
											assign node256 = (inp[7]) ? 1'b1 : node257;
												assign node257 = (inp[14]) ? 1'b1 : 1'b0;
								assign node263 = (inp[3]) ? node269 : node264;
									assign node264 = (inp[10]) ? 1'b0 : node265;
										assign node265 = (inp[9]) ? 1'b1 : 1'b0;
									assign node269 = (inp[7]) ? node275 : node270;
										assign node270 = (inp[9]) ? node272 : 1'b1;
											assign node272 = (inp[10]) ? 1'b1 : 1'b0;
										assign node275 = (inp[10]) ? 1'b0 : node276;
											assign node276 = (inp[9]) ? 1'b1 : 1'b0;
							assign node280 = (inp[15]) ? 1'b1 : node281;
								assign node281 = (inp[12]) ? node283 : 1'b1;
									assign node283 = (inp[9]) ? node285 : 1'b0;
										assign node285 = (inp[14]) ? 1'b0 : node286;
											assign node286 = (inp[3]) ? node288 : 1'b1;
												assign node288 = (inp[2]) ? node290 : 1'b0;
													assign node290 = (inp[7]) ? 1'b0 : 1'b1;
			assign node295 = (inp[11]) ? node541 : node296;
				assign node296 = (inp[13]) ? node424 : node297;
					assign node297 = (inp[14]) ? node365 : node298;
						assign node298 = (inp[0]) ? node326 : node299;
							assign node299 = (inp[5]) ? node319 : node300;
								assign node300 = (inp[6]) ? node308 : node301;
									assign node301 = (inp[12]) ? node303 : 1'b0;
										assign node303 = (inp[15]) ? 1'b0 : node304;
											assign node304 = (inp[9]) ? 1'b0 : 1'b1;
									assign node308 = (inp[15]) ? node314 : node309;
										assign node309 = (inp[12]) ? 1'b0 : node310;
											assign node310 = (inp[9]) ? 1'b0 : 1'b1;
										assign node314 = (inp[7]) ? node316 : 1'b1;
											assign node316 = (inp[9]) ? 1'b0 : 1'b1;
								assign node319 = (inp[12]) ? node321 : 1'b0;
									assign node321 = (inp[15]) ? 1'b0 : node322;
										assign node322 = (inp[2]) ? 1'b1 : 1'b0;
							assign node326 = (inp[4]) ? node346 : node327;
								assign node327 = (inp[6]) ? node329 : 1'b1;
									assign node329 = (inp[3]) ? node337 : node330;
										assign node330 = (inp[9]) ? 1'b1 : node331;
											assign node331 = (inp[15]) ? node333 : 1'b1;
												assign node333 = (inp[5]) ? 1'b1 : 1'b0;
										assign node337 = (inp[7]) ? 1'b0 : node338;
											assign node338 = (inp[9]) ? node340 : 1'b1;
												assign node340 = (inp[2]) ? 1'b0 : node341;
													assign node341 = (inp[5]) ? 1'b0 : 1'b1;
								assign node346 = (inp[5]) ? node360 : node347;
									assign node347 = (inp[6]) ? node355 : node348;
										assign node348 = (inp[12]) ? node350 : 1'b0;
											assign node350 = (inp[15]) ? 1'b0 : node351;
												assign node351 = (inp[10]) ? 1'b0 : 1'b1;
										assign node355 = (inp[15]) ? 1'b1 : node356;
											assign node356 = (inp[12]) ? 1'b0 : 1'b1;
									assign node360 = (inp[12]) ? node362 : 1'b0;
										assign node362 = (inp[15]) ? 1'b0 : 1'b1;
						assign node365 = (inp[2]) ? node395 : node366;
							assign node366 = (inp[9]) ? node386 : node367;
								assign node367 = (inp[4]) ? node375 : node368;
									assign node368 = (inp[12]) ? node370 : 1'b1;
										assign node370 = (inp[5]) ? 1'b0 : node371;
											assign node371 = (inp[0]) ? 1'b0 : 1'b1;
									assign node375 = (inp[5]) ? node381 : node376;
										assign node376 = (inp[0]) ? 1'b0 : node377;
											assign node377 = (inp[12]) ? 1'b1 : 1'b0;
										assign node381 = (inp[0]) ? 1'b1 : node382;
											assign node382 = (inp[7]) ? 1'b1 : 1'b0;
								assign node386 = (inp[4]) ? 1'b1 : node387;
									assign node387 = (inp[6]) ? node389 : 1'b1;
										assign node389 = (inp[12]) ? 1'b1 : node390;
											assign node390 = (inp[5]) ? 1'b1 : 1'b0;
							assign node395 = (inp[15]) ? node417 : node396;
								assign node396 = (inp[12]) ? node406 : node397;
									assign node397 = (inp[9]) ? 1'b0 : node398;
										assign node398 = (inp[3]) ? node400 : 1'b0;
											assign node400 = (inp[0]) ? 1'b1 : node401;
												assign node401 = (inp[10]) ? 1'b0 : 1'b1;
									assign node406 = (inp[5]) ? 1'b1 : node407;
										assign node407 = (inp[3]) ? 1'b0 : node408;
											assign node408 = (inp[6]) ? node412 : node409;
												assign node409 = (inp[9]) ? 1'b0 : 1'b1;
												assign node412 = (inp[9]) ? 1'b1 : 1'b0;
								assign node417 = (inp[4]) ? 1'b0 : node418;
									assign node418 = (inp[0]) ? node420 : 1'b0;
										assign node420 = (inp[6]) ? 1'b0 : 1'b1;
					assign node424 = (inp[9]) ? node498 : node425;
						assign node425 = (inp[0]) ? node463 : node426;
							assign node426 = (inp[2]) ? node444 : node427;
								assign node427 = (inp[14]) ? node437 : node428;
									assign node428 = (inp[10]) ? node430 : 1'b1;
										assign node430 = (inp[7]) ? 1'b0 : node431;
											assign node431 = (inp[4]) ? 1'b1 : node432;
												assign node432 = (inp[3]) ? 1'b1 : 1'b0;
									assign node437 = (inp[12]) ? node439 : 1'b0;
										assign node439 = (inp[15]) ? 1'b0 : node440;
											assign node440 = (inp[6]) ? 1'b0 : 1'b1;
								assign node444 = (inp[12]) ? node452 : node445;
									assign node445 = (inp[5]) ? 1'b1 : node446;
										assign node446 = (inp[6]) ? node448 : 1'b1;
											assign node448 = (inp[4]) ? 1'b1 : 1'b0;
									assign node452 = (inp[7]) ? node458 : node453;
										assign node453 = (inp[15]) ? 1'b1 : node454;
											assign node454 = (inp[10]) ? 1'b0 : 1'b1;
										assign node458 = (inp[15]) ? node460 : 1'b0;
											assign node460 = (inp[6]) ? 1'b0 : 1'b1;
							assign node463 = (inp[5]) ? node487 : node464;
								assign node464 = (inp[7]) ? node476 : node465;
									assign node465 = (inp[14]) ? node467 : 1'b1;
										assign node467 = (inp[3]) ? 1'b1 : node468;
											assign node468 = (inp[15]) ? node472 : node469;
												assign node469 = (inp[4]) ? 1'b0 : 1'b1;
												assign node472 = (inp[4]) ? 1'b1 : 1'b0;
									assign node476 = (inp[12]) ? 1'b0 : node477;
										assign node477 = (inp[3]) ? node479 : 1'b1;
											assign node479 = (inp[14]) ? node481 : 1'b0;
												assign node481 = (inp[4]) ? node483 : 1'b1;
													assign node483 = (inp[10]) ? 1'b0 : 1'b1;
								assign node487 = (inp[12]) ? node489 : 1'b1;
									assign node489 = (inp[4]) ? node495 : node490;
										assign node490 = (inp[15]) ? 1'b1 : node491;
											assign node491 = (inp[10]) ? 1'b0 : 1'b1;
										assign node495 = (inp[10]) ? 1'b1 : 1'b0;
						assign node498 = (inp[2]) ? node522 : node499;
							assign node499 = (inp[14]) ? node507 : node500;
								assign node500 = (inp[0]) ? node502 : 1'b1;
									assign node502 = (inp[5]) ? 1'b1 : node503;
										assign node503 = (inp[6]) ? 1'b0 : 1'b1;
								assign node507 = (inp[4]) ? node517 : node508;
									assign node508 = (inp[12]) ? node510 : 1'b1;
										assign node510 = (inp[10]) ? node512 : 1'b1;
											assign node512 = (inp[3]) ? node514 : 1'b0;
												assign node514 = (inp[6]) ? 1'b0 : 1'b1;
									assign node517 = (inp[6]) ? node519 : 1'b0;
										assign node519 = (inp[0]) ? 1'b0 : 1'b1;
							assign node522 = (inp[12]) ? node524 : 1'b1;
								assign node524 = (inp[14]) ? node526 : 1'b1;
									assign node526 = (inp[7]) ? 1'b1 : node527;
										assign node527 = (inp[0]) ? node535 : node528;
											assign node528 = (inp[15]) ? 1'b1 : node529;
												assign node529 = (inp[5]) ? node531 : 1'b0;
													assign node531 = (inp[6]) ? 1'b0 : 1'b1;
											assign node535 = (inp[15]) ? node537 : 1'b1;
												assign node537 = (inp[3]) ? 1'b0 : 1'b1;
				assign node541 = (inp[2]) ? node653 : node542;
					assign node542 = (inp[14]) ? node610 : node543;
						assign node543 = (inp[5]) ? node591 : node544;
							assign node544 = (inp[3]) ? node574 : node545;
								assign node545 = (inp[6]) ? node561 : node546;
									assign node546 = (inp[0]) ? node552 : node547;
										assign node547 = (inp[15]) ? 1'b0 : node548;
											assign node548 = (inp[7]) ? 1'b0 : 1'b1;
										assign node552 = (inp[13]) ? 1'b1 : node553;
											assign node553 = (inp[7]) ? 1'b0 : node554;
												assign node554 = (inp[15]) ? 1'b1 : node555;
													assign node555 = (inp[4]) ? 1'b1 : 1'b0;
									assign node561 = (inp[10]) ? 1'b1 : node562;
										assign node562 = (inp[0]) ? node566 : node563;
											assign node563 = (inp[9]) ? 1'b0 : 1'b1;
											assign node566 = (inp[13]) ? node570 : node567;
												assign node567 = (inp[12]) ? 1'b0 : 1'b1;
												assign node570 = (inp[9]) ? 1'b1 : 1'b0;
								assign node574 = (inp[13]) ? node584 : node575;
									assign node575 = (inp[7]) ? node577 : 1'b0;
										assign node577 = (inp[0]) ? node579 : 1'b0;
											assign node579 = (inp[6]) ? node581 : 1'b1;
												assign node581 = (inp[4]) ? 1'b1 : 1'b0;
									assign node584 = (inp[15]) ? 1'b0 : node585;
										assign node585 = (inp[0]) ? 1'b1 : node586;
											assign node586 = (inp[12]) ? 1'b1 : 1'b0;
							assign node591 = (inp[4]) ? node603 : node592;
								assign node592 = (inp[0]) ? node600 : node593;
									assign node593 = (inp[3]) ? 1'b0 : node594;
										assign node594 = (inp[12]) ? node596 : 1'b0;
											assign node596 = (inp[15]) ? 1'b0 : 1'b1;
									assign node600 = (inp[15]) ? 1'b1 : 1'b0;
								assign node603 = (inp[15]) ? 1'b0 : node604;
									assign node604 = (inp[12]) ? node606 : 1'b0;
										assign node606 = (inp[13]) ? 1'b0 : 1'b1;
						assign node610 = (inp[12]) ? node624 : node611;
							assign node611 = (inp[6]) ? node613 : 1'b1;
								assign node613 = (inp[5]) ? 1'b1 : node614;
									assign node614 = (inp[10]) ? 1'b0 : node615;
										assign node615 = (inp[15]) ? 1'b1 : node616;
											assign node616 = (inp[7]) ? node618 : 1'b0;
												assign node618 = (inp[3]) ? 1'b1 : 1'b0;
							assign node624 = (inp[15]) ? node638 : node625;
								assign node625 = (inp[7]) ? node633 : node626;
									assign node626 = (inp[6]) ? 1'b1 : node627;
										assign node627 = (inp[5]) ? 1'b0 : node628;
											assign node628 = (inp[10]) ? 1'b0 : 1'b1;
									assign node633 = (inp[9]) ? node635 : 1'b0;
										assign node635 = (inp[10]) ? 1'b0 : 1'b1;
								assign node638 = (inp[5]) ? 1'b1 : node639;
									assign node639 = (inp[6]) ? node641 : 1'b1;
										assign node641 = (inp[10]) ? 1'b0 : node642;
											assign node642 = (inp[4]) ? 1'b1 : node643;
												assign node643 = (inp[13]) ? 1'b0 : node644;
													assign node644 = (inp[0]) ? 1'b1 : node645;
														assign node645 = (inp[3]) ? 1'b1 : 1'b0;
					assign node653 = (inp[4]) ? node705 : node654;
						assign node654 = (inp[0]) ? node680 : node655;
							assign node655 = (inp[3]) ? node673 : node656;
								assign node656 = (inp[10]) ? node666 : node657;
									assign node657 = (inp[6]) ? node659 : 1'b0;
										assign node659 = (inp[5]) ? 1'b0 : node660;
											assign node660 = (inp[15]) ? 1'b1 : node661;
												assign node661 = (inp[12]) ? 1'b0 : 1'b1;
									assign node666 = (inp[7]) ? 1'b1 : node667;
										assign node667 = (inp[9]) ? node669 : 1'b0;
											assign node669 = (inp[15]) ? 1'b0 : 1'b1;
								assign node673 = (inp[12]) ? node675 : 1'b0;
									assign node675 = (inp[13]) ? node677 : 1'b0;
										assign node677 = (inp[5]) ? 1'b1 : 1'b0;
							assign node680 = (inp[15]) ? node696 : node681;
								assign node681 = (inp[12]) ? node687 : node682;
									assign node682 = (inp[3]) ? 1'b1 : node683;
										assign node683 = (inp[14]) ? 1'b1 : 1'b0;
									assign node687 = (inp[13]) ? node691 : node688;
										assign node688 = (inp[7]) ? 1'b0 : 1'b1;
										assign node691 = (inp[6]) ? node693 : 1'b0;
											assign node693 = (inp[3]) ? 1'b1 : 1'b0;
								assign node696 = (inp[6]) ? node698 : 1'b1;
									assign node698 = (inp[5]) ? 1'b1 : node699;
										assign node699 = (inp[10]) ? 1'b0 : node700;
											assign node700 = (inp[9]) ? 1'b1 : 1'b0;
						assign node705 = (inp[15]) ? node723 : node706;
							assign node706 = (inp[12]) ? node716 : node707;
								assign node707 = (inp[6]) ? node709 : 1'b0;
									assign node709 = (inp[5]) ? 1'b0 : node710;
										assign node710 = (inp[3]) ? node712 : 1'b1;
											assign node712 = (inp[7]) ? 1'b1 : 1'b0;
								assign node716 = (inp[5]) ? 1'b1 : node717;
									assign node717 = (inp[10]) ? node719 : 1'b0;
										assign node719 = (inp[13]) ? 1'b1 : 1'b0;
							assign node723 = (inp[6]) ? node725 : 1'b0;
								assign node725 = (inp[5]) ? 1'b0 : node726;
									assign node726 = (inp[7]) ? 1'b1 : node727;
										assign node727 = (inp[3]) ? 1'b0 : node728;
											assign node728 = (inp[10]) ? 1'b1 : 1'b0;
		assign node734 = (inp[4]) ? node1044 : node735;
			assign node735 = (inp[0]) ? node827 : node736;
				assign node736 = (inp[6]) ? node758 : node737;
					assign node737 = (inp[12]) ? node739 : 1'b1;
						assign node739 = (inp[15]) ? 1'b1 : node740;
							assign node740 = (inp[9]) ? node746 : node741;
								assign node741 = (inp[7]) ? 1'b0 : node742;
									assign node742 = (inp[3]) ? 1'b1 : 1'b0;
								assign node746 = (inp[10]) ? node752 : node747;
									assign node747 = (inp[7]) ? 1'b1 : node748;
										assign node748 = (inp[3]) ? 1'b0 : 1'b1;
									assign node752 = (inp[7]) ? 1'b0 : node753;
										assign node753 = (inp[3]) ? 1'b1 : 1'b0;
					assign node758 = (inp[5]) ? node800 : node759;
						assign node759 = (inp[3]) ? node777 : node760;
							assign node760 = (inp[10]) ? node772 : node761;
								assign node761 = (inp[9]) ? 1'b1 : node762;
									assign node762 = (inp[14]) ? node764 : 1'b0;
										assign node764 = (inp[7]) ? 1'b1 : node765;
											assign node765 = (inp[1]) ? node767 : 1'b0;
												assign node767 = (inp[15]) ? 1'b0 : 1'b1;
								assign node772 = (inp[12]) ? node774 : 1'b0;
									assign node774 = (inp[15]) ? 1'b0 : 1'b1;
							assign node777 = (inp[7]) ? node789 : node778;
								assign node778 = (inp[2]) ? 1'b1 : node779;
									assign node779 = (inp[10]) ? 1'b1 : node780;
										assign node780 = (inp[12]) ? node782 : 1'b0;
											assign node782 = (inp[11]) ? 1'b1 : node783;
												assign node783 = (inp[13]) ? 1'b1 : 1'b0;
								assign node789 = (inp[10]) ? node795 : node790;
									assign node790 = (inp[9]) ? 1'b1 : node791;
										assign node791 = (inp[13]) ? 1'b1 : 1'b0;
									assign node795 = (inp[12]) ? node797 : 1'b0;
										assign node797 = (inp[11]) ? 1'b1 : 1'b0;
						assign node800 = (inp[15]) ? 1'b1 : node801;
							assign node801 = (inp[12]) ? node803 : 1'b1;
								assign node803 = (inp[1]) ? node819 : node804;
									assign node804 = (inp[11]) ? node816 : node805;
										assign node805 = (inp[13]) ? node811 : node806;
											assign node806 = (inp[9]) ? node808 : 1'b0;
												assign node808 = (inp[14]) ? 1'b0 : 1'b1;
											assign node811 = (inp[9]) ? 1'b1 : node812;
												assign node812 = (inp[14]) ? 1'b1 : 1'b0;
										assign node816 = (inp[14]) ? 1'b1 : 1'b0;
									assign node819 = (inp[13]) ? 1'b0 : node820;
										assign node820 = (inp[3]) ? 1'b0 : node821;
											assign node821 = (inp[7]) ? 1'b0 : 1'b1;
				assign node827 = (inp[11]) ? node949 : node828;
					assign node828 = (inp[13]) ? node890 : node829;
						assign node829 = (inp[14]) ? node857 : node830;
							assign node830 = (inp[9]) ? node846 : node831;
								assign node831 = (inp[3]) ? node837 : node832;
									assign node832 = (inp[6]) ? 1'b1 : node833;
										assign node833 = (inp[15]) ? 1'b0 : 1'b1;
									assign node837 = (inp[7]) ? node839 : 1'b0;
										assign node839 = (inp[1]) ? node841 : 1'b0;
											assign node841 = (inp[15]) ? node843 : 1'b1;
												assign node843 = (inp[2]) ? 1'b0 : 1'b1;
								assign node846 = (inp[3]) ? node848 : 1'b0;
									assign node848 = (inp[6]) ? node854 : node849;
										assign node849 = (inp[1]) ? 1'b0 : node850;
											assign node850 = (inp[5]) ? 1'b1 : 1'b0;
										assign node854 = (inp[5]) ? 1'b0 : 1'b1;
							assign node857 = (inp[2]) ? node877 : node858;
								assign node858 = (inp[5]) ? node870 : node859;
									assign node859 = (inp[3]) ? 1'b1 : node860;
										assign node860 = (inp[15]) ? 1'b0 : node861;
											assign node861 = (inp[1]) ? 1'b1 : node862;
												assign node862 = (inp[6]) ? 1'b1 : node863;
													assign node863 = (inp[10]) ? 1'b0 : 1'b1;
									assign node870 = (inp[15]) ? 1'b1 : node871;
										assign node871 = (inp[3]) ? node873 : 1'b1;
											assign node873 = (inp[12]) ? 1'b0 : 1'b1;
								assign node877 = (inp[9]) ? 1'b0 : node878;
									assign node878 = (inp[5]) ? node884 : node879;
										assign node879 = (inp[12]) ? 1'b1 : node880;
											assign node880 = (inp[1]) ? 1'b1 : 1'b0;
										assign node884 = (inp[3]) ? 1'b0 : node885;
											assign node885 = (inp[15]) ? 1'b0 : 1'b1;
						assign node890 = (inp[2]) ? node920 : node891;
							assign node891 = (inp[14]) ? node909 : node892;
								assign node892 = (inp[9]) ? node904 : node893;
									assign node893 = (inp[5]) ? node901 : node894;
										assign node894 = (inp[12]) ? node896 : 1'b0;
											assign node896 = (inp[15]) ? node898 : 1'b1;
												assign node898 = (inp[3]) ? 1'b0 : 1'b1;
										assign node901 = (inp[15]) ? 1'b1 : 1'b0;
									assign node904 = (inp[10]) ? node906 : 1'b1;
										assign node906 = (inp[1]) ? 1'b0 : 1'b1;
								assign node909 = (inp[15]) ? 1'b0 : node910;
									assign node910 = (inp[6]) ? 1'b1 : node911;
										assign node911 = (inp[3]) ? 1'b0 : node912;
											assign node912 = (inp[12]) ? node914 : 1'b0;
												assign node914 = (inp[9]) ? 1'b0 : 1'b1;
							assign node920 = (inp[12]) ? node930 : node921;
								assign node921 = (inp[6]) ? node923 : 1'b1;
									assign node923 = (inp[5]) ? 1'b1 : node924;
										assign node924 = (inp[9]) ? 1'b1 : node925;
											assign node925 = (inp[3]) ? 1'b1 : 1'b0;
								assign node930 = (inp[15]) ? node944 : node931;
									assign node931 = (inp[6]) ? node939 : node932;
										assign node932 = (inp[3]) ? node934 : 1'b0;
											assign node934 = (inp[9]) ? 1'b0 : node935;
												assign node935 = (inp[7]) ? 1'b0 : 1'b1;
										assign node939 = (inp[5]) ? node941 : 1'b1;
											assign node941 = (inp[1]) ? 1'b1 : 1'b0;
									assign node944 = (inp[6]) ? node946 : 1'b1;
										assign node946 = (inp[5]) ? 1'b1 : 1'b0;
					assign node949 = (inp[14]) ? node997 : node950;
						assign node950 = (inp[6]) ? node964 : node951;
							assign node951 = (inp[12]) ? node953 : 1'b0;
								assign node953 = (inp[15]) ? 1'b0 : node954;
									assign node954 = (inp[1]) ? node956 : 1'b0;
										assign node956 = (inp[13]) ? node958 : 1'b1;
											assign node958 = (inp[5]) ? node960 : 1'b1;
												assign node960 = (inp[2]) ? 1'b1 : 1'b0;
							assign node964 = (inp[9]) ? node978 : node965;
								assign node965 = (inp[3]) ? node971 : node966;
									assign node966 = (inp[13]) ? node968 : 1'b1;
										assign node968 = (inp[2]) ? 1'b0 : 1'b1;
									assign node971 = (inp[7]) ? node973 : 1'b0;
										assign node973 = (inp[10]) ? node975 : 1'b1;
											assign node975 = (inp[1]) ? 1'b1 : 1'b0;
								assign node978 = (inp[10]) ? node986 : node979;
									assign node979 = (inp[12]) ? 1'b0 : node980;
										assign node980 = (inp[7]) ? 1'b0 : node981;
											assign node981 = (inp[13]) ? 1'b1 : 1'b0;
									assign node986 = (inp[13]) ? node988 : 1'b1;
										assign node988 = (inp[5]) ? 1'b0 : node989;
											assign node989 = (inp[2]) ? node991 : 1'b1;
												assign node991 = (inp[12]) ? 1'b0 : node992;
													assign node992 = (inp[15]) ? 1'b0 : 1'b1;
						assign node997 = (inp[2]) ? node1021 : node998;
							assign node998 = (inp[12]) ? node1008 : node999;
								assign node999 = (inp[5]) ? 1'b1 : node1000;
									assign node1000 = (inp[6]) ? node1002 : 1'b1;
										assign node1002 = (inp[1]) ? 1'b0 : node1003;
											assign node1003 = (inp[10]) ? 1'b0 : 1'b1;
								assign node1008 = (inp[3]) ? node1014 : node1009;
									assign node1009 = (inp[9]) ? node1011 : 1'b0;
										assign node1011 = (inp[1]) ? 1'b1 : 1'b0;
									assign node1014 = (inp[7]) ? node1016 : 1'b1;
										assign node1016 = (inp[9]) ? node1018 : 1'b0;
											assign node1018 = (inp[6]) ? 1'b0 : 1'b1;
							assign node1021 = (inp[12]) ? node1031 : node1022;
								assign node1022 = (inp[1]) ? node1024 : 1'b0;
									assign node1024 = (inp[6]) ? node1026 : 1'b0;
										assign node1026 = (inp[9]) ? 1'b0 : node1027;
											assign node1027 = (inp[5]) ? 1'b0 : 1'b1;
								assign node1031 = (inp[15]) ? node1039 : node1032;
									assign node1032 = (inp[5]) ? 1'b1 : node1033;
										assign node1033 = (inp[10]) ? node1035 : 1'b0;
											assign node1035 = (inp[7]) ? 1'b1 : 1'b0;
									assign node1039 = (inp[5]) ? 1'b0 : node1040;
										assign node1040 = (inp[6]) ? 1'b1 : 1'b0;
			assign node1044 = (inp[12]) ? node1066 : node1045;
				assign node1045 = (inp[5]) ? 1'b1 : node1046;
					assign node1046 = (inp[6]) ? node1048 : 1'b1;
						assign node1048 = (inp[10]) ? node1060 : node1049;
							assign node1049 = (inp[9]) ? node1055 : node1050;
								assign node1050 = (inp[3]) ? node1052 : 1'b0;
									assign node1052 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1055 = (inp[7]) ? 1'b1 : node1056;
									assign node1056 = (inp[3]) ? 1'b0 : 1'b1;
							assign node1060 = (inp[3]) ? node1062 : 1'b0;
								assign node1062 = (inp[7]) ? 1'b0 : 1'b1;
				assign node1066 = (inp[15]) ? node1104 : node1067;
					assign node1067 = (inp[5]) ? node1087 : node1068;
						assign node1068 = (inp[6]) ? 1'b1 : node1069;
							assign node1069 = (inp[9]) ? node1075 : node1070;
								assign node1070 = (inp[3]) ? node1072 : 1'b0;
									assign node1072 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1075 = (inp[10]) ? node1081 : node1076;
									assign node1076 = (inp[7]) ? 1'b1 : node1077;
										assign node1077 = (inp[0]) ? 1'b1 : 1'b0;
									assign node1081 = (inp[3]) ? node1083 : 1'b0;
										assign node1083 = (inp[0]) ? 1'b0 : 1'b1;
						assign node1087 = (inp[7]) ? node1099 : node1088;
							assign node1088 = (inp[3]) ? node1094 : node1089;
								assign node1089 = (inp[9]) ? node1091 : 1'b0;
									assign node1091 = (inp[10]) ? 1'b0 : 1'b1;
								assign node1094 = (inp[9]) ? node1096 : 1'b1;
									assign node1096 = (inp[10]) ? 1'b1 : 1'b0;
							assign node1099 = (inp[10]) ? 1'b0 : node1100;
								assign node1100 = (inp[9]) ? 1'b1 : 1'b0;
					assign node1104 = (inp[5]) ? 1'b1 : node1105;
						assign node1105 = (inp[6]) ? node1107 : 1'b1;
							assign node1107 = (inp[7]) ? node1119 : node1108;
								assign node1108 = (inp[3]) ? node1114 : node1109;
									assign node1109 = (inp[9]) ? node1111 : 1'b0;
										assign node1111 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1114 = (inp[10]) ? 1'b1 : node1115;
										assign node1115 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1119 = (inp[10]) ? 1'b0 : node1120;
									assign node1120 = (inp[9]) ? 1'b1 : 1'b0;

endmodule