module dtc_split875_bm45 (
	input  wire [16-1:0] inp,
	output wire [46-1:0] outp
);

	wire [46-1:0] node1;
	wire [46-1:0] node2;
	wire [46-1:0] node3;
	wire [46-1:0] node5;
	wire [46-1:0] node7;
	wire [46-1:0] node9;
	wire [46-1:0] node11;
	wire [46-1:0] node12;
	wire [46-1:0] node14;
	wire [46-1:0] node16;
	wire [46-1:0] node18;
	wire [46-1:0] node20;
	wire [46-1:0] node22;
	wire [46-1:0] node25;
	wire [46-1:0] node27;
	wire [46-1:0] node29;
	wire [46-1:0] node31;
	wire [46-1:0] node33;
	wire [46-1:0] node35;
	wire [46-1:0] node38;
	wire [46-1:0] node40;
	wire [46-1:0] node41;
	wire [46-1:0] node43;
	wire [46-1:0] node45;
	wire [46-1:0] node47;
	wire [46-1:0] node49;
	wire [46-1:0] node50;
	wire [46-1:0] node51;
	wire [46-1:0] node54;
	wire [46-1:0] node56;
	wire [46-1:0] node58;
	wire [46-1:0] node61;
	wire [46-1:0] node63;
	wire [46-1:0] node65;
	wire [46-1:0] node67;
	wire [46-1:0] node71;
	wire [46-1:0] node73;
	wire [46-1:0] node74;
	wire [46-1:0] node75;
	wire [46-1:0] node76;
	wire [46-1:0] node77;
	wire [46-1:0] node80;
	wire [46-1:0] node82;
	wire [46-1:0] node84;
	wire [46-1:0] node85;
	wire [46-1:0] node87;
	wire [46-1:0] node88;
	wire [46-1:0] node90;
	wire [46-1:0] node93;
	wire [46-1:0] node94;
	wire [46-1:0] node97;
	wire [46-1:0] node101;
	wire [46-1:0] node103;
	wire [46-1:0] node105;
	wire [46-1:0] node107;
	wire [46-1:0] node109;
	wire [46-1:0] node110;
	wire [46-1:0] node111;
	wire [46-1:0] node113;
	wire [46-1:0] node116;
	wire [46-1:0] node117;
	wire [46-1:0] node120;
	wire [46-1:0] node124;
	wire [46-1:0] node125;
	wire [46-1:0] node126;
	wire [46-1:0] node130;
	wire [46-1:0] node131;
	wire [46-1:0] node134;
	wire [46-1:0] node137;
	wire [46-1:0] node138;
	wire [46-1:0] node139;
	wire [46-1:0] node140;
	wire [46-1:0] node143;
	wire [46-1:0] node145;
	wire [46-1:0] node147;
	wire [46-1:0] node148;
	wire [46-1:0] node150;
	wire [46-1:0] node152;
	wire [46-1:0] node154;
	wire [46-1:0] node157;
	wire [46-1:0] node158;
	wire [46-1:0] node160;
	wire [46-1:0] node162;
	wire [46-1:0] node165;
	wire [46-1:0] node166;
	wire [46-1:0] node167;
	wire [46-1:0] node170;
	wire [46-1:0] node173;
	wire [46-1:0] node174;
	wire [46-1:0] node178;
	wire [46-1:0] node179;
	wire [46-1:0] node181;
	wire [46-1:0] node183;
	wire [46-1:0] node185;
	wire [46-1:0] node187;
	wire [46-1:0] node188;
	wire [46-1:0] node190;
	wire [46-1:0] node193;
	wire [46-1:0] node194;
	wire [46-1:0] node197;
	wire [46-1:0] node200;
	wire [46-1:0] node202;
	wire [46-1:0] node204;
	wire [46-1:0] node206;
	wire [46-1:0] node207;
	wire [46-1:0] node209;
	wire [46-1:0] node211;
	wire [46-1:0] node214;
	wire [46-1:0] node215;
	wire [46-1:0] node217;
	wire [46-1:0] node220;
	wire [46-1:0] node221;
	wire [46-1:0] node224;
	wire [46-1:0] node227;
	wire [46-1:0] node229;
	wire [46-1:0] node231;
	wire [46-1:0] node233;
	wire [46-1:0] node234;
	wire [46-1:0] node236;
	wire [46-1:0] node238;
	wire [46-1:0] node240;
	wire [46-1:0] node242;
	wire [46-1:0] node245;
	wire [46-1:0] node246;
	wire [46-1:0] node247;
	wire [46-1:0] node248;
	wire [46-1:0] node250;
	wire [46-1:0] node253;
	wire [46-1:0] node254;
	wire [46-1:0] node257;
	wire [46-1:0] node261;
	wire [46-1:0] node262;
	wire [46-1:0] node264;
	wire [46-1:0] node266;
	wire [46-1:0] node269;
	wire [46-1:0] node270;
	wire [46-1:0] node271;
	wire [46-1:0] node274;
	wire [46-1:0] node277;
	wire [46-1:0] node278;
	wire [46-1:0] node282;
	wire [46-1:0] node283;
	wire [46-1:0] node284;
	wire [46-1:0] node287;
	wire [46-1:0] node288;
	wire [46-1:0] node289;
	wire [46-1:0] node290;
	wire [46-1:0] node291;
	wire [46-1:0] node294;
	wire [46-1:0] node297;
	wire [46-1:0] node298;
	wire [46-1:0] node301;
	wire [46-1:0] node304;
	wire [46-1:0] node305;
	wire [46-1:0] node306;
	wire [46-1:0] node309;
	wire [46-1:0] node312;
	wire [46-1:0] node313;
	wire [46-1:0] node316;
	wire [46-1:0] node319;
	wire [46-1:0] node320;
	wire [46-1:0] node321;
	wire [46-1:0] node322;
	wire [46-1:0] node325;
	wire [46-1:0] node328;
	wire [46-1:0] node329;
	wire [46-1:0] node332;
	wire [46-1:0] node335;
	wire [46-1:0] node336;
	wire [46-1:0] node337;
	wire [46-1:0] node340;
	wire [46-1:0] node343;
	wire [46-1:0] node344;
	wire [46-1:0] node347;
	wire [46-1:0] node350;
	wire [46-1:0] node351;
	wire [46-1:0] node354;
	wire [46-1:0] node356;
	wire [46-1:0] node357;
	wire [46-1:0] node358;
	wire [46-1:0] node359;
	wire [46-1:0] node360;
	wire [46-1:0] node361;
	wire [46-1:0] node362;
	wire [46-1:0] node363;
	wire [46-1:0] node364;
	wire [46-1:0] node365;
	wire [46-1:0] node368;
	wire [46-1:0] node371;
	wire [46-1:0] node372;
	wire [46-1:0] node375;
	wire [46-1:0] node378;
	wire [46-1:0] node379;
	wire [46-1:0] node380;
	wire [46-1:0] node383;
	wire [46-1:0] node386;
	wire [46-1:0] node387;
	wire [46-1:0] node390;
	wire [46-1:0] node393;
	wire [46-1:0] node394;
	wire [46-1:0] node395;
	wire [46-1:0] node396;
	wire [46-1:0] node399;
	wire [46-1:0] node402;
	wire [46-1:0] node403;
	wire [46-1:0] node406;
	wire [46-1:0] node409;
	wire [46-1:0] node410;
	wire [46-1:0] node411;
	wire [46-1:0] node414;
	wire [46-1:0] node417;
	wire [46-1:0] node418;
	wire [46-1:0] node421;
	wire [46-1:0] node424;
	wire [46-1:0] node425;
	wire [46-1:0] node426;
	wire [46-1:0] node427;
	wire [46-1:0] node428;
	wire [46-1:0] node431;
	wire [46-1:0] node434;
	wire [46-1:0] node435;
	wire [46-1:0] node438;
	wire [46-1:0] node441;
	wire [46-1:0] node442;
	wire [46-1:0] node443;
	wire [46-1:0] node446;
	wire [46-1:0] node449;
	wire [46-1:0] node450;
	wire [46-1:0] node453;
	wire [46-1:0] node456;
	wire [46-1:0] node457;
	wire [46-1:0] node458;
	wire [46-1:0] node459;
	wire [46-1:0] node462;
	wire [46-1:0] node465;
	wire [46-1:0] node466;
	wire [46-1:0] node469;
	wire [46-1:0] node472;
	wire [46-1:0] node473;
	wire [46-1:0] node474;
	wire [46-1:0] node477;
	wire [46-1:0] node480;
	wire [46-1:0] node481;
	wire [46-1:0] node484;
	wire [46-1:0] node487;
	wire [46-1:0] node488;
	wire [46-1:0] node489;
	wire [46-1:0] node490;
	wire [46-1:0] node491;
	wire [46-1:0] node492;
	wire [46-1:0] node495;
	wire [46-1:0] node498;
	wire [46-1:0] node499;
	wire [46-1:0] node502;
	wire [46-1:0] node505;
	wire [46-1:0] node506;
	wire [46-1:0] node507;
	wire [46-1:0] node510;
	wire [46-1:0] node513;
	wire [46-1:0] node514;
	wire [46-1:0] node517;
	wire [46-1:0] node520;
	wire [46-1:0] node521;
	wire [46-1:0] node522;
	wire [46-1:0] node523;
	wire [46-1:0] node526;
	wire [46-1:0] node529;
	wire [46-1:0] node530;
	wire [46-1:0] node533;
	wire [46-1:0] node536;
	wire [46-1:0] node537;
	wire [46-1:0] node538;
	wire [46-1:0] node541;
	wire [46-1:0] node544;
	wire [46-1:0] node545;
	wire [46-1:0] node548;
	wire [46-1:0] node551;
	wire [46-1:0] node552;
	wire [46-1:0] node553;
	wire [46-1:0] node554;
	wire [46-1:0] node555;
	wire [46-1:0] node558;
	wire [46-1:0] node561;
	wire [46-1:0] node562;
	wire [46-1:0] node565;
	wire [46-1:0] node568;
	wire [46-1:0] node569;
	wire [46-1:0] node570;
	wire [46-1:0] node573;
	wire [46-1:0] node576;
	wire [46-1:0] node577;
	wire [46-1:0] node580;
	wire [46-1:0] node583;
	wire [46-1:0] node584;
	wire [46-1:0] node585;
	wire [46-1:0] node586;
	wire [46-1:0] node589;
	wire [46-1:0] node592;
	wire [46-1:0] node593;
	wire [46-1:0] node596;
	wire [46-1:0] node599;
	wire [46-1:0] node600;
	wire [46-1:0] node601;
	wire [46-1:0] node604;
	wire [46-1:0] node607;
	wire [46-1:0] node608;
	wire [46-1:0] node611;
	wire [46-1:0] node614;
	wire [46-1:0] node615;
	wire [46-1:0] node617;
	wire [46-1:0] node619;
	wire [46-1:0] node620;
	wire [46-1:0] node622;
	wire [46-1:0] node623;
	wire [46-1:0] node626;
	wire [46-1:0] node629;
	wire [46-1:0] node630;
	wire [46-1:0] node631;
	wire [46-1:0] node634;
	wire [46-1:0] node638;
	wire [46-1:0] node639;
	wire [46-1:0] node640;
	wire [46-1:0] node641;
	wire [46-1:0] node642;
	wire [46-1:0] node643;
	wire [46-1:0] node646;
	wire [46-1:0] node649;
	wire [46-1:0] node650;
	wire [46-1:0] node653;
	wire [46-1:0] node656;
	wire [46-1:0] node657;
	wire [46-1:0] node658;
	wire [46-1:0] node661;
	wire [46-1:0] node664;
	wire [46-1:0] node665;
	wire [46-1:0] node668;
	wire [46-1:0] node671;
	wire [46-1:0] node672;
	wire [46-1:0] node673;
	wire [46-1:0] node674;
	wire [46-1:0] node677;
	wire [46-1:0] node680;
	wire [46-1:0] node681;
	wire [46-1:0] node684;
	wire [46-1:0] node687;
	wire [46-1:0] node688;
	wire [46-1:0] node689;
	wire [46-1:0] node692;
	wire [46-1:0] node695;
	wire [46-1:0] node696;
	wire [46-1:0] node699;
	wire [46-1:0] node702;
	wire [46-1:0] node703;
	wire [46-1:0] node704;
	wire [46-1:0] node705;
	wire [46-1:0] node706;
	wire [46-1:0] node709;
	wire [46-1:0] node712;
	wire [46-1:0] node713;
	wire [46-1:0] node716;
	wire [46-1:0] node719;
	wire [46-1:0] node720;
	wire [46-1:0] node721;
	wire [46-1:0] node724;
	wire [46-1:0] node727;
	wire [46-1:0] node728;
	wire [46-1:0] node731;
	wire [46-1:0] node734;
	wire [46-1:0] node735;
	wire [46-1:0] node736;
	wire [46-1:0] node737;
	wire [46-1:0] node740;
	wire [46-1:0] node743;
	wire [46-1:0] node744;
	wire [46-1:0] node747;
	wire [46-1:0] node750;
	wire [46-1:0] node751;
	wire [46-1:0] node752;
	wire [46-1:0] node755;
	wire [46-1:0] node758;
	wire [46-1:0] node759;
	wire [46-1:0] node762;
	wire [46-1:0] node765;
	wire [46-1:0] node766;
	wire [46-1:0] node767;
	wire [46-1:0] node768;
	wire [46-1:0] node769;
	wire [46-1:0] node771;
	wire [46-1:0] node772;
	wire [46-1:0] node773;
	wire [46-1:0] node776;
	wire [46-1:0] node779;
	wire [46-1:0] node780;
	wire [46-1:0] node784;
	wire [46-1:0] node785;
	wire [46-1:0] node786;
	wire [46-1:0] node787;
	wire [46-1:0] node791;
	wire [46-1:0] node792;
	wire [46-1:0] node795;
	wire [46-1:0] node799;
	wire [46-1:0] node800;
	wire [46-1:0] node801;
	wire [46-1:0] node803;
	wire [46-1:0] node804;
	wire [46-1:0] node808;
	wire [46-1:0] node810;
	wire [46-1:0] node811;
	wire [46-1:0] node817;
	wire [46-1:0] node818;
	wire [46-1:0] node819;
	wire [46-1:0] node820;
	wire [46-1:0] node821;
	wire [46-1:0] node822;
	wire [46-1:0] node823;
	wire [46-1:0] node826;
	wire [46-1:0] node829;
	wire [46-1:0] node830;
	wire [46-1:0] node833;
	wire [46-1:0] node836;
	wire [46-1:0] node837;
	wire [46-1:0] node838;
	wire [46-1:0] node841;
	wire [46-1:0] node844;
	wire [46-1:0] node845;
	wire [46-1:0] node848;
	wire [46-1:0] node851;
	wire [46-1:0] node852;
	wire [46-1:0] node853;
	wire [46-1:0] node854;
	wire [46-1:0] node857;
	wire [46-1:0] node860;
	wire [46-1:0] node861;
	wire [46-1:0] node864;
	wire [46-1:0] node867;
	wire [46-1:0] node868;
	wire [46-1:0] node869;
	wire [46-1:0] node872;
	wire [46-1:0] node875;
	wire [46-1:0] node876;
	wire [46-1:0] node879;
	wire [46-1:0] node882;
	wire [46-1:0] node883;
	wire [46-1:0] node884;
	wire [46-1:0] node885;
	wire [46-1:0] node886;
	wire [46-1:0] node889;
	wire [46-1:0] node892;
	wire [46-1:0] node893;
	wire [46-1:0] node896;
	wire [46-1:0] node899;
	wire [46-1:0] node900;
	wire [46-1:0] node901;
	wire [46-1:0] node904;
	wire [46-1:0] node907;
	wire [46-1:0] node908;
	wire [46-1:0] node911;
	wire [46-1:0] node914;
	wire [46-1:0] node915;
	wire [46-1:0] node916;
	wire [46-1:0] node917;
	wire [46-1:0] node920;
	wire [46-1:0] node923;
	wire [46-1:0] node924;
	wire [46-1:0] node927;
	wire [46-1:0] node930;
	wire [46-1:0] node931;
	wire [46-1:0] node932;
	wire [46-1:0] node935;
	wire [46-1:0] node938;
	wire [46-1:0] node939;
	wire [46-1:0] node942;
	wire [46-1:0] node945;
	wire [46-1:0] node946;
	wire [46-1:0] node947;
	wire [46-1:0] node948;
	wire [46-1:0] node949;
	wire [46-1:0] node950;
	wire [46-1:0] node953;
	wire [46-1:0] node956;
	wire [46-1:0] node957;
	wire [46-1:0] node960;
	wire [46-1:0] node963;
	wire [46-1:0] node964;
	wire [46-1:0] node965;
	wire [46-1:0] node968;
	wire [46-1:0] node971;
	wire [46-1:0] node972;
	wire [46-1:0] node975;
	wire [46-1:0] node978;
	wire [46-1:0] node979;
	wire [46-1:0] node980;
	wire [46-1:0] node981;
	wire [46-1:0] node984;
	wire [46-1:0] node987;
	wire [46-1:0] node988;
	wire [46-1:0] node991;
	wire [46-1:0] node994;
	wire [46-1:0] node995;
	wire [46-1:0] node996;
	wire [46-1:0] node999;
	wire [46-1:0] node1002;
	wire [46-1:0] node1003;
	wire [46-1:0] node1006;
	wire [46-1:0] node1009;
	wire [46-1:0] node1010;
	wire [46-1:0] node1011;
	wire [46-1:0] node1012;
	wire [46-1:0] node1013;
	wire [46-1:0] node1016;
	wire [46-1:0] node1019;
	wire [46-1:0] node1020;
	wire [46-1:0] node1023;
	wire [46-1:0] node1026;
	wire [46-1:0] node1027;
	wire [46-1:0] node1028;
	wire [46-1:0] node1031;
	wire [46-1:0] node1034;
	wire [46-1:0] node1035;
	wire [46-1:0] node1038;
	wire [46-1:0] node1041;
	wire [46-1:0] node1042;
	wire [46-1:0] node1043;
	wire [46-1:0] node1044;
	wire [46-1:0] node1047;
	wire [46-1:0] node1050;
	wire [46-1:0] node1051;
	wire [46-1:0] node1054;
	wire [46-1:0] node1057;
	wire [46-1:0] node1058;
	wire [46-1:0] node1059;
	wire [46-1:0] node1062;
	wire [46-1:0] node1065;
	wire [46-1:0] node1066;
	wire [46-1:0] node1069;
	wire [46-1:0] node1072;
	wire [46-1:0] node1073;
	wire [46-1:0] node1074;
	wire [46-1:0] node1075;
	wire [46-1:0] node1077;
	wire [46-1:0] node1079;
	wire [46-1:0] node1081;
	wire [46-1:0] node1083;
	wire [46-1:0] node1084;
	wire [46-1:0] node1087;
	wire [46-1:0] node1090;
	wire [46-1:0] node1091;
	wire [46-1:0] node1093;
	wire [46-1:0] node1095;
	wire [46-1:0] node1097;
	wire [46-1:0] node1098;
	wire [46-1:0] node1101;
	wire [46-1:0] node1104;
	wire [46-1:0] node1105;
	wire [46-1:0] node1106;
	wire [46-1:0] node1107;
	wire [46-1:0] node1108;
	wire [46-1:0] node1111;
	wire [46-1:0] node1114;
	wire [46-1:0] node1115;
	wire [46-1:0] node1118;
	wire [46-1:0] node1121;
	wire [46-1:0] node1122;
	wire [46-1:0] node1123;
	wire [46-1:0] node1126;
	wire [46-1:0] node1129;
	wire [46-1:0] node1130;
	wire [46-1:0] node1133;
	wire [46-1:0] node1136;
	wire [46-1:0] node1137;
	wire [46-1:0] node1139;
	wire [46-1:0] node1140;
	wire [46-1:0] node1143;
	wire [46-1:0] node1146;
	wire [46-1:0] node1147;
	wire [46-1:0] node1148;
	wire [46-1:0] node1151;
	wire [46-1:0] node1155;
	wire [46-1:0] node1156;
	wire [46-1:0] node1157;
	wire [46-1:0] node1158;
	wire [46-1:0] node1159;
	wire [46-1:0] node1160;
	wire [46-1:0] node1161;
	wire [46-1:0] node1164;
	wire [46-1:0] node1167;
	wire [46-1:0] node1168;
	wire [46-1:0] node1171;
	wire [46-1:0] node1174;
	wire [46-1:0] node1175;
	wire [46-1:0] node1176;
	wire [46-1:0] node1179;
	wire [46-1:0] node1182;
	wire [46-1:0] node1183;
	wire [46-1:0] node1186;
	wire [46-1:0] node1189;
	wire [46-1:0] node1190;
	wire [46-1:0] node1191;
	wire [46-1:0] node1192;
	wire [46-1:0] node1195;
	wire [46-1:0] node1198;
	wire [46-1:0] node1199;
	wire [46-1:0] node1202;
	wire [46-1:0] node1205;
	wire [46-1:0] node1206;
	wire [46-1:0] node1207;
	wire [46-1:0] node1210;
	wire [46-1:0] node1213;
	wire [46-1:0] node1214;
	wire [46-1:0] node1217;
	wire [46-1:0] node1220;
	wire [46-1:0] node1221;
	wire [46-1:0] node1222;
	wire [46-1:0] node1223;
	wire [46-1:0] node1224;
	wire [46-1:0] node1227;
	wire [46-1:0] node1230;
	wire [46-1:0] node1231;
	wire [46-1:0] node1234;
	wire [46-1:0] node1237;
	wire [46-1:0] node1238;
	wire [46-1:0] node1239;
	wire [46-1:0] node1242;
	wire [46-1:0] node1245;
	wire [46-1:0] node1246;
	wire [46-1:0] node1249;
	wire [46-1:0] node1252;
	wire [46-1:0] node1253;
	wire [46-1:0] node1254;
	wire [46-1:0] node1255;
	wire [46-1:0] node1258;
	wire [46-1:0] node1261;
	wire [46-1:0] node1262;
	wire [46-1:0] node1265;
	wire [46-1:0] node1268;
	wire [46-1:0] node1269;
	wire [46-1:0] node1270;
	wire [46-1:0] node1273;
	wire [46-1:0] node1276;
	wire [46-1:0] node1277;
	wire [46-1:0] node1280;
	wire [46-1:0] node1283;
	wire [46-1:0] node1284;
	wire [46-1:0] node1285;
	wire [46-1:0] node1286;
	wire [46-1:0] node1287;
	wire [46-1:0] node1288;
	wire [46-1:0] node1291;
	wire [46-1:0] node1294;
	wire [46-1:0] node1295;
	wire [46-1:0] node1298;
	wire [46-1:0] node1301;
	wire [46-1:0] node1302;
	wire [46-1:0] node1303;
	wire [46-1:0] node1306;
	wire [46-1:0] node1309;
	wire [46-1:0] node1310;
	wire [46-1:0] node1313;
	wire [46-1:0] node1316;
	wire [46-1:0] node1317;
	wire [46-1:0] node1318;
	wire [46-1:0] node1319;
	wire [46-1:0] node1322;
	wire [46-1:0] node1325;
	wire [46-1:0] node1326;
	wire [46-1:0] node1329;
	wire [46-1:0] node1332;
	wire [46-1:0] node1333;
	wire [46-1:0] node1334;
	wire [46-1:0] node1337;
	wire [46-1:0] node1340;
	wire [46-1:0] node1341;
	wire [46-1:0] node1344;
	wire [46-1:0] node1347;
	wire [46-1:0] node1348;
	wire [46-1:0] node1349;
	wire [46-1:0] node1350;
	wire [46-1:0] node1351;
	wire [46-1:0] node1354;
	wire [46-1:0] node1357;
	wire [46-1:0] node1358;
	wire [46-1:0] node1361;
	wire [46-1:0] node1364;
	wire [46-1:0] node1365;
	wire [46-1:0] node1366;
	wire [46-1:0] node1369;
	wire [46-1:0] node1372;
	wire [46-1:0] node1373;
	wire [46-1:0] node1376;
	wire [46-1:0] node1379;
	wire [46-1:0] node1380;
	wire [46-1:0] node1381;
	wire [46-1:0] node1382;
	wire [46-1:0] node1385;
	wire [46-1:0] node1388;
	wire [46-1:0] node1389;
	wire [46-1:0] node1392;
	wire [46-1:0] node1395;
	wire [46-1:0] node1396;
	wire [46-1:0] node1397;
	wire [46-1:0] node1400;
	wire [46-1:0] node1403;
	wire [46-1:0] node1404;
	wire [46-1:0] node1407;
	wire [46-1:0] node1410;
	wire [46-1:0] node1411;
	wire [46-1:0] node1412;
	wire [46-1:0] node1413;
	wire [46-1:0] node1414;
	wire [46-1:0] node1415;
	wire [46-1:0] node1418;
	wire [46-1:0] node1423;
	wire [46-1:0] node1424;
	wire [46-1:0] node1425;
	wire [46-1:0] node1426;
	wire [46-1:0] node1429;
	wire [46-1:0] node1432;
	wire [46-1:0] node1433;
	wire [46-1:0] node1436;
	wire [46-1:0] node1439;
	wire [46-1:0] node1440;
	wire [46-1:0] node1441;
	wire [46-1:0] node1444;
	wire [46-1:0] node1448;
	wire [46-1:0] node1449;
	wire [46-1:0] node1450;
	wire [46-1:0] node1451;
	wire [46-1:0] node1452;
	wire [46-1:0] node1455;
	wire [46-1:0] node1458;
	wire [46-1:0] node1459;
	wire [46-1:0] node1462;
	wire [46-1:0] node1465;
	wire [46-1:0] node1466;
	wire [46-1:0] node1467;
	wire [46-1:0] node1470;
	wire [46-1:0] node1474;
	wire [46-1:0] node1475;
	wire [46-1:0] node1476;
	wire [46-1:0] node1477;
	wire [46-1:0] node1480;

	assign outp = (inp[1]) ? node282 : node1;
		assign node1 = (inp[15]) ? node71 : node2;
			assign node2 = (inp[13]) ? node38 : node3;
				assign node3 = (inp[0]) ? node5 : 46'b0000000000000000000000000000000000000000000000;
					assign node5 = (inp[10]) ? node7 : 46'b0000000000000000000000000000000000000000000000;
						assign node7 = (inp[9]) ? node9 : 46'b0000000000000000000000000000000000000000000000;
							assign node9 = (inp[8]) ? node11 : 46'b0000000000000000000000000000000000000000000000;
								assign node11 = (inp[11]) ? node25 : node12;
									assign node12 = (inp[7]) ? node14 : 46'b0000000000000000000000000000000000000000000000;
										assign node14 = (inp[2]) ? node16 : 46'b0000000000000000000000000000000000000000000000;
											assign node16 = (inp[5]) ? node18 : 46'b0000000000000000000000000000000000000000000000;
												assign node18 = (inp[14]) ? node20 : 46'b0000000000000000000000000000000000000000000000;
													assign node20 = (inp[12]) ? node22 : 46'b0000000000000000000000000000000000000000000000;
														assign node22 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
									assign node25 = (inp[3]) ? node27 : 46'b0000000000000000000000000000000000000000000000;
										assign node27 = (inp[7]) ? node29 : 46'b0000000000000000000000000000000000000000000000;
											assign node29 = (inp[12]) ? node31 : 46'b0000000000000000000000000000000000000000000000;
												assign node31 = (inp[4]) ? node33 : 46'b0000000000000000000000000000000000000000000000;
													assign node33 = (inp[14]) ? node35 : 46'b0000000000000000000000000000000000000000000000;
														assign node35 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
				assign node38 = (inp[2]) ? node40 : 46'b0000000000000000000000000000000000000000000000;
					assign node40 = (inp[11]) ? 46'b0000000000000000000000000000000000000000000000 : node41;
						assign node41 = (inp[7]) ? node43 : 46'b0000000000000000000000000000000000000000000000;
							assign node43 = (inp[6]) ? node45 : 46'b0000000000000000000000000000000000000000000000;
								assign node45 = (inp[5]) ? node47 : 46'b0000000000000000000000000000000000000000000000;
									assign node47 = (inp[12]) ? node49 : 46'b0000000000000000000000000000000000000000000000;
										assign node49 = (inp[9]) ? node61 : node50;
											assign node50 = (inp[0]) ? node54 : node51;
												assign node51 = (inp[3]) ? 46'b0000000000000000000000000000000000000100000000 : 46'b0000000000000000000000000000000000000000000000;
												assign node54 = (inp[8]) ? node56 : 46'b0000000000000000000000000000000000000000000000;
													assign node56 = (inp[10]) ? node58 : 46'b0000000000000000000000000000000000000000000000;
														assign node58 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
											assign node61 = (inp[4]) ? node63 : 46'b0000000000000000000000000000000000000000000000;
												assign node63 = (inp[0]) ? node65 : 46'b0000000000000000000000000000000000000000000000;
													assign node65 = (inp[8]) ? node67 : 46'b0000000000000000000000000000000000000000000000;
														assign node67 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
			assign node71 = (inp[3]) ? node73 : 46'b0000000000000000000000000000001000000000000000;
				assign node73 = (inp[9]) ? node137 : node74;
					assign node74 = (inp[11]) ? node124 : node75;
						assign node75 = (inp[2]) ? node101 : node76;
							assign node76 = (inp[13]) ? node80 : node77;
								assign node77 = (inp[0]) ? 46'b0000000000001000000000000010000000000000000000 : 46'b0000001000001000000000000000000000000000000000;
								assign node80 = (inp[5]) ? node82 : 46'b0000000000000000000000000000000000000000000000;
									assign node82 = (inp[6]) ? node84 : 46'b0000000000000000000000000000000000000000000000;
										assign node84 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node85;
											assign node85 = (inp[14]) ? node87 : 46'b0000000000000000000000000000000000000000000000;
												assign node87 = (inp[4]) ? node93 : node88;
													assign node88 = (inp[10]) ? node90 : 46'b0000000000000000000000000000000000000000000000;
														assign node90 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
													assign node93 = (inp[7]) ? node97 : node94;
														assign node94 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
														assign node97 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000001000010100000000000000000000010000;
							assign node101 = (inp[14]) ? node103 : 46'b0000000000000000000000000000000000000000000000;
								assign node103 = (inp[13]) ? node105 : 46'b0000000000000000000000000000000000000000000000;
									assign node105 = (inp[6]) ? node107 : 46'b0000000000000000000000000000000000000000000000;
										assign node107 = (inp[5]) ? node109 : 46'b0000000000000000000000000000000000000000000000;
											assign node109 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node110;
												assign node110 = (inp[8]) ? node116 : node111;
													assign node111 = (inp[10]) ? node113 : 46'b0000000000000000000000000000000000000000000000;
														assign node113 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
													assign node116 = (inp[10]) ? node120 : node117;
														assign node117 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
														assign node120 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
						assign node124 = (inp[13]) ? node130 : node125;
							assign node125 = (inp[2]) ? 46'b0000000000000000000000000000000000000000000000 : node126;
								assign node126 = (inp[0]) ? 46'b0000010000000000000000000010000000000000000000 : 46'b0000011000000000000000000000000000000000000000;
							assign node130 = (inp[2]) ? node134 : node131;
								assign node131 = (inp[0]) ? 46'b0000001000000000011000000100000000000000010000 : 46'b0000001000000000010000000100000000000000010010;
								assign node134 = (inp[0]) ? 46'b0000001000000000010010000000010000000010000000 : 46'b0000001000000000010010100000000000000010000000;
					assign node137 = (inp[2]) ? node227 : node138;
						assign node138 = (inp[0]) ? node178 : node139;
							assign node139 = (inp[13]) ? node143 : node140;
								assign node140 = (inp[11]) ? 46'b0000010100000000000000000000000000000000000000 : 46'b0000000100001000000000000000000000000000000000;
								assign node143 = (inp[5]) ? node145 : 46'b0000000000000000000000000000000000000000000000;
									assign node145 = (inp[14]) ? node147 : 46'b0000000000000000000000000000000000000000000000;
										assign node147 = (inp[6]) ? node157 : node148;
											assign node148 = (inp[11]) ? node150 : 46'b0000000000000000000000000000000000000000000000;
												assign node150 = (inp[10]) ? node152 : 46'b0000000000000000000000000000000000000000000000;
													assign node152 = (inp[4]) ? node154 : 46'b0000000000000000000000000000000000000000000000;
														assign node154 = (inp[8]) ? 46'b0000000000000000000000000100000000000000000010 : 46'b0000000000000000000000000000000000000000000000;
											assign node157 = (inp[4]) ? node165 : node158;
												assign node158 = (inp[10]) ? node160 : 46'b0000000000000000000000000000000000000000000000;
													assign node160 = (inp[8]) ? node162 : 46'b0000000000000000000000000000000000000000000000;
														assign node162 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000010000000000000000010000;
												assign node165 = (inp[7]) ? node173 : node166;
													assign node166 = (inp[12]) ? node170 : node167;
														assign node167 = (inp[11]) ? 46'b0010000000000000000000000100000000000000010010 : 46'b0010000000000000000000000000000000000000010000;
														assign node170 = (inp[10]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
													assign node173 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node174;
														assign node174 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
							assign node178 = (inp[11]) ? node200 : node179;
								assign node179 = (inp[13]) ? node181 : 46'b0010001000000000000000000000000000000000010000;
									assign node181 = (inp[14]) ? node183 : 46'b0000000000000000000000000000000000000000000000;
										assign node183 = (inp[6]) ? node185 : 46'b0000000000000000000000000000000000000000000000;
											assign node185 = (inp[5]) ? node187 : 46'b0000000000000000000000000000000000000000000000;
												assign node187 = (inp[8]) ? node193 : node188;
													assign node188 = (inp[10]) ? node190 : 46'b0000000000000000000000000000000000000000000000;
														assign node190 = (inp[4]) ? 46'b0000000000010000010000000000000000000000010100 : 46'b0000000000000000000000000000000000000000000000;
													assign node193 = (inp[12]) ? node197 : node194;
														assign node194 = (inp[7]) ? 46'b0000000000001000010000000000000000000000010100 : 46'b0000000000000000000000000000000000000000000000;
														assign node197 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000010000000000010000000000000000000000010100;
								assign node200 = (inp[5]) ? node202 : 46'b0000000000000000000000000000000000000000000000;
									assign node202 = (inp[14]) ? node204 : 46'b0000000000000000000000000000000000000000000000;
										assign node204 = (inp[13]) ? node206 : 46'b0000000000000000000000000000000000000000000000;
											assign node206 = (inp[6]) ? node214 : node207;
												assign node207 = (inp[4]) ? node209 : 46'b0000000000000000000000000000000000000000000000;
													assign node209 = (inp[10]) ? node211 : 46'b0000000000000000000000000000000000000000000000;
														assign node211 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
												assign node214 = (inp[10]) ? node220 : node215;
													assign node215 = (inp[4]) ? node217 : 46'b0000000000000000000000000000000000000000000000;
														assign node217 = (inp[8]) ? 46'b0000000000000000001000000100000100000000010000 : 46'b0000000000000000000000000000000000000000000000;
													assign node220 = (inp[8]) ? node224 : node221;
														assign node221 = (inp[4]) ? 46'b0000000000010000001000000100000000000000010000 : 46'b0000000000000000000000000000000000000000000000;
														assign node224 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000011000010100000000000000010000;
						assign node227 = (inp[14]) ? node229 : 46'b0000000000000000000000000000000000000000000000;
							assign node229 = (inp[13]) ? node231 : 46'b0000000000000000000000000000000000000000000000;
								assign node231 = (inp[5]) ? node233 : 46'b0000000000000000000000000000000000000000000000;
									assign node233 = (inp[6]) ? node245 : node234;
										assign node234 = (inp[11]) ? node236 : 46'b0000000000000000000000000000000000000000000000;
											assign node236 = (inp[4]) ? node238 : 46'b0000000000000000000000000000000000000000000000;
												assign node238 = (inp[10]) ? node240 : 46'b0000000000000000000000000000000000000000000000;
													assign node240 = (inp[8]) ? node242 : 46'b0000000000000000000000000000000000000000000000;
														assign node242 = (inp[0]) ? 46'b0000000000000000000010000000010000000000000000 : 46'b0000000000000000000010100000000000000000000000;
										assign node245 = (inp[11]) ? node261 : node246;
											assign node246 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node247;
												assign node247 = (inp[10]) ? node253 : node248;
													assign node248 = (inp[8]) ? node250 : 46'b0000000000000000000000000000000000000000000000;
														assign node250 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
													assign node253 = (inp[7]) ? node257 : node254;
														assign node254 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000010000000000000010000000;
														assign node257 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
											assign node261 = (inp[4]) ? node269 : node262;
												assign node262 = (inp[10]) ? node264 : 46'b0000000000000000000000000000000000000000000000;
													assign node264 = (inp[8]) ? node266 : 46'b0000000000000000000000000000000000000000000000;
														assign node266 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000001000010010010000010000000010000000;
												assign node269 = (inp[12]) ? node277 : node270;
													assign node270 = (inp[7]) ? node274 : node271;
														assign node271 = (inp[10]) ? 46'b0010000000010000000010000000000000000010000000 : 46'b0000000000000000000000000000000000000000000000;
														assign node274 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
													assign node277 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node278;
														assign node278 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
		assign node282 = (inp[15]) ? node350 : node283;
			assign node283 = (inp[13]) ? node287 : node284;
				assign node284 = (inp[3]) ? 46'b0000100000000000000000000000001000000000000000 : 46'b0000100000000000000000000000000000000000000000;
				assign node287 = (inp[2]) ? node319 : node288;
					assign node288 = (inp[11]) ? node304 : node289;
						assign node289 = (inp[0]) ? node297 : node290;
							assign node290 = (inp[9]) ? node294 : node291;
								assign node291 = (inp[3]) ? 46'b0000100000001000010000010100001000000000010010 : 46'b0000100000001000010000010100000000000000010010;
								assign node294 = (inp[3]) ? 46'b0000110000000000010000010100001000000000010010 : 46'b0000110000000000010000010100000000000000010010;
							assign node297 = (inp[9]) ? node301 : node298;
								assign node298 = (inp[3]) ? 46'b0000100000001000010000000100001100000000010010 : 46'b0000100000001000010000000100000100000000010010;
								assign node301 = (inp[3]) ? 46'b0000110000000000010000000100001100000000010010 : 46'b0000110000000000010000000100000100000000010010;
						assign node304 = (inp[0]) ? node312 : node305;
							assign node305 = (inp[9]) ? node309 : node306;
								assign node306 = (inp[3]) ? 46'b0000100000001000011000010100001000000000010000 : 46'b0000100000001000011000010100000000000000010000;
								assign node309 = (inp[3]) ? 46'b0000110000000000011000010100001000000000010000 : 46'b0000110000000000011000010100000000000000010000;
							assign node312 = (inp[9]) ? node316 : node313;
								assign node313 = (inp[3]) ? 46'b0000100000001000011000000100001100000000010000 : 46'b0000100000001000011000000100000100000000010000;
								assign node316 = (inp[3]) ? 46'b0000110000000000011000000100001100000000010000 : 46'b0000110000000000011000000100000100000000010000;
					assign node319 = (inp[9]) ? node335 : node320;
						assign node320 = (inp[0]) ? node328 : node321;
							assign node321 = (inp[11]) ? node325 : node322;
								assign node322 = (inp[3]) ? 46'b0000100000001000010010110000001000000010000000 : 46'b0000100000001000010010110000000000000010000000;
								assign node325 = (inp[3]) ? 46'b0000100000001000010010010000011000000010000000 : 46'b0000100000001000010010010000010000000010000000;
							assign node328 = (inp[11]) ? node332 : node329;
								assign node329 = (inp[3]) ? 46'b0000100000001000010010100000001100000010000000 : 46'b0000100000001000010010100000000100000010000000;
								assign node332 = (inp[3]) ? 46'b0000100000001000010010000000011100000010000000 : 46'b0000100000001000010010000000010100000010000000;
						assign node335 = (inp[11]) ? node343 : node336;
							assign node336 = (inp[0]) ? node340 : node337;
								assign node337 = (inp[3]) ? 46'b0000110000000000010010110000001000000010000000 : 46'b0000110000000000010010110000000000000010000000;
								assign node340 = (inp[3]) ? 46'b0000110000000000010010100000001100000010000000 : 46'b0000110000000000010010100000000100000010000000;
							assign node343 = (inp[0]) ? node347 : node344;
								assign node344 = (inp[3]) ? 46'b0000110000000000010010010000011000000010000000 : 46'b0000110000000000010010010000010000000010000000;
								assign node347 = (inp[3]) ? 46'b0000110000000000010010000000011100000010000000 : 46'b0000110000000000010010000000010100000010000000;
			assign node350 = (inp[13]) ? node354 : node351;
				assign node351 = (inp[3]) ? 46'b0000000000000000000000000000000000000000001000 : 46'b0000000000000000000000000000001000000000001000;
				assign node354 = (inp[3]) ? node356 : 46'b0000000000000000000000000000001000000000000000;
					assign node356 = (inp[2]) ? node1072 : node357;
						assign node357 = (inp[9]) ? node765 : node358;
							assign node358 = (inp[11]) ? node614 : node359;
								assign node359 = (inp[7]) ? node487 : node360;
									assign node360 = (inp[6]) ? node424 : node361;
										assign node361 = (inp[12]) ? node393 : node362;
											assign node362 = (inp[0]) ? node378 : node363;
												assign node363 = (inp[5]) ? node371 : node364;
													assign node364 = (inp[8]) ? node368 : node365;
														assign node365 = (inp[14]) ? 46'b0011000000000000001000010001100010110001010000 : 46'b0011000000000100000000010000100010110001010000;
														assign node368 = (inp[14]) ? 46'b0011000000000010000000010000100010110001010000 : 46'b0011000000000000000000010001100010110001010010;
													assign node371 = (inp[8]) ? node375 : node372;
														assign node372 = (inp[14]) ? 46'b0010000000000000001000010001100010110001010000 : 46'b0010000000000100000000010000100010110001010000;
														assign node375 = (inp[14]) ? 46'b0010000000000010000000010001100010110001010000 : 46'b0010000000000000000000010001100010110001010010;
												assign node378 = (inp[5]) ? node386 : node379;
													assign node379 = (inp[4]) ? node383 : node380;
														assign node380 = (inp[10]) ? 46'b0011000000000000000000010001100010110000010010 : 46'b0011000000000100000000010000100010110000010000;
														assign node383 = (inp[10]) ? 46'b0011000000000010000000010000100010110000010000 : 46'b0011000000000000001000010001100010110000010000;
													assign node386 = (inp[14]) ? node390 : node387;
														assign node387 = (inp[8]) ? 46'b0010000000000000000000010001100010110000010010 : 46'b0010000000000100000000010000100010110000010000;
														assign node390 = (inp[4]) ? 46'b0010000000000010001000010001100010110000010000 : 46'b0010000000000000000000010001100010110000010010;
											assign node393 = (inp[5]) ? node409 : node394;
												assign node394 = (inp[0]) ? node402 : node395;
													assign node395 = (inp[4]) ? node399 : node396;
														assign node396 = (inp[10]) ? 46'b0011000000000000000000010001100000110001010010 : 46'b0011000000000100000000010001100000110001010000;
														assign node399 = (inp[10]) ? 46'b0011000000000010000000010000100000110001010000 : 46'b0011000000000000001000010001100000110001010000;
													assign node402 = (inp[4]) ? node406 : node403;
														assign node403 = (inp[10]) ? 46'b0011000000000000000000010001100000110000010010 : 46'b0011000000000100000000010001100000110000010000;
														assign node406 = (inp[10]) ? 46'b0011000000000010000000010000100000110000010000 : 46'b0011000000000000001000010001100000110000010000;
												assign node409 = (inp[0]) ? node417 : node410;
													assign node410 = (inp[8]) ? node414 : node411;
														assign node411 = (inp[14]) ? 46'b0010000000000000001000010001100000110001010000 : 46'b0010000000000100000000010000100000110001010000;
														assign node414 = (inp[10]) ? 46'b0010000000000010000000010001100000110001010010 : 46'b0010000000000000001000010001100000110001010010;
													assign node417 = (inp[14]) ? node421 : node418;
														assign node418 = (inp[8]) ? 46'b0010000000000000000000010001100000110000010010 : 46'b0010000000000100000000010000100000110000010000;
														assign node421 = (inp[8]) ? 46'b0010000000000010000000010000100000110000010000 : 46'b0010000000000000001000010001100000110000010000;
										assign node424 = (inp[5]) ? node456 : node425;
											assign node425 = (inp[0]) ? node441 : node426;
												assign node426 = (inp[12]) ? node434 : node427;
													assign node427 = (inp[14]) ? node431 : node428;
														assign node428 = (inp[8]) ? 46'b0011000000000000000000010001100010010001010010 : 46'b0011000000000100000000010000100010010001010000;
														assign node431 = (inp[8]) ? 46'b0011000000000010000000010000100010010001010000 : 46'b0011000000000000001000010001100010010001010000;
													assign node434 = (inp[8]) ? node438 : node435;
														assign node435 = (inp[14]) ? 46'b0011000000000000001000010001100000010001010000 : 46'b0011000000000100000000010001100000010001010000;
														assign node438 = (inp[14]) ? 46'b0011000000000010000000010000100000010001010000 : 46'b0011000000000000000000010001100000010001010010;
												assign node441 = (inp[12]) ? node449 : node442;
													assign node442 = (inp[8]) ? node446 : node443;
														assign node443 = (inp[14]) ? 46'b0011000000000000001000010001100010010000010000 : 46'b0011000000000100000000010000100010010000010000;
														assign node446 = (inp[14]) ? 46'b0011000000000010000000010000100010010000010000 : 46'b0011000000000000000000010001100010010000010010;
													assign node449 = (inp[14]) ? node453 : node450;
														assign node450 = (inp[8]) ? 46'b0011000000000000000000010001100000010000010010 : 46'b0011000000000100000000010000100000010000010000;
														assign node453 = (inp[8]) ? 46'b0011000000000010000000010000100000010000010000 : 46'b0011000000000000001000010001100000010000010000;
											assign node456 = (inp[12]) ? node472 : node457;
												assign node457 = (inp[0]) ? node465 : node458;
													assign node458 = (inp[4]) ? node462 : node459;
														assign node459 = (inp[10]) ? 46'b0010000000000000000000010001100010010001010010 : 46'b0010000000000100000000010000100010010001010000;
														assign node462 = (inp[10]) ? 46'b0010000000000010000000010000100010010001010000 : 46'b0010000000000000001000010001100010010001010000;
													assign node465 = (inp[4]) ? node469 : node466;
														assign node466 = (inp[10]) ? 46'b0010000000000000000000010001100010010000010010 : 46'b0010000000000100000000010000100010010000010000;
														assign node469 = (inp[10]) ? 46'b0010000000000010000000010000100010010000010000 : 46'b0010000000000000001000010001100010010000010000;
												assign node472 = (inp[0]) ? node480 : node473;
													assign node473 = (inp[10]) ? node477 : node474;
														assign node474 = (inp[4]) ? 46'b0010000000000000001000010001100000010001010000 : 46'b0010000000000100000000010000100000010001010000;
														assign node477 = (inp[4]) ? 46'b0010000000000010000000010000100000010001010000 : 46'b0010000000000000000000010001100000010001010010;
													assign node480 = (inp[8]) ? node484 : node481;
														assign node481 = (inp[14]) ? 46'b0010000000000000001000010001100000010000010000 : 46'b0010000000000100000000010000100000010000010000;
														assign node484 = (inp[14]) ? 46'b0010000000000010000000010000100000010000010000 : 46'b0010000000000000000000010001100000010000010010;
									assign node487 = (inp[12]) ? node551 : node488;
										assign node488 = (inp[6]) ? node520 : node489;
											assign node489 = (inp[5]) ? node505 : node490;
												assign node490 = (inp[0]) ? node498 : node491;
													assign node491 = (inp[4]) ? node495 : node492;
														assign node492 = (inp[10]) ? 46'b0011000000000000000000010001000010110001010010 : 46'b0011000000000100000000010000000010110001010000;
														assign node495 = (inp[10]) ? 46'b0011000000000010000000010000000010110001010000 : 46'b0011000000000000001000010001000010110001010000;
													assign node498 = (inp[8]) ? node502 : node499;
														assign node499 = (inp[14]) ? 46'b0011000000000000001000010001000010110000010000 : 46'b0011000000000100000000010001000010110000010000;
														assign node502 = (inp[10]) ? 46'b0011000000000010000000010001000010110000010010 : 46'b0011000000000110000000010000000010110000010000;
												assign node505 = (inp[0]) ? node513 : node506;
													assign node506 = (inp[8]) ? node510 : node507;
														assign node507 = (inp[14]) ? 46'b0010000000000000001000010001000010110001010000 : 46'b0010000000000100000000010000000010110001010000;
														assign node510 = (inp[14]) ? 46'b0010000000000010000000010000000010110001010000 : 46'b0010000000000000000000010001000010110001010010;
													assign node513 = (inp[14]) ? node517 : node514;
														assign node514 = (inp[8]) ? 46'b0010000000000000000000010001000010110000010010 : 46'b0010000000000100000000010000000010110000010000;
														assign node517 = (inp[8]) ? 46'b0010000000000010000000010000000010110000010000 : 46'b0010000000000000001000010001000010110000010000;
											assign node520 = (inp[5]) ? node536 : node521;
												assign node521 = (inp[0]) ? node529 : node522;
													assign node522 = (inp[14]) ? node526 : node523;
														assign node523 = (inp[8]) ? 46'b0011000000000000000000010001000010010001010010 : 46'b0011000000000100000000010000000010010001010000;
														assign node526 = (inp[8]) ? 46'b0011000000000010000000010000000010010001010000 : 46'b0011000000000000001000010001000010010001010000;
													assign node529 = (inp[8]) ? node533 : node530;
														assign node530 = (inp[14]) ? 46'b0011000000000000001000010001000010010000010000 : 46'b0011000000000100000000010000000010010000010000;
														assign node533 = (inp[14]) ? 46'b0011000000000010000000010001000010010000010000 : 46'b0011000000000000000000010001000010010000010010;
												assign node536 = (inp[0]) ? node544 : node537;
													assign node537 = (inp[8]) ? node541 : node538;
														assign node538 = (inp[14]) ? 46'b0010000000000000001000010001000010010001010000 : 46'b0010000000000100000000010000000010010001010000;
														assign node541 = (inp[14]) ? 46'b0010000000000010000000010000000010010001010000 : 46'b0010000000000000000000010001000010010001010010;
													assign node544 = (inp[14]) ? node548 : node545;
														assign node545 = (inp[8]) ? 46'b0010000000000000000000010001000010010000010010 : 46'b0010000000000100000000010000000010010000010000;
														assign node548 = (inp[8]) ? 46'b0010000000000010000000010001000010010000010000 : 46'b0010000000000000001000010001000010010000010000;
										assign node551 = (inp[0]) ? node583 : node552;
											assign node552 = (inp[5]) ? node568 : node553;
												assign node553 = (inp[6]) ? node561 : node554;
													assign node554 = (inp[4]) ? node558 : node555;
														assign node555 = (inp[10]) ? 46'b0011000000000000000000010001000000110001010010 : 46'b0011000000000100000000010000000000110001010000;
														assign node558 = (inp[10]) ? 46'b0011000000000010000000010000000000110001010000 : 46'b0011000000000000001000010001000000110001010000;
													assign node561 = (inp[14]) ? node565 : node562;
														assign node562 = (inp[8]) ? 46'b0011000000000000000000010001000000010001010010 : 46'b0011000000000100000000010000000000010001010000;
														assign node565 = (inp[8]) ? 46'b0011000000000010000000010000000000010001010000 : 46'b0011000000000000001000010001000000010001010000;
												assign node568 = (inp[6]) ? node576 : node569;
													assign node569 = (inp[14]) ? node573 : node570;
														assign node570 = (inp[8]) ? 46'b0010000000000000000000010001000000110001010010 : 46'b0010000000000100000000010000000000110001010000;
														assign node573 = (inp[8]) ? 46'b0010000000000010000000010000000000110001010000 : 46'b0010000000000000001000010001000000110001010000;
													assign node576 = (inp[8]) ? node580 : node577;
														assign node577 = (inp[14]) ? 46'b0010000000000000001000010001000000010001010000 : 46'b0010000000000100000000010000000000010001010000;
														assign node580 = (inp[14]) ? 46'b0010000000000010000000010000000000010001010000 : 46'b0010000000000000000000010001000000010001010010;
											assign node583 = (inp[6]) ? node599 : node584;
												assign node584 = (inp[5]) ? node592 : node585;
													assign node585 = (inp[4]) ? node589 : node586;
														assign node586 = (inp[10]) ? 46'b0011000000000000000000010001000000110000010010 : 46'b0011000000000100000000010000000000110000010000;
														assign node589 = (inp[10]) ? 46'b0011000000000010000000010000000000110000010000 : 46'b0011000000000000001000010001000000110000010000;
													assign node592 = (inp[4]) ? node596 : node593;
														assign node593 = (inp[10]) ? 46'b0010000000000000000000010001000000110000010010 : 46'b0010000000000100000000010000000000110000010000;
														assign node596 = (inp[10]) ? 46'b0010000000000010000000010000000000110000010000 : 46'b0010000000000000001000010001000000110000010000;
												assign node599 = (inp[5]) ? node607 : node600;
													assign node600 = (inp[10]) ? node604 : node601;
														assign node601 = (inp[4]) ? 46'b0011000000000000001000010001000000010000010000 : 46'b0011000000000100000000010000000000010000010000;
														assign node604 = (inp[8]) ? 46'b0011000000000010000000010001000000010000010010 : 46'b0011000000000000001000010001000000010000010010;
													assign node607 = (inp[14]) ? node611 : node608;
														assign node608 = (inp[8]) ? 46'b0010000000000000000000010001000000010000010010 : 46'b0010000000000100000000010000000000010000010000;
														assign node611 = (inp[8]) ? 46'b0010000000000010000000010000000000010000010000 : 46'b0010000000000000001000010001000000010000010000;
								assign node614 = (inp[0]) ? node638 : node615;
									assign node615 = (inp[5]) ? node617 : 46'b0000000000000000000000000000000000000000000000;
										assign node617 = (inp[7]) ? node619 : 46'b0000000000000000000000000000000000000000000000;
											assign node619 = (inp[6]) ? node629 : node620;
												assign node620 = (inp[12]) ? node622 : 46'b0000000000000000000000000000000000000000000000;
													assign node622 = (inp[4]) ? node626 : node623;
														assign node623 = (inp[10]) ? 46'b0000000000000000000001000001000000100000000010 : 46'b0000000000000100000001000000000000100000000000;
														assign node626 = (inp[10]) ? 46'b0000000000000010000001000000000000100000000000 : 46'b0000000000000000001001000001000000100000000000;
												assign node629 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node630;
													assign node630 = (inp[10]) ? node634 : node631;
														assign node631 = (inp[4]) ? 46'b0000000000000000001001000001000010000000000000 : 46'b0000000000000100000001000000000010000000000000;
														assign node634 = (inp[4]) ? 46'b0000000000000010000001000000000010000000000000 : 46'b0000000000000000000001000001000010000000000010;
									assign node638 = (inp[6]) ? node702 : node639;
										assign node639 = (inp[7]) ? node671 : node640;
											assign node640 = (inp[5]) ? node656 : node641;
												assign node641 = (inp[12]) ? node649 : node642;
													assign node642 = (inp[8]) ? node646 : node643;
														assign node643 = (inp[14]) ? 46'b0101000000000000001000000001100010100000000000 : 46'b0101000000000100000000000000100010100000000000;
														assign node646 = (inp[14]) ? 46'b0101000000000010000000000000100010100000000000 : 46'b0101000000000000000000000001100010100000000010;
													assign node649 = (inp[8]) ? node653 : node650;
														assign node650 = (inp[14]) ? 46'b0101000000000000001000000001100000100000000000 : 46'b0101000000000100000000000001100000100000000000;
														assign node653 = (inp[14]) ? 46'b0101000000000010000000000000100000100000000000 : 46'b0101000000000000000000000001100000100000000010;
												assign node656 = (inp[12]) ? node664 : node657;
													assign node657 = (inp[4]) ? node661 : node658;
														assign node658 = (inp[10]) ? 46'b0100000000000000000000000001100010100000000010 : 46'b0100000000000100000000000000100010100000000000;
														assign node661 = (inp[10]) ? 46'b0100000000000010000000000000100010100000000000 : 46'b0100000000000000001000000001100010100000000000;
													assign node664 = (inp[8]) ? node668 : node665;
														assign node665 = (inp[14]) ? 46'b0100000000000000001000000001100000100000000000 : 46'b0100000000000100000000000001100000100000000000;
														assign node668 = (inp[14]) ? 46'b0100000000000010000000000000100000100000000000 : 46'b0100000000000000000000000001100000100000000010;
											assign node671 = (inp[5]) ? node687 : node672;
												assign node672 = (inp[12]) ? node680 : node673;
													assign node673 = (inp[14]) ? node677 : node674;
														assign node674 = (inp[8]) ? 46'b0101000000000000000000000001000010100000000010 : 46'b0101000000000100000000000000000010100000000000;
														assign node677 = (inp[8]) ? 46'b0101000000000010000000000000000010100000000000 : 46'b0101000000000000001000000001000010100000000000;
													assign node680 = (inp[8]) ? node684 : node681;
														assign node681 = (inp[14]) ? 46'b0101000000000000001000000001000000100000000000 : 46'b0101000000000100000000000000000000100000000000;
														assign node684 = (inp[14]) ? 46'b0101000000000010000000000000000000100000000000 : 46'b0101000000000000000000000001000000100000000010;
												assign node687 = (inp[12]) ? node695 : node688;
													assign node688 = (inp[8]) ? node692 : node689;
														assign node689 = (inp[14]) ? 46'b0100000000000000001000000001000010100000000000 : 46'b0100000000000100000000000001000010100000000000;
														assign node692 = (inp[14]) ? 46'b0100000000000010000000000000000010100000000000 : 46'b0100000000000000000000000001000010100000000010;
													assign node695 = (inp[8]) ? node699 : node696;
														assign node696 = (inp[14]) ? 46'b0100000000000000001000000001000000100000000000 : 46'b0100000000000100000000000000000000100000000000;
														assign node699 = (inp[14]) ? 46'b0100000000000010000000000000000000100000000000 : 46'b0100000000000000000000000001000000100000000010;
										assign node702 = (inp[5]) ? node734 : node703;
											assign node703 = (inp[7]) ? node719 : node704;
												assign node704 = (inp[12]) ? node712 : node705;
													assign node705 = (inp[4]) ? node709 : node706;
														assign node706 = (inp[10]) ? 46'b0101000000000000000000000001100010000000000010 : 46'b0101000000000100000000000000100010000000000000;
														assign node709 = (inp[10]) ? 46'b0101000000000010000000000001100010000000000000 : 46'b0101000000000000001000000001100010000000000000;
													assign node712 = (inp[8]) ? node716 : node713;
														assign node713 = (inp[14]) ? 46'b0101000000000000001000000001100000000000000000 : 46'b0101000000000100000000000000100000000000000000;
														assign node716 = (inp[14]) ? 46'b0101000000000010000000000000100000000000000000 : 46'b0101000000000000000000000001100000000000000010;
												assign node719 = (inp[12]) ? node727 : node720;
													assign node720 = (inp[14]) ? node724 : node721;
														assign node721 = (inp[8]) ? 46'b0101000000000000000000000001000010000000000010 : 46'b0101000000000100000000000000000010000000000000;
														assign node724 = (inp[8]) ? 46'b0101000000000010000000000000000010000000000000 : 46'b0101000000000000001000000001000010000000000000;
													assign node727 = (inp[4]) ? node731 : node728;
														assign node728 = (inp[14]) ? 46'b0101000000000000001000000001000000000000000000 : 46'b0101000000000100000000000001000000000000000010;
														assign node731 = (inp[10]) ? 46'b0101000000000010000000000000000000000000000000 : 46'b0101000000000000001000000001000000000000000000;
											assign node734 = (inp[12]) ? node750 : node735;
												assign node735 = (inp[7]) ? node743 : node736;
													assign node736 = (inp[8]) ? node740 : node737;
														assign node737 = (inp[14]) ? 46'b0100000000000000001000000001100010000000000000 : 46'b0100000000000100000000000000100010000000000000;
														assign node740 = (inp[14]) ? 46'b0100000000000010000000000000100010000000000000 : 46'b0100000000000000000000000001100010000000000010;
													assign node743 = (inp[4]) ? node747 : node744;
														assign node744 = (inp[10]) ? 46'b0100000000000000000000000001000010000000000010 : 46'b0100000000000100000000000000000010000000000000;
														assign node747 = (inp[14]) ? 46'b0100000000000010001000000001000010000000000000 : 46'b0100000000000100000000000000000010000000000000;
												assign node750 = (inp[7]) ? node758 : node751;
													assign node751 = (inp[14]) ? node755 : node752;
														assign node752 = (inp[8]) ? 46'b0100000000000000000000000001100000000000000010 : 46'b0100000000000100000000000000100000000000000000;
														assign node755 = (inp[8]) ? 46'b0100000000000010000000000000100000000000000000 : 46'b0100000000000000001000000001100000000000000000;
													assign node758 = (inp[10]) ? node762 : node759;
														assign node759 = (inp[4]) ? 46'b0100000000000000001000000001000000000000000000 : 46'b0100000000000100000000000001000000000000000000;
														assign node762 = (inp[4]) ? 46'b0100000000000010000000000000000000000000000000 : 46'b0100000000000000000000000001000000000000000010;
							assign node765 = (inp[11]) ? node817 : node766;
								assign node766 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node767;
									assign node767 = (inp[4]) ? node799 : node768;
										assign node768 = (inp[5]) ? node784 : node769;
											assign node769 = (inp[7]) ? node771 : 46'b0000000000000000000000000000000000000000000000;
												assign node771 = (inp[10]) ? node779 : node772;
													assign node772 = (inp[6]) ? node776 : node773;
														assign node773 = (inp[12]) ? 46'b0001000000000100000000001000000000100000000000 : 46'b0001000000000100000000001000000010100000000000;
														assign node776 = (inp[12]) ? 46'b0001000000000100000000001000000000000000000000 : 46'b0001000000000100000000001000000010000000000000;
													assign node779 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : node780;
														assign node780 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000000100000000001001000000000000000010;
											assign node784 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node785;
												assign node785 = (inp[10]) ? node791 : node786;
													assign node786 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : node787;
														assign node787 = (inp[8]) ? 46'b0000000000000100000000001001100000000000000010 : 46'b0000000000000000000000000000000000000000000000;
													assign node791 = (inp[6]) ? node795 : node792;
														assign node792 = (inp[12]) ? 46'b0000000000000000000000001001100000100000000010 : 46'b0000000000000000000000001001100010100000000010;
														assign node795 = (inp[12]) ? 46'b0000000000000000000000001001100000000000000010 : 46'b0000000000000000000000001001100010000000000010;
										assign node799 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : node800;
											assign node800 = (inp[8]) ? node808 : node801;
												assign node801 = (inp[7]) ? node803 : 46'b0000000000000000000000000000000000000000000000;
													assign node803 = (inp[5]) ? 46'b0000000000000000000000000000000000000000000000 : node804;
														assign node804 = (inp[10]) ? 46'b0001000000000110000000001000000000000000000000 : 46'b0001000000000100001000001001000000000000000000;
												assign node808 = (inp[5]) ? node810 : 46'b0000000000000000000000000000000000000000000000;
													assign node810 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node811;
														assign node811 = (inp[10]) ? 46'b0000000000000010000000001001100000000000000010 : 46'b0000000000000000001000001001100000000000000010;
								assign node817 = (inp[0]) ? node945 : node818;
									assign node818 = (inp[12]) ? node882 : node819;
										assign node819 = (inp[7]) ? node851 : node820;
											assign node820 = (inp[5]) ? node836 : node821;
												assign node821 = (inp[6]) ? node829 : node822;
													assign node822 = (inp[10]) ? node826 : node823;
														assign node823 = (inp[4]) ? 46'b1001000000000000001000000001100010100000000000 : 46'b1001000000000100000000000000100010100000000000;
														assign node826 = (inp[4]) ? 46'b1001000000000010000000000000100010100000000000 : 46'b1001000000000000000000000001100010100000000010;
													assign node829 = (inp[10]) ? node833 : node830;
														assign node830 = (inp[4]) ? 46'b1001000000000000001000000001100010000000000000 : 46'b1001000000000100000000000000100010000000000000;
														assign node833 = (inp[4]) ? 46'b1001000000000010000000000001100010000000000000 : 46'b1001000000000000000000000001100010000000000010;
												assign node836 = (inp[6]) ? node844 : node837;
													assign node837 = (inp[8]) ? node841 : node838;
														assign node838 = (inp[14]) ? 46'b1000000000000000001000000001100010100000000000 : 46'b1000000000000100000000000000100010100000000000;
														assign node841 = (inp[14]) ? 46'b1000000000000010000000000001100010100000000000 : 46'b1000000000000000000000000001100010100000000010;
													assign node844 = (inp[14]) ? node848 : node845;
														assign node845 = (inp[8]) ? 46'b1000000000000000000000000001100010000000000010 : 46'b1000000000000100000000000000100010000000000000;
														assign node848 = (inp[8]) ? 46'b1000000000000010000000000000100010000000000000 : 46'b1000000000000000001000000001100010000000000000;
											assign node851 = (inp[5]) ? node867 : node852;
												assign node852 = (inp[6]) ? node860 : node853;
													assign node853 = (inp[4]) ? node857 : node854;
														assign node854 = (inp[10]) ? 46'b1001000000000000000000000001000010100000000010 : 46'b1001000000000100000000000001000010100000000000;
														assign node857 = (inp[10]) ? 46'b1001000000000010000000000000000010100000000000 : 46'b1001000000000000001000000001000010100000000000;
													assign node860 = (inp[8]) ? node864 : node861;
														assign node861 = (inp[14]) ? 46'b1001000000000000001000000001000010000000000000 : 46'b1001000000000100000000000000000010000000000000;
														assign node864 = (inp[14]) ? 46'b1001000000000010000000000001000010000000000000 : 46'b1001000000000000000000000001000010000000000010;
												assign node867 = (inp[6]) ? node875 : node868;
													assign node868 = (inp[4]) ? node872 : node869;
														assign node869 = (inp[10]) ? 46'b1000000000000000000000000001000010100000000010 : 46'b1000000000000100000000000000000010100000000000;
														assign node872 = (inp[10]) ? 46'b1000000000000010000000000000000010100000000000 : 46'b1000000000000000001000000001000010100000000000;
													assign node875 = (inp[14]) ? node879 : node876;
														assign node876 = (inp[8]) ? 46'b1000000000000000000000000001000010000000000010 : 46'b1000000000000100000000000000000010000000000000;
														assign node879 = (inp[8]) ? 46'b1000000000000010000000000000000010000000000000 : 46'b1000000000000000001000000001000010000000000000;
										assign node882 = (inp[7]) ? node914 : node883;
											assign node883 = (inp[6]) ? node899 : node884;
												assign node884 = (inp[5]) ? node892 : node885;
													assign node885 = (inp[4]) ? node889 : node886;
														assign node886 = (inp[14]) ? 46'b1001000000000000000000000001100000100000000010 : 46'b1001000000000100000000000001100000100000000010;
														assign node889 = (inp[10]) ? 46'b1001000000000010000000000001100000100000000000 : 46'b1001000000000000001000000001100000100000000000;
													assign node892 = (inp[10]) ? node896 : node893;
														assign node893 = (inp[8]) ? 46'b1000000000000000001000000001100000100000000010 : 46'b1000000000000100001000000001100000100000000000;
														assign node896 = (inp[4]) ? 46'b1000000000000010000000000000100000100000000000 : 46'b1000000000000000000000000001100000100000000010;
												assign node899 = (inp[5]) ? node907 : node900;
													assign node900 = (inp[8]) ? node904 : node901;
														assign node901 = (inp[14]) ? 46'b1001000000000000001000000001100000000000000000 : 46'b1001000000000100000000000000100000000000000000;
														assign node904 = (inp[14]) ? 46'b1001000000000010000000000000100000000000000000 : 46'b1001000000000000000000000001100000000000000010;
													assign node907 = (inp[14]) ? node911 : node908;
														assign node908 = (inp[8]) ? 46'b1000000000000000000000000001100000000000000010 : 46'b1000000000000100000000000000100000000000000000;
														assign node911 = (inp[8]) ? 46'b1000000000000010000000000000100000000000000000 : 46'b1000000000000000001000000001100000000000000000;
											assign node914 = (inp[5]) ? node930 : node915;
												assign node915 = (inp[6]) ? node923 : node916;
													assign node916 = (inp[4]) ? node920 : node917;
														assign node917 = (inp[10]) ? 46'b1001000000000000000000000001000000100000000010 : 46'b1001000000000100000000000000000000100000000000;
														assign node920 = (inp[10]) ? 46'b1001000000000010000000000000000000100000000000 : 46'b1001000000000000001000000001000000100000000000;
													assign node923 = (inp[10]) ? node927 : node924;
														assign node924 = (inp[8]) ? 46'b1001000000000000000000000001000000000000000010 : 46'b1001000000000100001000000001000000000000000000;
														assign node927 = (inp[4]) ? 46'b1001000000000010000000000000000000000000000000 : 46'b1001000000000000000000000001000000000000000010;
												assign node930 = (inp[6]) ? node938 : node931;
													assign node931 = (inp[10]) ? node935 : node932;
														assign node932 = (inp[4]) ? 46'b1000000000000000001000000001000000100000000000 : 46'b1000000000000100000000000000000000100000000000;
														assign node935 = (inp[4]) ? 46'b1000000000000010000000000000000000100000000000 : 46'b1000000000000000000000000001000000100000000010;
													assign node938 = (inp[10]) ? node942 : node939;
														assign node939 = (inp[4]) ? 46'b1000000000000000001000000001000000000000000000 : 46'b1000000000000100000000000000000000000000000000;
														assign node942 = (inp[4]) ? 46'b1000000000000010000000000000000000000000000000 : 46'b1000000000000000000000000001000000000000000010;
									assign node945 = (inp[12]) ? node1009 : node946;
										assign node946 = (inp[5]) ? node978 : node947;
											assign node947 = (inp[6]) ? node963 : node948;
												assign node948 = (inp[7]) ? node956 : node949;
													assign node949 = (inp[4]) ? node953 : node950;
														assign node950 = (inp[10]) ? 46'b0001000000000000000000000001100010101000000010 : 46'b0001000000000100000000000000100010101000000000;
														assign node953 = (inp[10]) ? 46'b0001000000000010000000000000100010101000000000 : 46'b0001000000000000001000000001100010101000000000;
													assign node956 = (inp[14]) ? node960 : node957;
														assign node957 = (inp[8]) ? 46'b0001000000000000000000000001000010101000000010 : 46'b0001000000000100000000000000000010101000000000;
														assign node960 = (inp[8]) ? 46'b0001000000000010000000000000000010101000000000 : 46'b0001000000000000001000000001000010101000000000;
												assign node963 = (inp[7]) ? node971 : node964;
													assign node964 = (inp[4]) ? node968 : node965;
														assign node965 = (inp[10]) ? 46'b0001000000000000000000000001100010001000000010 : 46'b0001000000000100000000000001100010001000000000;
														assign node968 = (inp[10]) ? 46'b0001000000000010000000000000100010001000000000 : 46'b0001000000000000001000000001100010001000000000;
													assign node971 = (inp[4]) ? node975 : node972;
														assign node972 = (inp[10]) ? 46'b0001000000000000000000000001000010001000000010 : 46'b0001000000000100000000000000000010001000000000;
														assign node975 = (inp[10]) ? 46'b0001000000000010000000000000000010001000000000 : 46'b0001000000000000001000000001000010001000000000;
											assign node978 = (inp[7]) ? node994 : node979;
												assign node979 = (inp[6]) ? node987 : node980;
													assign node980 = (inp[10]) ? node984 : node981;
														assign node981 = (inp[4]) ? 46'b0000000000000000001000000001100010101000000000 : 46'b0000000000000100000000000000100010101000000000;
														assign node984 = (inp[4]) ? 46'b0000000000000010000000000001100010101000000000 : 46'b0000000000000000000000000001100010101000000010;
													assign node987 = (inp[8]) ? node991 : node988;
														assign node988 = (inp[14]) ? 46'b0000000000000000001000000001100010001000000000 : 46'b0000000000000100000000000000100010001000000000;
														assign node991 = (inp[14]) ? 46'b0000000000000010000000000000100010001000000000 : 46'b0000000000000000000000000001100010001000000010;
												assign node994 = (inp[6]) ? node1002 : node995;
													assign node995 = (inp[14]) ? node999 : node996;
														assign node996 = (inp[8]) ? 46'b0000000000000000000000000001000010101000000010 : 46'b0000000000000100000000000000000010101000000000;
														assign node999 = (inp[8]) ? 46'b0000000000000010000000000000000010101000000000 : 46'b0000000000000000001000000001000010101000000000;
													assign node1002 = (inp[4]) ? node1006 : node1003;
														assign node1003 = (inp[14]) ? 46'b0000000000000100000000000000000010001000000000 : 46'b0000000000000100000000000001000010001000000010;
														assign node1006 = (inp[10]) ? 46'b0000000000000010000000000000000010001000000000 : 46'b0000000000000000001000000001000010001000000000;
										assign node1009 = (inp[7]) ? node1041 : node1010;
											assign node1010 = (inp[6]) ? node1026 : node1011;
												assign node1011 = (inp[5]) ? node1019 : node1012;
													assign node1012 = (inp[8]) ? node1016 : node1013;
														assign node1013 = (inp[14]) ? 46'b0001000000000000001000000001100000101000000000 : 46'b0001000000000100000000000000100000101000000000;
														assign node1016 = (inp[14]) ? 46'b0001000000000010000000000000100000101000000000 : 46'b0001000000000000000000000001100000101000000010;
													assign node1019 = (inp[10]) ? node1023 : node1020;
														assign node1020 = (inp[4]) ? 46'b0000000000000000001000000001100000101000000000 : 46'b0000000000000110000000000000100000101000000000;
														assign node1023 = (inp[4]) ? 46'b0000000000000010000000000000100000101000000000 : 46'b0000000000000000000000000001100000101000000010;
												assign node1026 = (inp[5]) ? node1034 : node1027;
													assign node1027 = (inp[8]) ? node1031 : node1028;
														assign node1028 = (inp[14]) ? 46'b0001000000000000001000000001100000001000000000 : 46'b0001000000000100000000000000100000001000000000;
														assign node1031 = (inp[14]) ? 46'b0001000000000010000000000000100000001000000000 : 46'b0001000000000000000000000001100000001000000010;
													assign node1034 = (inp[8]) ? node1038 : node1035;
														assign node1035 = (inp[14]) ? 46'b0000000000000000001000000001100000001000000000 : 46'b0000000000000100000000000000100000001000000000;
														assign node1038 = (inp[14]) ? 46'b0000000000000010000000000000100000001000000000 : 46'b0000000000000000000000000001100000001000000010;
											assign node1041 = (inp[6]) ? node1057 : node1042;
												assign node1042 = (inp[5]) ? node1050 : node1043;
													assign node1043 = (inp[4]) ? node1047 : node1044;
														assign node1044 = (inp[10]) ? 46'b0001000000000000000000000001000000101000000010 : 46'b0001000000000100000000000000000000101000000000;
														assign node1047 = (inp[10]) ? 46'b0001000000000010000000000000000000101000000000 : 46'b0001000000000000001000000001000000101000000000;
													assign node1050 = (inp[8]) ? node1054 : node1051;
														assign node1051 = (inp[14]) ? 46'b0000000000000000001000000001000000101000000000 : 46'b0000000000000100000000000000000000101000000000;
														assign node1054 = (inp[14]) ? 46'b0000000000000010000000000000000000101000000000 : 46'b0000000000000000000000000001000000101000000010;
												assign node1057 = (inp[5]) ? node1065 : node1058;
													assign node1058 = (inp[8]) ? node1062 : node1059;
														assign node1059 = (inp[14]) ? 46'b0001000000000000001000000001000000001000000000 : 46'b0001000000000100000000000000000000001000000000;
														assign node1062 = (inp[14]) ? 46'b0001000000000010000000000000000000001000000000 : 46'b0001000000000000000000000001000000001000000010;
													assign node1065 = (inp[8]) ? node1069 : node1066;
														assign node1066 = (inp[14]) ? 46'b0000000000000000001000000001000000001000000000 : 46'b0000000000000100000000000000000000001000000000;
														assign node1069 = (inp[14]) ? 46'b0000000000000010000000000000000000001000000000 : 46'b0000000000000000000000000001000000001000000010;
						assign node1072 = (inp[11]) ? node1410 : node1073;
							assign node1073 = (inp[9]) ? node1155 : node1074;
								assign node1074 = (inp[5]) ? node1090 : node1075;
									assign node1075 = (inp[0]) ? node1077 : 46'b0000000000000000000000000000000000000000000000;
										assign node1077 = (inp[7]) ? node1079 : 46'b0000000000000000000000000000000000000000000000;
											assign node1079 = (inp[12]) ? node1081 : 46'b0000000000000000000000000000000000000000000000;
												assign node1081 = (inp[6]) ? node1083 : 46'b0000000000000000000000000000000000000000000000;
													assign node1083 = (inp[8]) ? node1087 : node1084;
														assign node1084 = (inp[14]) ? 46'b0001000000000001001000000001000000000000100000 : 46'b0001000000000101000000000000000000000000100000;
														assign node1087 = (inp[10]) ? 46'b0001000000000011000000000001000000000000100010 : 46'b0001000000000001001000000001000000000000100000;
									assign node1090 = (inp[7]) ? node1104 : node1091;
										assign node1091 = (inp[0]) ? node1093 : 46'b0000000000000000000000000000000000000000000000;
											assign node1093 = (inp[12]) ? node1095 : 46'b0000000000000000000000000000000000000000000000;
												assign node1095 = (inp[6]) ? node1097 : 46'b0000000000000000000000000000000000000000000000;
													assign node1097 = (inp[14]) ? node1101 : node1098;
														assign node1098 = (inp[8]) ? 46'b0000000000000001000000000001100000000000100010 : 46'b0000000000000101000000000001100000000000100000;
														assign node1101 = (inp[8]) ? 46'b0000000000000011000000000000100000000000100000 : 46'b0000000000000001001000000001100000000000100000;
										assign node1104 = (inp[0]) ? node1136 : node1105;
											assign node1105 = (inp[12]) ? node1121 : node1106;
												assign node1106 = (inp[6]) ? node1114 : node1107;
													assign node1107 = (inp[8]) ? node1111 : node1108;
														assign node1108 = (inp[14]) ? 46'b0000000000100000001001000001000010100000000000 : 46'b0000000000100100000001000000000010100000000000;
														assign node1111 = (inp[14]) ? 46'b0000000000100010000001000000000010100000000000 : 46'b0000000000100000000001000001000010100000000010;
													assign node1114 = (inp[8]) ? node1118 : node1115;
														assign node1115 = (inp[14]) ? 46'b0000000000100000001001000001000010000000000000 : 46'b0000000000100100000001000000000010000000000000;
														assign node1118 = (inp[14]) ? 46'b0000000000100010000001000000000010000000000000 : 46'b0000000000100000000001000001000010000000000010;
												assign node1121 = (inp[6]) ? node1129 : node1122;
													assign node1122 = (inp[8]) ? node1126 : node1123;
														assign node1123 = (inp[14]) ? 46'b0000000000100000001001000001000000100000000000 : 46'b0000000000100100000001000000000000100000000000;
														assign node1126 = (inp[14]) ? 46'b0000000000100010000001000001000000100000000000 : 46'b0000000000100000000001000001000000100000000010;
													assign node1129 = (inp[4]) ? node1133 : node1130;
														assign node1130 = (inp[10]) ? 46'b0000000000100000000001000001000000000000000010 : 46'b0000000000100100000001000000000000000000000000;
														assign node1133 = (inp[14]) ? 46'b0000000000100010001001000001000000000000000000 : 46'b0000000000100000000001000001000000000000000010;
											assign node1136 = (inp[6]) ? node1146 : node1137;
												assign node1137 = (inp[12]) ? node1139 : 46'b0000000000000000000000000000000000000000000000;
													assign node1139 = (inp[10]) ? node1143 : node1140;
														assign node1140 = (inp[4]) ? 46'b0000000000000001001000000001000000100000100000 : 46'b0000000000000101000000000000000000100000100000;
														assign node1143 = (inp[4]) ? 46'b0000000000000011000000000000000000100000100000 : 46'b0000000000000001000000000001000000100000100010;
												assign node1146 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node1147;
													assign node1147 = (inp[8]) ? node1151 : node1148;
														assign node1148 = (inp[14]) ? 46'b0000000000000001001000000001000010000000100000 : 46'b0000000000000101000000000000000010000000100000;
														assign node1151 = (inp[14]) ? 46'b0000000000000011000000000000000010000000100000 : 46'b0000000000000001000000000001000010000000100010;
								assign node1155 = (inp[6]) ? node1283 : node1156;
									assign node1156 = (inp[0]) ? node1220 : node1157;
										assign node1157 = (inp[12]) ? node1189 : node1158;
											assign node1158 = (inp[5]) ? node1174 : node1159;
												assign node1159 = (inp[7]) ? node1167 : node1160;
													assign node1160 = (inp[14]) ? node1164 : node1161;
														assign node1161 = (inp[8]) ? 46'b0001000000100000000000000001100010100000100010 : 46'b0001000000100100000000000000100010100000100000;
														assign node1164 = (inp[8]) ? 46'b0001000000100010000000000000100010100000100000 : 46'b0001000000100000001000000001100010100000100000;
													assign node1167 = (inp[4]) ? node1171 : node1168;
														assign node1168 = (inp[10]) ? 46'b0001000000100000000000000001000010100000100010 : 46'b0001000000100100000000000000000010100000100000;
														assign node1171 = (inp[10]) ? 46'b0001000000100010000000000001000010100000100000 : 46'b0001000000100000001000000001000010100000100000;
												assign node1174 = (inp[7]) ? node1182 : node1175;
													assign node1175 = (inp[4]) ? node1179 : node1176;
														assign node1176 = (inp[14]) ? 46'b0000000000100100001000000001100010100000100000 : 46'b0000000000100100000000000001100010100000100010;
														assign node1179 = (inp[10]) ? 46'b0000000000100010000000000000100010100000100000 : 46'b0000000000100000001000000001100010100000100000;
													assign node1182 = (inp[14]) ? node1186 : node1183;
														assign node1183 = (inp[8]) ? 46'b0000000000100000000000000001000010100000100010 : 46'b0000000000100100000000000000000010100000100000;
														assign node1186 = (inp[8]) ? 46'b0000000000100010000000000000000010100000100000 : 46'b0000000000100000001000000001000010100000100000;
											assign node1189 = (inp[7]) ? node1205 : node1190;
												assign node1190 = (inp[5]) ? node1198 : node1191;
													assign node1191 = (inp[14]) ? node1195 : node1192;
														assign node1192 = (inp[8]) ? 46'b0001000000100000000000000001100000100000100010 : 46'b0001000000100100000000000000100000100000100000;
														assign node1195 = (inp[8]) ? 46'b0001000000100010000000000000100000100000100000 : 46'b0001000000100000001000000001100000100000100000;
													assign node1198 = (inp[8]) ? node1202 : node1199;
														assign node1199 = (inp[14]) ? 46'b0000000000100000001000000001100000100000100000 : 46'b0000000000100100000000000001100000100000100000;
														assign node1202 = (inp[14]) ? 46'b0000000000100010000000000000100000100000100000 : 46'b0000000000100000000000000001100000100000100010;
												assign node1205 = (inp[5]) ? node1213 : node1206;
													assign node1206 = (inp[8]) ? node1210 : node1207;
														assign node1207 = (inp[14]) ? 46'b0001000000100000001000000001000000100000100000 : 46'b0001000000100100000000000000000000100000100000;
														assign node1210 = (inp[14]) ? 46'b0001000000100010000000000000000000100000100000 : 46'b0001000000100000000000000001000000100000100010;
													assign node1213 = (inp[4]) ? node1217 : node1214;
														assign node1214 = (inp[10]) ? 46'b0000000000100000000000000001000000100000100010 : 46'b0000000000100100000000000000000000100000100000;
														assign node1217 = (inp[10]) ? 46'b0000000000100010000000000000000000100000100000 : 46'b0000000000100000001000000001000000100000100000;
										assign node1220 = (inp[7]) ? node1252 : node1221;
											assign node1221 = (inp[12]) ? node1237 : node1222;
												assign node1222 = (inp[5]) ? node1230 : node1223;
													assign node1223 = (inp[14]) ? node1227 : node1224;
														assign node1224 = (inp[8]) ? 46'b0001000000000000000000000001100010100000100010 : 46'b0001000000000100000000000000100010100000100000;
														assign node1227 = (inp[8]) ? 46'b0001000000000010000000000000100010100000100000 : 46'b0001000000000000001000000001100010100000100010;
													assign node1230 = (inp[10]) ? node1234 : node1231;
														assign node1231 = (inp[4]) ? 46'b0000000000000000001000000001100010100000100000 : 46'b0000000000000100000000000000100010100000100000;
														assign node1234 = (inp[4]) ? 46'b0000000000000010000000000000100010100000100000 : 46'b0000000000000000000000000001100010100000100010;
												assign node1237 = (inp[5]) ? node1245 : node1238;
													assign node1238 = (inp[8]) ? node1242 : node1239;
														assign node1239 = (inp[14]) ? 46'b0001000000000000001000000001100000100000100000 : 46'b0001000000000100000000000000100000100000100000;
														assign node1242 = (inp[14]) ? 46'b0001000000000010000000000001100000100000100000 : 46'b0001000000000000000000000001100000100000100010;
													assign node1245 = (inp[14]) ? node1249 : node1246;
														assign node1246 = (inp[8]) ? 46'b0000000000000000000000000001100000100000100010 : 46'b0000000000000100000000000000100000100000100000;
														assign node1249 = (inp[4]) ? 46'b0000000000000010001000000001100000100000100000 : 46'b0000000000000000001000000001100000100000100000;
											assign node1252 = (inp[5]) ? node1268 : node1253;
												assign node1253 = (inp[12]) ? node1261 : node1254;
													assign node1254 = (inp[4]) ? node1258 : node1255;
														assign node1255 = (inp[10]) ? 46'b0001000000000000000000000001000010100000100010 : 46'b0001000000000100000000000001000010100000100000;
														assign node1258 = (inp[10]) ? 46'b0001000000000010000000000000000010100000100000 : 46'b0001000000000000001000000001000010100000100000;
													assign node1261 = (inp[4]) ? node1265 : node1262;
														assign node1262 = (inp[10]) ? 46'b0001000000000000000000000001000000100000100010 : 46'b0001000000000100000000000000000000100000100000;
														assign node1265 = (inp[10]) ? 46'b0001000000000010000000000000000000100000100000 : 46'b0001000000000000001000000001000000100000100000;
												assign node1268 = (inp[12]) ? node1276 : node1269;
													assign node1269 = (inp[10]) ? node1273 : node1270;
														assign node1270 = (inp[4]) ? 46'b0000000000000000001000000001000010100000100000 : 46'b0000000000000100000000000001000010100000100000;
														assign node1273 = (inp[4]) ? 46'b0000000000000010000000000000000010100000100000 : 46'b0000000000000000000000000001000010100000100010;
													assign node1276 = (inp[4]) ? node1280 : node1277;
														assign node1277 = (inp[10]) ? 46'b0000000000000000000000000001000000100000100010 : 46'b0000000000000100000000000000000000100000100000;
														assign node1280 = (inp[10]) ? 46'b0000000000000010000000000000000000100000100000 : 46'b0000000000000000001000000001000000100000100000;
									assign node1283 = (inp[0]) ? node1347 : node1284;
										assign node1284 = (inp[12]) ? node1316 : node1285;
											assign node1285 = (inp[7]) ? node1301 : node1286;
												assign node1286 = (inp[5]) ? node1294 : node1287;
													assign node1287 = (inp[4]) ? node1291 : node1288;
														assign node1288 = (inp[10]) ? 46'b0001000000100000000000000001100010000000100010 : 46'b0001000000100100000000000001100010000000100000;
														assign node1291 = (inp[10]) ? 46'b0001000000100010000000000000100010000000100000 : 46'b0001000000100000001000000001100010000000100000;
													assign node1294 = (inp[8]) ? node1298 : node1295;
														assign node1295 = (inp[14]) ? 46'b0000000000100000001000000001100010000000100000 : 46'b0000000000100100000000000001100010000000100000;
														assign node1298 = (inp[14]) ? 46'b0000000000100010000000000000100010000000100000 : 46'b0000000000100000000000000001100010000000100010;
												assign node1301 = (inp[5]) ? node1309 : node1302;
													assign node1302 = (inp[10]) ? node1306 : node1303;
														assign node1303 = (inp[4]) ? 46'b0001000000100000001000000001000010000000100000 : 46'b0001000000100100000000000000000010000000100000;
														assign node1306 = (inp[4]) ? 46'b0001000000100010000000000000000010000000100000 : 46'b0001000000100000000000000001000010000000100010;
													assign node1309 = (inp[4]) ? node1313 : node1310;
														assign node1310 = (inp[10]) ? 46'b0000000000100000000000000001000010000000100010 : 46'b0000000000100100000000000000000010000000100000;
														assign node1313 = (inp[10]) ? 46'b0000000000100010000000000000000010000000100000 : 46'b0000000000100000001000000001000010000000100000;
											assign node1316 = (inp[5]) ? node1332 : node1317;
												assign node1317 = (inp[7]) ? node1325 : node1318;
													assign node1318 = (inp[10]) ? node1322 : node1319;
														assign node1319 = (inp[4]) ? 46'b0001000000100000001000000001100000000000100000 : 46'b0001000000100100000000000000100000000000100000;
														assign node1322 = (inp[4]) ? 46'b0001000000100010000000000000100000000000100000 : 46'b0001000000100000000000000001100000000000100010;
													assign node1325 = (inp[8]) ? node1329 : node1326;
														assign node1326 = (inp[14]) ? 46'b0001000000100000001000000001000000000000100000 : 46'b0001000000100100000000000000000000000000100000;
														assign node1329 = (inp[14]) ? 46'b0001000000100010000000000000000000000000100000 : 46'b0001000000100000000000000001000000000000100010;
												assign node1332 = (inp[7]) ? node1340 : node1333;
													assign node1333 = (inp[14]) ? node1337 : node1334;
														assign node1334 = (inp[8]) ? 46'b0000000000100000000000000001100000000000100010 : 46'b0000000000100100000000000001100000000000100000;
														assign node1337 = (inp[8]) ? 46'b0000000000100010000000000000100000000000100000 : 46'b0000000000100000001000000001100000000000100000;
													assign node1340 = (inp[4]) ? node1344 : node1341;
														assign node1341 = (inp[10]) ? 46'b0000000000100000000000000001000000000000100010 : 46'b0000000000100100000000000000000000000000100000;
														assign node1344 = (inp[10]) ? 46'b0000000000100010000000000000000000000000100000 : 46'b0000000000100000001000000001000000000000100000;
										assign node1347 = (inp[5]) ? node1379 : node1348;
											assign node1348 = (inp[7]) ? node1364 : node1349;
												assign node1349 = (inp[12]) ? node1357 : node1350;
													assign node1350 = (inp[4]) ? node1354 : node1351;
														assign node1351 = (inp[10]) ? 46'b0001000000000000000000000001100010000000100010 : 46'b0001000000000100000000000000100010000000100000;
														assign node1354 = (inp[10]) ? 46'b0001000000000010000000000000100010000000100000 : 46'b0001000000000000001000000001100010000000100000;
													assign node1357 = (inp[4]) ? node1361 : node1358;
														assign node1358 = (inp[10]) ? 46'b0001000000000000000000000001100000000000100010 : 46'b0001000000000100000000000000100000000000100000;
														assign node1361 = (inp[10]) ? 46'b0001000000000010000000000000100000000000100000 : 46'b0001000000000000001000000001100000000000100000;
												assign node1364 = (inp[12]) ? node1372 : node1365;
													assign node1365 = (inp[4]) ? node1369 : node1366;
														assign node1366 = (inp[10]) ? 46'b0001000000000000000000000001000010000000100010 : 46'b0001000000000100000000000001000010000000100000;
														assign node1369 = (inp[14]) ? 46'b0001000000000010001000000001000010000000100000 : 46'b0001000000000100001000000001000010000000100000;
													assign node1372 = (inp[8]) ? node1376 : node1373;
														assign node1373 = (inp[14]) ? 46'b0001000000000000001000000001000000000000100000 : 46'b0001000000000100000000000000000000000000100000;
														assign node1376 = (inp[14]) ? 46'b0001000000000010000000000000000000000000100000 : 46'b0001000000000000000000000001000000000000100010;
											assign node1379 = (inp[12]) ? node1395 : node1380;
												assign node1380 = (inp[7]) ? node1388 : node1381;
													assign node1381 = (inp[10]) ? node1385 : node1382;
														assign node1382 = (inp[4]) ? 46'b0000000000000000001000000001100010000000100000 : 46'b0000000000000100000000000000100010000000100000;
														assign node1385 = (inp[4]) ? 46'b0000000000000010000000000000100010000000100000 : 46'b0000000000000000000000000001100010000000100010;
													assign node1388 = (inp[14]) ? node1392 : node1389;
														assign node1389 = (inp[8]) ? 46'b0000000000000000000000000001000010000000100010 : 46'b0000000000000100000000000000000010000000100000;
														assign node1392 = (inp[8]) ? 46'b0000000000000010000000000000000010000000100000 : 46'b0000000000000000001000000001000010000000100000;
												assign node1395 = (inp[7]) ? node1403 : node1396;
													assign node1396 = (inp[4]) ? node1400 : node1397;
														assign node1397 = (inp[10]) ? 46'b0000000000000000000000000001100000000000100010 : 46'b0000000000000100000000000000100000000000100000;
														assign node1400 = (inp[10]) ? 46'b0000000000000010000000000000100000000000100000 : 46'b0000000000000000001000000001100000000000100000;
													assign node1403 = (inp[8]) ? node1407 : node1404;
														assign node1404 = (inp[14]) ? 46'b0000000000000000001000000001000000000000100000 : 46'b0000000000000100000000000000000000000000100000;
														assign node1407 = (inp[14]) ? 46'b0000000000000010000000000000000000000000100000 : 46'b0000000000000000000000000001000000000000100010;
							assign node1410 = (inp[7]) ? node1448 : node1411;
								assign node1411 = (inp[5]) ? node1423 : node1412;
									assign node1412 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1413;
										assign node1413 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1414;
											assign node1414 = (inp[12]) ? node1418 : node1415;
												assign node1415 = (inp[6]) ? 46'b0001000000100010000000000000100010000000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1418 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000100000001000000001100000100000100000;
									assign node1423 = (inp[0]) ? node1439 : node1424;
										assign node1424 = (inp[9]) ? node1432 : node1425;
											assign node1425 = (inp[6]) ? node1429 : node1426;
												assign node1426 = (inp[12]) ? 46'b0000000000100000001000000001100000100000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1429 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000100010000000000000100010000000100000;
											assign node1432 = (inp[12]) ? node1436 : node1433;
												assign node1433 = (inp[6]) ? 46'b0000000010000000000000000001100010000001000010 : 46'b0000000010000000000000000001100010100001000010;
												assign node1436 = (inp[6]) ? 46'b0000000010000000000000000001100000000001000010 : 46'b0000000010000000000000000001100000100001000010;
										assign node1439 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1440;
											assign node1440 = (inp[6]) ? node1444 : node1441;
												assign node1441 = (inp[12]) ? 46'b0000000010000000000000000001100000100000000010 : 46'b0000000010000000000000000001100010100000000010;
												assign node1444 = (inp[12]) ? 46'b0000000010000000000000000001100000000000000010 : 46'b0000000010000000000000000001100010000000000010;
								assign node1448 = (inp[5]) ? node1474 : node1449;
									assign node1449 = (inp[9]) ? node1465 : node1450;
										assign node1450 = (inp[0]) ? node1458 : node1451;
											assign node1451 = (inp[6]) ? node1455 : node1452;
												assign node1452 = (inp[12]) ? 46'b0001000000100000001000000001000000100000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1455 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000100010000000000000000010000000100000;
											assign node1458 = (inp[12]) ? node1462 : node1459;
												assign node1459 = (inp[6]) ? 46'b0001000010000100000000000000000010000000000000 : 46'b0001000010000100000000000000000010100000000000;
												assign node1462 = (inp[6]) ? 46'b0001000010000100000000000000000000000000000000 : 46'b0001000010000100000000000000000000100000000000;
										assign node1465 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1466;
											assign node1466 = (inp[12]) ? node1470 : node1467;
												assign node1467 = (inp[6]) ? 46'b0001000010000100000000000000000010000001000000 : 46'b0001000010000100000000000000000010100001000000;
												assign node1470 = (inp[6]) ? 46'b0001000010000100000000000000000000000001000000 : 46'b0001000010000100000000000000000000100001000000;
									assign node1474 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node1475;
										assign node1475 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node1476;
											assign node1476 = (inp[12]) ? node1480 : node1477;
												assign node1477 = (inp[6]) ? 46'b0000000000100010000000000000000010000000100000 : 46'b0000000000000000000000000000000000000000000000;
												assign node1480 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000100000001000000001000000100000100000;

endmodule