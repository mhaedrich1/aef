module dtc_split25_bm64 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node14;
	wire [4-1:0] node18;
	wire [4-1:0] node19;
	wire [4-1:0] node21;
	wire [4-1:0] node26;
	wire [4-1:0] node28;
	wire [4-1:0] node29;
	wire [4-1:0] node31;
	wire [4-1:0] node36;
	wire [4-1:0] node38;
	wire [4-1:0] node39;
	wire [4-1:0] node40;
	wire [4-1:0] node44;
	wire [4-1:0] node46;
	wire [4-1:0] node48;
	wire [4-1:0] node52;
	wire [4-1:0] node54;
	wire [4-1:0] node55;
	wire [4-1:0] node56;
	wire [4-1:0] node57;
	wire [4-1:0] node58;
	wire [4-1:0] node62;
	wire [4-1:0] node64;
	wire [4-1:0] node66;
	wire [4-1:0] node70;
	wire [4-1:0] node72;
	wire [4-1:0] node73;
	wire [4-1:0] node75;
	wire [4-1:0] node78;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node86;
	wire [4-1:0] node87;
	wire [4-1:0] node88;
	wire [4-1:0] node89;
	wire [4-1:0] node90;
	wire [4-1:0] node91;
	wire [4-1:0] node93;
	wire [4-1:0] node94;
	wire [4-1:0] node99;
	wire [4-1:0] node101;
	wire [4-1:0] node102;
	wire [4-1:0] node103;
	wire [4-1:0] node104;
	wire [4-1:0] node106;
	wire [4-1:0] node112;
	wire [4-1:0] node113;
	wire [4-1:0] node114;
	wire [4-1:0] node116;
	wire [4-1:0] node120;
	wire [4-1:0] node122;
	wire [4-1:0] node123;
	wire [4-1:0] node125;
	wire [4-1:0] node126;
	wire [4-1:0] node130;
	wire [4-1:0] node132;
	wire [4-1:0] node133;
	wire [4-1:0] node135;
	wire [4-1:0] node136;
	wire [4-1:0] node141;
	wire [4-1:0] node142;
	wire [4-1:0] node143;
	wire [4-1:0] node144;
	wire [4-1:0] node146;
	wire [4-1:0] node147;
	wire [4-1:0] node148;
	wire [4-1:0] node149;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node160;
	wire [4-1:0] node162;
	wire [4-1:0] node164;
	wire [4-1:0] node166;
	wire [4-1:0] node169;
	wire [4-1:0] node171;
	wire [4-1:0] node172;
	wire [4-1:0] node173;
	wire [4-1:0] node174;
	wire [4-1:0] node179;
	wire [4-1:0] node180;
	wire [4-1:0] node182;
	wire [4-1:0] node184;
	wire [4-1:0] node187;
	wire [4-1:0] node188;
	wire [4-1:0] node190;
	wire [4-1:0] node192;
	wire [4-1:0] node193;
	wire [4-1:0] node198;
	wire [4-1:0] node200;
	wire [4-1:0] node201;
	wire [4-1:0] node202;
	wire [4-1:0] node203;
	wire [4-1:0] node204;
	wire [4-1:0] node205;
	wire [4-1:0] node208;
	wire [4-1:0] node209;
	wire [4-1:0] node214;
	wire [4-1:0] node216;
	wire [4-1:0] node218;
	wire [4-1:0] node220;
	wire [4-1:0] node222;
	wire [4-1:0] node226;
	wire [4-1:0] node228;
	wire [4-1:0] node229;
	wire [4-1:0] node230;
	wire [4-1:0] node232;
	wire [4-1:0] node236;
	wire [4-1:0] node238;
	wire [4-1:0] node239;
	wire [4-1:0] node240;
	wire [4-1:0] node245;
	wire [4-1:0] node246;
	wire [4-1:0] node248;
	wire [4-1:0] node249;
	wire [4-1:0] node250;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node253;
	wire [4-1:0] node254;
	wire [4-1:0] node255;
	wire [4-1:0] node260;
	wire [4-1:0] node262;
	wire [4-1:0] node266;
	wire [4-1:0] node268;
	wire [4-1:0] node269;
	wire [4-1:0] node270;
	wire [4-1:0] node271;
	wire [4-1:0] node272;
	wire [4-1:0] node277;
	wire [4-1:0] node279;
	wire [4-1:0] node282;
	wire [4-1:0] node284;
	wire [4-1:0] node288;
	wire [4-1:0] node290;
	wire [4-1:0] node291;
	wire [4-1:0] node292;
	wire [4-1:0] node293;
	wire [4-1:0] node295;
	wire [4-1:0] node296;
	wire [4-1:0] node300;
	wire [4-1:0] node302;
	wire [4-1:0] node303;
	wire [4-1:0] node308;
	wire [4-1:0] node310;
	wire [4-1:0] node311;
	wire [4-1:0] node313;
	wire [4-1:0] node315;
	wire [4-1:0] node317;
	wire [4-1:0] node320;
	wire [4-1:0] node321;
	wire [4-1:0] node323;
	wire [4-1:0] node327;
	wire [4-1:0] node328;
	wire [4-1:0] node329;
	wire [4-1:0] node330;
	wire [4-1:0] node331;
	wire [4-1:0] node332;
	wire [4-1:0] node333;
	wire [4-1:0] node334;
	wire [4-1:0] node335;
	wire [4-1:0] node341;
	wire [4-1:0] node342;
	wire [4-1:0] node344;
	wire [4-1:0] node345;
	wire [4-1:0] node349;
	wire [4-1:0] node350;
	wire [4-1:0] node351;
	wire [4-1:0] node352;
	wire [4-1:0] node358;
	wire [4-1:0] node360;
	wire [4-1:0] node361;
	wire [4-1:0] node362;
	wire [4-1:0] node364;
	wire [4-1:0] node368;
	wire [4-1:0] node370;
	wire [4-1:0] node371;
	wire [4-1:0] node375;
	wire [4-1:0] node376;
	wire [4-1:0] node377;
	wire [4-1:0] node378;
	wire [4-1:0] node379;
	wire [4-1:0] node380;
	wire [4-1:0] node381;
	wire [4-1:0] node387;
	wire [4-1:0] node388;
	wire [4-1:0] node389;
	wire [4-1:0] node390;
	wire [4-1:0] node397;
	wire [4-1:0] node399;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node403;
	wire [4-1:0] node408;
	wire [4-1:0] node409;
	wire [4-1:0] node410;
	wire [4-1:0] node411;
	wire [4-1:0] node412;
	wire [4-1:0] node413;
	wire [4-1:0] node414;
	wire [4-1:0] node415;
	wire [4-1:0] node419;
	wire [4-1:0] node423;
	wire [4-1:0] node424;
	wire [4-1:0] node426;
	wire [4-1:0] node427;
	wire [4-1:0] node431;
	wire [4-1:0] node433;
	wire [4-1:0] node435;
	wire [4-1:0] node438;
	wire [4-1:0] node439;
	wire [4-1:0] node440;
	wire [4-1:0] node441;
	wire [4-1:0] node444;
	wire [4-1:0] node445;
	wire [4-1:0] node449;
	wire [4-1:0] node450;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node456;
	wire [4-1:0] node457;
	wire [4-1:0] node458;
	wire [4-1:0] node464;
	wire [4-1:0] node466;
	wire [4-1:0] node468;
	wire [4-1:0] node469;
	wire [4-1:0] node473;
	wire [4-1:0] node474;
	wire [4-1:0] node475;
	wire [4-1:0] node476;
	wire [4-1:0] node478;
	wire [4-1:0] node479;
	wire [4-1:0] node483;
	wire [4-1:0] node486;
	wire [4-1:0] node487;
	wire [4-1:0] node488;
	wire [4-1:0] node489;
	wire [4-1:0] node490;
	wire [4-1:0] node497;
	wire [4-1:0] node498;
	wire [4-1:0] node499;
	wire [4-1:0] node500;
	wire [4-1:0] node502;
	wire [4-1:0] node505;
	wire [4-1:0] node509;
	wire [4-1:0] node510;
	wire [4-1:0] node512;
	wire [4-1:0] node516;
	wire [4-1:0] node517;
	wire [4-1:0] node518;
	wire [4-1:0] node519;
	wire [4-1:0] node520;
	wire [4-1:0] node522;
	wire [4-1:0] node525;
	wire [4-1:0] node527;
	wire [4-1:0] node528;
	wire [4-1:0] node531;
	wire [4-1:0] node534;
	wire [4-1:0] node535;
	wire [4-1:0] node536;
	wire [4-1:0] node541;
	wire [4-1:0] node542;
	wire [4-1:0] node543;
	wire [4-1:0] node544;
	wire [4-1:0] node548;
	wire [4-1:0] node550;
	wire [4-1:0] node551;
	wire [4-1:0] node555;
	wire [4-1:0] node556;
	wire [4-1:0] node560;
	wire [4-1:0] node561;
	wire [4-1:0] node562;
	wire [4-1:0] node563;
	wire [4-1:0] node565;
	wire [4-1:0] node567;
	wire [4-1:0] node570;
	wire [4-1:0] node572;
	wire [4-1:0] node575;
	wire [4-1:0] node576;
	wire [4-1:0] node577;
	wire [4-1:0] node578;
	wire [4-1:0] node582;
	wire [4-1:0] node585;
	wire [4-1:0] node586;
	wire [4-1:0] node590;
	wire [4-1:0] node591;
	wire [4-1:0] node592;
	wire [4-1:0] node593;
	wire [4-1:0] node594;
	wire [4-1:0] node599;
	wire [4-1:0] node600;
	wire [4-1:0] node601;
	wire [4-1:0] node602;
	wire [4-1:0] node605;
	wire [4-1:0] node607;
	wire [4-1:0] node610;
	wire [4-1:0] node612;
	wire [4-1:0] node616;
	wire [4-1:0] node617;
	wire [4-1:0] node620;
	wire [4-1:0] node623;
	wire [4-1:0] node624;
	wire [4-1:0] node625;
	wire [4-1:0] node626;
	wire [4-1:0] node627;
	wire [4-1:0] node628;
	wire [4-1:0] node629;
	wire [4-1:0] node631;
	wire [4-1:0] node635;
	wire [4-1:0] node636;
	wire [4-1:0] node637;
	wire [4-1:0] node639;
	wire [4-1:0] node643;
	wire [4-1:0] node646;
	wire [4-1:0] node647;
	wire [4-1:0] node648;
	wire [4-1:0] node651;
	wire [4-1:0] node653;
	wire [4-1:0] node654;
	wire [4-1:0] node658;
	wire [4-1:0] node660;
	wire [4-1:0] node661;
	wire [4-1:0] node662;
	wire [4-1:0] node667;
	wire [4-1:0] node668;
	wire [4-1:0] node669;
	wire [4-1:0] node671;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node678;
	wire [4-1:0] node680;
	wire [4-1:0] node683;
	wire [4-1:0] node684;
	wire [4-1:0] node685;
	wire [4-1:0] node687;
	wire [4-1:0] node691;
	wire [4-1:0] node692;
	wire [4-1:0] node696;
	wire [4-1:0] node697;
	wire [4-1:0] node698;
	wire [4-1:0] node699;
	wire [4-1:0] node700;
	wire [4-1:0] node701;
	wire [4-1:0] node706;
	wire [4-1:0] node708;
	wire [4-1:0] node709;
	wire [4-1:0] node713;
	wire [4-1:0] node714;
	wire [4-1:0] node715;
	wire [4-1:0] node720;
	wire [4-1:0] node721;
	wire [4-1:0] node722;
	wire [4-1:0] node724;
	wire [4-1:0] node725;
	wire [4-1:0] node727;
	wire [4-1:0] node731;
	wire [4-1:0] node733;
	wire [4-1:0] node736;
	wire [4-1:0] node737;
	wire [4-1:0] node739;
	wire [4-1:0] node740;
	wire [4-1:0] node744;
	wire [4-1:0] node746;
	wire [4-1:0] node747;
	wire [4-1:0] node751;
	wire [4-1:0] node752;
	wire [4-1:0] node753;
	wire [4-1:0] node754;
	wire [4-1:0] node755;
	wire [4-1:0] node756;
	wire [4-1:0] node758;
	wire [4-1:0] node761;
	wire [4-1:0] node762;
	wire [4-1:0] node764;
	wire [4-1:0] node767;
	wire [4-1:0] node768;
	wire [4-1:0] node772;
	wire [4-1:0] node773;
	wire [4-1:0] node774;
	wire [4-1:0] node777;
	wire [4-1:0] node780;
	wire [4-1:0] node783;
	wire [4-1:0] node784;
	wire [4-1:0] node785;
	wire [4-1:0] node786;
	wire [4-1:0] node788;
	wire [4-1:0] node791;
	wire [4-1:0] node794;
	wire [4-1:0] node795;
	wire [4-1:0] node798;
	wire [4-1:0] node801;
	wire [4-1:0] node802;
	wire [4-1:0] node803;
	wire [4-1:0] node805;
	wire [4-1:0] node809;
	wire [4-1:0] node810;
	wire [4-1:0] node811;
	wire [4-1:0] node815;
	wire [4-1:0] node816;
	wire [4-1:0] node820;
	wire [4-1:0] node821;
	wire [4-1:0] node822;
	wire [4-1:0] node823;
	wire [4-1:0] node826;
	wire [4-1:0] node827;
	wire [4-1:0] node831;
	wire [4-1:0] node832;
	wire [4-1:0] node834;
	wire [4-1:0] node837;
	wire [4-1:0] node839;
	wire [4-1:0] node842;
	wire [4-1:0] node843;
	wire [4-1:0] node844;
	wire [4-1:0] node845;
	wire [4-1:0] node849;
	wire [4-1:0] node850;
	wire [4-1:0] node854;
	wire [4-1:0] node855;
	wire [4-1:0] node856;
	wire [4-1:0] node859;
	wire [4-1:0] node861;
	wire [4-1:0] node863;
	wire [4-1:0] node866;
	wire [4-1:0] node869;
	wire [4-1:0] node870;
	wire [4-1:0] node871;
	wire [4-1:0] node872;
	wire [4-1:0] node873;
	wire [4-1:0] node874;
	wire [4-1:0] node875;
	wire [4-1:0] node878;
	wire [4-1:0] node881;
	wire [4-1:0] node882;
	wire [4-1:0] node883;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node891;
	wire [4-1:0] node893;
	wire [4-1:0] node895;
	wire [4-1:0] node898;
	wire [4-1:0] node901;
	wire [4-1:0] node902;
	wire [4-1:0] node903;
	wire [4-1:0] node904;
	wire [4-1:0] node907;
	wire [4-1:0] node910;
	wire [4-1:0] node913;
	wire [4-1:0] node914;
	wire [4-1:0] node915;
	wire [4-1:0] node916;
	wire [4-1:0] node918;
	wire [4-1:0] node921;
	wire [4-1:0] node922;
	wire [4-1:0] node928;
	wire [4-1:0] node929;
	wire [4-1:0] node930;
	wire [4-1:0] node933;
	wire [4-1:0] node936;
	wire [4-1:0] node937;
	wire [4-1:0] node940;
	wire [4-1:0] node943;
	wire [4-1:0] node944;
	wire [4-1:0] node945;
	wire [4-1:0] node946;
	wire [4-1:0] node949;
	wire [4-1:0] node952;
	wire [4-1:0] node953;
	wire [4-1:0] node956;
	wire [4-1:0] node960;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node964;
	wire [4-1:0] node965;
	wire [4-1:0] node966;
	wire [4-1:0] node967;
	wire [4-1:0] node968;
	wire [4-1:0] node970;
	wire [4-1:0] node974;
	wire [4-1:0] node976;
	wire [4-1:0] node977;
	wire [4-1:0] node978;
	wire [4-1:0] node982;
	wire [4-1:0] node984;
	wire [4-1:0] node988;
	wire [4-1:0] node989;
	wire [4-1:0] node990;
	wire [4-1:0] node991;
	wire [4-1:0] node992;
	wire [4-1:0] node993;
	wire [4-1:0] node998;
	wire [4-1:0] node1000;
	wire [4-1:0] node1001;
	wire [4-1:0] node1002;
	wire [4-1:0] node1003;
	wire [4-1:0] node1008;
	wire [4-1:0] node1010;
	wire [4-1:0] node1012;
	wire [4-1:0] node1016;
	wire [4-1:0] node1017;
	wire [4-1:0] node1018;
	wire [4-1:0] node1019;
	wire [4-1:0] node1021;
	wire [4-1:0] node1022;
	wire [4-1:0] node1024;
	wire [4-1:0] node1029;
	wire [4-1:0] node1030;
	wire [4-1:0] node1031;
	wire [4-1:0] node1032;
	wire [4-1:0] node1033;
	wire [4-1:0] node1039;
	wire [4-1:0] node1040;
	wire [4-1:0] node1042;
	wire [4-1:0] node1046;
	wire [4-1:0] node1047;
	wire [4-1:0] node1048;
	wire [4-1:0] node1049;
	wire [4-1:0] node1050;
	wire [4-1:0] node1051;
	wire [4-1:0] node1057;
	wire [4-1:0] node1058;
	wire [4-1:0] node1060;
	wire [4-1:0] node1061;
	wire [4-1:0] node1066;
	wire [4-1:0] node1067;
	wire [4-1:0] node1068;
	wire [4-1:0] node1070;
	wire [4-1:0] node1075;
	wire [4-1:0] node1076;
	wire [4-1:0] node1078;
	wire [4-1:0] node1079;
	wire [4-1:0] node1080;
	wire [4-1:0] node1081;
	wire [4-1:0] node1082;
	wire [4-1:0] node1086;
	wire [4-1:0] node1087;
	wire [4-1:0] node1089;
	wire [4-1:0] node1092;
	wire [4-1:0] node1093;
	wire [4-1:0] node1094;
	wire [4-1:0] node1100;
	wire [4-1:0] node1102;
	wire [4-1:0] node1103;
	wire [4-1:0] node1105;
	wire [4-1:0] node1106;
	wire [4-1:0] node1108;
	wire [4-1:0] node1112;
	wire [4-1:0] node1114;
	wire [4-1:0] node1115;
	wire [4-1:0] node1116;
	wire [4-1:0] node1118;
	wire [4-1:0] node1123;
	wire [4-1:0] node1124;
	wire [4-1:0] node1125;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1128;
	wire [4-1:0] node1129;
	wire [4-1:0] node1133;
	wire [4-1:0] node1135;
	wire [4-1:0] node1137;
	wire [4-1:0] node1140;
	wire [4-1:0] node1143;
	wire [4-1:0] node1144;
	wire [4-1:0] node1145;
	wire [4-1:0] node1148;
	wire [4-1:0] node1149;
	wire [4-1:0] node1150;
	wire [4-1:0] node1153;
	wire [4-1:0] node1155;
	wire [4-1:0] node1158;
	wire [4-1:0] node1160;
	wire [4-1:0] node1163;
	wire [4-1:0] node1164;
	wire [4-1:0] node1165;
	wire [4-1:0] node1168;
	wire [4-1:0] node1171;
	wire [4-1:0] node1174;
	wire [4-1:0] node1175;
	wire [4-1:0] node1176;
	wire [4-1:0] node1177;
	wire [4-1:0] node1178;
	wire [4-1:0] node1179;
	wire [4-1:0] node1183;
	wire [4-1:0] node1185;
	wire [4-1:0] node1188;
	wire [4-1:0] node1190;
	wire [4-1:0] node1192;
	wire [4-1:0] node1195;
	wire [4-1:0] node1196;
	wire [4-1:0] node1198;
	wire [4-1:0] node1201;
	wire [4-1:0] node1202;
	wire [4-1:0] node1203;
	wire [4-1:0] node1206;
	wire [4-1:0] node1209;
	wire [4-1:0] node1212;
	wire [4-1:0] node1213;
	wire [4-1:0] node1215;
	wire [4-1:0] node1216;
	wire [4-1:0] node1220;
	wire [4-1:0] node1221;
	wire [4-1:0] node1222;
	wire [4-1:0] node1223;
	wire [4-1:0] node1224;
	wire [4-1:0] node1230;
	wire [4-1:0] node1231;
	wire [4-1:0] node1235;
	wire [4-1:0] node1236;
	wire [4-1:0] node1237;
	wire [4-1:0] node1238;
	wire [4-1:0] node1240;
	wire [4-1:0] node1241;
	wire [4-1:0] node1245;
	wire [4-1:0] node1246;
	wire [4-1:0] node1247;
	wire [4-1:0] node1248;
	wire [4-1:0] node1249;
	wire [4-1:0] node1255;
	wire [4-1:0] node1257;
	wire [4-1:0] node1258;
	wire [4-1:0] node1260;
	wire [4-1:0] node1263;
	wire [4-1:0] node1266;
	wire [4-1:0] node1267;
	wire [4-1:0] node1268;
	wire [4-1:0] node1270;
	wire [4-1:0] node1273;
	wire [4-1:0] node1275;
	wire [4-1:0] node1278;
	wire [4-1:0] node1280;
	wire [4-1:0] node1281;
	wire [4-1:0] node1285;
	wire [4-1:0] node1286;
	wire [4-1:0] node1287;
	wire [4-1:0] node1288;
	wire [4-1:0] node1289;
	wire [4-1:0] node1290;
	wire [4-1:0] node1294;
	wire [4-1:0] node1297;
	wire [4-1:0] node1300;
	wire [4-1:0] node1301;
	wire [4-1:0] node1302;
	wire [4-1:0] node1305;
	wire [4-1:0] node1306;
	wire [4-1:0] node1310;
	wire [4-1:0] node1313;
	wire [4-1:0] node1314;
	wire [4-1:0] node1315;
	wire [4-1:0] node1316;
	wire [4-1:0] node1319;
	wire [4-1:0] node1322;
	wire [4-1:0] node1323;
	wire [4-1:0] node1326;
	wire [4-1:0] node1330;
	wire [4-1:0] node1332;
	wire [4-1:0] node1333;
	wire [4-1:0] node1334;
	wire [4-1:0] node1335;
	wire [4-1:0] node1336;
	wire [4-1:0] node1337;
	wire [4-1:0] node1338;
	wire [4-1:0] node1339;
	wire [4-1:0] node1344;
	wire [4-1:0] node1346;
	wire [4-1:0] node1347;
	wire [4-1:0] node1349;
	wire [4-1:0] node1354;
	wire [4-1:0] node1355;
	wire [4-1:0] node1356;
	wire [4-1:0] node1358;
	wire [4-1:0] node1359;
	wire [4-1:0] node1363;
	wire [4-1:0] node1364;
	wire [4-1:0] node1366;
	wire [4-1:0] node1367;
	wire [4-1:0] node1370;
	wire [4-1:0] node1373;
	wire [4-1:0] node1375;
	wire [4-1:0] node1377;
	wire [4-1:0] node1378;
	wire [4-1:0] node1381;
	wire [4-1:0] node1384;
	wire [4-1:0] node1386;
	wire [4-1:0] node1387;
	wire [4-1:0] node1389;
	wire [4-1:0] node1390;
	wire [4-1:0] node1394;
	wire [4-1:0] node1396;
	wire [4-1:0] node1397;
	wire [4-1:0] node1401;
	wire [4-1:0] node1402;
	wire [4-1:0] node1404;
	wire [4-1:0] node1405;
	wire [4-1:0] node1406;
	wire [4-1:0] node1407;
	wire [4-1:0] node1409;
	wire [4-1:0] node1413;
	wire [4-1:0] node1416;
	wire [4-1:0] node1418;
	wire [4-1:0] node1421;
	wire [4-1:0] node1422;
	wire [4-1:0] node1423;
	wire [4-1:0] node1424;
	wire [4-1:0] node1425;
	wire [4-1:0] node1426;
	wire [4-1:0] node1430;
	wire [4-1:0] node1431;
	wire [4-1:0] node1435;
	wire [4-1:0] node1436;
	wire [4-1:0] node1440;
	wire [4-1:0] node1441;
	wire [4-1:0] node1442;
	wire [4-1:0] node1443;
	wire [4-1:0] node1444;
	wire [4-1:0] node1448;
	wire [4-1:0] node1451;
	wire [4-1:0] node1454;
	wire [4-1:0] node1455;
	wire [4-1:0] node1459;
	wire [4-1:0] node1460;
	wire [4-1:0] node1461;
	wire [4-1:0] node1464;
	wire [4-1:0] node1467;
	wire [4-1:0] node1468;
	wire [4-1:0] node1470;
	wire [4-1:0] node1471;
	wire [4-1:0] node1475;
	wire [4-1:0] node1477;
	wire [4-1:0] node1480;
	wire [4-1:0] node1482;
	wire [4-1:0] node1483;
	wire [4-1:0] node1484;
	wire [4-1:0] node1485;
	wire [4-1:0] node1488;
	wire [4-1:0] node1490;
	wire [4-1:0] node1493;
	wire [4-1:0] node1494;
	wire [4-1:0] node1495;
	wire [4-1:0] node1497;
	wire [4-1:0] node1501;
	wire [4-1:0] node1502;
	wire [4-1:0] node1503;
	wire [4-1:0] node1506;
	wire [4-1:0] node1510;
	wire [4-1:0] node1512;
	wire [4-1:0] node1513;
	wire [4-1:0] node1514;
	wire [4-1:0] node1516;
	wire [4-1:0] node1519;
	wire [4-1:0] node1520;
	wire [4-1:0] node1521;
	wire [4-1:0] node1526;
	wire [4-1:0] node1527;

	assign outp = (inp[14]) ? node2 : 4'b0000;
		assign node2 = (inp[12]) ? node960 : node3;
			assign node3 = (inp[3]) ? node245 : node4;
				assign node4 = (inp[0]) ? node86 : node5;
					assign node5 = (inp[4]) ? 4'b0000 : node6;
						assign node6 = (inp[7]) ? node52 : node7;
							assign node7 = (inp[11]) ? 4'b0000 : node8;
								assign node8 = (inp[5]) ? node36 : node9;
									assign node9 = (inp[9]) ? 4'b0010 : node10;
										assign node10 = (inp[15]) ? node26 : node11;
											assign node11 = (inp[13]) ? 4'b0010 : node12;
												assign node12 = (inp[1]) ? node18 : node13;
													assign node13 = (inp[8]) ? 4'b0000 : node14;
														assign node14 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node18 = (inp[6]) ? 4'b0010 : node19;
														assign node19 = (inp[8]) ? node21 : 4'b0010;
															assign node21 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node26 = (inp[13]) ? node28 : 4'b0000;
												assign node28 = (inp[10]) ? 4'b0000 : node29;
													assign node29 = (inp[8]) ? node31 : 4'b0010;
														assign node31 = (inp[6]) ? 4'b0010 : 4'b0000;
									assign node36 = (inp[9]) ? node38 : 4'b0000;
										assign node38 = (inp[13]) ? node44 : node39;
											assign node39 = (inp[15]) ? 4'b0000 : node40;
												assign node40 = (inp[1]) ? 4'b0010 : 4'b0000;
											assign node44 = (inp[15]) ? node46 : 4'b0010;
												assign node46 = (inp[10]) ? node48 : 4'b0010;
													assign node48 = (inp[8]) ? 4'b0000 : 4'b0010;
							assign node52 = (inp[11]) ? node54 : 4'b0010;
								assign node54 = (inp[9]) ? node70 : node55;
									assign node55 = (inp[5]) ? 4'b0000 : node56;
										assign node56 = (inp[13]) ? node62 : node57;
											assign node57 = (inp[8]) ? 4'b0000 : node58;
												assign node58 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node62 = (inp[8]) ? node64 : 4'b0010;
												assign node64 = (inp[15]) ? node66 : 4'b0010;
													assign node66 = (inp[2]) ? 4'b0000 : 4'b0010;
									assign node70 = (inp[5]) ? node72 : 4'b0010;
										assign node72 = (inp[15]) ? node78 : node73;
											assign node73 = (inp[8]) ? node75 : 4'b0010;
												assign node75 = (inp[1]) ? 4'b0010 : 4'b0000;
											assign node78 = (inp[13]) ? node80 : 4'b0000;
												assign node80 = (inp[1]) ? 4'b0010 : node81;
													assign node81 = (inp[8]) ? 4'b0000 : 4'b0010;
					assign node86 = (inp[4]) ? node198 : node87;
						assign node87 = (inp[5]) ? node141 : node88;
							assign node88 = (inp[7]) ? node112 : node89;
								assign node89 = (inp[11]) ? node99 : node90;
									assign node90 = (inp[9]) ? 4'b0000 : node91;
										assign node91 = (inp[15]) ? node93 : 4'b0000;
											assign node93 = (inp[13]) ? 4'b0000 : node94;
												assign node94 = (inp[2]) ? 4'b0010 : 4'b0000;
									assign node99 = (inp[9]) ? node101 : 4'b0010;
										assign node101 = (inp[13]) ? 4'b0000 : node102;
											assign node102 = (inp[1]) ? 4'b0000 : node103;
												assign node103 = (inp[15]) ? 4'b0010 : node104;
													assign node104 = (inp[8]) ? node106 : 4'b0000;
														assign node106 = (inp[6]) ? 4'b0000 : 4'b0010;
								assign node112 = (inp[9]) ? node120 : node113;
									assign node113 = (inp[11]) ? 4'b0000 : node114;
										assign node114 = (inp[13]) ? node116 : 4'b0000;
											assign node116 = (inp[15]) ? 4'b0000 : 4'b0010;
									assign node120 = (inp[11]) ? node122 : 4'b0010;
										assign node122 = (inp[13]) ? node130 : node123;
											assign node123 = (inp[1]) ? node125 : 4'b0000;
												assign node125 = (inp[15]) ? 4'b0000 : node126;
													assign node126 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node130 = (inp[15]) ? node132 : 4'b0010;
												assign node132 = (inp[2]) ? 4'b0010 : node133;
													assign node133 = (inp[8]) ? node135 : 4'b0010;
														assign node135 = (inp[1]) ? 4'b0010 : node136;
															assign node136 = (inp[6]) ? 4'b0010 : 4'b0000;
							assign node141 = (inp[7]) ? node169 : node142;
								assign node142 = (inp[11]) ? node160 : node143;
									assign node143 = (inp[9]) ? 4'b0000 : node144;
										assign node144 = (inp[13]) ? node146 : 4'b0010;
											assign node146 = (inp[8]) ? node154 : node147;
												assign node147 = (inp[10]) ? 4'b0000 : node148;
													assign node148 = (inp[2]) ? 4'b0000 : node149;
														assign node149 = (inp[1]) ? 4'b0000 : 4'b0010;
												assign node154 = (inp[15]) ? 4'b0010 : node155;
													assign node155 = (inp[6]) ? 4'b0000 : 4'b0010;
									assign node160 = (inp[13]) ? node162 : 4'b0010;
										assign node162 = (inp[9]) ? node164 : 4'b0010;
											assign node164 = (inp[15]) ? node166 : 4'b0000;
												assign node166 = (inp[10]) ? 4'b0000 : 4'b0010;
								assign node169 = (inp[9]) ? node171 : 4'b0000;
									assign node171 = (inp[13]) ? node179 : node172;
										assign node172 = (inp[11]) ? 4'b0000 : node173;
											assign node173 = (inp[1]) ? 4'b0010 : node174;
												assign node174 = (inp[8]) ? 4'b0000 : 4'b0010;
										assign node179 = (inp[1]) ? node187 : node180;
											assign node180 = (inp[11]) ? node182 : 4'b0010;
												assign node182 = (inp[6]) ? node184 : 4'b0000;
													assign node184 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node187 = (inp[10]) ? 4'b0010 : node188;
												assign node188 = (inp[8]) ? node190 : 4'b0010;
													assign node190 = (inp[15]) ? node192 : 4'b0010;
														assign node192 = (inp[6]) ? 4'b0010 : node193;
															assign node193 = (inp[11]) ? 4'b0000 : 4'b0010;
						assign node198 = (inp[7]) ? node200 : 4'b0010;
							assign node200 = (inp[9]) ? node226 : node201;
								assign node201 = (inp[11]) ? 4'b0010 : node202;
									assign node202 = (inp[13]) ? node214 : node203;
										assign node203 = (inp[5]) ? 4'b0010 : node204;
											assign node204 = (inp[1]) ? node208 : node205;
												assign node205 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node208 = (inp[6]) ? 4'b0000 : node209;
													assign node209 = (inp[2]) ? 4'b0000 : 4'b0010;
										assign node214 = (inp[15]) ? node216 : 4'b0000;
											assign node216 = (inp[5]) ? node218 : 4'b0000;
												assign node218 = (inp[1]) ? node220 : 4'b0010;
													assign node220 = (inp[8]) ? node222 : 4'b0000;
														assign node222 = (inp[10]) ? 4'b0000 : 4'b0010;
								assign node226 = (inp[11]) ? node228 : 4'b0000;
									assign node228 = (inp[5]) ? node236 : node229;
										assign node229 = (inp[13]) ? 4'b0000 : node230;
											assign node230 = (inp[15]) ? node232 : 4'b0000;
												assign node232 = (inp[1]) ? 4'b0000 : 4'b0010;
										assign node236 = (inp[13]) ? node238 : 4'b0010;
											assign node238 = (inp[1]) ? 4'b0000 : node239;
												assign node239 = (inp[15]) ? 4'b0010 : node240;
													assign node240 = (inp[6]) ? 4'b0000 : 4'b0010;
				assign node245 = (inp[0]) ? node327 : node246;
					assign node246 = (inp[4]) ? node248 : 4'b0010;
						assign node248 = (inp[7]) ? node288 : node249;
							assign node249 = (inp[11]) ? 4'b0000 : node250;
								assign node250 = (inp[9]) ? node266 : node251;
									assign node251 = (inp[5]) ? 4'b0000 : node252;
										assign node252 = (inp[15]) ? node260 : node253;
											assign node253 = (inp[13]) ? 4'b0010 : node254;
												assign node254 = (inp[2]) ? 4'b0010 : node255;
													assign node255 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node260 = (inp[13]) ? node262 : 4'b0000;
												assign node262 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node266 = (inp[5]) ? node268 : 4'b0010;
										assign node268 = (inp[1]) ? node282 : node269;
											assign node269 = (inp[13]) ? node277 : node270;
												assign node270 = (inp[10]) ? 4'b0000 : node271;
													assign node271 = (inp[8]) ? 4'b0000 : node272;
														assign node272 = (inp[2]) ? 4'b0010 : 4'b0000;
												assign node277 = (inp[8]) ? node279 : 4'b0010;
													assign node279 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node282 = (inp[2]) ? node284 : 4'b0010;
												assign node284 = (inp[15]) ? 4'b0000 : 4'b0010;
							assign node288 = (inp[11]) ? node290 : 4'b0010;
								assign node290 = (inp[5]) ? node308 : node291;
									assign node291 = (inp[9]) ? 4'b0010 : node292;
										assign node292 = (inp[15]) ? node300 : node293;
											assign node293 = (inp[8]) ? node295 : 4'b0010;
												assign node295 = (inp[1]) ? 4'b0010 : node296;
													assign node296 = (inp[13]) ? 4'b0010 : 4'b0000;
											assign node300 = (inp[13]) ? node302 : 4'b0000;
												assign node302 = (inp[1]) ? 4'b0010 : node303;
													assign node303 = (inp[10]) ? 4'b0010 : 4'b0000;
									assign node308 = (inp[9]) ? node310 : 4'b0000;
										assign node310 = (inp[15]) ? node320 : node311;
											assign node311 = (inp[10]) ? node313 : 4'b0010;
												assign node313 = (inp[1]) ? node315 : 4'b0000;
													assign node315 = (inp[2]) ? node317 : 4'b0010;
														assign node317 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node320 = (inp[8]) ? 4'b0000 : node321;
												assign node321 = (inp[13]) ? node323 : 4'b0000;
													assign node323 = (inp[1]) ? 4'b0010 : 4'b0000;
					assign node327 = (inp[9]) ? node623 : node328;
						assign node328 = (inp[7]) ? node408 : node329;
							assign node329 = (inp[4]) ? node375 : node330;
								assign node330 = (inp[11]) ? node358 : node331;
									assign node331 = (inp[1]) ? node341 : node332;
										assign node332 = (inp[13]) ? 4'b1000 : node333;
											assign node333 = (inp[5]) ? 4'b0010 : node334;
												assign node334 = (inp[6]) ? 4'b1000 : node335;
													assign node335 = (inp[15]) ? 4'b0010 : 4'b1000;
										assign node341 = (inp[13]) ? node349 : node342;
											assign node342 = (inp[15]) ? node344 : 4'b1000;
												assign node344 = (inp[6]) ? 4'b1000 : node345;
													assign node345 = (inp[5]) ? 4'b0010 : 4'b1000;
											assign node349 = (inp[5]) ? 4'b1000 : node350;
												assign node350 = (inp[6]) ? 4'b1010 : node351;
													assign node351 = (inp[15]) ? 4'b1000 : node352;
														assign node352 = (inp[2]) ? 4'b1010 : 4'b1000;
									assign node358 = (inp[13]) ? node360 : 4'b0010;
										assign node360 = (inp[1]) ? node368 : node361;
											assign node361 = (inp[5]) ? 4'b0010 : node362;
												assign node362 = (inp[15]) ? node364 : 4'b1000;
													assign node364 = (inp[6]) ? 4'b1000 : 4'b0010;
											assign node368 = (inp[5]) ? node370 : 4'b1000;
												assign node370 = (inp[6]) ? 4'b1000 : node371;
													assign node371 = (inp[15]) ? 4'b0010 : 4'b1000;
								assign node375 = (inp[11]) ? node397 : node376;
									assign node376 = (inp[13]) ? 4'b0010 : node377;
										assign node377 = (inp[5]) ? node387 : node378;
											assign node378 = (inp[1]) ? 4'b0010 : node379;
												assign node379 = (inp[2]) ? 4'b0000 : node380;
													assign node380 = (inp[6]) ? 4'b0010 : node381;
														assign node381 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node387 = (inp[15]) ? 4'b0000 : node388;
												assign node388 = (inp[10]) ? 4'b0000 : node389;
													assign node389 = (inp[6]) ? 4'b0000 : node390;
														assign node390 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node397 = (inp[1]) ? node399 : 4'b0000;
										assign node399 = (inp[13]) ? node401 : 4'b0000;
											assign node401 = (inp[5]) ? 4'b0000 : node402;
												assign node402 = (inp[6]) ? 4'b0010 : node403;
													assign node403 = (inp[15]) ? 4'b0000 : 4'b0010;
							assign node408 = (inp[13]) ? node516 : node409;
								assign node409 = (inp[4]) ? node473 : node410;
									assign node410 = (inp[1]) ? node438 : node411;
										assign node411 = (inp[11]) ? node423 : node412;
											assign node412 = (inp[2]) ? 4'b0000 : node413;
												assign node413 = (inp[8]) ? node419 : node414;
													assign node414 = (inp[10]) ? 4'b0000 : node415;
														assign node415 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node419 = (inp[5]) ? 4'b1010 : 4'b0000;
											assign node423 = (inp[5]) ? node431 : node424;
												assign node424 = (inp[8]) ? node426 : 4'b1010;
													assign node426 = (inp[6]) ? 4'b1010 : node427;
														assign node427 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node431 = (inp[6]) ? node433 : 4'b1000;
													assign node433 = (inp[10]) ? node435 : 4'b1010;
														assign node435 = (inp[8]) ? 4'b1000 : 4'b1010;
										assign node438 = (inp[8]) ? node454 : node439;
											assign node439 = (inp[6]) ? node449 : node440;
												assign node440 = (inp[5]) ? node444 : node441;
													assign node441 = (inp[11]) ? 4'b0000 : 4'b0010;
													assign node444 = (inp[11]) ? 4'b1010 : node445;
														assign node445 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node449 = (inp[15]) ? 4'b0000 : node450;
													assign node450 = (inp[11]) ? 4'b0000 : 4'b0010;
											assign node454 = (inp[15]) ? node464 : node455;
												assign node455 = (inp[11]) ? 4'b0000 : node456;
													assign node456 = (inp[2]) ? 4'b0010 : node457;
														assign node457 = (inp[5]) ? 4'b0000 : node458;
															assign node458 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node464 = (inp[2]) ? node466 : 4'b0000;
													assign node466 = (inp[10]) ? node468 : 4'b0000;
														assign node468 = (inp[6]) ? 4'b0000 : node469;
															assign node469 = (inp[5]) ? 4'b1010 : 4'b0000;
									assign node473 = (inp[1]) ? node497 : node474;
										assign node474 = (inp[8]) ? node486 : node475;
											assign node475 = (inp[11]) ? node483 : node476;
												assign node476 = (inp[5]) ? node478 : 4'b1000;
													assign node478 = (inp[15]) ? 4'b1010 : node479;
														assign node479 = (inp[6]) ? 4'b1000 : 4'b1010;
												assign node483 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node486 = (inp[5]) ? 4'b1000 : node487;
												assign node487 = (inp[6]) ? 4'b1010 : node488;
													assign node488 = (inp[10]) ? 4'b1000 : node489;
														assign node489 = (inp[11]) ? 4'b1010 : node490;
															assign node490 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node497 = (inp[15]) ? node509 : node498;
											assign node498 = (inp[8]) ? 4'b1010 : node499;
												assign node499 = (inp[11]) ? node505 : node500;
													assign node500 = (inp[5]) ? node502 : 4'b1010;
														assign node502 = (inp[6]) ? 4'b1010 : 4'b1000;
													assign node505 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node509 = (inp[11]) ? 4'b1010 : node510;
												assign node510 = (inp[2]) ? node512 : 4'b1000;
													assign node512 = (inp[5]) ? 4'b1000 : 4'b1010;
								assign node516 = (inp[11]) ? node560 : node517;
									assign node517 = (inp[4]) ? node541 : node518;
										assign node518 = (inp[1]) ? node534 : node519;
											assign node519 = (inp[8]) ? node525 : node520;
												assign node520 = (inp[5]) ? node522 : 4'b1000;
													assign node522 = (inp[6]) ? 4'b0010 : 4'b0000;
												assign node525 = (inp[10]) ? node527 : 4'b0010;
													assign node527 = (inp[5]) ? node531 : node528;
														assign node528 = (inp[6]) ? 4'b1000 : 4'b0010;
														assign node531 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node534 = (inp[5]) ? 4'b1000 : node535;
												assign node535 = (inp[15]) ? 4'b1010 : node536;
													assign node536 = (inp[8]) ? 4'b1010 : 4'b1000;
										assign node541 = (inp[5]) ? node555 : node542;
											assign node542 = (inp[6]) ? node548 : node543;
												assign node543 = (inp[2]) ? 4'b0000 : node544;
													assign node544 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node548 = (inp[8]) ? node550 : 4'b0010;
													assign node550 = (inp[1]) ? 4'b0010 : node551;
														assign node551 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node555 = (inp[6]) ? 4'b0000 : node556;
												assign node556 = (inp[1]) ? 4'b0010 : 4'b1010;
									assign node560 = (inp[4]) ? node590 : node561;
										assign node561 = (inp[1]) ? node575 : node562;
											assign node562 = (inp[6]) ? node570 : node563;
												assign node563 = (inp[2]) ? node565 : 4'b0010;
													assign node565 = (inp[5]) ? node567 : 4'b0010;
														assign node567 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node570 = (inp[2]) ? node572 : 4'b0000;
													assign node572 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node575 = (inp[2]) ? node585 : node576;
												assign node576 = (inp[15]) ? node582 : node577;
													assign node577 = (inp[5]) ? 4'b1000 : node578;
														assign node578 = (inp[6]) ? 4'b1010 : 4'b1000;
													assign node582 = (inp[6]) ? 4'b1010 : 4'b0010;
												assign node585 = (inp[6]) ? 4'b1000 : node586;
													assign node586 = (inp[5]) ? 4'b0010 : 4'b1000;
										assign node590 = (inp[1]) ? node616 : node591;
											assign node591 = (inp[5]) ? node599 : node592;
												assign node592 = (inp[6]) ? 4'b1010 : node593;
													assign node593 = (inp[8]) ? 4'b1000 : node594;
														assign node594 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node599 = (inp[2]) ? 4'b1000 : node600;
													assign node600 = (inp[10]) ? node610 : node601;
														assign node601 = (inp[8]) ? node605 : node602;
															assign node602 = (inp[6]) ? 4'b1010 : 4'b1000;
															assign node605 = (inp[15]) ? node607 : 4'b1000;
																assign node607 = (inp[6]) ? 4'b1000 : 4'b1010;
														assign node610 = (inp[8]) ? node612 : 4'b1010;
															assign node612 = (inp[6]) ? 4'b1000 : 4'b1010;
											assign node616 = (inp[5]) ? node620 : node617;
												assign node617 = (inp[6]) ? 4'b0010 : 4'b0000;
												assign node620 = (inp[6]) ? 4'b0000 : 4'b1010;
						assign node623 = (inp[7]) ? node751 : node624;
							assign node624 = (inp[4]) ? node696 : node625;
								assign node625 = (inp[11]) ? node667 : node626;
									assign node626 = (inp[13]) ? node646 : node627;
										assign node627 = (inp[2]) ? node635 : node628;
											assign node628 = (inp[5]) ? 4'b1010 : node629;
												assign node629 = (inp[1]) ? node631 : 4'b1010;
													assign node631 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node635 = (inp[1]) ? node643 : node636;
												assign node636 = (inp[6]) ? 4'b1010 : node637;
													assign node637 = (inp[5]) ? node639 : 4'b1010;
														assign node639 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node643 = (inp[5]) ? 4'b1010 : 4'b1000;
										assign node646 = (inp[1]) ? node658 : node647;
											assign node647 = (inp[8]) ? node651 : node648;
												assign node648 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node651 = (inp[15]) ? node653 : 4'b1000;
													assign node653 = (inp[6]) ? 4'b1000 : node654;
														assign node654 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node658 = (inp[5]) ? node660 : 4'b1010;
												assign node660 = (inp[6]) ? 4'b1010 : node661;
													assign node661 = (inp[8]) ? 4'b1000 : node662;
														assign node662 = (inp[2]) ? 4'b1000 : 4'b1010;
									assign node667 = (inp[13]) ? node683 : node668;
										assign node668 = (inp[1]) ? node678 : node669;
											assign node669 = (inp[2]) ? node671 : 4'b1000;
												assign node671 = (inp[8]) ? 4'b1000 : node672;
													assign node672 = (inp[15]) ? 4'b1000 : node673;
														assign node673 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node678 = (inp[15]) ? node680 : 4'b1010;
												assign node680 = (inp[5]) ? 4'b1000 : 4'b1010;
										assign node683 = (inp[1]) ? node691 : node684;
											assign node684 = (inp[15]) ? 4'b1010 : node685;
												assign node685 = (inp[6]) ? node687 : 4'b1010;
													assign node687 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node691 = (inp[6]) ? 4'b1000 : node692;
												assign node692 = (inp[5]) ? 4'b1010 : 4'b1000;
								assign node696 = (inp[13]) ? node720 : node697;
									assign node697 = (inp[11]) ? node713 : node698;
										assign node698 = (inp[5]) ? node706 : node699;
											assign node699 = (inp[1]) ? 4'b1000 : node700;
												assign node700 = (inp[6]) ? 4'b1000 : node701;
													assign node701 = (inp[15]) ? 4'b0010 : 4'b1000;
											assign node706 = (inp[1]) ? node708 : 4'b0010;
												assign node708 = (inp[6]) ? 4'b1000 : node709;
													assign node709 = (inp[15]) ? 4'b0010 : 4'b1000;
										assign node713 = (inp[1]) ? 4'b0010 : node714;
											assign node714 = (inp[6]) ? 4'b0010 : node715;
												assign node715 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node720 = (inp[11]) ? node736 : node721;
										assign node721 = (inp[1]) ? node731 : node722;
											assign node722 = (inp[6]) ? node724 : 4'b1000;
												assign node724 = (inp[5]) ? 4'b1000 : node725;
													assign node725 = (inp[10]) ? node727 : 4'b1010;
														assign node727 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node731 = (inp[5]) ? node733 : 4'b1010;
												assign node733 = (inp[6]) ? 4'b1010 : 4'b1000;
										assign node736 = (inp[5]) ? node744 : node737;
											assign node737 = (inp[15]) ? node739 : 4'b1000;
												assign node739 = (inp[1]) ? 4'b1000 : node740;
													assign node740 = (inp[10]) ? 4'b1000 : 4'b0010;
											assign node744 = (inp[1]) ? node746 : 4'b0010;
												assign node746 = (inp[6]) ? 4'b1000 : node747;
													assign node747 = (inp[15]) ? 4'b0010 : 4'b1000;
							assign node751 = (inp[13]) ? node869 : node752;
								assign node752 = (inp[4]) ? node820 : node753;
									assign node753 = (inp[15]) ? node783 : node754;
										assign node754 = (inp[1]) ? node772 : node755;
											assign node755 = (inp[6]) ? node761 : node756;
												assign node756 = (inp[11]) ? node758 : 4'b0001;
													assign node758 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node761 = (inp[11]) ? node767 : node762;
													assign node762 = (inp[2]) ? node764 : 4'b0011;
														assign node764 = (inp[8]) ? 4'b1001 : 4'b1011;
													assign node767 = (inp[2]) ? 4'b0001 : node768;
														assign node768 = (inp[5]) ? 4'b0011 : 4'b0001;
											assign node772 = (inp[6]) ? node780 : node773;
												assign node773 = (inp[5]) ? node777 : node774;
													assign node774 = (inp[11]) ? 4'b1011 : 4'b0011;
													assign node777 = (inp[11]) ? 4'b1001 : 4'b1011;
												assign node780 = (inp[11]) ? 4'b0011 : 4'b1011;
										assign node783 = (inp[8]) ? node801 : node784;
											assign node784 = (inp[1]) ? node794 : node785;
												assign node785 = (inp[11]) ? node791 : node786;
													assign node786 = (inp[10]) ? node788 : 4'b0011;
														assign node788 = (inp[6]) ? 4'b0011 : 4'b0001;
													assign node791 = (inp[6]) ? 4'b0001 : 4'b1000;
												assign node794 = (inp[6]) ? node798 : node795;
													assign node795 = (inp[11]) ? 4'b0011 : 4'b0001;
													assign node798 = (inp[11]) ? 4'b0001 : 4'b1001;
											assign node801 = (inp[11]) ? node809 : node802;
												assign node802 = (inp[6]) ? 4'b1001 : node803;
													assign node803 = (inp[10]) ? node805 : 4'b0001;
														assign node805 = (inp[1]) ? 4'b0001 : 4'b0011;
												assign node809 = (inp[6]) ? node815 : node810;
													assign node810 = (inp[2]) ? 4'b1010 : node811;
														assign node811 = (inp[10]) ? 4'b1001 : 4'b1011;
													assign node815 = (inp[1]) ? 4'b0001 : node816;
														assign node816 = (inp[5]) ? 4'b0001 : 4'b0011;
									assign node820 = (inp[1]) ? node842 : node821;
										assign node821 = (inp[11]) ? node831 : node822;
											assign node822 = (inp[15]) ? node826 : node823;
												assign node823 = (inp[10]) ? 4'b1010 : 4'b1000;
												assign node826 = (inp[6]) ? 4'b1010 : node827;
													assign node827 = (inp[5]) ? 4'b0010 : 4'b1000;
											assign node831 = (inp[5]) ? node837 : node832;
												assign node832 = (inp[6]) ? node834 : 4'b0000;
													assign node834 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node837 = (inp[15]) ? node839 : 4'b0010;
													assign node839 = (inp[6]) ? 4'b0000 : 4'b0010;
										assign node842 = (inp[15]) ? node854 : node843;
											assign node843 = (inp[2]) ? node849 : node844;
												assign node844 = (inp[11]) ? 4'b0011 : node845;
													assign node845 = (inp[6]) ? 4'b1011 : 4'b0011;
												assign node849 = (inp[11]) ? 4'b1010 : node850;
													assign node850 = (inp[6]) ? 4'b1011 : 4'b0001;
											assign node854 = (inp[6]) ? node866 : node855;
												assign node855 = (inp[11]) ? node859 : node856;
													assign node856 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node859 = (inp[5]) ? node861 : 4'b1000;
														assign node861 = (inp[8]) ? node863 : 4'b1010;
															assign node863 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node866 = (inp[11]) ? 4'b0001 : 4'b1001;
								assign node869 = (inp[6]) ? node943 : node870;
									assign node870 = (inp[1]) ? node928 : node871;
										assign node871 = (inp[4]) ? node901 : node872;
											assign node872 = (inp[2]) ? node888 : node873;
												assign node873 = (inp[10]) ? node881 : node874;
													assign node874 = (inp[11]) ? node878 : node875;
														assign node875 = (inp[8]) ? 4'b1010 : 4'b1000;
														assign node878 = (inp[15]) ? 4'b0000 : 4'b1000;
													assign node881 = (inp[15]) ? 4'b0010 : node882;
														assign node882 = (inp[11]) ? 4'b1000 : node883;
															assign node883 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node888 = (inp[10]) ? node898 : node889;
													assign node889 = (inp[11]) ? node891 : 4'b0000;
														assign node891 = (inp[15]) ? node893 : 4'b1010;
															assign node893 = (inp[8]) ? node895 : 4'b0010;
																assign node895 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node898 = (inp[11]) ? 4'b0000 : 4'b1000;
											assign node901 = (inp[11]) ? node913 : node902;
												assign node902 = (inp[8]) ? node910 : node903;
													assign node903 = (inp[15]) ? node907 : node904;
														assign node904 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node907 = (inp[10]) ? 4'b0011 : 4'b1001;
													assign node910 = (inp[5]) ? 4'b0011 : 4'b1011;
												assign node913 = (inp[5]) ? 4'b1011 : node914;
													assign node914 = (inp[10]) ? 4'b0001 : node915;
														assign node915 = (inp[2]) ? node921 : node916;
															assign node916 = (inp[15]) ? node918 : 4'b0001;
																assign node918 = (inp[8]) ? 4'b0001 : 4'b0011;
															assign node921 = (inp[15]) ? 4'b0001 : node922;
																assign node922 = (inp[8]) ? 4'b0011 : 4'b0001;
										assign node928 = (inp[15]) ? node936 : node929;
											assign node929 = (inp[10]) ? node933 : node930;
												assign node930 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node933 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node936 = (inp[10]) ? node940 : node937;
												assign node937 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node940 = (inp[11]) ? 4'b0100 : 4'b0101;
									assign node943 = (inp[1]) ? 4'b0000 : node944;
										assign node944 = (inp[8]) ? node952 : node945;
											assign node945 = (inp[4]) ? node949 : node946;
												assign node946 = (inp[5]) ? 4'b0011 : 4'b1011;
												assign node949 = (inp[5]) ? 4'b0010 : 4'b1010;
											assign node952 = (inp[5]) ? node956 : node953;
												assign node953 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node956 = (inp[4]) ? 4'b0000 : 4'b0001;
			assign node960 = (inp[0]) ? node962 : 4'b0000;
				assign node962 = (inp[4]) ? node1330 : node963;
					assign node963 = (inp[7]) ? node1075 : node964;
						assign node964 = (inp[3]) ? node988 : node965;
							assign node965 = (inp[11]) ? 4'b0000 : node966;
								assign node966 = (inp[5]) ? node974 : node967;
									assign node967 = (inp[9]) ? 4'b0010 : node968;
										assign node968 = (inp[15]) ? node970 : 4'b0010;
											assign node970 = (inp[13]) ? 4'b0010 : 4'b0000;
									assign node974 = (inp[9]) ? node976 : 4'b0000;
										assign node976 = (inp[15]) ? node982 : node977;
											assign node977 = (inp[13]) ? 4'b0010 : node978;
												assign node978 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node982 = (inp[13]) ? node984 : 4'b0000;
												assign node984 = (inp[10]) ? 4'b0000 : 4'b0010;
							assign node988 = (inp[9]) ? node1016 : node989;
								assign node989 = (inp[11]) ? 4'b0010 : node990;
									assign node990 = (inp[5]) ? node998 : node991;
										assign node991 = (inp[6]) ? 4'b0000 : node992;
											assign node992 = (inp[13]) ? 4'b0000 : node993;
												assign node993 = (inp[1]) ? 4'b0000 : 4'b0010;
										assign node998 = (inp[13]) ? node1000 : 4'b0010;
											assign node1000 = (inp[15]) ? node1008 : node1001;
												assign node1001 = (inp[6]) ? 4'b0000 : node1002;
													assign node1002 = (inp[1]) ? 4'b0000 : node1003;
														assign node1003 = (inp[8]) ? 4'b0010 : 4'b0000;
												assign node1008 = (inp[1]) ? node1010 : 4'b0010;
													assign node1010 = (inp[8]) ? node1012 : 4'b0000;
														assign node1012 = (inp[6]) ? 4'b0000 : 4'b0010;
								assign node1016 = (inp[1]) ? node1046 : node1017;
									assign node1017 = (inp[11]) ? node1029 : node1018;
										assign node1018 = (inp[5]) ? 4'b0000 : node1019;
											assign node1019 = (inp[13]) ? node1021 : 4'b0000;
												assign node1021 = (inp[6]) ? 4'b0010 : node1022;
													assign node1022 = (inp[15]) ? node1024 : 4'b0010;
														assign node1024 = (inp[8]) ? 4'b0000 : 4'b0010;
										assign node1029 = (inp[13]) ? node1039 : node1030;
											assign node1030 = (inp[5]) ? 4'b0010 : node1031;
												assign node1031 = (inp[6]) ? 4'b0000 : node1032;
													assign node1032 = (inp[8]) ? 4'b0010 : node1033;
														assign node1033 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node1039 = (inp[6]) ? 4'b0000 : node1040;
												assign node1040 = (inp[5]) ? node1042 : 4'b0000;
													assign node1042 = (inp[8]) ? 4'b0010 : 4'b0000;
									assign node1046 = (inp[11]) ? node1066 : node1047;
										assign node1047 = (inp[13]) ? node1057 : node1048;
											assign node1048 = (inp[8]) ? 4'b0000 : node1049;
												assign node1049 = (inp[15]) ? 4'b0000 : node1050;
													assign node1050 = (inp[6]) ? 4'b0010 : node1051;
														assign node1051 = (inp[10]) ? 4'b0000 : 4'b0010;
											assign node1057 = (inp[6]) ? 4'b0010 : node1058;
												assign node1058 = (inp[8]) ? node1060 : 4'b0010;
													assign node1060 = (inp[2]) ? 4'b0010 : node1061;
														assign node1061 = (inp[10]) ? 4'b0000 : 4'b0010;
										assign node1066 = (inp[13]) ? 4'b0000 : node1067;
											assign node1067 = (inp[5]) ? 4'b0010 : node1068;
												assign node1068 = (inp[8]) ? node1070 : 4'b0000;
													assign node1070 = (inp[10]) ? 4'b0010 : 4'b0000;
						assign node1075 = (inp[3]) ? node1123 : node1076;
							assign node1076 = (inp[11]) ? node1078 : 4'b0010;
								assign node1078 = (inp[5]) ? node1100 : node1079;
									assign node1079 = (inp[9]) ? 4'b0010 : node1080;
										assign node1080 = (inp[8]) ? node1086 : node1081;
											assign node1081 = (inp[13]) ? 4'b0010 : node1082;
												assign node1082 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node1086 = (inp[1]) ? node1092 : node1087;
												assign node1087 = (inp[13]) ? node1089 : 4'b0000;
													assign node1089 = (inp[10]) ? 4'b0010 : 4'b0000;
												assign node1092 = (inp[6]) ? 4'b0010 : node1093;
													assign node1093 = (inp[2]) ? 4'b0000 : node1094;
														assign node1094 = (inp[13]) ? 4'b0010 : 4'b0000;
									assign node1100 = (inp[9]) ? node1102 : 4'b0000;
										assign node1102 = (inp[15]) ? node1112 : node1103;
											assign node1103 = (inp[2]) ? node1105 : 4'b0010;
												assign node1105 = (inp[6]) ? 4'b0010 : node1106;
													assign node1106 = (inp[8]) ? node1108 : 4'b0010;
														assign node1108 = (inp[13]) ? 4'b0010 : 4'b0000;
											assign node1112 = (inp[13]) ? node1114 : 4'b0000;
												assign node1114 = (inp[1]) ? 4'b0010 : node1115;
													assign node1115 = (inp[8]) ? 4'b0000 : node1116;
														assign node1116 = (inp[10]) ? node1118 : 4'b0010;
															assign node1118 = (inp[6]) ? 4'b0010 : 4'b0000;
							assign node1123 = (inp[13]) ? node1235 : node1124;
								assign node1124 = (inp[10]) ? node1174 : node1125;
									assign node1125 = (inp[9]) ? node1143 : node1126;
										assign node1126 = (inp[11]) ? node1140 : node1127;
											assign node1127 = (inp[1]) ? node1133 : node1128;
												assign node1128 = (inp[5]) ? 4'b0010 : node1129;
													assign node1129 = (inp[15]) ? 4'b0010 : 4'b1000;
												assign node1133 = (inp[8]) ? node1135 : 4'b1000;
													assign node1135 = (inp[6]) ? node1137 : 4'b0010;
														assign node1137 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node1140 = (inp[5]) ? 4'b0000 : 4'b0010;
										assign node1143 = (inp[1]) ? node1163 : node1144;
											assign node1144 = (inp[11]) ? node1148 : node1145;
												assign node1145 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node1148 = (inp[8]) ? node1158 : node1149;
													assign node1149 = (inp[5]) ? node1153 : node1150;
														assign node1150 = (inp[6]) ? 4'b1010 : 4'b1000;
														assign node1153 = (inp[6]) ? node1155 : 4'b1010;
															assign node1155 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node1158 = (inp[2]) ? node1160 : 4'b1000;
														assign node1160 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node1163 = (inp[15]) ? node1171 : node1164;
												assign node1164 = (inp[11]) ? node1168 : node1165;
													assign node1165 = (inp[6]) ? 4'b1010 : 4'b0010;
													assign node1168 = (inp[5]) ? 4'b1010 : 4'b0010;
												assign node1171 = (inp[11]) ? 4'b0000 : 4'b1000;
									assign node1174 = (inp[11]) ? node1212 : node1175;
										assign node1175 = (inp[1]) ? node1195 : node1176;
											assign node1176 = (inp[5]) ? node1188 : node1177;
												assign node1177 = (inp[9]) ? node1183 : node1178;
													assign node1178 = (inp[6]) ? 4'b1000 : node1179;
														assign node1179 = (inp[2]) ? 4'b1000 : 4'b0010;
													assign node1183 = (inp[15]) ? node1185 : 4'b0000;
														assign node1185 = (inp[2]) ? 4'b0000 : 4'b0010;
												assign node1188 = (inp[9]) ? node1190 : 4'b0010;
													assign node1190 = (inp[15]) ? node1192 : 4'b0010;
														assign node1192 = (inp[2]) ? 4'b0000 : 4'b1000;
											assign node1195 = (inp[9]) ? node1201 : node1196;
												assign node1196 = (inp[6]) ? node1198 : 4'b1000;
													assign node1198 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node1201 = (inp[6]) ? node1209 : node1202;
													assign node1202 = (inp[15]) ? node1206 : node1203;
														assign node1203 = (inp[5]) ? 4'b0000 : 4'b1000;
														assign node1206 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node1209 = (inp[8]) ? 4'b1010 : 4'b1000;
										assign node1212 = (inp[1]) ? node1220 : node1213;
											assign node1213 = (inp[9]) ? node1215 : 4'b0000;
												assign node1215 = (inp[6]) ? 4'b1010 : node1216;
													assign node1216 = (inp[2]) ? 4'b1010 : 4'b1000;
											assign node1220 = (inp[15]) ? node1230 : node1221;
												assign node1221 = (inp[6]) ? 4'b0010 : node1222;
													assign node1222 = (inp[2]) ? 4'b0000 : node1223;
														assign node1223 = (inp[9]) ? 4'b1010 : node1224;
															assign node1224 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node1230 = (inp[5]) ? 4'b0000 : node1231;
													assign node1231 = (inp[9]) ? 4'b0000 : 4'b0010;
								assign node1235 = (inp[9]) ? node1285 : node1236;
									assign node1236 = (inp[11]) ? node1266 : node1237;
										assign node1237 = (inp[2]) ? node1245 : node1238;
											assign node1238 = (inp[6]) ? node1240 : 4'b1010;
												assign node1240 = (inp[8]) ? 4'b1010 : node1241;
													assign node1241 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node1245 = (inp[8]) ? node1255 : node1246;
												assign node1246 = (inp[15]) ? 4'b1010 : node1247;
													assign node1247 = (inp[5]) ? 4'b1000 : node1248;
														assign node1248 = (inp[10]) ? 4'b1000 : node1249;
															assign node1249 = (inp[1]) ? 4'b1010 : 4'b1000;
												assign node1255 = (inp[15]) ? node1257 : 4'b1010;
													assign node1257 = (inp[6]) ? node1263 : node1258;
														assign node1258 = (inp[5]) ? node1260 : 4'b1000;
															assign node1260 = (inp[1]) ? 4'b1010 : 4'b1000;
														assign node1263 = (inp[5]) ? 4'b1000 : 4'b1010;
										assign node1266 = (inp[5]) ? node1278 : node1267;
											assign node1267 = (inp[1]) ? node1273 : node1268;
												assign node1268 = (inp[15]) ? node1270 : 4'b1000;
													assign node1270 = (inp[10]) ? 4'b0010 : 4'b1000;
												assign node1273 = (inp[15]) ? node1275 : 4'b1010;
													assign node1275 = (inp[6]) ? 4'b1010 : 4'b1000;
											assign node1278 = (inp[1]) ? node1280 : 4'b0010;
												assign node1280 = (inp[6]) ? 4'b1000 : node1281;
													assign node1281 = (inp[15]) ? 4'b0010 : 4'b1000;
									assign node1285 = (inp[1]) ? node1313 : node1286;
										assign node1286 = (inp[5]) ? node1300 : node1287;
											assign node1287 = (inp[6]) ? node1297 : node1288;
												assign node1288 = (inp[11]) ? node1294 : node1289;
													assign node1289 = (inp[15]) ? 4'b0001 : node1290;
														assign node1290 = (inp[10]) ? 4'b1001 : 4'b1011;
													assign node1294 = (inp[2]) ? 4'b1000 : 4'b1010;
												assign node1297 = (inp[8]) ? 4'b1001 : 4'b1011;
											assign node1300 = (inp[6]) ? node1310 : node1301;
												assign node1301 = (inp[11]) ? node1305 : node1302;
													assign node1302 = (inp[10]) ? 4'b0001 : 4'b0011;
													assign node1305 = (inp[10]) ? 4'b1000 : node1306;
														assign node1306 = (inp[15]) ? 4'b0010 : 4'b1010;
												assign node1310 = (inp[8]) ? 4'b0001 : 4'b0011;
										assign node1313 = (inp[6]) ? 4'b0000 : node1314;
											assign node1314 = (inp[15]) ? node1322 : node1315;
												assign node1315 = (inp[11]) ? node1319 : node1316;
													assign node1316 = (inp[10]) ? 4'b1001 : 4'b1011;
													assign node1319 = (inp[10]) ? 4'b1000 : 4'b1010;
												assign node1322 = (inp[11]) ? node1326 : node1323;
													assign node1323 = (inp[10]) ? 4'b0001 : 4'b0011;
													assign node1326 = (inp[10]) ? 4'b0000 : 4'b0010;
					assign node1330 = (inp[3]) ? node1332 : 4'b0000;
						assign node1332 = (inp[11]) ? node1480 : node1333;
							assign node1333 = (inp[9]) ? node1401 : node1334;
								assign node1334 = (inp[7]) ? node1354 : node1335;
									assign node1335 = (inp[5]) ? 4'b0000 : node1336;
										assign node1336 = (inp[13]) ? node1344 : node1337;
											assign node1337 = (inp[8]) ? 4'b0000 : node1338;
												assign node1338 = (inp[15]) ? 4'b0000 : node1339;
													assign node1339 = (inp[1]) ? 4'b0010 : 4'b0000;
											assign node1344 = (inp[15]) ? node1346 : 4'b0010;
												assign node1346 = (inp[1]) ? 4'b0010 : node1347;
													assign node1347 = (inp[6]) ? node1349 : 4'b0000;
														assign node1349 = (inp[8]) ? 4'b0000 : 4'b0010;
									assign node1354 = (inp[5]) ? node1384 : node1355;
										assign node1355 = (inp[15]) ? node1363 : node1356;
											assign node1356 = (inp[13]) ? node1358 : 4'b0000;
												assign node1358 = (inp[1]) ? 4'b0010 : node1359;
													assign node1359 = (inp[8]) ? 4'b0000 : 4'b0010;
											assign node1363 = (inp[10]) ? node1373 : node1364;
												assign node1364 = (inp[2]) ? node1366 : 4'b0010;
													assign node1366 = (inp[6]) ? node1370 : node1367;
														assign node1367 = (inp[13]) ? 4'b0010 : 4'b0000;
														assign node1370 = (inp[13]) ? 4'b0000 : 4'b0010;
												assign node1373 = (inp[6]) ? node1375 : 4'b0010;
													assign node1375 = (inp[2]) ? node1377 : 4'b0000;
														assign node1377 = (inp[13]) ? node1381 : node1378;
															assign node1378 = (inp[1]) ? 4'b0000 : 4'b0010;
															assign node1381 = (inp[1]) ? 4'b0010 : 4'b0000;
										assign node1384 = (inp[13]) ? node1386 : 4'b0010;
											assign node1386 = (inp[15]) ? node1394 : node1387;
												assign node1387 = (inp[2]) ? node1389 : 4'b0000;
													assign node1389 = (inp[1]) ? 4'b0000 : node1390;
														assign node1390 = (inp[6]) ? 4'b0000 : 4'b0010;
												assign node1394 = (inp[1]) ? node1396 : 4'b0010;
													assign node1396 = (inp[10]) ? 4'b0000 : node1397;
														assign node1397 = (inp[6]) ? 4'b0000 : 4'b0010;
								assign node1401 = (inp[7]) ? node1421 : node1402;
									assign node1402 = (inp[5]) ? node1404 : 4'b0010;
										assign node1404 = (inp[1]) ? node1416 : node1405;
											assign node1405 = (inp[13]) ? node1413 : node1406;
												assign node1406 = (inp[8]) ? 4'b0000 : node1407;
													assign node1407 = (inp[6]) ? node1409 : 4'b0000;
														assign node1409 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node1413 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node1416 = (inp[15]) ? node1418 : 4'b0010;
												assign node1418 = (inp[13]) ? 4'b0010 : 4'b0000;
									assign node1421 = (inp[15]) ? node1459 : node1422;
										assign node1422 = (inp[13]) ? node1440 : node1423;
											assign node1423 = (inp[1]) ? node1435 : node1424;
												assign node1424 = (inp[5]) ? node1430 : node1425;
													assign node1425 = (inp[8]) ? 4'b1000 : node1426;
														assign node1426 = (inp[6]) ? 4'b1010 : 4'b1000;
													assign node1430 = (inp[6]) ? 4'b0010 : node1431;
														assign node1431 = (inp[10]) ? 4'b0000 : 4'b0010;
												assign node1435 = (inp[6]) ? 4'b1010 : node1436;
													assign node1436 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node1440 = (inp[1]) ? node1454 : node1441;
												assign node1441 = (inp[8]) ? node1451 : node1442;
													assign node1442 = (inp[2]) ? node1448 : node1443;
														assign node1443 = (inp[10]) ? 4'b1010 : node1444;
															assign node1444 = (inp[5]) ? 4'b1010 : 4'b0000;
														assign node1448 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node1451 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node1454 = (inp[6]) ? 4'b0000 : node1455;
													assign node1455 = (inp[2]) ? 4'b1001 : 4'b1011;
										assign node1459 = (inp[6]) ? node1467 : node1460;
											assign node1460 = (inp[13]) ? node1464 : node1461;
												assign node1461 = (inp[1]) ? 4'b0010 : 4'b0000;
												assign node1464 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node1467 = (inp[5]) ? node1475 : node1468;
												assign node1468 = (inp[13]) ? node1470 : 4'b1000;
													assign node1470 = (inp[1]) ? 4'b0000 : node1471;
														assign node1471 = (inp[8]) ? 4'b1000 : 4'b1010;
												assign node1475 = (inp[8]) ? node1477 : 4'b0010;
													assign node1477 = (inp[1]) ? 4'b1000 : 4'b0000;
							assign node1480 = (inp[7]) ? node1482 : 4'b0000;
								assign node1482 = (inp[5]) ? node1510 : node1483;
									assign node1483 = (inp[13]) ? node1493 : node1484;
										assign node1484 = (inp[15]) ? node1488 : node1485;
											assign node1485 = (inp[1]) ? 4'b0010 : 4'b0000;
											assign node1488 = (inp[9]) ? node1490 : 4'b0000;
												assign node1490 = (inp[10]) ? 4'b0010 : 4'b0000;
										assign node1493 = (inp[9]) ? node1501 : node1494;
											assign node1494 = (inp[1]) ? 4'b0010 : node1495;
												assign node1495 = (inp[15]) ? node1497 : 4'b0010;
													assign node1497 = (inp[6]) ? 4'b0010 : 4'b0000;
											assign node1501 = (inp[1]) ? 4'b0000 : node1502;
												assign node1502 = (inp[6]) ? node1506 : node1503;
													assign node1503 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node1506 = (inp[2]) ? 4'b1010 : 4'b1000;
									assign node1510 = (inp[9]) ? node1512 : 4'b0000;
										assign node1512 = (inp[15]) ? node1526 : node1513;
											assign node1513 = (inp[13]) ? node1519 : node1514;
												assign node1514 = (inp[8]) ? node1516 : 4'b0010;
													assign node1516 = (inp[1]) ? 4'b0010 : 4'b0000;
												assign node1519 = (inp[1]) ? 4'b1000 : node1520;
													assign node1520 = (inp[6]) ? 4'b0000 : node1521;
														assign node1521 = (inp[8]) ? 4'b0010 : 4'b0000;
											assign node1526 = (inp[10]) ? 4'b0000 : node1527;
												assign node1527 = (inp[1]) ? 4'b0010 : 4'b0000;

endmodule