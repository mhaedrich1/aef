module dtc_split66_bm56 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node215;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node232;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node243;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node317;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node333;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node344;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node354;
	wire [3-1:0] node357;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node363;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node376;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node392;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node401;
	wire [3-1:0] node403;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node409;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node425;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node433;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node443;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node450;
	wire [3-1:0] node454;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node486;
	wire [3-1:0] node488;
	wire [3-1:0] node490;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node501;
	wire [3-1:0] node503;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node510;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node537;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node544;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node551;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node561;
	wire [3-1:0] node564;
	wire [3-1:0] node566;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node573;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node591;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node597;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node604;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node620;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node628;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node635;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node644;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node652;
	wire [3-1:0] node655;
	wire [3-1:0] node657;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node664;
	wire [3-1:0] node666;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node676;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node684;
	wire [3-1:0] node686;
	wire [3-1:0] node689;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node696;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node703;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node716;
	wire [3-1:0] node719;
	wire [3-1:0] node721;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node736;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node743;
	wire [3-1:0] node746;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node766;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node774;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node785;
	wire [3-1:0] node788;
	wire [3-1:0] node790;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node796;
	wire [3-1:0] node799;
	wire [3-1:0] node801;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node809;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node814;
	wire [3-1:0] node815;
	wire [3-1:0] node818;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node825;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node831;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node840;
	wire [3-1:0] node843;
	wire [3-1:0] node845;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node851;
	wire [3-1:0] node854;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node864;
	wire [3-1:0] node867;
	wire [3-1:0] node868;
	wire [3-1:0] node869;
	wire [3-1:0] node871;
	wire [3-1:0] node874;
	wire [3-1:0] node876;
	wire [3-1:0] node879;
	wire [3-1:0] node881;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node897;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node904;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node911;
	wire [3-1:0] node914;
	wire [3-1:0] node916;
	wire [3-1:0] node919;
	wire [3-1:0] node921;
	wire [3-1:0] node923;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node931;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node938;
	wire [3-1:0] node941;
	wire [3-1:0] node943;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node950;
	wire [3-1:0] node953;
	wire [3-1:0] node955;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node961;
	wire [3-1:0] node964;
	wire [3-1:0] node967;
	wire [3-1:0] node968;
	wire [3-1:0] node969;
	wire [3-1:0] node970;
	wire [3-1:0] node971;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node976;
	wire [3-1:0] node979;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node985;
	wire [3-1:0] node988;
	wire [3-1:0] node990;
	wire [3-1:0] node993;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node1000;
	wire [3-1:0] node1001;
	wire [3-1:0] node1002;
	wire [3-1:0] node1007;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1012;
	wire [3-1:0] node1015;
	wire [3-1:0] node1016;
	wire [3-1:0] node1017;
	wire [3-1:0] node1020;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1031;
	wire [3-1:0] node1034;
	wire [3-1:0] node1035;
	wire [3-1:0] node1036;
	wire [3-1:0] node1039;
	wire [3-1:0] node1043;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1048;
	wire [3-1:0] node1051;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1056;
	wire [3-1:0] node1060;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1064;
	wire [3-1:0] node1065;
	wire [3-1:0] node1069;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1074;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1081;
	wire [3-1:0] node1084;
	wire [3-1:0] node1085;
	wire [3-1:0] node1088;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1095;
	wire [3-1:0] node1098;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1104;
	wire [3-1:0] node1105;
	wire [3-1:0] node1108;
	wire [3-1:0] node1111;
	wire [3-1:0] node1112;
	wire [3-1:0] node1113;
	wire [3-1:0] node1116;
	wire [3-1:0] node1119;
	wire [3-1:0] node1121;
	wire [3-1:0] node1124;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1131;
	wire [3-1:0] node1132;
	wire [3-1:0] node1135;
	wire [3-1:0] node1137;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1142;
	wire [3-1:0] node1146;
	wire [3-1:0] node1147;
	wire [3-1:0] node1148;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1155;
	wire [3-1:0] node1156;
	wire [3-1:0] node1157;
	wire [3-1:0] node1158;
	wire [3-1:0] node1161;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1167;
	wire [3-1:0] node1171;
	wire [3-1:0] node1174;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1179;
	wire [3-1:0] node1180;
	wire [3-1:0] node1184;
	wire [3-1:0] node1186;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1191;
	wire [3-1:0] node1193;
	wire [3-1:0] node1196;
	wire [3-1:0] node1197;
	wire [3-1:0] node1201;
	wire [3-1:0] node1202;
	wire [3-1:0] node1203;
	wire [3-1:0] node1207;
	wire [3-1:0] node1208;
	wire [3-1:0] node1209;
	wire [3-1:0] node1214;
	wire [3-1:0] node1215;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1219;
	wire [3-1:0] node1220;
	wire [3-1:0] node1222;
	wire [3-1:0] node1226;
	wire [3-1:0] node1227;
	wire [3-1:0] node1230;
	wire [3-1:0] node1233;
	wire [3-1:0] node1235;
	wire [3-1:0] node1237;
	wire [3-1:0] node1238;
	wire [3-1:0] node1242;
	wire [3-1:0] node1243;
	wire [3-1:0] node1244;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1250;
	wire [3-1:0] node1253;
	wire [3-1:0] node1254;
	wire [3-1:0] node1255;
	wire [3-1:0] node1259;
	wire [3-1:0] node1260;
	wire [3-1:0] node1264;
	wire [3-1:0] node1265;
	wire [3-1:0] node1266;
	wire [3-1:0] node1268;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1277;
	wire [3-1:0] node1278;
	wire [3-1:0] node1279;
	wire [3-1:0] node1280;
	wire [3-1:0] node1282;
	wire [3-1:0] node1285;
	wire [3-1:0] node1286;
	wire [3-1:0] node1287;
	wire [3-1:0] node1291;
	wire [3-1:0] node1294;
	wire [3-1:0] node1295;
	wire [3-1:0] node1297;
	wire [3-1:0] node1298;
	wire [3-1:0] node1302;
	wire [3-1:0] node1303;
	wire [3-1:0] node1304;
	wire [3-1:0] node1307;
	wire [3-1:0] node1311;
	wire [3-1:0] node1312;
	wire [3-1:0] node1313;
	wire [3-1:0] node1314;
	wire [3-1:0] node1318;
	wire [3-1:0] node1321;
	wire [3-1:0] node1322;
	wire [3-1:0] node1323;
	wire [3-1:0] node1324;
	wire [3-1:0] node1328;
	wire [3-1:0] node1329;
	wire [3-1:0] node1333;
	wire [3-1:0] node1335;
	wire [3-1:0] node1338;
	wire [3-1:0] node1339;
	wire [3-1:0] node1340;
	wire [3-1:0] node1341;
	wire [3-1:0] node1342;
	wire [3-1:0] node1344;
	wire [3-1:0] node1345;
	wire [3-1:0] node1348;
	wire [3-1:0] node1351;
	wire [3-1:0] node1353;
	wire [3-1:0] node1354;
	wire [3-1:0] node1358;
	wire [3-1:0] node1359;
	wire [3-1:0] node1360;
	wire [3-1:0] node1361;
	wire [3-1:0] node1364;
	wire [3-1:0] node1368;
	wire [3-1:0] node1369;
	wire [3-1:0] node1370;
	wire [3-1:0] node1374;
	wire [3-1:0] node1377;
	wire [3-1:0] node1378;
	wire [3-1:0] node1379;
	wire [3-1:0] node1381;
	wire [3-1:0] node1383;
	wire [3-1:0] node1386;
	wire [3-1:0] node1387;
	wire [3-1:0] node1388;
	wire [3-1:0] node1392;
	wire [3-1:0] node1393;
	wire [3-1:0] node1397;
	wire [3-1:0] node1398;
	wire [3-1:0] node1400;
	wire [3-1:0] node1401;
	wire [3-1:0] node1405;
	wire [3-1:0] node1408;
	wire [3-1:0] node1409;
	wire [3-1:0] node1410;
	wire [3-1:0] node1412;
	wire [3-1:0] node1413;
	wire [3-1:0] node1417;
	wire [3-1:0] node1418;
	wire [3-1:0] node1419;
	wire [3-1:0] node1422;
	wire [3-1:0] node1425;
	wire [3-1:0] node1427;
	wire [3-1:0] node1430;
	wire [3-1:0] node1431;
	wire [3-1:0] node1432;
	wire [3-1:0] node1434;
	wire [3-1:0] node1437;
	wire [3-1:0] node1438;
	wire [3-1:0] node1442;
	wire [3-1:0] node1443;
	wire [3-1:0] node1444;
	wire [3-1:0] node1449;
	wire [3-1:0] node1450;
	wire [3-1:0] node1451;
	wire [3-1:0] node1452;
	wire [3-1:0] node1453;
	wire [3-1:0] node1454;
	wire [3-1:0] node1455;
	wire [3-1:0] node1458;
	wire [3-1:0] node1459;
	wire [3-1:0] node1461;
	wire [3-1:0] node1464;
	wire [3-1:0] node1465;
	wire [3-1:0] node1469;
	wire [3-1:0] node1470;
	wire [3-1:0] node1472;
	wire [3-1:0] node1475;
	wire [3-1:0] node1476;
	wire [3-1:0] node1477;
	wire [3-1:0] node1482;
	wire [3-1:0] node1483;
	wire [3-1:0] node1484;
	wire [3-1:0] node1485;
	wire [3-1:0] node1488;
	wire [3-1:0] node1489;
	wire [3-1:0] node1492;
	wire [3-1:0] node1495;
	wire [3-1:0] node1496;
	wire [3-1:0] node1498;
	wire [3-1:0] node1501;
	wire [3-1:0] node1502;
	wire [3-1:0] node1506;
	wire [3-1:0] node1507;
	wire [3-1:0] node1509;
	wire [3-1:0] node1512;
	wire [3-1:0] node1513;
	wire [3-1:0] node1516;
	wire [3-1:0] node1517;
	wire [3-1:0] node1521;
	wire [3-1:0] node1522;
	wire [3-1:0] node1523;
	wire [3-1:0] node1524;
	wire [3-1:0] node1525;
	wire [3-1:0] node1528;
	wire [3-1:0] node1531;
	wire [3-1:0] node1532;
	wire [3-1:0] node1535;
	wire [3-1:0] node1536;
	wire [3-1:0] node1540;
	wire [3-1:0] node1541;
	wire [3-1:0] node1542;
	wire [3-1:0] node1545;
	wire [3-1:0] node1548;
	wire [3-1:0] node1550;
	wire [3-1:0] node1553;
	wire [3-1:0] node1554;
	wire [3-1:0] node1555;
	wire [3-1:0] node1556;
	wire [3-1:0] node1559;
	wire [3-1:0] node1563;
	wire [3-1:0] node1564;
	wire [3-1:0] node1565;
	wire [3-1:0] node1566;
	wire [3-1:0] node1569;
	wire [3-1:0] node1572;
	wire [3-1:0] node1573;
	wire [3-1:0] node1576;
	wire [3-1:0] node1579;
	wire [3-1:0] node1580;
	wire [3-1:0] node1581;
	wire [3-1:0] node1586;
	wire [3-1:0] node1587;
	wire [3-1:0] node1588;
	wire [3-1:0] node1589;
	wire [3-1:0] node1591;
	wire [3-1:0] node1592;
	wire [3-1:0] node1593;
	wire [3-1:0] node1596;
	wire [3-1:0] node1599;
	wire [3-1:0] node1601;
	wire [3-1:0] node1604;
	wire [3-1:0] node1605;
	wire [3-1:0] node1606;
	wire [3-1:0] node1607;
	wire [3-1:0] node1612;
	wire [3-1:0] node1614;
	wire [3-1:0] node1617;
	wire [3-1:0] node1618;
	wire [3-1:0] node1619;
	wire [3-1:0] node1621;
	wire [3-1:0] node1624;
	wire [3-1:0] node1626;
	wire [3-1:0] node1629;
	wire [3-1:0] node1630;
	wire [3-1:0] node1631;
	wire [3-1:0] node1634;
	wire [3-1:0] node1637;
	wire [3-1:0] node1638;
	wire [3-1:0] node1639;
	wire [3-1:0] node1643;
	wire [3-1:0] node1644;
	wire [3-1:0] node1648;
	wire [3-1:0] node1649;
	wire [3-1:0] node1650;
	wire [3-1:0] node1651;
	wire [3-1:0] node1652;
	wire [3-1:0] node1655;
	wire [3-1:0] node1658;
	wire [3-1:0] node1659;
	wire [3-1:0] node1662;
	wire [3-1:0] node1665;
	wire [3-1:0] node1666;
	wire [3-1:0] node1667;
	wire [3-1:0] node1668;
	wire [3-1:0] node1671;
	wire [3-1:0] node1674;
	wire [3-1:0] node1675;
	wire [3-1:0] node1679;
	wire [3-1:0] node1681;
	wire [3-1:0] node1682;
	wire [3-1:0] node1685;
	wire [3-1:0] node1688;
	wire [3-1:0] node1689;
	wire [3-1:0] node1690;
	wire [3-1:0] node1692;
	wire [3-1:0] node1695;
	wire [3-1:0] node1696;
	wire [3-1:0] node1697;
	wire [3-1:0] node1701;
	wire [3-1:0] node1703;
	wire [3-1:0] node1706;
	wire [3-1:0] node1707;
	wire [3-1:0] node1709;
	wire [3-1:0] node1710;
	wire [3-1:0] node1714;
	wire [3-1:0] node1715;
	wire [3-1:0] node1716;
	wire [3-1:0] node1719;
	wire [3-1:0] node1723;
	wire [3-1:0] node1724;
	wire [3-1:0] node1725;
	wire [3-1:0] node1726;
	wire [3-1:0] node1727;
	wire [3-1:0] node1728;
	wire [3-1:0] node1729;
	wire [3-1:0] node1731;
	wire [3-1:0] node1734;
	wire [3-1:0] node1736;
	wire [3-1:0] node1739;
	wire [3-1:0] node1741;
	wire [3-1:0] node1744;
	wire [3-1:0] node1745;
	wire [3-1:0] node1747;
	wire [3-1:0] node1748;
	wire [3-1:0] node1752;
	wire [3-1:0] node1753;
	wire [3-1:0] node1754;
	wire [3-1:0] node1757;
	wire [3-1:0] node1761;
	wire [3-1:0] node1762;
	wire [3-1:0] node1763;
	wire [3-1:0] node1764;
	wire [3-1:0] node1766;
	wire [3-1:0] node1769;
	wire [3-1:0] node1771;
	wire [3-1:0] node1774;
	wire [3-1:0] node1775;
	wire [3-1:0] node1778;
	wire [3-1:0] node1781;
	wire [3-1:0] node1782;
	wire [3-1:0] node1784;
	wire [3-1:0] node1785;
	wire [3-1:0] node1789;
	wire [3-1:0] node1792;
	wire [3-1:0] node1793;
	wire [3-1:0] node1794;
	wire [3-1:0] node1795;
	wire [3-1:0] node1796;
	wire [3-1:0] node1797;
	wire [3-1:0] node1800;
	wire [3-1:0] node1803;
	wire [3-1:0] node1805;
	wire [3-1:0] node1808;
	wire [3-1:0] node1810;
	wire [3-1:0] node1813;
	wire [3-1:0] node1814;
	wire [3-1:0] node1815;
	wire [3-1:0] node1818;
	wire [3-1:0] node1821;
	wire [3-1:0] node1822;
	wire [3-1:0] node1825;
	wire [3-1:0] node1828;
	wire [3-1:0] node1829;
	wire [3-1:0] node1830;
	wire [3-1:0] node1832;
	wire [3-1:0] node1835;
	wire [3-1:0] node1836;
	wire [3-1:0] node1839;
	wire [3-1:0] node1842;
	wire [3-1:0] node1843;
	wire [3-1:0] node1844;
	wire [3-1:0] node1848;
	wire [3-1:0] node1851;
	wire [3-1:0] node1852;
	wire [3-1:0] node1853;
	wire [3-1:0] node1854;
	wire [3-1:0] node1855;
	wire [3-1:0] node1856;
	wire [3-1:0] node1859;
	wire [3-1:0] node1862;
	wire [3-1:0] node1863;
	wire [3-1:0] node1866;
	wire [3-1:0] node1869;
	wire [3-1:0] node1870;
	wire [3-1:0] node1873;
	wire [3-1:0] node1876;
	wire [3-1:0] node1877;
	wire [3-1:0] node1878;
	wire [3-1:0] node1879;
	wire [3-1:0] node1882;
	wire [3-1:0] node1885;
	wire [3-1:0] node1887;
	wire [3-1:0] node1890;
	wire [3-1:0] node1891;
	wire [3-1:0] node1892;
	wire [3-1:0] node1895;
	wire [3-1:0] node1898;
	wire [3-1:0] node1899;
	wire [3-1:0] node1900;
	wire [3-1:0] node1903;
	wire [3-1:0] node1907;
	wire [3-1:0] node1908;
	wire [3-1:0] node1909;
	wire [3-1:0] node1910;
	wire [3-1:0] node1912;
	wire [3-1:0] node1913;
	wire [3-1:0] node1916;
	wire [3-1:0] node1919;
	wire [3-1:0] node1920;
	wire [3-1:0] node1923;
	wire [3-1:0] node1926;
	wire [3-1:0] node1927;
	wire [3-1:0] node1928;
	wire [3-1:0] node1930;
	wire [3-1:0] node1933;
	wire [3-1:0] node1934;
	wire [3-1:0] node1937;
	wire [3-1:0] node1940;
	wire [3-1:0] node1941;
	wire [3-1:0] node1942;
	wire [3-1:0] node1945;
	wire [3-1:0] node1949;
	wire [3-1:0] node1950;
	wire [3-1:0] node1951;
	wire [3-1:0] node1952;
	wire [3-1:0] node1955;
	wire [3-1:0] node1958;
	wire [3-1:0] node1960;
	wire [3-1:0] node1963;
	wire [3-1:0] node1964;
	wire [3-1:0] node1967;
	wire [3-1:0] node1970;
	wire [3-1:0] node1971;
	wire [3-1:0] node1972;
	wire [3-1:0] node1973;
	wire [3-1:0] node1974;
	wire [3-1:0] node1975;
	wire [3-1:0] node1976;
	wire [3-1:0] node1977;
	wire [3-1:0] node1978;
	wire [3-1:0] node1980;
	wire [3-1:0] node1983;
	wire [3-1:0] node1984;
	wire [3-1:0] node1985;
	wire [3-1:0] node1989;
	wire [3-1:0] node1990;
	wire [3-1:0] node1993;
	wire [3-1:0] node1996;
	wire [3-1:0] node1998;
	wire [3-1:0] node1999;
	wire [3-1:0] node2000;
	wire [3-1:0] node2003;
	wire [3-1:0] node2006;
	wire [3-1:0] node2007;
	wire [3-1:0] node2010;
	wire [3-1:0] node2013;
	wire [3-1:0] node2014;
	wire [3-1:0] node2015;
	wire [3-1:0] node2018;
	wire [3-1:0] node2020;
	wire [3-1:0] node2023;
	wire [3-1:0] node2024;
	wire [3-1:0] node2026;
	wire [3-1:0] node2029;
	wire [3-1:0] node2032;
	wire [3-1:0] node2033;
	wire [3-1:0] node2034;
	wire [3-1:0] node2035;
	wire [3-1:0] node2037;
	wire [3-1:0] node2040;
	wire [3-1:0] node2042;
	wire [3-1:0] node2045;
	wire [3-1:0] node2046;
	wire [3-1:0] node2048;
	wire [3-1:0] node2051;
	wire [3-1:0] node2053;
	wire [3-1:0] node2056;
	wire [3-1:0] node2057;
	wire [3-1:0] node2058;
	wire [3-1:0] node2060;
	wire [3-1:0] node2063;
	wire [3-1:0] node2065;
	wire [3-1:0] node2066;
	wire [3-1:0] node2070;
	wire [3-1:0] node2072;
	wire [3-1:0] node2075;
	wire [3-1:0] node2076;
	wire [3-1:0] node2077;
	wire [3-1:0] node2078;
	wire [3-1:0] node2079;
	wire [3-1:0] node2080;
	wire [3-1:0] node2083;
	wire [3-1:0] node2085;
	wire [3-1:0] node2088;
	wire [3-1:0] node2089;
	wire [3-1:0] node2091;
	wire [3-1:0] node2095;
	wire [3-1:0] node2096;
	wire [3-1:0] node2098;
	wire [3-1:0] node2101;
	wire [3-1:0] node2103;
	wire [3-1:0] node2104;
	wire [3-1:0] node2108;
	wire [3-1:0] node2109;
	wire [3-1:0] node2110;
	wire [3-1:0] node2112;
	wire [3-1:0] node2115;
	wire [3-1:0] node2116;
	wire [3-1:0] node2120;
	wire [3-1:0] node2121;
	wire [3-1:0] node2123;
	wire [3-1:0] node2127;
	wire [3-1:0] node2128;
	wire [3-1:0] node2129;
	wire [3-1:0] node2130;
	wire [3-1:0] node2131;
	wire [3-1:0] node2134;
	wire [3-1:0] node2137;
	wire [3-1:0] node2139;
	wire [3-1:0] node2140;
	wire [3-1:0] node2143;
	wire [3-1:0] node2146;
	wire [3-1:0] node2147;
	wire [3-1:0] node2148;
	wire [3-1:0] node2149;
	wire [3-1:0] node2154;
	wire [3-1:0] node2155;
	wire [3-1:0] node2156;
	wire [3-1:0] node2159;
	wire [3-1:0] node2163;
	wire [3-1:0] node2164;
	wire [3-1:0] node2165;
	wire [3-1:0] node2166;
	wire [3-1:0] node2168;
	wire [3-1:0] node2171;
	wire [3-1:0] node2173;
	wire [3-1:0] node2176;
	wire [3-1:0] node2177;
	wire [3-1:0] node2179;
	wire [3-1:0] node2183;
	wire [3-1:0] node2184;
	wire [3-1:0] node2185;
	wire [3-1:0] node2186;
	wire [3-1:0] node2189;
	wire [3-1:0] node2193;
	wire [3-1:0] node2194;
	wire [3-1:0] node2195;
	wire [3-1:0] node2198;
	wire [3-1:0] node2202;
	wire [3-1:0] node2203;
	wire [3-1:0] node2204;
	wire [3-1:0] node2205;
	wire [3-1:0] node2206;
	wire [3-1:0] node2207;
	wire [3-1:0] node2208;
	wire [3-1:0] node2210;
	wire [3-1:0] node2213;
	wire [3-1:0] node2214;
	wire [3-1:0] node2217;
	wire [3-1:0] node2220;
	wire [3-1:0] node2222;
	wire [3-1:0] node2225;
	wire [3-1:0] node2226;
	wire [3-1:0] node2227;
	wire [3-1:0] node2231;
	wire [3-1:0] node2233;
	wire [3-1:0] node2235;
	wire [3-1:0] node2238;
	wire [3-1:0] node2239;
	wire [3-1:0] node2240;
	wire [3-1:0] node2241;
	wire [3-1:0] node2244;
	wire [3-1:0] node2246;
	wire [3-1:0] node2249;
	wire [3-1:0] node2250;
	wire [3-1:0] node2253;
	wire [3-1:0] node2256;
	wire [3-1:0] node2257;
	wire [3-1:0] node2258;
	wire [3-1:0] node2261;
	wire [3-1:0] node2263;
	wire [3-1:0] node2266;
	wire [3-1:0] node2267;
	wire [3-1:0] node2271;
	wire [3-1:0] node2272;
	wire [3-1:0] node2273;
	wire [3-1:0] node2274;
	wire [3-1:0] node2276;
	wire [3-1:0] node2279;
	wire [3-1:0] node2280;
	wire [3-1:0] node2281;
	wire [3-1:0] node2286;
	wire [3-1:0] node2287;
	wire [3-1:0] node2288;
	wire [3-1:0] node2292;
	wire [3-1:0] node2294;
	wire [3-1:0] node2297;
	wire [3-1:0] node2298;
	wire [3-1:0] node2299;
	wire [3-1:0] node2300;
	wire [3-1:0] node2301;
	wire [3-1:0] node2305;
	wire [3-1:0] node2308;
	wire [3-1:0] node2310;
	wire [3-1:0] node2313;
	wire [3-1:0] node2314;
	wire [3-1:0] node2315;
	wire [3-1:0] node2319;
	wire [3-1:0] node2322;
	wire [3-1:0] node2323;
	wire [3-1:0] node2324;
	wire [3-1:0] node2325;
	wire [3-1:0] node2326;
	wire [3-1:0] node2328;
	wire [3-1:0] node2331;
	wire [3-1:0] node2332;
	wire [3-1:0] node2333;
	wire [3-1:0] node2336;
	wire [3-1:0] node2340;
	wire [3-1:0] node2341;
	wire [3-1:0] node2342;
	wire [3-1:0] node2347;
	wire [3-1:0] node2348;
	wire [3-1:0] node2349;
	wire [3-1:0] node2350;
	wire [3-1:0] node2354;
	wire [3-1:0] node2355;
	wire [3-1:0] node2359;
	wire [3-1:0] node2360;
	wire [3-1:0] node2361;
	wire [3-1:0] node2365;
	wire [3-1:0] node2366;
	wire [3-1:0] node2370;
	wire [3-1:0] node2371;
	wire [3-1:0] node2372;
	wire [3-1:0] node2373;
	wire [3-1:0] node2375;
	wire [3-1:0] node2378;
	wire [3-1:0] node2379;
	wire [3-1:0] node2380;
	wire [3-1:0] node2384;
	wire [3-1:0] node2385;
	wire [3-1:0] node2388;
	wire [3-1:0] node2391;
	wire [3-1:0] node2392;
	wire [3-1:0] node2394;
	wire [3-1:0] node2397;
	wire [3-1:0] node2399;
	wire [3-1:0] node2402;
	wire [3-1:0] node2403;
	wire [3-1:0] node2405;
	wire [3-1:0] node2406;
	wire [3-1:0] node2407;
	wire [3-1:0] node2410;
	wire [3-1:0] node2414;
	wire [3-1:0] node2415;
	wire [3-1:0] node2416;
	wire [3-1:0] node2417;
	wire [3-1:0] node2420;
	wire [3-1:0] node2424;
	wire [3-1:0] node2425;
	wire [3-1:0] node2426;
	wire [3-1:0] node2430;
	wire [3-1:0] node2432;
	wire [3-1:0] node2435;
	wire [3-1:0] node2436;
	wire [3-1:0] node2437;
	wire [3-1:0] node2438;
	wire [3-1:0] node2439;
	wire [3-1:0] node2440;
	wire [3-1:0] node2441;
	wire [3-1:0] node2442;
	wire [3-1:0] node2445;
	wire [3-1:0] node2448;
	wire [3-1:0] node2449;
	wire [3-1:0] node2452;
	wire [3-1:0] node2455;
	wire [3-1:0] node2456;
	wire [3-1:0] node2457;
	wire [3-1:0] node2460;
	wire [3-1:0] node2463;
	wire [3-1:0] node2465;
	wire [3-1:0] node2468;
	wire [3-1:0] node2469;
	wire [3-1:0] node2470;
	wire [3-1:0] node2473;
	wire [3-1:0] node2475;
	wire [3-1:0] node2478;
	wire [3-1:0] node2479;
	wire [3-1:0] node2481;
	wire [3-1:0] node2484;
	wire [3-1:0] node2486;
	wire [3-1:0] node2489;
	wire [3-1:0] node2490;
	wire [3-1:0] node2491;
	wire [3-1:0] node2492;
	wire [3-1:0] node2493;
	wire [3-1:0] node2496;
	wire [3-1:0] node2499;
	wire [3-1:0] node2500;
	wire [3-1:0] node2504;
	wire [3-1:0] node2505;
	wire [3-1:0] node2506;
	wire [3-1:0] node2507;
	wire [3-1:0] node2511;
	wire [3-1:0] node2512;
	wire [3-1:0] node2516;
	wire [3-1:0] node2517;
	wire [3-1:0] node2519;
	wire [3-1:0] node2523;
	wire [3-1:0] node2524;
	wire [3-1:0] node2525;
	wire [3-1:0] node2526;
	wire [3-1:0] node2528;
	wire [3-1:0] node2531;
	wire [3-1:0] node2532;
	wire [3-1:0] node2536;
	wire [3-1:0] node2538;
	wire [3-1:0] node2540;
	wire [3-1:0] node2543;
	wire [3-1:0] node2544;
	wire [3-1:0] node2545;
	wire [3-1:0] node2546;
	wire [3-1:0] node2551;
	wire [3-1:0] node2552;
	wire [3-1:0] node2555;
	wire [3-1:0] node2558;
	wire [3-1:0] node2559;
	wire [3-1:0] node2560;
	wire [3-1:0] node2561;
	wire [3-1:0] node2562;
	wire [3-1:0] node2563;
	wire [3-1:0] node2566;
	wire [3-1:0] node2569;
	wire [3-1:0] node2570;
	wire [3-1:0] node2573;
	wire [3-1:0] node2576;
	wire [3-1:0] node2577;
	wire [3-1:0] node2578;
	wire [3-1:0] node2581;
	wire [3-1:0] node2584;
	wire [3-1:0] node2585;
	wire [3-1:0] node2586;
	wire [3-1:0] node2590;
	wire [3-1:0] node2593;
	wire [3-1:0] node2594;
	wire [3-1:0] node2595;
	wire [3-1:0] node2596;
	wire [3-1:0] node2597;
	wire [3-1:0] node2600;
	wire [3-1:0] node2604;
	wire [3-1:0] node2605;
	wire [3-1:0] node2609;
	wire [3-1:0] node2610;
	wire [3-1:0] node2611;
	wire [3-1:0] node2615;
	wire [3-1:0] node2618;
	wire [3-1:0] node2619;
	wire [3-1:0] node2620;
	wire [3-1:0] node2621;
	wire [3-1:0] node2623;
	wire [3-1:0] node2626;
	wire [3-1:0] node2627;
	wire [3-1:0] node2631;
	wire [3-1:0] node2632;
	wire [3-1:0] node2633;
	wire [3-1:0] node2637;
	wire [3-1:0] node2640;
	wire [3-1:0] node2641;
	wire [3-1:0] node2643;
	wire [3-1:0] node2644;
	wire [3-1:0] node2648;
	wire [3-1:0] node2649;
	wire [3-1:0] node2650;
	wire [3-1:0] node2655;
	wire [3-1:0] node2656;
	wire [3-1:0] node2657;
	wire [3-1:0] node2658;
	wire [3-1:0] node2659;
	wire [3-1:0] node2660;
	wire [3-1:0] node2661;
	wire [3-1:0] node2664;
	wire [3-1:0] node2667;
	wire [3-1:0] node2668;
	wire [3-1:0] node2671;
	wire [3-1:0] node2674;
	wire [3-1:0] node2675;
	wire [3-1:0] node2678;
	wire [3-1:0] node2681;
	wire [3-1:0] node2682;
	wire [3-1:0] node2683;
	wire [3-1:0] node2685;
	wire [3-1:0] node2686;
	wire [3-1:0] node2689;
	wire [3-1:0] node2692;
	wire [3-1:0] node2693;
	wire [3-1:0] node2694;
	wire [3-1:0] node2697;
	wire [3-1:0] node2701;
	wire [3-1:0] node2702;
	wire [3-1:0] node2703;
	wire [3-1:0] node2706;
	wire [3-1:0] node2708;
	wire [3-1:0] node2712;
	wire [3-1:0] node2713;
	wire [3-1:0] node2714;
	wire [3-1:0] node2715;
	wire [3-1:0] node2716;
	wire [3-1:0] node2720;
	wire [3-1:0] node2722;
	wire [3-1:0] node2725;
	wire [3-1:0] node2726;
	wire [3-1:0] node2727;
	wire [3-1:0] node2730;
	wire [3-1:0] node2733;
	wire [3-1:0] node2734;
	wire [3-1:0] node2737;
	wire [3-1:0] node2740;
	wire [3-1:0] node2741;
	wire [3-1:0] node2742;
	wire [3-1:0] node2743;
	wire [3-1:0] node2746;
	wire [3-1:0] node2749;
	wire [3-1:0] node2750;
	wire [3-1:0] node2753;
	wire [3-1:0] node2756;
	wire [3-1:0] node2757;
	wire [3-1:0] node2758;
	wire [3-1:0] node2762;
	wire [3-1:0] node2765;
	wire [3-1:0] node2766;
	wire [3-1:0] node2767;
	wire [3-1:0] node2768;
	wire [3-1:0] node2769;
	wire [3-1:0] node2770;
	wire [3-1:0] node2773;
	wire [3-1:0] node2775;
	wire [3-1:0] node2778;
	wire [3-1:0] node2779;
	wire [3-1:0] node2782;
	wire [3-1:0] node2785;
	wire [3-1:0] node2786;
	wire [3-1:0] node2787;
	wire [3-1:0] node2791;
	wire [3-1:0] node2794;
	wire [3-1:0] node2795;
	wire [3-1:0] node2796;
	wire [3-1:0] node2798;
	wire [3-1:0] node2801;
	wire [3-1:0] node2802;
	wire [3-1:0] node2805;
	wire [3-1:0] node2808;
	wire [3-1:0] node2810;
	wire [3-1:0] node2811;
	wire [3-1:0] node2814;
	wire [3-1:0] node2817;
	wire [3-1:0] node2818;
	wire [3-1:0] node2819;
	wire [3-1:0] node2820;
	wire [3-1:0] node2821;
	wire [3-1:0] node2823;
	wire [3-1:0] node2827;
	wire [3-1:0] node2830;
	wire [3-1:0] node2831;
	wire [3-1:0] node2832;
	wire [3-1:0] node2833;
	wire [3-1:0] node2836;
	wire [3-1:0] node2839;
	wire [3-1:0] node2842;
	wire [3-1:0] node2843;
	wire [3-1:0] node2846;
	wire [3-1:0] node2848;
	wire [3-1:0] node2851;
	wire [3-1:0] node2852;
	wire [3-1:0] node2853;
	wire [3-1:0] node2854;
	wire [3-1:0] node2857;
	wire [3-1:0] node2858;
	wire [3-1:0] node2862;
	wire [3-1:0] node2864;
	wire [3-1:0] node2866;
	wire [3-1:0] node2869;
	wire [3-1:0] node2870;
	wire [3-1:0] node2872;
	wire [3-1:0] node2875;
	wire [3-1:0] node2876;
	wire [3-1:0] node2880;
	wire [3-1:0] node2881;
	wire [3-1:0] node2882;
	wire [3-1:0] node2883;
	wire [3-1:0] node2884;
	wire [3-1:0] node2885;
	wire [3-1:0] node2886;
	wire [3-1:0] node2887;
	wire [3-1:0] node2888;
	wire [3-1:0] node2891;
	wire [3-1:0] node2894;
	wire [3-1:0] node2896;
	wire [3-1:0] node2897;
	wire [3-1:0] node2900;
	wire [3-1:0] node2903;
	wire [3-1:0] node2904;
	wire [3-1:0] node2905;
	wire [3-1:0] node2908;
	wire [3-1:0] node2911;
	wire [3-1:0] node2912;
	wire [3-1:0] node2915;
	wire [3-1:0] node2918;
	wire [3-1:0] node2919;
	wire [3-1:0] node2920;
	wire [3-1:0] node2922;
	wire [3-1:0] node2923;
	wire [3-1:0] node2926;
	wire [3-1:0] node2929;
	wire [3-1:0] node2930;
	wire [3-1:0] node2931;
	wire [3-1:0] node2934;
	wire [3-1:0] node2938;
	wire [3-1:0] node2939;
	wire [3-1:0] node2940;
	wire [3-1:0] node2941;
	wire [3-1:0] node2945;
	wire [3-1:0] node2946;
	wire [3-1:0] node2950;
	wire [3-1:0] node2951;
	wire [3-1:0] node2953;
	wire [3-1:0] node2957;
	wire [3-1:0] node2958;
	wire [3-1:0] node2959;
	wire [3-1:0] node2960;
	wire [3-1:0] node2961;
	wire [3-1:0] node2964;
	wire [3-1:0] node2967;
	wire [3-1:0] node2968;
	wire [3-1:0] node2969;
	wire [3-1:0] node2972;
	wire [3-1:0] node2976;
	wire [3-1:0] node2977;
	wire [3-1:0] node2979;
	wire [3-1:0] node2983;
	wire [3-1:0] node2984;
	wire [3-1:0] node2985;
	wire [3-1:0] node2986;
	wire [3-1:0] node2987;
	wire [3-1:0] node2990;
	wire [3-1:0] node2993;
	wire [3-1:0] node2995;
	wire [3-1:0] node2998;
	wire [3-1:0] node2999;
	wire [3-1:0] node3000;
	wire [3-1:0] node3003;
	wire [3-1:0] node3006;
	wire [3-1:0] node3008;
	wire [3-1:0] node3011;
	wire [3-1:0] node3012;
	wire [3-1:0] node3013;
	wire [3-1:0] node3016;
	wire [3-1:0] node3019;
	wire [3-1:0] node3020;
	wire [3-1:0] node3021;
	wire [3-1:0] node3024;
	wire [3-1:0] node3027;
	wire [3-1:0] node3029;
	wire [3-1:0] node3032;
	wire [3-1:0] node3033;
	wire [3-1:0] node3034;
	wire [3-1:0] node3035;
	wire [3-1:0] node3036;
	wire [3-1:0] node3037;
	wire [3-1:0] node3038;
	wire [3-1:0] node3043;
	wire [3-1:0] node3044;
	wire [3-1:0] node3047;
	wire [3-1:0] node3048;
	wire [3-1:0] node3051;
	wire [3-1:0] node3054;
	wire [3-1:0] node3055;
	wire [3-1:0] node3058;
	wire [3-1:0] node3059;
	wire [3-1:0] node3061;
	wire [3-1:0] node3065;
	wire [3-1:0] node3066;
	wire [3-1:0] node3067;
	wire [3-1:0] node3068;
	wire [3-1:0] node3070;
	wire [3-1:0] node3073;
	wire [3-1:0] node3074;
	wire [3-1:0] node3077;
	wire [3-1:0] node3080;
	wire [3-1:0] node3081;
	wire [3-1:0] node3082;
	wire [3-1:0] node3085;
	wire [3-1:0] node3088;
	wire [3-1:0] node3091;
	wire [3-1:0] node3092;
	wire [3-1:0] node3094;
	wire [3-1:0] node3095;
	wire [3-1:0] node3098;
	wire [3-1:0] node3101;
	wire [3-1:0] node3103;
	wire [3-1:0] node3106;
	wire [3-1:0] node3107;
	wire [3-1:0] node3108;
	wire [3-1:0] node3109;
	wire [3-1:0] node3110;
	wire [3-1:0] node3113;
	wire [3-1:0] node3116;
	wire [3-1:0] node3117;
	wire [3-1:0] node3120;
	wire [3-1:0] node3123;
	wire [3-1:0] node3124;
	wire [3-1:0] node3127;
	wire [3-1:0] node3129;
	wire [3-1:0] node3132;
	wire [3-1:0] node3133;
	wire [3-1:0] node3134;
	wire [3-1:0] node3136;
	wire [3-1:0] node3137;
	wire [3-1:0] node3141;
	wire [3-1:0] node3142;
	wire [3-1:0] node3145;
	wire [3-1:0] node3148;
	wire [3-1:0] node3149;
	wire [3-1:0] node3150;
	wire [3-1:0] node3152;
	wire [3-1:0] node3155;
	wire [3-1:0] node3158;
	wire [3-1:0] node3159;
	wire [3-1:0] node3162;
	wire [3-1:0] node3165;
	wire [3-1:0] node3166;
	wire [3-1:0] node3167;
	wire [3-1:0] node3168;
	wire [3-1:0] node3169;
	wire [3-1:0] node3170;
	wire [3-1:0] node3171;
	wire [3-1:0] node3172;
	wire [3-1:0] node3176;
	wire [3-1:0] node3177;
	wire [3-1:0] node3181;
	wire [3-1:0] node3182;
	wire [3-1:0] node3186;
	wire [3-1:0] node3187;
	wire [3-1:0] node3188;
	wire [3-1:0] node3191;
	wire [3-1:0] node3194;
	wire [3-1:0] node3195;
	wire [3-1:0] node3199;
	wire [3-1:0] node3200;
	wire [3-1:0] node3201;
	wire [3-1:0] node3202;
	wire [3-1:0] node3206;
	wire [3-1:0] node3207;
	wire [3-1:0] node3208;
	wire [3-1:0] node3211;
	wire [3-1:0] node3215;
	wire [3-1:0] node3216;
	wire [3-1:0] node3217;
	wire [3-1:0] node3220;
	wire [3-1:0] node3223;
	wire [3-1:0] node3224;
	wire [3-1:0] node3228;
	wire [3-1:0] node3229;
	wire [3-1:0] node3230;
	wire [3-1:0] node3231;
	wire [3-1:0] node3232;
	wire [3-1:0] node3235;
	wire [3-1:0] node3238;
	wire [3-1:0] node3240;
	wire [3-1:0] node3241;
	wire [3-1:0] node3244;
	wire [3-1:0] node3247;
	wire [3-1:0] node3248;
	wire [3-1:0] node3249;
	wire [3-1:0] node3251;
	wire [3-1:0] node3254;
	wire [3-1:0] node3255;
	wire [3-1:0] node3258;
	wire [3-1:0] node3261;
	wire [3-1:0] node3262;
	wire [3-1:0] node3266;
	wire [3-1:0] node3267;
	wire [3-1:0] node3268;
	wire [3-1:0] node3269;
	wire [3-1:0] node3270;
	wire [3-1:0] node3274;
	wire [3-1:0] node3275;
	wire [3-1:0] node3278;
	wire [3-1:0] node3281;
	wire [3-1:0] node3282;
	wire [3-1:0] node3284;
	wire [3-1:0] node3287;
	wire [3-1:0] node3289;
	wire [3-1:0] node3292;
	wire [3-1:0] node3294;
	wire [3-1:0] node3295;
	wire [3-1:0] node3296;
	wire [3-1:0] node3299;
	wire [3-1:0] node3302;
	wire [3-1:0] node3303;
	wire [3-1:0] node3306;
	wire [3-1:0] node3309;
	wire [3-1:0] node3310;
	wire [3-1:0] node3311;
	wire [3-1:0] node3312;
	wire [3-1:0] node3313;
	wire [3-1:0] node3315;
	wire [3-1:0] node3316;
	wire [3-1:0] node3320;
	wire [3-1:0] node3321;
	wire [3-1:0] node3323;
	wire [3-1:0] node3326;
	wire [3-1:0] node3327;
	wire [3-1:0] node3331;
	wire [3-1:0] node3332;
	wire [3-1:0] node3333;
	wire [3-1:0] node3334;
	wire [3-1:0] node3339;
	wire [3-1:0] node3340;
	wire [3-1:0] node3341;
	wire [3-1:0] node3344;
	wire [3-1:0] node3347;
	wire [3-1:0] node3348;
	wire [3-1:0] node3351;
	wire [3-1:0] node3354;
	wire [3-1:0] node3355;
	wire [3-1:0] node3356;
	wire [3-1:0] node3357;
	wire [3-1:0] node3361;
	wire [3-1:0] node3364;
	wire [3-1:0] node3365;
	wire [3-1:0] node3366;
	wire [3-1:0] node3367;
	wire [3-1:0] node3370;
	wire [3-1:0] node3373;
	wire [3-1:0] node3375;
	wire [3-1:0] node3378;
	wire [3-1:0] node3381;
	wire [3-1:0] node3382;
	wire [3-1:0] node3383;
	wire [3-1:0] node3385;
	wire [3-1:0] node3387;
	wire [3-1:0] node3388;
	wire [3-1:0] node3391;
	wire [3-1:0] node3394;
	wire [3-1:0] node3395;
	wire [3-1:0] node3396;
	wire [3-1:0] node3399;
	wire [3-1:0] node3401;
	wire [3-1:0] node3404;
	wire [3-1:0] node3406;
	wire [3-1:0] node3409;
	wire [3-1:0] node3410;
	wire [3-1:0] node3411;
	wire [3-1:0] node3414;
	wire [3-1:0] node3417;
	wire [3-1:0] node3418;
	wire [3-1:0] node3419;
	wire [3-1:0] node3422;
	wire [3-1:0] node3425;
	wire [3-1:0] node3426;
	wire [3-1:0] node3430;
	wire [3-1:0] node3431;
	wire [3-1:0] node3432;
	wire [3-1:0] node3433;
	wire [3-1:0] node3434;
	wire [3-1:0] node3435;
	wire [3-1:0] node3436;
	wire [3-1:0] node3437;
	wire [3-1:0] node3440;
	wire [3-1:0] node3443;
	wire [3-1:0] node3445;
	wire [3-1:0] node3448;
	wire [3-1:0] node3449;
	wire [3-1:0] node3450;
	wire [3-1:0] node3453;
	wire [3-1:0] node3457;
	wire [3-1:0] node3458;
	wire [3-1:0] node3459;
	wire [3-1:0] node3460;
	wire [3-1:0] node3463;
	wire [3-1:0] node3466;
	wire [3-1:0] node3468;
	wire [3-1:0] node3471;
	wire [3-1:0] node3472;
	wire [3-1:0] node3475;
	wire [3-1:0] node3478;
	wire [3-1:0] node3479;
	wire [3-1:0] node3480;
	wire [3-1:0] node3481;
	wire [3-1:0] node3482;
	wire [3-1:0] node3483;
	wire [3-1:0] node3487;
	wire [3-1:0] node3488;
	wire [3-1:0] node3491;
	wire [3-1:0] node3494;
	wire [3-1:0] node3495;
	wire [3-1:0] node3499;
	wire [3-1:0] node3500;
	wire [3-1:0] node3503;
	wire [3-1:0] node3506;
	wire [3-1:0] node3507;
	wire [3-1:0] node3508;
	wire [3-1:0] node3509;
	wire [3-1:0] node3513;
	wire [3-1:0] node3515;
	wire [3-1:0] node3516;
	wire [3-1:0] node3519;
	wire [3-1:0] node3522;
	wire [3-1:0] node3523;
	wire [3-1:0] node3524;
	wire [3-1:0] node3527;
	wire [3-1:0] node3530;
	wire [3-1:0] node3531;
	wire [3-1:0] node3532;
	wire [3-1:0] node3535;
	wire [3-1:0] node3538;
	wire [3-1:0] node3539;
	wire [3-1:0] node3542;
	wire [3-1:0] node3545;
	wire [3-1:0] node3546;
	wire [3-1:0] node3547;
	wire [3-1:0] node3548;
	wire [3-1:0] node3549;
	wire [3-1:0] node3550;
	wire [3-1:0] node3554;
	wire [3-1:0] node3555;
	wire [3-1:0] node3558;
	wire [3-1:0] node3561;
	wire [3-1:0] node3562;
	wire [3-1:0] node3564;
	wire [3-1:0] node3566;
	wire [3-1:0] node3569;
	wire [3-1:0] node3570;
	wire [3-1:0] node3571;
	wire [3-1:0] node3574;
	wire [3-1:0] node3577;
	wire [3-1:0] node3578;
	wire [3-1:0] node3581;
	wire [3-1:0] node3584;
	wire [3-1:0] node3585;
	wire [3-1:0] node3586;
	wire [3-1:0] node3587;
	wire [3-1:0] node3590;
	wire [3-1:0] node3593;
	wire [3-1:0] node3594;
	wire [3-1:0] node3597;
	wire [3-1:0] node3600;
	wire [3-1:0] node3601;
	wire [3-1:0] node3602;
	wire [3-1:0] node3606;
	wire [3-1:0] node3608;
	wire [3-1:0] node3611;
	wire [3-1:0] node3612;
	wire [3-1:0] node3613;
	wire [3-1:0] node3614;
	wire [3-1:0] node3617;
	wire [3-1:0] node3620;
	wire [3-1:0] node3621;
	wire [3-1:0] node3624;
	wire [3-1:0] node3627;
	wire [3-1:0] node3628;
	wire [3-1:0] node3629;
	wire [3-1:0] node3632;
	wire [3-1:0] node3635;
	wire [3-1:0] node3636;
	wire [3-1:0] node3639;
	wire [3-1:0] node3642;
	wire [3-1:0] node3643;
	wire [3-1:0] node3644;
	wire [3-1:0] node3645;
	wire [3-1:0] node3646;
	wire [3-1:0] node3647;
	wire [3-1:0] node3649;
	wire [3-1:0] node3652;
	wire [3-1:0] node3653;
	wire [3-1:0] node3656;
	wire [3-1:0] node3659;
	wire [3-1:0] node3660;
	wire [3-1:0] node3661;
	wire [3-1:0] node3662;
	wire [3-1:0] node3665;
	wire [3-1:0] node3669;
	wire [3-1:0] node3670;
	wire [3-1:0] node3674;
	wire [3-1:0] node3675;
	wire [3-1:0] node3676;
	wire [3-1:0] node3677;
	wire [3-1:0] node3679;
	wire [3-1:0] node3683;
	wire [3-1:0] node3684;
	wire [3-1:0] node3687;
	wire [3-1:0] node3690;
	wire [3-1:0] node3691;
	wire [3-1:0] node3692;
	wire [3-1:0] node3695;
	wire [3-1:0] node3698;
	wire [3-1:0] node3699;
	wire [3-1:0] node3702;
	wire [3-1:0] node3705;
	wire [3-1:0] node3706;
	wire [3-1:0] node3707;
	wire [3-1:0] node3708;
	wire [3-1:0] node3709;
	wire [3-1:0] node3713;
	wire [3-1:0] node3714;
	wire [3-1:0] node3717;
	wire [3-1:0] node3720;
	wire [3-1:0] node3721;
	wire [3-1:0] node3723;
	wire [3-1:0] node3726;
	wire [3-1:0] node3729;
	wire [3-1:0] node3730;
	wire [3-1:0] node3731;
	wire [3-1:0] node3732;
	wire [3-1:0] node3735;
	wire [3-1:0] node3738;
	wire [3-1:0] node3739;
	wire [3-1:0] node3742;
	wire [3-1:0] node3745;
	wire [3-1:0] node3747;
	wire [3-1:0] node3748;
	wire [3-1:0] node3750;
	wire [3-1:0] node3753;
	wire [3-1:0] node3754;
	wire [3-1:0] node3757;
	wire [3-1:0] node3760;
	wire [3-1:0] node3761;
	wire [3-1:0] node3762;
	wire [3-1:0] node3763;
	wire [3-1:0] node3765;
	wire [3-1:0] node3767;
	wire [3-1:0] node3770;
	wire [3-1:0] node3771;
	wire [3-1:0] node3772;
	wire [3-1:0] node3776;
	wire [3-1:0] node3777;
	wire [3-1:0] node3778;
	wire [3-1:0] node3783;
	wire [3-1:0] node3784;
	wire [3-1:0] node3785;
	wire [3-1:0] node3786;
	wire [3-1:0] node3789;
	wire [3-1:0] node3792;
	wire [3-1:0] node3794;
	wire [3-1:0] node3797;
	wire [3-1:0] node3798;
	wire [3-1:0] node3799;
	wire [3-1:0] node3800;
	wire [3-1:0] node3803;
	wire [3-1:0] node3806;
	wire [3-1:0] node3808;
	wire [3-1:0] node3811;
	wire [3-1:0] node3813;
	wire [3-1:0] node3814;
	wire [3-1:0] node3817;
	wire [3-1:0] node3820;
	wire [3-1:0] node3821;
	wire [3-1:0] node3822;
	wire [3-1:0] node3823;
	wire [3-1:0] node3826;
	wire [3-1:0] node3829;
	wire [3-1:0] node3830;
	wire [3-1:0] node3833;
	wire [3-1:0] node3836;
	wire [3-1:0] node3837;
	wire [3-1:0] node3840;

	assign outp = (inp[10]) ? node1970 : node1;
		assign node1 = (inp[6]) ? node967 : node2;
			assign node2 = (inp[1]) ? node528 : node3;
				assign node3 = (inp[11]) ? node261 : node4;
					assign node4 = (inp[5]) ? node118 : node5;
						assign node5 = (inp[8]) ? node59 : node6;
							assign node6 = (inp[4]) ? node34 : node7;
								assign node7 = (inp[2]) ? node15 : node8;
									assign node8 = (inp[7]) ? node12 : node9;
										assign node9 = (inp[9]) ? 3'b110 : 3'b111;
										assign node12 = (inp[9]) ? 3'b111 : 3'b110;
									assign node15 = (inp[3]) ? node29 : node16;
										assign node16 = (inp[0]) ? node24 : node17;
											assign node17 = (inp[9]) ? node21 : node18;
												assign node18 = (inp[7]) ? 3'b110 : 3'b111;
												assign node21 = (inp[7]) ? 3'b111 : 3'b110;
											assign node24 = (inp[9]) ? 3'b111 : node25;
												assign node25 = (inp[7]) ? 3'b111 : 3'b110;
										assign node29 = (inp[7]) ? node31 : 3'b110;
											assign node31 = (inp[0]) ? 3'b110 : 3'b111;
								assign node34 = (inp[9]) ? node46 : node35;
									assign node35 = (inp[7]) ? node41 : node36;
										assign node36 = (inp[0]) ? node38 : 3'b101;
											assign node38 = (inp[2]) ? 3'b100 : 3'b101;
										assign node41 = (inp[2]) ? node43 : 3'b100;
											assign node43 = (inp[0]) ? 3'b101 : 3'b100;
									assign node46 = (inp[2]) ? node48 : 3'b101;
										assign node48 = (inp[3]) ? node54 : node49;
											assign node49 = (inp[7]) ? node51 : 3'b101;
												assign node51 = (inp[0]) ? 3'b100 : 3'b101;
											assign node54 = (inp[7]) ? 3'b101 : node55;
												assign node55 = (inp[0]) ? 3'b101 : 3'b100;
							assign node59 = (inp[4]) ? node91 : node60;
								assign node60 = (inp[3]) ? node74 : node61;
									assign node61 = (inp[7]) ? node69 : node62;
										assign node62 = (inp[9]) ? node64 : 3'b101;
											assign node64 = (inp[0]) ? node66 : 3'b100;
												assign node66 = (inp[2]) ? 3'b101 : 3'b100;
										assign node69 = (inp[9]) ? node71 : 3'b100;
											assign node71 = (inp[2]) ? 3'b100 : 3'b101;
									assign node74 = (inp[7]) ? node86 : node75;
										assign node75 = (inp[9]) ? node81 : node76;
											assign node76 = (inp[2]) ? node78 : 3'b101;
												assign node78 = (inp[0]) ? 3'b100 : 3'b101;
											assign node81 = (inp[2]) ? node83 : 3'b100;
												assign node83 = (inp[0]) ? 3'b101 : 3'b100;
										assign node86 = (inp[9]) ? 3'b101 : node87;
											assign node87 = (inp[2]) ? 3'b101 : 3'b100;
								assign node91 = (inp[2]) ? node111 : node92;
									assign node92 = (inp[3]) ? node100 : node93;
										assign node93 = (inp[9]) ? node95 : 3'b110;
											assign node95 = (inp[0]) ? 3'b110 : node96;
												assign node96 = (inp[7]) ? 3'b111 : 3'b110;
										assign node100 = (inp[7]) ? node106 : node101;
											assign node101 = (inp[0]) ? 3'b111 : node102;
												assign node102 = (inp[9]) ? 3'b110 : 3'b111;
											assign node106 = (inp[0]) ? 3'b110 : node107;
												assign node107 = (inp[9]) ? 3'b111 : 3'b110;
									assign node111 = (inp[9]) ? node115 : node112;
										assign node112 = (inp[7]) ? 3'b111 : 3'b110;
										assign node115 = (inp[7]) ? 3'b110 : 3'b111;
						assign node118 = (inp[9]) ? node186 : node119;
							assign node119 = (inp[3]) ? node151 : node120;
								assign node120 = (inp[7]) ? node138 : node121;
									assign node121 = (inp[0]) ? node135 : node122;
										assign node122 = (inp[2]) ? node130 : node123;
											assign node123 = (inp[4]) ? node127 : node124;
												assign node124 = (inp[8]) ? 3'b101 : 3'b111;
												assign node127 = (inp[8]) ? 3'b111 : 3'b101;
											assign node130 = (inp[4]) ? node132 : 3'b101;
												assign node132 = (inp[8]) ? 3'b110 : 3'b101;
										assign node135 = (inp[2]) ? 3'b100 : 3'b110;
									assign node138 = (inp[2]) ? node140 : 3'b100;
										assign node140 = (inp[0]) ? node148 : node141;
											assign node141 = (inp[8]) ? node145 : node142;
												assign node142 = (inp[4]) ? 3'b100 : 3'b110;
												assign node145 = (inp[4]) ? 3'b111 : 3'b100;
											assign node148 = (inp[4]) ? 3'b101 : 3'b111;
								assign node151 = (inp[2]) ? node171 : node152;
									assign node152 = (inp[8]) ? node162 : node153;
										assign node153 = (inp[4]) ? node155 : 3'b100;
											assign node155 = (inp[0]) ? node159 : node156;
												assign node156 = (inp[7]) ? 3'b110 : 3'b111;
												assign node159 = (inp[7]) ? 3'b111 : 3'b110;
										assign node162 = (inp[4]) ? node164 : 3'b111;
											assign node164 = (inp[7]) ? node168 : node165;
												assign node165 = (inp[0]) ? 3'b100 : 3'b101;
												assign node168 = (inp[0]) ? 3'b101 : 3'b100;
									assign node171 = (inp[0]) ? node183 : node172;
										assign node172 = (inp[4]) ? node180 : node173;
											assign node173 = (inp[8]) ? node177 : node174;
												assign node174 = (inp[7]) ? 3'b100 : 3'b101;
												assign node177 = (inp[7]) ? 3'b111 : 3'b110;
											assign node180 = (inp[7]) ? 3'b111 : 3'b110;
										assign node183 = (inp[4]) ? 3'b100 : 3'b110;
							assign node186 = (inp[3]) ? node222 : node187;
								assign node187 = (inp[7]) ? node205 : node188;
									assign node188 = (inp[2]) ? node198 : node189;
										assign node189 = (inp[4]) ? node193 : node190;
											assign node190 = (inp[8]) ? 3'b100 : 3'b110;
											assign node193 = (inp[0]) ? 3'b111 : node194;
												assign node194 = (inp[8]) ? 3'b110 : 3'b100;
										assign node198 = (inp[0]) ? 3'b101 : node199;
											assign node199 = (inp[4]) ? 3'b111 : node200;
												assign node200 = (inp[8]) ? 3'b100 : 3'b110;
									assign node205 = (inp[2]) ? node215 : node206;
										assign node206 = (inp[4]) ? node210 : node207;
											assign node207 = (inp[8]) ? 3'b101 : 3'b111;
											assign node210 = (inp[0]) ? 3'b110 : node211;
												assign node211 = (inp[8]) ? 3'b111 : 3'b101;
										assign node215 = (inp[0]) ? node217 : 3'b110;
											assign node217 = (inp[4]) ? 3'b100 : node218;
												assign node218 = (inp[8]) ? 3'b100 : 3'b110;
								assign node222 = (inp[2]) ? node246 : node223;
									assign node223 = (inp[7]) ? node237 : node224;
										assign node224 = (inp[0]) ? node232 : node225;
											assign node225 = (inp[4]) ? node229 : node226;
												assign node226 = (inp[8]) ? 3'b110 : 3'b100;
												assign node229 = (inp[8]) ? 3'b100 : 3'b110;
											assign node232 = (inp[8]) ? node234 : 3'b100;
												assign node234 = (inp[4]) ? 3'b101 : 3'b111;
										assign node237 = (inp[8]) ? node241 : node238;
											assign node238 = (inp[4]) ? 3'b111 : 3'b101;
											assign node241 = (inp[4]) ? node243 : 3'b110;
												assign node243 = (inp[0]) ? 3'b100 : 3'b101;
									assign node246 = (inp[7]) ? node254 : node247;
										assign node247 = (inp[4]) ? node251 : node248;
											assign node248 = (inp[8]) ? 3'b111 : 3'b101;
											assign node251 = (inp[8]) ? 3'b101 : 3'b111;
										assign node254 = (inp[4]) ? node258 : node255;
											assign node255 = (inp[8]) ? 3'b110 : 3'b101;
											assign node258 = (inp[8]) ? 3'b100 : 3'b110;
					assign node261 = (inp[3]) ? node395 : node262;
						assign node262 = (inp[5]) ? node336 : node263;
							assign node263 = (inp[7]) ? node303 : node264;
								assign node264 = (inp[0]) ? node284 : node265;
									assign node265 = (inp[9]) ? node275 : node266;
										assign node266 = (inp[8]) ? node270 : node267;
											assign node267 = (inp[4]) ? 3'b001 : 3'b011;
											assign node270 = (inp[4]) ? node272 : 3'b001;
												assign node272 = (inp[2]) ? 3'b010 : 3'b011;
										assign node275 = (inp[4]) ? node279 : node276;
											assign node276 = (inp[8]) ? 3'b000 : 3'b010;
											assign node279 = (inp[2]) ? 3'b011 : node280;
												assign node280 = (inp[8]) ? 3'b010 : 3'b000;
									assign node284 = (inp[2]) ? node294 : node285;
										assign node285 = (inp[8]) ? node289 : node286;
											assign node286 = (inp[9]) ? 3'b010 : 3'b011;
											assign node289 = (inp[4]) ? node291 : 3'b001;
												assign node291 = (inp[9]) ? 3'b011 : 3'b010;
										assign node294 = (inp[9]) ? node296 : 3'b000;
											assign node296 = (inp[4]) ? node300 : node297;
												assign node297 = (inp[8]) ? 3'b001 : 3'b011;
												assign node300 = (inp[8]) ? 3'b011 : 3'b001;
								assign node303 = (inp[9]) ? node323 : node304;
									assign node304 = (inp[2]) ? node314 : node305;
										assign node305 = (inp[8]) ? node309 : node306;
											assign node306 = (inp[4]) ? 3'b000 : 3'b010;
											assign node309 = (inp[4]) ? node311 : 3'b000;
												assign node311 = (inp[0]) ? 3'b011 : 3'b010;
										assign node314 = (inp[8]) ? node320 : node315;
											assign node315 = (inp[4]) ? node317 : 3'b011;
												assign node317 = (inp[0]) ? 3'b001 : 3'b000;
											assign node320 = (inp[4]) ? 3'b011 : 3'b001;
									assign node323 = (inp[2]) ? node331 : node324;
										assign node324 = (inp[4]) ? node328 : node325;
											assign node325 = (inp[8]) ? 3'b001 : 3'b011;
											assign node328 = (inp[8]) ? 3'b011 : 3'b001;
										assign node331 = (inp[0]) ? node333 : 3'b001;
											assign node333 = (inp[4]) ? 3'b010 : 3'b000;
							assign node336 = (inp[8]) ? node366 : node337;
								assign node337 = (inp[4]) ? node349 : node338;
									assign node338 = (inp[9]) ? node340 : 3'b011;
										assign node340 = (inp[2]) ? node344 : node341;
											assign node341 = (inp[7]) ? 3'b011 : 3'b010;
											assign node344 = (inp[0]) ? node346 : 3'b010;
												assign node346 = (inp[7]) ? 3'b010 : 3'b011;
									assign node349 = (inp[0]) ? node357 : node350;
										assign node350 = (inp[7]) ? node354 : node351;
											assign node351 = (inp[9]) ? 3'b000 : 3'b001;
											assign node354 = (inp[9]) ? 3'b001 : 3'b000;
										assign node357 = (inp[9]) ? node359 : 3'b000;
											assign node359 = (inp[7]) ? node363 : node360;
												assign node360 = (inp[2]) ? 3'b001 : 3'b000;
												assign node363 = (inp[2]) ? 3'b000 : 3'b001;
								assign node366 = (inp[4]) ? node380 : node367;
									assign node367 = (inp[7]) ? node373 : node368;
										assign node368 = (inp[9]) ? 3'b000 : node369;
											assign node369 = (inp[0]) ? 3'b000 : 3'b001;
										assign node373 = (inp[9]) ? 3'b001 : node374;
											assign node374 = (inp[0]) ? node376 : 3'b000;
												assign node376 = (inp[2]) ? 3'b001 : 3'b000;
									assign node380 = (inp[7]) ? node386 : node381;
										assign node381 = (inp[9]) ? 3'b011 : node382;
											assign node382 = (inp[2]) ? 3'b010 : 3'b011;
										assign node386 = (inp[2]) ? node392 : node387;
											assign node387 = (inp[0]) ? 3'b010 : node388;
												assign node388 = (inp[9]) ? 3'b011 : 3'b010;
											assign node392 = (inp[9]) ? 3'b010 : 3'b011;
						assign node395 = (inp[9]) ? node461 : node396;
							assign node396 = (inp[5]) ? node428 : node397;
								assign node397 = (inp[7]) ? node419 : node398;
									assign node398 = (inp[2]) ? node406 : node399;
										assign node399 = (inp[8]) ? node401 : 3'b001;
											assign node401 = (inp[4]) ? node403 : 3'b001;
												assign node403 = (inp[0]) ? 3'b010 : 3'b011;
										assign node406 = (inp[0]) ? node412 : node407;
											assign node407 = (inp[4]) ? node409 : 3'b001;
												assign node409 = (inp[8]) ? 3'b010 : 3'b001;
											assign node412 = (inp[8]) ? node416 : node413;
												assign node413 = (inp[4]) ? 3'b000 : 3'b010;
												assign node416 = (inp[4]) ? 3'b010 : 3'b000;
									assign node419 = (inp[2]) ? node425 : node420;
										assign node420 = (inp[8]) ? 3'b000 : node421;
											assign node421 = (inp[4]) ? 3'b000 : 3'b010;
										assign node425 = (inp[0]) ? 3'b001 : 3'b000;
								assign node428 = (inp[8]) ? node446 : node429;
									assign node429 = (inp[4]) ? node437 : node430;
										assign node430 = (inp[7]) ? 3'b000 : node431;
											assign node431 = (inp[0]) ? node433 : 3'b001;
												assign node433 = (inp[2]) ? 3'b000 : 3'b001;
										assign node437 = (inp[7]) ? node443 : node438;
											assign node438 = (inp[2]) ? 3'b010 : node439;
												assign node439 = (inp[0]) ? 3'b010 : 3'b011;
											assign node443 = (inp[0]) ? 3'b011 : 3'b010;
									assign node446 = (inp[4]) ? node454 : node447;
										assign node447 = (inp[0]) ? 3'b010 : node448;
											assign node448 = (inp[7]) ? node450 : 3'b011;
												assign node450 = (inp[2]) ? 3'b011 : 3'b010;
										assign node454 = (inp[7]) ? node456 : 3'b000;
											assign node456 = (inp[0]) ? 3'b001 : node457;
												assign node457 = (inp[2]) ? 3'b001 : 3'b000;
							assign node461 = (inp[0]) ? node493 : node462;
								assign node462 = (inp[7]) ? node480 : node463;
									assign node463 = (inp[8]) ? node469 : node464;
										assign node464 = (inp[5]) ? 3'b000 : node465;
											assign node465 = (inp[4]) ? 3'b000 : 3'b010;
										assign node469 = (inp[2]) ? node475 : node470;
											assign node470 = (inp[5]) ? 3'b010 : node471;
												assign node471 = (inp[4]) ? 3'b010 : 3'b000;
											assign node475 = (inp[4]) ? 3'b011 : node476;
												assign node476 = (inp[5]) ? 3'b011 : 3'b000;
									assign node480 = (inp[2]) ? node486 : node481;
										assign node481 = (inp[8]) ? 3'b011 : node482;
											assign node482 = (inp[5]) ? 3'b001 : 3'b011;
										assign node486 = (inp[5]) ? node488 : 3'b011;
											assign node488 = (inp[8]) ? node490 : 3'b010;
												assign node490 = (inp[4]) ? 3'b000 : 3'b010;
								assign node493 = (inp[7]) ? node513 : node494;
									assign node494 = (inp[8]) ? node506 : node495;
										assign node495 = (inp[2]) ? node501 : node496;
											assign node496 = (inp[4]) ? 3'b000 : node497;
												assign node497 = (inp[5]) ? 3'b000 : 3'b010;
											assign node501 = (inp[5]) ? node503 : 3'b001;
												assign node503 = (inp[4]) ? 3'b011 : 3'b001;
										assign node506 = (inp[4]) ? node510 : node507;
											assign node507 = (inp[5]) ? 3'b011 : 3'b001;
											assign node510 = (inp[5]) ? 3'b001 : 3'b011;
									assign node513 = (inp[4]) ? node521 : node514;
										assign node514 = (inp[5]) ? 3'b010 : node515;
											assign node515 = (inp[8]) ? 3'b001 : node516;
												assign node516 = (inp[2]) ? 3'b010 : 3'b011;
										assign node521 = (inp[5]) ? node525 : node522;
											assign node522 = (inp[2]) ? 3'b000 : 3'b001;
											assign node525 = (inp[8]) ? 3'b000 : 3'b010;
				assign node528 = (inp[0]) ? node778 : node529;
					assign node529 = (inp[4]) ? node669 : node530;
						assign node530 = (inp[8]) ? node584 : node531;
							assign node531 = (inp[3]) ? node569 : node532;
								assign node532 = (inp[11]) ? node554 : node533;
									assign node533 = (inp[5]) ? node547 : node534;
										assign node534 = (inp[2]) ? node540 : node535;
											assign node535 = (inp[7]) ? node537 : 3'b011;
												assign node537 = (inp[9]) ? 3'b011 : 3'b010;
											assign node540 = (inp[9]) ? node544 : node541;
												assign node541 = (inp[7]) ? 3'b010 : 3'b011;
												assign node544 = (inp[7]) ? 3'b011 : 3'b010;
										assign node547 = (inp[7]) ? node551 : node548;
											assign node548 = (inp[9]) ? 3'b010 : 3'b011;
											assign node551 = (inp[9]) ? 3'b011 : 3'b010;
									assign node554 = (inp[5]) ? node564 : node555;
										assign node555 = (inp[2]) ? node557 : 3'b011;
											assign node557 = (inp[9]) ? node561 : node558;
												assign node558 = (inp[7]) ? 3'b010 : 3'b011;
												assign node561 = (inp[7]) ? 3'b011 : 3'b010;
										assign node564 = (inp[9]) ? node566 : 3'b011;
											assign node566 = (inp[7]) ? 3'b011 : 3'b010;
								assign node569 = (inp[5]) ? node577 : node570;
									assign node570 = (inp[2]) ? 3'b011 : node571;
										assign node571 = (inp[9]) ? node573 : 3'b010;
											assign node573 = (inp[7]) ? 3'b011 : 3'b010;
									assign node577 = (inp[7]) ? node581 : node578;
										assign node578 = (inp[9]) ? 3'b000 : 3'b001;
										assign node581 = (inp[9]) ? 3'b001 : 3'b000;
							assign node584 = (inp[5]) ? node638 : node585;
								assign node585 = (inp[11]) ? node607 : node586;
									assign node586 = (inp[2]) ? node594 : node587;
										assign node587 = (inp[9]) ? node591 : node588;
											assign node588 = (inp[7]) ? 3'b000 : 3'b001;
											assign node591 = (inp[7]) ? 3'b001 : 3'b000;
										assign node594 = (inp[3]) ? node600 : node595;
											assign node595 = (inp[9]) ? node597 : 3'b001;
												assign node597 = (inp[7]) ? 3'b001 : 3'b000;
											assign node600 = (inp[7]) ? node604 : node601;
												assign node601 = (inp[9]) ? 3'b000 : 3'b001;
												assign node604 = (inp[9]) ? 3'b001 : 3'b000;
									assign node607 = (inp[3]) ? node623 : node608;
										assign node608 = (inp[2]) ? node616 : node609;
											assign node609 = (inp[9]) ? node613 : node610;
												assign node610 = (inp[7]) ? 3'b000 : 3'b001;
												assign node613 = (inp[7]) ? 3'b001 : 3'b000;
											assign node616 = (inp[7]) ? node620 : node617;
												assign node617 = (inp[9]) ? 3'b000 : 3'b001;
												assign node620 = (inp[9]) ? 3'b001 : 3'b000;
										assign node623 = (inp[2]) ? node631 : node624;
											assign node624 = (inp[9]) ? node628 : node625;
												assign node625 = (inp[7]) ? 3'b000 : 3'b001;
												assign node628 = (inp[7]) ? 3'b001 : 3'b000;
											assign node631 = (inp[9]) ? node635 : node632;
												assign node632 = (inp[7]) ? 3'b000 : 3'b001;
												assign node635 = (inp[7]) ? 3'b001 : 3'b000;
								assign node638 = (inp[3]) ? node648 : node639;
									assign node639 = (inp[11]) ? 3'b001 : node640;
										assign node640 = (inp[7]) ? node644 : node641;
											assign node641 = (inp[9]) ? 3'b000 : 3'b001;
											assign node644 = (inp[9]) ? 3'b001 : 3'b000;
									assign node648 = (inp[9]) ? node660 : node649;
										assign node649 = (inp[11]) ? node655 : node650;
											assign node650 = (inp[7]) ? node652 : 3'b011;
												assign node652 = (inp[2]) ? 3'b011 : 3'b010;
											assign node655 = (inp[2]) ? node657 : 3'b011;
												assign node657 = (inp[7]) ? 3'b011 : 3'b010;
										assign node660 = (inp[11]) ? node664 : node661;
											assign node661 = (inp[7]) ? 3'b011 : 3'b010;
											assign node664 = (inp[2]) ? node666 : 3'b010;
												assign node666 = (inp[7]) ? 3'b010 : 3'b011;
						assign node669 = (inp[8]) ? node729 : node670;
							assign node670 = (inp[3]) ? node706 : node671;
								assign node671 = (inp[5]) ? node689 : node672;
									assign node672 = (inp[11]) ? node684 : node673;
										assign node673 = (inp[2]) ? node679 : node674;
											assign node674 = (inp[7]) ? node676 : 3'b000;
												assign node676 = (inp[9]) ? 3'b001 : 3'b000;
											assign node679 = (inp[7]) ? 3'b000 : node680;
												assign node680 = (inp[9]) ? 3'b000 : 3'b001;
										assign node684 = (inp[9]) ? node686 : 3'b001;
											assign node686 = (inp[7]) ? 3'b001 : 3'b000;
									assign node689 = (inp[11]) ? node691 : 3'b001;
										assign node691 = (inp[2]) ? node699 : node692;
											assign node692 = (inp[7]) ? node696 : node693;
												assign node693 = (inp[9]) ? 3'b000 : 3'b001;
												assign node696 = (inp[9]) ? 3'b001 : 3'b000;
											assign node699 = (inp[7]) ? node703 : node700;
												assign node700 = (inp[9]) ? 3'b000 : 3'b001;
												assign node703 = (inp[9]) ? 3'b001 : 3'b000;
								assign node706 = (inp[5]) ? node712 : node707;
									assign node707 = (inp[9]) ? 3'b001 : node708;
										assign node708 = (inp[7]) ? 3'b000 : 3'b001;
									assign node712 = (inp[11]) ? node724 : node713;
										assign node713 = (inp[9]) ? node719 : node714;
											assign node714 = (inp[2]) ? node716 : 3'b010;
												assign node716 = (inp[7]) ? 3'b011 : 3'b010;
											assign node719 = (inp[2]) ? node721 : 3'b011;
												assign node721 = (inp[7]) ? 3'b010 : 3'b011;
										assign node724 = (inp[9]) ? 3'b010 : node725;
											assign node725 = (inp[7]) ? 3'b010 : 3'b011;
							assign node729 = (inp[5]) ? node755 : node730;
								assign node730 = (inp[11]) ? node746 : node731;
									assign node731 = (inp[2]) ? node739 : node732;
										assign node732 = (inp[9]) ? node736 : node733;
											assign node733 = (inp[7]) ? 3'b010 : 3'b011;
											assign node736 = (inp[7]) ? 3'b011 : 3'b010;
										assign node739 = (inp[7]) ? node743 : node740;
											assign node740 = (inp[9]) ? 3'b011 : 3'b010;
											assign node743 = (inp[9]) ? 3'b010 : 3'b011;
									assign node746 = (inp[7]) ? node748 : 3'b010;
										assign node748 = (inp[2]) ? node752 : node749;
											assign node749 = (inp[9]) ? 3'b011 : 3'b010;
											assign node752 = (inp[9]) ? 3'b010 : 3'b011;
								assign node755 = (inp[3]) ? node769 : node756;
									assign node756 = (inp[7]) ? node762 : node757;
										assign node757 = (inp[9]) ? 3'b010 : node758;
											assign node758 = (inp[2]) ? 3'b010 : 3'b011;
										assign node762 = (inp[9]) ? node766 : node763;
											assign node763 = (inp[2]) ? 3'b011 : 3'b010;
											assign node766 = (inp[2]) ? 3'b010 : 3'b011;
									assign node769 = (inp[7]) ? 3'b000 : node770;
										assign node770 = (inp[2]) ? node774 : node771;
											assign node771 = (inp[9]) ? 3'b000 : 3'b001;
											assign node774 = (inp[9]) ? 3'b001 : 3'b000;
					assign node778 = (inp[7]) ? node884 : node779;
						assign node779 = (inp[9]) ? node835 : node780;
							assign node780 = (inp[2]) ? node804 : node781;
								assign node781 = (inp[8]) ? node793 : node782;
									assign node782 = (inp[4]) ? node788 : node783;
										assign node783 = (inp[5]) ? node785 : 3'b011;
											assign node785 = (inp[3]) ? 3'b001 : 3'b011;
										assign node788 = (inp[5]) ? node790 : 3'b001;
											assign node790 = (inp[3]) ? 3'b010 : 3'b001;
									assign node793 = (inp[4]) ? node799 : node794;
										assign node794 = (inp[3]) ? node796 : 3'b001;
											assign node796 = (inp[5]) ? 3'b010 : 3'b001;
										assign node799 = (inp[5]) ? node801 : 3'b010;
											assign node801 = (inp[3]) ? 3'b000 : 3'b010;
								assign node804 = (inp[3]) ? node812 : node805;
									assign node805 = (inp[8]) ? node809 : node806;
										assign node806 = (inp[4]) ? 3'b000 : 3'b010;
										assign node809 = (inp[4]) ? 3'b010 : 3'b000;
									assign node812 = (inp[11]) ? node828 : node813;
										assign node813 = (inp[5]) ? node821 : node814;
											assign node814 = (inp[8]) ? node818 : node815;
												assign node815 = (inp[4]) ? 3'b000 : 3'b010;
												assign node818 = (inp[4]) ? 3'b010 : 3'b000;
											assign node821 = (inp[8]) ? node825 : node822;
												assign node822 = (inp[4]) ? 3'b010 : 3'b000;
												assign node825 = (inp[4]) ? 3'b000 : 3'b010;
										assign node828 = (inp[4]) ? 3'b010 : node829;
											assign node829 = (inp[8]) ? node831 : 3'b010;
												assign node831 = (inp[5]) ? 3'b010 : 3'b000;
							assign node835 = (inp[2]) ? node859 : node836;
								assign node836 = (inp[4]) ? node848 : node837;
									assign node837 = (inp[8]) ? node843 : node838;
										assign node838 = (inp[3]) ? node840 : 3'b010;
											assign node840 = (inp[5]) ? 3'b000 : 3'b010;
										assign node843 = (inp[5]) ? node845 : 3'b000;
											assign node845 = (inp[3]) ? 3'b011 : 3'b000;
									assign node848 = (inp[8]) ? node854 : node849;
										assign node849 = (inp[3]) ? node851 : 3'b000;
											assign node851 = (inp[5]) ? 3'b011 : 3'b000;
										assign node854 = (inp[5]) ? node856 : 3'b011;
											assign node856 = (inp[3]) ? 3'b001 : 3'b011;
								assign node859 = (inp[3]) ? node867 : node860;
									assign node860 = (inp[4]) ? node864 : node861;
										assign node861 = (inp[8]) ? 3'b001 : 3'b011;
										assign node864 = (inp[8]) ? 3'b011 : 3'b001;
									assign node867 = (inp[5]) ? node879 : node868;
										assign node868 = (inp[11]) ? node874 : node869;
											assign node869 = (inp[8]) ? node871 : 3'b001;
												assign node871 = (inp[4]) ? 3'b011 : 3'b001;
											assign node874 = (inp[4]) ? node876 : 3'b011;
												assign node876 = (inp[8]) ? 3'b011 : 3'b001;
										assign node879 = (inp[8]) ? node881 : 3'b011;
											assign node881 = (inp[4]) ? 3'b001 : 3'b011;
						assign node884 = (inp[9]) ? node926 : node885;
							assign node885 = (inp[2]) ? node907 : node886;
								assign node886 = (inp[3]) ? node892 : node887;
									assign node887 = (inp[8]) ? 3'b000 : node888;
										assign node888 = (inp[4]) ? 3'b000 : 3'b010;
									assign node892 = (inp[8]) ? node900 : node893;
										assign node893 = (inp[5]) ? node897 : node894;
											assign node894 = (inp[4]) ? 3'b000 : 3'b010;
											assign node897 = (inp[4]) ? 3'b011 : 3'b000;
										assign node900 = (inp[4]) ? node904 : node901;
											assign node901 = (inp[5]) ? 3'b011 : 3'b000;
											assign node904 = (inp[5]) ? 3'b001 : 3'b011;
								assign node907 = (inp[8]) ? node919 : node908;
									assign node908 = (inp[4]) ? node914 : node909;
										assign node909 = (inp[5]) ? node911 : 3'b011;
											assign node911 = (inp[3]) ? 3'b001 : 3'b011;
										assign node914 = (inp[5]) ? node916 : 3'b001;
											assign node916 = (inp[3]) ? 3'b011 : 3'b001;
									assign node919 = (inp[4]) ? node921 : 3'b001;
										assign node921 = (inp[3]) ? node923 : 3'b011;
											assign node923 = (inp[5]) ? 3'b001 : 3'b011;
							assign node926 = (inp[2]) ? node946 : node927;
								assign node927 = (inp[4]) ? node935 : node928;
									assign node928 = (inp[8]) ? 3'b001 : node929;
										assign node929 = (inp[3]) ? node931 : 3'b011;
											assign node931 = (inp[5]) ? 3'b001 : 3'b011;
									assign node935 = (inp[8]) ? node941 : node936;
										assign node936 = (inp[3]) ? node938 : 3'b001;
											assign node938 = (inp[5]) ? 3'b010 : 3'b001;
										assign node941 = (inp[5]) ? node943 : 3'b010;
											assign node943 = (inp[3]) ? 3'b000 : 3'b010;
								assign node946 = (inp[4]) ? node958 : node947;
									assign node947 = (inp[8]) ? node953 : node948;
										assign node948 = (inp[3]) ? node950 : 3'b010;
											assign node950 = (inp[5]) ? 3'b000 : 3'b010;
										assign node953 = (inp[3]) ? node955 : 3'b000;
											assign node955 = (inp[5]) ? 3'b010 : 3'b000;
									assign node958 = (inp[8]) ? node964 : node959;
										assign node959 = (inp[3]) ? node961 : 3'b000;
											assign node961 = (inp[5]) ? 3'b010 : 3'b000;
										assign node964 = (inp[3]) ? 3'b000 : 3'b010;
			assign node967 = (inp[11]) ? node1449 : node968;
				assign node968 = (inp[1]) ? node1214 : node969;
					assign node969 = (inp[8]) ? node1091 : node970;
						assign node970 = (inp[4]) ? node1024 : node971;
							assign node971 = (inp[3]) ? node993 : node972;
								assign node972 = (inp[9]) ? node982 : node973;
									assign node973 = (inp[7]) ? node979 : node974;
										assign node974 = (inp[2]) ? node976 : 3'b011;
											assign node976 = (inp[0]) ? 3'b010 : 3'b011;
										assign node979 = (inp[2]) ? 3'b011 : 3'b010;
									assign node982 = (inp[7]) ? node988 : node983;
										assign node983 = (inp[0]) ? node985 : 3'b010;
											assign node985 = (inp[2]) ? 3'b011 : 3'b010;
										assign node988 = (inp[0]) ? node990 : 3'b011;
											assign node990 = (inp[2]) ? 3'b010 : 3'b011;
								assign node993 = (inp[5]) ? node1007 : node994;
									assign node994 = (inp[2]) ? node1000 : node995;
										assign node995 = (inp[9]) ? 3'b011 : node996;
											assign node996 = (inp[7]) ? 3'b010 : 3'b011;
										assign node1000 = (inp[9]) ? 3'b010 : node1001;
											assign node1001 = (inp[7]) ? 3'b010 : node1002;
												assign node1002 = (inp[0]) ? 3'b010 : 3'b011;
									assign node1007 = (inp[2]) ? node1015 : node1008;
										assign node1008 = (inp[9]) ? node1012 : node1009;
											assign node1009 = (inp[7]) ? 3'b000 : 3'b001;
											assign node1012 = (inp[7]) ? 3'b001 : 3'b000;
										assign node1015 = (inp[0]) ? 3'b000 : node1016;
											assign node1016 = (inp[7]) ? node1020 : node1017;
												assign node1017 = (inp[9]) ? 3'b000 : 3'b001;
												assign node1020 = (inp[9]) ? 3'b001 : 3'b000;
							assign node1024 = (inp[3]) ? node1060 : node1025;
								assign node1025 = (inp[5]) ? node1043 : node1026;
									assign node1026 = (inp[2]) ? node1034 : node1027;
										assign node1027 = (inp[7]) ? node1031 : node1028;
											assign node1028 = (inp[9]) ? 3'b000 : 3'b001;
											assign node1031 = (inp[9]) ? 3'b001 : 3'b000;
										assign node1034 = (inp[0]) ? 3'b001 : node1035;
											assign node1035 = (inp[7]) ? node1039 : node1036;
												assign node1036 = (inp[9]) ? 3'b000 : 3'b001;
												assign node1039 = (inp[9]) ? 3'b001 : 3'b000;
									assign node1043 = (inp[0]) ? node1051 : node1044;
										assign node1044 = (inp[7]) ? node1048 : node1045;
											assign node1045 = (inp[9]) ? 3'b000 : 3'b001;
											assign node1048 = (inp[9]) ? 3'b001 : 3'b000;
										assign node1051 = (inp[2]) ? 3'b000 : node1052;
											assign node1052 = (inp[7]) ? node1056 : node1053;
												assign node1053 = (inp[9]) ? 3'b000 : 3'b001;
												assign node1056 = (inp[9]) ? 3'b001 : 3'b000;
								assign node1060 = (inp[5]) ? node1078 : node1061;
									assign node1061 = (inp[0]) ? node1069 : node1062;
										assign node1062 = (inp[2]) ? node1064 : 3'b000;
											assign node1064 = (inp[7]) ? 3'b000 : node1065;
												assign node1065 = (inp[9]) ? 3'b000 : 3'b001;
										assign node1069 = (inp[9]) ? 3'b001 : node1070;
											assign node1070 = (inp[2]) ? node1074 : node1071;
												assign node1071 = (inp[7]) ? 3'b000 : 3'b001;
												assign node1074 = (inp[7]) ? 3'b001 : 3'b000;
									assign node1078 = (inp[9]) ? node1084 : node1079;
										assign node1079 = (inp[7]) ? node1081 : 3'b010;
											assign node1081 = (inp[2]) ? 3'b011 : 3'b010;
										assign node1084 = (inp[7]) ? node1088 : node1085;
											assign node1085 = (inp[0]) ? 3'b011 : 3'b010;
											assign node1088 = (inp[2]) ? 3'b010 : 3'b011;
						assign node1091 = (inp[4]) ? node1153 : node1092;
							assign node1092 = (inp[3]) ? node1124 : node1093;
								assign node1093 = (inp[2]) ? node1101 : node1094;
									assign node1094 = (inp[7]) ? node1098 : node1095;
										assign node1095 = (inp[9]) ? 3'b000 : 3'b001;
										assign node1098 = (inp[9]) ? 3'b001 : 3'b000;
									assign node1101 = (inp[5]) ? node1111 : node1102;
										assign node1102 = (inp[7]) ? node1104 : 3'b001;
											assign node1104 = (inp[9]) ? node1108 : node1105;
												assign node1105 = (inp[0]) ? 3'b001 : 3'b000;
												assign node1108 = (inp[0]) ? 3'b000 : 3'b001;
										assign node1111 = (inp[7]) ? node1119 : node1112;
											assign node1112 = (inp[0]) ? node1116 : node1113;
												assign node1113 = (inp[9]) ? 3'b000 : 3'b001;
												assign node1116 = (inp[9]) ? 3'b001 : 3'b000;
											assign node1119 = (inp[9]) ? node1121 : 3'b001;
												assign node1121 = (inp[0]) ? 3'b000 : 3'b001;
								assign node1124 = (inp[5]) ? node1140 : node1125;
									assign node1125 = (inp[9]) ? node1131 : node1126;
										assign node1126 = (inp[7]) ? 3'b000 : node1127;
											assign node1127 = (inp[2]) ? 3'b000 : 3'b001;
										assign node1131 = (inp[0]) ? node1135 : node1132;
											assign node1132 = (inp[2]) ? 3'b001 : 3'b000;
											assign node1135 = (inp[2]) ? node1137 : 3'b001;
												assign node1137 = (inp[7]) ? 3'b000 : 3'b001;
									assign node1140 = (inp[9]) ? node1146 : node1141;
										assign node1141 = (inp[7]) ? 3'b011 : node1142;
											assign node1142 = (inp[2]) ? 3'b010 : 3'b011;
										assign node1146 = (inp[2]) ? 3'b011 : node1147;
											assign node1147 = (inp[0]) ? 3'b010 : node1148;
												assign node1148 = (inp[7]) ? 3'b011 : 3'b010;
							assign node1153 = (inp[5]) ? node1189 : node1154;
								assign node1154 = (inp[3]) ? node1174 : node1155;
									assign node1155 = (inp[7]) ? node1165 : node1156;
										assign node1156 = (inp[2]) ? 3'b010 : node1157;
											assign node1157 = (inp[9]) ? node1161 : node1158;
												assign node1158 = (inp[0]) ? 3'b010 : 3'b011;
												assign node1161 = (inp[0]) ? 3'b011 : 3'b010;
										assign node1165 = (inp[9]) ? node1171 : node1166;
											assign node1166 = (inp[0]) ? 3'b011 : node1167;
												assign node1167 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1171 = (inp[0]) ? 3'b010 : 3'b011;
									assign node1174 = (inp[7]) ? node1184 : node1175;
										assign node1175 = (inp[9]) ? node1179 : node1176;
											assign node1176 = (inp[0]) ? 3'b010 : 3'b011;
											assign node1179 = (inp[0]) ? 3'b011 : node1180;
												assign node1180 = (inp[2]) ? 3'b011 : 3'b010;
										assign node1184 = (inp[0]) ? node1186 : 3'b010;
											assign node1186 = (inp[9]) ? 3'b010 : 3'b011;
								assign node1189 = (inp[3]) ? node1201 : node1190;
									assign node1190 = (inp[0]) ? node1196 : node1191;
										assign node1191 = (inp[2]) ? node1193 : 3'b010;
											assign node1193 = (inp[7]) ? 3'b010 : 3'b011;
										assign node1196 = (inp[7]) ? 3'b011 : node1197;
											assign node1197 = (inp[9]) ? 3'b011 : 3'b010;
									assign node1201 = (inp[7]) ? node1207 : node1202;
										assign node1202 = (inp[9]) ? 3'b001 : node1203;
											assign node1203 = (inp[2]) ? 3'b000 : 3'b001;
										assign node1207 = (inp[9]) ? 3'b000 : node1208;
											assign node1208 = (inp[2]) ? 3'b001 : node1209;
												assign node1209 = (inp[0]) ? 3'b001 : 3'b000;
					assign node1214 = (inp[7]) ? node1338 : node1215;
						assign node1215 = (inp[9]) ? node1277 : node1216;
							assign node1216 = (inp[2]) ? node1242 : node1217;
								assign node1217 = (inp[0]) ? node1233 : node1218;
									assign node1218 = (inp[3]) ? node1226 : node1219;
										assign node1219 = (inp[4]) ? 3'b101 : node1220;
											assign node1220 = (inp[8]) ? node1222 : 3'b101;
												assign node1222 = (inp[5]) ? 3'b111 : 3'b101;
										assign node1226 = (inp[8]) ? node1230 : node1227;
											assign node1227 = (inp[4]) ? 3'b111 : 3'b101;
											assign node1230 = (inp[4]) ? 3'b101 : 3'b111;
									assign node1233 = (inp[4]) ? node1235 : 3'b101;
										assign node1235 = (inp[8]) ? node1237 : 3'b110;
											assign node1237 = (inp[5]) ? 3'b100 : node1238;
												assign node1238 = (inp[3]) ? 3'b100 : 3'b110;
								assign node1242 = (inp[0]) ? node1264 : node1243;
									assign node1243 = (inp[4]) ? node1253 : node1244;
										assign node1244 = (inp[8]) ? node1250 : node1245;
											assign node1245 = (inp[5]) ? 3'b101 : node1246;
												assign node1246 = (inp[3]) ? 3'b101 : 3'b111;
											assign node1250 = (inp[3]) ? 3'b110 : 3'b101;
										assign node1253 = (inp[8]) ? node1259 : node1254;
											assign node1254 = (inp[5]) ? 3'b110 : node1255;
												assign node1255 = (inp[3]) ? 3'b110 : 3'b101;
											assign node1259 = (inp[5]) ? 3'b100 : node1260;
												assign node1260 = (inp[3]) ? 3'b100 : 3'b110;
									assign node1264 = (inp[3]) ? node1272 : node1265;
										assign node1265 = (inp[4]) ? 3'b110 : node1266;
											assign node1266 = (inp[5]) ? node1268 : 3'b110;
												assign node1268 = (inp[8]) ? 3'b110 : 3'b100;
										assign node1272 = (inp[5]) ? 3'b100 : node1273;
											assign node1273 = (inp[8]) ? 3'b110 : 3'b100;
							assign node1277 = (inp[0]) ? node1311 : node1278;
								assign node1278 = (inp[2]) ? node1294 : node1279;
									assign node1279 = (inp[4]) ? node1285 : node1280;
										assign node1280 = (inp[5]) ? node1282 : 3'b100;
											assign node1282 = (inp[8]) ? 3'b110 : 3'b100;
										assign node1285 = (inp[8]) ? node1291 : node1286;
											assign node1286 = (inp[5]) ? 3'b110 : node1287;
												assign node1287 = (inp[3]) ? 3'b110 : 3'b100;
											assign node1291 = (inp[3]) ? 3'b100 : 3'b110;
									assign node1294 = (inp[8]) ? node1302 : node1295;
										assign node1295 = (inp[4]) ? node1297 : 3'b100;
											assign node1297 = (inp[5]) ? 3'b111 : node1298;
												assign node1298 = (inp[3]) ? 3'b111 : 3'b100;
										assign node1302 = (inp[3]) ? 3'b111 : node1303;
											assign node1303 = (inp[4]) ? node1307 : node1304;
												assign node1304 = (inp[5]) ? 3'b111 : 3'b100;
												assign node1307 = (inp[5]) ? 3'b101 : 3'b111;
								assign node1311 = (inp[2]) ? node1321 : node1312;
									assign node1312 = (inp[4]) ? node1318 : node1313;
										assign node1313 = (inp[8]) ? 3'b111 : node1314;
											assign node1314 = (inp[3]) ? 3'b100 : 3'b110;
										assign node1318 = (inp[8]) ? 3'b101 : 3'b111;
									assign node1321 = (inp[8]) ? node1333 : node1322;
										assign node1322 = (inp[4]) ? node1328 : node1323;
											assign node1323 = (inp[5]) ? 3'b101 : node1324;
												assign node1324 = (inp[3]) ? 3'b101 : 3'b111;
											assign node1328 = (inp[3]) ? 3'b111 : node1329;
												assign node1329 = (inp[5]) ? 3'b111 : 3'b101;
										assign node1333 = (inp[4]) ? node1335 : 3'b111;
											assign node1335 = (inp[5]) ? 3'b101 : 3'b111;
						assign node1338 = (inp[3]) ? node1408 : node1339;
							assign node1339 = (inp[0]) ? node1377 : node1340;
								assign node1340 = (inp[9]) ? node1358 : node1341;
									assign node1341 = (inp[2]) ? node1351 : node1342;
										assign node1342 = (inp[8]) ? node1344 : 3'b110;
											assign node1344 = (inp[5]) ? node1348 : node1345;
												assign node1345 = (inp[4]) ? 3'b110 : 3'b100;
												assign node1348 = (inp[4]) ? 3'b100 : 3'b110;
										assign node1351 = (inp[5]) ? node1353 : 3'b100;
											assign node1353 = (inp[8]) ? 3'b111 : node1354;
												assign node1354 = (inp[4]) ? 3'b111 : 3'b100;
									assign node1358 = (inp[2]) ? node1368 : node1359;
										assign node1359 = (inp[5]) ? 3'b111 : node1360;
											assign node1360 = (inp[8]) ? node1364 : node1361;
												assign node1361 = (inp[4]) ? 3'b101 : 3'b111;
												assign node1364 = (inp[4]) ? 3'b111 : 3'b101;
										assign node1368 = (inp[8]) ? node1374 : node1369;
											assign node1369 = (inp[4]) ? 3'b101 : node1370;
												assign node1370 = (inp[5]) ? 3'b101 : 3'b111;
											assign node1374 = (inp[4]) ? 3'b100 : 3'b110;
								assign node1377 = (inp[9]) ? node1397 : node1378;
									assign node1378 = (inp[2]) ? node1386 : node1379;
										assign node1379 = (inp[8]) ? node1381 : 3'b100;
											assign node1381 = (inp[4]) ? node1383 : 3'b100;
												assign node1383 = (inp[5]) ? 3'b101 : 3'b111;
										assign node1386 = (inp[8]) ? node1392 : node1387;
											assign node1387 = (inp[5]) ? 3'b111 : node1388;
												assign node1388 = (inp[4]) ? 3'b101 : 3'b111;
											assign node1392 = (inp[5]) ? 3'b101 : node1393;
												assign node1393 = (inp[4]) ? 3'b111 : 3'b101;
									assign node1397 = (inp[4]) ? node1405 : node1398;
										assign node1398 = (inp[2]) ? node1400 : 3'b110;
											assign node1400 = (inp[8]) ? 3'b100 : node1401;
												assign node1401 = (inp[5]) ? 3'b100 : 3'b110;
										assign node1405 = (inp[5]) ? 3'b100 : 3'b101;
							assign node1408 = (inp[9]) ? node1430 : node1409;
								assign node1409 = (inp[2]) ? node1417 : node1410;
									assign node1410 = (inp[0]) ? node1412 : 3'b110;
										assign node1412 = (inp[8]) ? 3'b111 : node1413;
											assign node1413 = (inp[4]) ? 3'b111 : 3'b100;
									assign node1417 = (inp[5]) ? node1425 : node1418;
										assign node1418 = (inp[4]) ? node1422 : node1419;
											assign node1419 = (inp[8]) ? 3'b111 : 3'b101;
											assign node1422 = (inp[0]) ? 3'b111 : 3'b101;
										assign node1425 = (inp[4]) ? node1427 : 3'b111;
											assign node1427 = (inp[8]) ? 3'b101 : 3'b111;
								assign node1430 = (inp[2]) ? node1442 : node1431;
									assign node1431 = (inp[0]) ? node1437 : node1432;
										assign node1432 = (inp[8]) ? node1434 : 3'b111;
											assign node1434 = (inp[4]) ? 3'b101 : 3'b111;
										assign node1437 = (inp[4]) ? 3'b110 : node1438;
											assign node1438 = (inp[8]) ? 3'b110 : 3'b101;
									assign node1442 = (inp[8]) ? 3'b110 : node1443;
										assign node1443 = (inp[4]) ? 3'b110 : node1444;
											assign node1444 = (inp[0]) ? 3'b100 : 3'b101;
				assign node1449 = (inp[3]) ? node1723 : node1450;
					assign node1450 = (inp[0]) ? node1586 : node1451;
						assign node1451 = (inp[1]) ? node1521 : node1452;
							assign node1452 = (inp[2]) ? node1482 : node1453;
								assign node1453 = (inp[4]) ? node1469 : node1454;
									assign node1454 = (inp[8]) ? node1458 : node1455;
										assign node1455 = (inp[5]) ? 3'b100 : 3'b110;
										assign node1458 = (inp[5]) ? node1464 : node1459;
											assign node1459 = (inp[7]) ? node1461 : 3'b100;
												assign node1461 = (inp[9]) ? 3'b101 : 3'b100;
											assign node1464 = (inp[7]) ? 3'b110 : node1465;
												assign node1465 = (inp[9]) ? 3'b110 : 3'b111;
									assign node1469 = (inp[8]) ? node1475 : node1470;
										assign node1470 = (inp[9]) ? node1472 : 3'b110;
											assign node1472 = (inp[7]) ? 3'b111 : 3'b110;
										assign node1475 = (inp[5]) ? 3'b101 : node1476;
											assign node1476 = (inp[7]) ? 3'b111 : node1477;
												assign node1477 = (inp[9]) ? 3'b110 : 3'b111;
								assign node1482 = (inp[9]) ? node1506 : node1483;
									assign node1483 = (inp[4]) ? node1495 : node1484;
										assign node1484 = (inp[5]) ? node1488 : node1485;
											assign node1485 = (inp[8]) ? 3'b101 : 3'b111;
											assign node1488 = (inp[8]) ? node1492 : node1489;
												assign node1489 = (inp[7]) ? 3'b100 : 3'b101;
												assign node1492 = (inp[7]) ? 3'b111 : 3'b110;
										assign node1495 = (inp[7]) ? node1501 : node1496;
											assign node1496 = (inp[8]) ? node1498 : 3'b110;
												assign node1498 = (inp[5]) ? 3'b100 : 3'b110;
											assign node1501 = (inp[5]) ? 3'b111 : node1502;
												assign node1502 = (inp[8]) ? 3'b111 : 3'b100;
									assign node1506 = (inp[8]) ? node1512 : node1507;
										assign node1507 = (inp[7]) ? node1509 : 3'b111;
											assign node1509 = (inp[5]) ? 3'b101 : 3'b111;
										assign node1512 = (inp[4]) ? node1516 : node1513;
											assign node1513 = (inp[7]) ? 3'b101 : 3'b100;
											assign node1516 = (inp[7]) ? 3'b100 : node1517;
												assign node1517 = (inp[5]) ? 3'b101 : 3'b111;
							assign node1521 = (inp[5]) ? node1553 : node1522;
								assign node1522 = (inp[9]) ? node1540 : node1523;
									assign node1523 = (inp[7]) ? node1531 : node1524;
										assign node1524 = (inp[4]) ? node1528 : node1525;
											assign node1525 = (inp[8]) ? 3'b101 : 3'b111;
											assign node1528 = (inp[8]) ? 3'b110 : 3'b101;
										assign node1531 = (inp[8]) ? node1535 : node1532;
											assign node1532 = (inp[4]) ? 3'b100 : 3'b110;
											assign node1535 = (inp[2]) ? 3'b111 : node1536;
												assign node1536 = (inp[4]) ? 3'b110 : 3'b100;
									assign node1540 = (inp[7]) ? node1548 : node1541;
										assign node1541 = (inp[8]) ? node1545 : node1542;
											assign node1542 = (inp[4]) ? 3'b100 : 3'b110;
											assign node1545 = (inp[4]) ? 3'b110 : 3'b100;
										assign node1548 = (inp[4]) ? node1550 : 3'b101;
											assign node1550 = (inp[8]) ? 3'b110 : 3'b101;
								assign node1553 = (inp[8]) ? node1563 : node1554;
									assign node1554 = (inp[4]) ? 3'b111 : node1555;
										assign node1555 = (inp[9]) ? node1559 : node1556;
											assign node1556 = (inp[7]) ? 3'b100 : 3'b101;
											assign node1559 = (inp[7]) ? 3'b101 : 3'b100;
									assign node1563 = (inp[4]) ? node1579 : node1564;
										assign node1564 = (inp[7]) ? node1572 : node1565;
											assign node1565 = (inp[2]) ? node1569 : node1566;
												assign node1566 = (inp[9]) ? 3'b110 : 3'b111;
												assign node1569 = (inp[9]) ? 3'b111 : 3'b110;
											assign node1572 = (inp[2]) ? node1576 : node1573;
												assign node1573 = (inp[9]) ? 3'b111 : 3'b110;
												assign node1576 = (inp[9]) ? 3'b110 : 3'b111;
										assign node1579 = (inp[2]) ? 3'b100 : node1580;
											assign node1580 = (inp[9]) ? 3'b101 : node1581;
												assign node1581 = (inp[7]) ? 3'b100 : 3'b101;
						assign node1586 = (inp[7]) ? node1648 : node1587;
							assign node1587 = (inp[9]) ? node1617 : node1588;
								assign node1588 = (inp[2]) ? node1604 : node1589;
									assign node1589 = (inp[1]) ? node1591 : 3'b101;
										assign node1591 = (inp[4]) ? node1599 : node1592;
											assign node1592 = (inp[8]) ? node1596 : node1593;
												assign node1593 = (inp[5]) ? 3'b101 : 3'b111;
												assign node1596 = (inp[5]) ? 3'b110 : 3'b101;
											assign node1599 = (inp[5]) ? node1601 : 3'b110;
												assign node1601 = (inp[8]) ? 3'b100 : 3'b110;
									assign node1604 = (inp[4]) ? node1612 : node1605;
										assign node1605 = (inp[1]) ? 3'b100 : node1606;
											assign node1606 = (inp[5]) ? 3'b110 : node1607;
												assign node1607 = (inp[8]) ? 3'b100 : 3'b110;
										assign node1612 = (inp[5]) ? node1614 : 3'b110;
											assign node1614 = (inp[8]) ? 3'b100 : 3'b110;
								assign node1617 = (inp[2]) ? node1629 : node1618;
									assign node1618 = (inp[5]) ? node1624 : node1619;
										assign node1619 = (inp[1]) ? node1621 : 3'b100;
											assign node1621 = (inp[8]) ? 3'b111 : 3'b110;
										assign node1624 = (inp[8]) ? node1626 : 3'b111;
											assign node1626 = (inp[4]) ? 3'b101 : 3'b111;
									assign node1629 = (inp[4]) ? node1637 : node1630;
										assign node1630 = (inp[5]) ? node1634 : node1631;
											assign node1631 = (inp[8]) ? 3'b101 : 3'b111;
											assign node1634 = (inp[8]) ? 3'b111 : 3'b101;
										assign node1637 = (inp[1]) ? node1643 : node1638;
											assign node1638 = (inp[5]) ? 3'b101 : node1639;
												assign node1639 = (inp[8]) ? 3'b111 : 3'b101;
											assign node1643 = (inp[8]) ? 3'b101 : node1644;
												assign node1644 = (inp[5]) ? 3'b111 : 3'b101;
							assign node1648 = (inp[9]) ? node1688 : node1649;
								assign node1649 = (inp[2]) ? node1665 : node1650;
									assign node1650 = (inp[4]) ? node1658 : node1651;
										assign node1651 = (inp[5]) ? node1655 : node1652;
											assign node1652 = (inp[8]) ? 3'b100 : 3'b110;
											assign node1655 = (inp[8]) ? 3'b111 : 3'b100;
										assign node1658 = (inp[5]) ? node1662 : node1659;
											assign node1659 = (inp[8]) ? 3'b111 : 3'b100;
											assign node1662 = (inp[8]) ? 3'b101 : 3'b111;
									assign node1665 = (inp[1]) ? node1679 : node1666;
										assign node1666 = (inp[4]) ? node1674 : node1667;
											assign node1667 = (inp[8]) ? node1671 : node1668;
												assign node1668 = (inp[5]) ? 3'b101 : 3'b111;
												assign node1671 = (inp[5]) ? 3'b111 : 3'b101;
											assign node1674 = (inp[5]) ? 3'b111 : node1675;
												assign node1675 = (inp[8]) ? 3'b111 : 3'b101;
										assign node1679 = (inp[8]) ? node1681 : 3'b111;
											assign node1681 = (inp[5]) ? node1685 : node1682;
												assign node1682 = (inp[4]) ? 3'b111 : 3'b101;
												assign node1685 = (inp[4]) ? 3'b101 : 3'b111;
								assign node1688 = (inp[2]) ? node1706 : node1689;
									assign node1689 = (inp[8]) ? node1695 : node1690;
										assign node1690 = (inp[5]) ? node1692 : 3'b101;
											assign node1692 = (inp[4]) ? 3'b110 : 3'b101;
										assign node1695 = (inp[1]) ? node1701 : node1696;
											assign node1696 = (inp[5]) ? 3'b110 : node1697;
												assign node1697 = (inp[4]) ? 3'b110 : 3'b101;
											assign node1701 = (inp[5]) ? node1703 : 3'b110;
												assign node1703 = (inp[4]) ? 3'b100 : 3'b110;
									assign node1706 = (inp[1]) ? node1714 : node1707;
										assign node1707 = (inp[8]) ? node1709 : 3'b110;
											assign node1709 = (inp[4]) ? 3'b110 : node1710;
												assign node1710 = (inp[5]) ? 3'b110 : 3'b100;
										assign node1714 = (inp[8]) ? 3'b100 : node1715;
											assign node1715 = (inp[4]) ? node1719 : node1716;
												assign node1716 = (inp[5]) ? 3'b100 : 3'b110;
												assign node1719 = (inp[5]) ? 3'b110 : 3'b100;
					assign node1723 = (inp[1]) ? node1851 : node1724;
						assign node1724 = (inp[7]) ? node1792 : node1725;
							assign node1725 = (inp[5]) ? node1761 : node1726;
								assign node1726 = (inp[8]) ? node1744 : node1727;
									assign node1727 = (inp[4]) ? node1739 : node1728;
										assign node1728 = (inp[9]) ? node1734 : node1729;
											assign node1729 = (inp[0]) ? node1731 : 3'b101;
												assign node1731 = (inp[2]) ? 3'b100 : 3'b101;
											assign node1734 = (inp[0]) ? node1736 : 3'b100;
												assign node1736 = (inp[2]) ? 3'b101 : 3'b100;
										assign node1739 = (inp[2]) ? node1741 : 3'b111;
											assign node1741 = (inp[9]) ? 3'b111 : 3'b110;
									assign node1744 = (inp[4]) ? node1752 : node1745;
										assign node1745 = (inp[9]) ? node1747 : 3'b110;
											assign node1747 = (inp[0]) ? 3'b111 : node1748;
												assign node1748 = (inp[2]) ? 3'b111 : 3'b110;
										assign node1752 = (inp[2]) ? 3'b100 : node1753;
											assign node1753 = (inp[0]) ? node1757 : node1754;
												assign node1754 = (inp[9]) ? 3'b100 : 3'b101;
												assign node1757 = (inp[9]) ? 3'b101 : 3'b100;
								assign node1761 = (inp[9]) ? node1781 : node1762;
									assign node1762 = (inp[0]) ? node1774 : node1763;
										assign node1763 = (inp[2]) ? node1769 : node1764;
											assign node1764 = (inp[8]) ? node1766 : 3'b111;
												assign node1766 = (inp[4]) ? 3'b101 : 3'b111;
											assign node1769 = (inp[4]) ? node1771 : 3'b101;
												assign node1771 = (inp[8]) ? 3'b100 : 3'b110;
										assign node1774 = (inp[8]) ? node1778 : node1775;
											assign node1775 = (inp[4]) ? 3'b110 : 3'b100;
											assign node1778 = (inp[4]) ? 3'b100 : 3'b110;
									assign node1781 = (inp[4]) ? node1789 : node1782;
										assign node1782 = (inp[8]) ? node1784 : 3'b100;
											assign node1784 = (inp[0]) ? 3'b111 : node1785;
												assign node1785 = (inp[2]) ? 3'b111 : 3'b110;
										assign node1789 = (inp[8]) ? 3'b101 : 3'b111;
							assign node1792 = (inp[9]) ? node1828 : node1793;
								assign node1793 = (inp[0]) ? node1813 : node1794;
									assign node1794 = (inp[2]) ? node1808 : node1795;
										assign node1795 = (inp[5]) ? node1803 : node1796;
											assign node1796 = (inp[8]) ? node1800 : node1797;
												assign node1797 = (inp[4]) ? 3'b110 : 3'b100;
												assign node1800 = (inp[4]) ? 3'b100 : 3'b110;
											assign node1803 = (inp[8]) ? node1805 : 3'b100;
												assign node1805 = (inp[4]) ? 3'b100 : 3'b110;
										assign node1808 = (inp[8]) ? node1810 : 3'b100;
											assign node1810 = (inp[4]) ? 3'b101 : 3'b111;
									assign node1813 = (inp[5]) ? node1821 : node1814;
										assign node1814 = (inp[8]) ? node1818 : node1815;
											assign node1815 = (inp[4]) ? 3'b111 : 3'b100;
											assign node1818 = (inp[4]) ? 3'b101 : 3'b111;
										assign node1821 = (inp[4]) ? node1825 : node1822;
											assign node1822 = (inp[2]) ? 3'b101 : 3'b100;
											assign node1825 = (inp[8]) ? 3'b101 : 3'b111;
								assign node1828 = (inp[2]) ? node1842 : node1829;
									assign node1829 = (inp[0]) ? node1835 : node1830;
										assign node1830 = (inp[4]) ? node1832 : 3'b101;
											assign node1832 = (inp[8]) ? 3'b101 : 3'b111;
										assign node1835 = (inp[4]) ? node1839 : node1836;
											assign node1836 = (inp[8]) ? 3'b110 : 3'b101;
											assign node1839 = (inp[8]) ? 3'b100 : 3'b110;
									assign node1842 = (inp[4]) ? node1848 : node1843;
										assign node1843 = (inp[8]) ? 3'b110 : node1844;
											assign node1844 = (inp[0]) ? 3'b100 : 3'b101;
										assign node1848 = (inp[8]) ? 3'b100 : 3'b110;
						assign node1851 = (inp[9]) ? node1907 : node1852;
							assign node1852 = (inp[7]) ? node1876 : node1853;
								assign node1853 = (inp[2]) ? node1869 : node1854;
									assign node1854 = (inp[0]) ? node1862 : node1855;
										assign node1855 = (inp[8]) ? node1859 : node1856;
											assign node1856 = (inp[4]) ? 3'b111 : 3'b101;
											assign node1859 = (inp[4]) ? 3'b101 : 3'b111;
										assign node1862 = (inp[4]) ? node1866 : node1863;
											assign node1863 = (inp[8]) ? 3'b110 : 3'b101;
											assign node1866 = (inp[8]) ? 3'b100 : 3'b110;
									assign node1869 = (inp[8]) ? node1873 : node1870;
										assign node1870 = (inp[4]) ? 3'b110 : 3'b100;
										assign node1873 = (inp[4]) ? 3'b100 : 3'b110;
								assign node1876 = (inp[0]) ? node1890 : node1877;
									assign node1877 = (inp[2]) ? node1885 : node1878;
										assign node1878 = (inp[4]) ? node1882 : node1879;
											assign node1879 = (inp[8]) ? 3'b110 : 3'b100;
											assign node1882 = (inp[8]) ? 3'b100 : 3'b110;
										assign node1885 = (inp[8]) ? node1887 : 3'b100;
											assign node1887 = (inp[4]) ? 3'b101 : 3'b111;
									assign node1890 = (inp[2]) ? node1898 : node1891;
										assign node1891 = (inp[4]) ? node1895 : node1892;
											assign node1892 = (inp[8]) ? 3'b111 : 3'b100;
											assign node1895 = (inp[8]) ? 3'b101 : 3'b111;
										assign node1898 = (inp[5]) ? 3'b101 : node1899;
											assign node1899 = (inp[8]) ? node1903 : node1900;
												assign node1900 = (inp[4]) ? 3'b111 : 3'b101;
												assign node1903 = (inp[4]) ? 3'b101 : 3'b111;
							assign node1907 = (inp[7]) ? node1949 : node1908;
								assign node1908 = (inp[0]) ? node1926 : node1909;
									assign node1909 = (inp[2]) ? node1919 : node1910;
										assign node1910 = (inp[5]) ? node1912 : 3'b100;
											assign node1912 = (inp[4]) ? node1916 : node1913;
												assign node1913 = (inp[8]) ? 3'b110 : 3'b100;
												assign node1916 = (inp[8]) ? 3'b100 : 3'b110;
										assign node1919 = (inp[4]) ? node1923 : node1920;
											assign node1920 = (inp[8]) ? 3'b111 : 3'b100;
											assign node1923 = (inp[8]) ? 3'b101 : 3'b111;
									assign node1926 = (inp[5]) ? node1940 : node1927;
										assign node1927 = (inp[2]) ? node1933 : node1928;
											assign node1928 = (inp[8]) ? node1930 : 3'b111;
												assign node1930 = (inp[4]) ? 3'b101 : 3'b111;
											assign node1933 = (inp[8]) ? node1937 : node1934;
												assign node1934 = (inp[4]) ? 3'b111 : 3'b101;
												assign node1937 = (inp[4]) ? 3'b101 : 3'b111;
										assign node1940 = (inp[2]) ? 3'b101 : node1941;
											assign node1941 = (inp[4]) ? node1945 : node1942;
												assign node1942 = (inp[8]) ? 3'b111 : 3'b100;
												assign node1945 = (inp[8]) ? 3'b101 : 3'b111;
								assign node1949 = (inp[2]) ? node1963 : node1950;
									assign node1950 = (inp[0]) ? node1958 : node1951;
										assign node1951 = (inp[8]) ? node1955 : node1952;
											assign node1952 = (inp[4]) ? 3'b111 : 3'b101;
											assign node1955 = (inp[4]) ? 3'b101 : 3'b111;
										assign node1958 = (inp[4]) ? node1960 : 3'b101;
											assign node1960 = (inp[8]) ? 3'b100 : 3'b110;
									assign node1963 = (inp[4]) ? node1967 : node1964;
										assign node1964 = (inp[8]) ? 3'b110 : 3'b100;
										assign node1967 = (inp[8]) ? 3'b100 : 3'b110;
		assign node1970 = (inp[6]) ? node2880 : node1971;
			assign node1971 = (inp[1]) ? node2435 : node1972;
				assign node1972 = (inp[11]) ? node2202 : node1973;
					assign node1973 = (inp[3]) ? node2075 : node1974;
						assign node1974 = (inp[4]) ? node2032 : node1975;
							assign node1975 = (inp[8]) ? node2013 : node1976;
								assign node1976 = (inp[0]) ? node1996 : node1977;
									assign node1977 = (inp[2]) ? node1983 : node1978;
										assign node1978 = (inp[5]) ? node1980 : 3'b011;
											assign node1980 = (inp[7]) ? 3'b010 : 3'b011;
										assign node1983 = (inp[5]) ? node1989 : node1984;
											assign node1984 = (inp[9]) ? 3'b010 : node1985;
												assign node1985 = (inp[7]) ? 3'b010 : 3'b011;
											assign node1989 = (inp[9]) ? node1993 : node1990;
												assign node1990 = (inp[7]) ? 3'b010 : 3'b011;
												assign node1993 = (inp[7]) ? 3'b011 : 3'b010;
									assign node1996 = (inp[2]) ? node1998 : 3'b010;
										assign node1998 = (inp[5]) ? node2006 : node1999;
											assign node1999 = (inp[7]) ? node2003 : node2000;
												assign node2000 = (inp[9]) ? 3'b011 : 3'b010;
												assign node2003 = (inp[9]) ? 3'b010 : 3'b011;
											assign node2006 = (inp[7]) ? node2010 : node2007;
												assign node2007 = (inp[9]) ? 3'b011 : 3'b010;
												assign node2010 = (inp[9]) ? 3'b010 : 3'b011;
								assign node2013 = (inp[7]) ? node2023 : node2014;
									assign node2014 = (inp[9]) ? node2018 : node2015;
										assign node2015 = (inp[0]) ? 3'b000 : 3'b001;
										assign node2018 = (inp[0]) ? node2020 : 3'b000;
											assign node2020 = (inp[2]) ? 3'b001 : 3'b000;
									assign node2023 = (inp[9]) ? node2029 : node2024;
										assign node2024 = (inp[0]) ? node2026 : 3'b000;
											assign node2026 = (inp[2]) ? 3'b001 : 3'b000;
										assign node2029 = (inp[2]) ? 3'b000 : 3'b001;
							assign node2032 = (inp[8]) ? node2056 : node2033;
								assign node2033 = (inp[9]) ? node2045 : node2034;
									assign node2034 = (inp[7]) ? node2040 : node2035;
										assign node2035 = (inp[0]) ? node2037 : 3'b001;
											assign node2037 = (inp[2]) ? 3'b000 : 3'b001;
										assign node2040 = (inp[0]) ? node2042 : 3'b000;
											assign node2042 = (inp[2]) ? 3'b001 : 3'b000;
									assign node2045 = (inp[7]) ? node2051 : node2046;
										assign node2046 = (inp[2]) ? node2048 : 3'b000;
											assign node2048 = (inp[0]) ? 3'b001 : 3'b000;
										assign node2051 = (inp[0]) ? node2053 : 3'b001;
											assign node2053 = (inp[2]) ? 3'b000 : 3'b001;
								assign node2056 = (inp[5]) ? node2070 : node2057;
									assign node2057 = (inp[7]) ? node2063 : node2058;
										assign node2058 = (inp[9]) ? node2060 : 3'b010;
											assign node2060 = (inp[2]) ? 3'b011 : 3'b010;
										assign node2063 = (inp[9]) ? node2065 : 3'b011;
											assign node2065 = (inp[2]) ? 3'b010 : node2066;
												assign node2066 = (inp[0]) ? 3'b010 : 3'b011;
									assign node2070 = (inp[9]) ? node2072 : 3'b011;
										assign node2072 = (inp[7]) ? 3'b011 : 3'b010;
						assign node2075 = (inp[8]) ? node2127 : node2076;
							assign node2076 = (inp[9]) ? node2108 : node2077;
								assign node2077 = (inp[5]) ? node2095 : node2078;
									assign node2078 = (inp[4]) ? node2088 : node2079;
										assign node2079 = (inp[7]) ? node2083 : node2080;
											assign node2080 = (inp[0]) ? 3'b010 : 3'b011;
											assign node2083 = (inp[0]) ? node2085 : 3'b010;
												assign node2085 = (inp[2]) ? 3'b011 : 3'b010;
										assign node2088 = (inp[7]) ? 3'b000 : node2089;
											assign node2089 = (inp[0]) ? node2091 : 3'b001;
												assign node2091 = (inp[2]) ? 3'b000 : 3'b001;
									assign node2095 = (inp[4]) ? node2101 : node2096;
										assign node2096 = (inp[7]) ? node2098 : 3'b001;
											assign node2098 = (inp[0]) ? 3'b001 : 3'b000;
										assign node2101 = (inp[7]) ? node2103 : 3'b010;
											assign node2103 = (inp[0]) ? 3'b011 : node2104;
												assign node2104 = (inp[2]) ? 3'b011 : 3'b010;
								assign node2108 = (inp[2]) ? node2120 : node2109;
									assign node2109 = (inp[7]) ? node2115 : node2110;
										assign node2110 = (inp[4]) ? node2112 : 3'b000;
											assign node2112 = (inp[0]) ? 3'b011 : 3'b010;
										assign node2115 = (inp[5]) ? 3'b001 : node2116;
											assign node2116 = (inp[4]) ? 3'b001 : 3'b011;
									assign node2120 = (inp[7]) ? 3'b010 : node2121;
										assign node2121 = (inp[4]) ? node2123 : 3'b010;
											assign node2123 = (inp[5]) ? 3'b011 : 3'b001;
							assign node2127 = (inp[4]) ? node2163 : node2128;
								assign node2128 = (inp[5]) ? node2146 : node2129;
									assign node2129 = (inp[9]) ? node2137 : node2130;
										assign node2130 = (inp[7]) ? node2134 : node2131;
											assign node2131 = (inp[0]) ? 3'b000 : 3'b001;
											assign node2134 = (inp[0]) ? 3'b001 : 3'b000;
										assign node2137 = (inp[0]) ? node2139 : 3'b000;
											assign node2139 = (inp[2]) ? node2143 : node2140;
												assign node2140 = (inp[7]) ? 3'b001 : 3'b000;
												assign node2143 = (inp[7]) ? 3'b000 : 3'b001;
									assign node2146 = (inp[9]) ? node2154 : node2147;
										assign node2147 = (inp[0]) ? 3'b011 : node2148;
											assign node2148 = (inp[2]) ? 3'b010 : node2149;
												assign node2149 = (inp[7]) ? 3'b010 : 3'b011;
										assign node2154 = (inp[0]) ? 3'b010 : node2155;
											assign node2155 = (inp[7]) ? node2159 : node2156;
												assign node2156 = (inp[2]) ? 3'b011 : 3'b010;
												assign node2159 = (inp[2]) ? 3'b010 : 3'b011;
								assign node2163 = (inp[5]) ? node2183 : node2164;
									assign node2164 = (inp[2]) ? node2176 : node2165;
										assign node2165 = (inp[0]) ? node2171 : node2166;
											assign node2166 = (inp[7]) ? node2168 : 3'b011;
												assign node2168 = (inp[9]) ? 3'b011 : 3'b010;
											assign node2171 = (inp[7]) ? node2173 : 3'b010;
												assign node2173 = (inp[9]) ? 3'b010 : 3'b011;
										assign node2176 = (inp[0]) ? 3'b011 : node2177;
											assign node2177 = (inp[9]) ? node2179 : 3'b011;
												assign node2179 = (inp[7]) ? 3'b010 : 3'b011;
									assign node2183 = (inp[2]) ? node2193 : node2184;
										assign node2184 = (inp[0]) ? 3'b001 : node2185;
											assign node2185 = (inp[7]) ? node2189 : node2186;
												assign node2186 = (inp[9]) ? 3'b000 : 3'b001;
												assign node2189 = (inp[9]) ? 3'b001 : 3'b000;
										assign node2193 = (inp[0]) ? 3'b000 : node2194;
											assign node2194 = (inp[7]) ? node2198 : node2195;
												assign node2195 = (inp[9]) ? 3'b001 : 3'b000;
												assign node2198 = (inp[9]) ? 3'b000 : 3'b001;
					assign node2202 = (inp[8]) ? node2322 : node2203;
						assign node2203 = (inp[4]) ? node2271 : node2204;
							assign node2204 = (inp[3]) ? node2238 : node2205;
								assign node2205 = (inp[5]) ? node2225 : node2206;
									assign node2206 = (inp[0]) ? node2220 : node2207;
										assign node2207 = (inp[2]) ? node2213 : node2208;
											assign node2208 = (inp[7]) ? node2210 : 3'b110;
												assign node2210 = (inp[9]) ? 3'b111 : 3'b110;
											assign node2213 = (inp[9]) ? node2217 : node2214;
												assign node2214 = (inp[7]) ? 3'b110 : 3'b111;
												assign node2217 = (inp[7]) ? 3'b111 : 3'b110;
										assign node2220 = (inp[7]) ? node2222 : 3'b111;
											assign node2222 = (inp[9]) ? 3'b110 : 3'b111;
									assign node2225 = (inp[9]) ? node2231 : node2226;
										assign node2226 = (inp[7]) ? 3'b100 : node2227;
											assign node2227 = (inp[0]) ? 3'b100 : 3'b101;
										assign node2231 = (inp[2]) ? node2233 : 3'b101;
											assign node2233 = (inp[7]) ? node2235 : 3'b100;
												assign node2235 = (inp[0]) ? 3'b100 : 3'b101;
								assign node2238 = (inp[5]) ? node2256 : node2239;
									assign node2239 = (inp[9]) ? node2249 : node2240;
										assign node2240 = (inp[7]) ? node2244 : node2241;
											assign node2241 = (inp[0]) ? 3'b100 : 3'b101;
											assign node2244 = (inp[2]) ? node2246 : 3'b100;
												assign node2246 = (inp[0]) ? 3'b101 : 3'b100;
										assign node2249 = (inp[7]) ? node2253 : node2250;
											assign node2250 = (inp[2]) ? 3'b101 : 3'b100;
											assign node2253 = (inp[2]) ? 3'b100 : 3'b101;
									assign node2256 = (inp[7]) ? node2266 : node2257;
										assign node2257 = (inp[0]) ? node2261 : node2258;
											assign node2258 = (inp[2]) ? 3'b101 : 3'b100;
											assign node2261 = (inp[2]) ? node2263 : 3'b101;
												assign node2263 = (inp[9]) ? 3'b101 : 3'b100;
										assign node2266 = (inp[9]) ? 3'b101 : node2267;
											assign node2267 = (inp[0]) ? 3'b101 : 3'b100;
							assign node2271 = (inp[5]) ? node2297 : node2272;
								assign node2272 = (inp[3]) ? node2286 : node2273;
									assign node2273 = (inp[0]) ? node2279 : node2274;
										assign node2274 = (inp[9]) ? node2276 : 3'b100;
											assign node2276 = (inp[7]) ? 3'b101 : 3'b100;
										assign node2279 = (inp[2]) ? 3'b101 : node2280;
											assign node2280 = (inp[7]) ? 3'b101 : node2281;
												assign node2281 = (inp[9]) ? 3'b100 : 3'b101;
									assign node2286 = (inp[0]) ? node2292 : node2287;
										assign node2287 = (inp[9]) ? 3'b111 : node2288;
											assign node2288 = (inp[7]) ? 3'b111 : 3'b110;
										assign node2292 = (inp[9]) ? node2294 : 3'b110;
											assign node2294 = (inp[7]) ? 3'b110 : 3'b111;
								assign node2297 = (inp[3]) ? node2313 : node2298;
									assign node2298 = (inp[7]) ? node2308 : node2299;
										assign node2299 = (inp[9]) ? node2305 : node2300;
											assign node2300 = (inp[0]) ? 3'b110 : node2301;
												assign node2301 = (inp[2]) ? 3'b110 : 3'b111;
											assign node2305 = (inp[0]) ? 3'b111 : 3'b110;
										assign node2308 = (inp[2]) ? node2310 : 3'b110;
											assign node2310 = (inp[0]) ? 3'b110 : 3'b111;
									assign node2313 = (inp[9]) ? node2319 : node2314;
										assign node2314 = (inp[7]) ? 3'b111 : node2315;
											assign node2315 = (inp[2]) ? 3'b110 : 3'b111;
										assign node2319 = (inp[7]) ? 3'b110 : 3'b111;
						assign node2322 = (inp[4]) ? node2370 : node2323;
							assign node2323 = (inp[3]) ? node2347 : node2324;
								assign node2324 = (inp[5]) ? node2340 : node2325;
									assign node2325 = (inp[2]) ? node2331 : node2326;
										assign node2326 = (inp[0]) ? node2328 : 3'b101;
											assign node2328 = (inp[9]) ? 3'b101 : 3'b100;
										assign node2331 = (inp[9]) ? 3'b100 : node2332;
											assign node2332 = (inp[0]) ? node2336 : node2333;
												assign node2333 = (inp[7]) ? 3'b100 : 3'b101;
												assign node2336 = (inp[7]) ? 3'b101 : 3'b100;
									assign node2340 = (inp[9]) ? 3'b110 : node2341;
										assign node2341 = (inp[0]) ? 3'b111 : node2342;
											assign node2342 = (inp[7]) ? 3'b110 : 3'b111;
								assign node2347 = (inp[9]) ? node2359 : node2348;
									assign node2348 = (inp[7]) ? node2354 : node2349;
										assign node2349 = (inp[0]) ? 3'b110 : node2350;
											assign node2350 = (inp[2]) ? 3'b110 : 3'b111;
										assign node2354 = (inp[0]) ? 3'b111 : node2355;
											assign node2355 = (inp[2]) ? 3'b111 : 3'b110;
									assign node2359 = (inp[7]) ? node2365 : node2360;
										assign node2360 = (inp[2]) ? 3'b111 : node2361;
											assign node2361 = (inp[0]) ? 3'b111 : 3'b110;
										assign node2365 = (inp[2]) ? 3'b110 : node2366;
											assign node2366 = (inp[0]) ? 3'b110 : 3'b111;
							assign node2370 = (inp[3]) ? node2402 : node2371;
								assign node2371 = (inp[5]) ? node2391 : node2372;
									assign node2372 = (inp[0]) ? node2378 : node2373;
										assign node2373 = (inp[9]) ? node2375 : 3'b111;
											assign node2375 = (inp[7]) ? 3'b110 : 3'b111;
										assign node2378 = (inp[2]) ? node2384 : node2379;
											assign node2379 = (inp[7]) ? 3'b110 : node2380;
												assign node2380 = (inp[9]) ? 3'b111 : 3'b110;
											assign node2384 = (inp[9]) ? node2388 : node2385;
												assign node2385 = (inp[7]) ? 3'b111 : 3'b110;
												assign node2388 = (inp[7]) ? 3'b110 : 3'b111;
									assign node2391 = (inp[0]) ? node2397 : node2392;
										assign node2392 = (inp[9]) ? node2394 : 3'b100;
											assign node2394 = (inp[7]) ? 3'b101 : 3'b100;
										assign node2397 = (inp[9]) ? node2399 : 3'b101;
											assign node2399 = (inp[7]) ? 3'b100 : 3'b101;
								assign node2402 = (inp[2]) ? node2414 : node2403;
									assign node2403 = (inp[5]) ? node2405 : 3'b100;
										assign node2405 = (inp[9]) ? 3'b100 : node2406;
											assign node2406 = (inp[0]) ? node2410 : node2407;
												assign node2407 = (inp[7]) ? 3'b100 : 3'b101;
												assign node2410 = (inp[7]) ? 3'b101 : 3'b100;
									assign node2414 = (inp[5]) ? node2424 : node2415;
										assign node2415 = (inp[0]) ? 3'b101 : node2416;
											assign node2416 = (inp[7]) ? node2420 : node2417;
												assign node2417 = (inp[9]) ? 3'b101 : 3'b100;
												assign node2420 = (inp[9]) ? 3'b100 : 3'b101;
										assign node2424 = (inp[0]) ? node2430 : node2425;
											assign node2425 = (inp[9]) ? 3'b100 : node2426;
												assign node2426 = (inp[7]) ? 3'b101 : 3'b100;
											assign node2430 = (inp[9]) ? node2432 : 3'b100;
												assign node2432 = (inp[7]) ? 3'b100 : 3'b101;
				assign node2435 = (inp[5]) ? node2655 : node2436;
					assign node2436 = (inp[8]) ? node2558 : node2437;
						assign node2437 = (inp[4]) ? node2489 : node2438;
							assign node2438 = (inp[3]) ? node2468 : node2439;
								assign node2439 = (inp[0]) ? node2455 : node2440;
									assign node2440 = (inp[2]) ? node2448 : node2441;
										assign node2441 = (inp[7]) ? node2445 : node2442;
											assign node2442 = (inp[9]) ? 3'b110 : 3'b111;
											assign node2445 = (inp[9]) ? 3'b111 : 3'b110;
										assign node2448 = (inp[7]) ? node2452 : node2449;
											assign node2449 = (inp[9]) ? 3'b110 : 3'b111;
											assign node2452 = (inp[9]) ? 3'b111 : 3'b110;
									assign node2455 = (inp[9]) ? node2463 : node2456;
										assign node2456 = (inp[2]) ? node2460 : node2457;
											assign node2457 = (inp[7]) ? 3'b110 : 3'b111;
											assign node2460 = (inp[7]) ? 3'b111 : 3'b110;
										assign node2463 = (inp[2]) ? node2465 : 3'b111;
											assign node2465 = (inp[7]) ? 3'b110 : 3'b111;
								assign node2468 = (inp[7]) ? node2478 : node2469;
									assign node2469 = (inp[9]) ? node2473 : node2470;
										assign node2470 = (inp[2]) ? 3'b100 : 3'b101;
										assign node2473 = (inp[2]) ? node2475 : 3'b100;
											assign node2475 = (inp[0]) ? 3'b101 : 3'b100;
									assign node2478 = (inp[9]) ? node2484 : node2479;
										assign node2479 = (inp[2]) ? node2481 : 3'b100;
											assign node2481 = (inp[11]) ? 3'b100 : 3'b101;
										assign node2484 = (inp[0]) ? node2486 : 3'b101;
											assign node2486 = (inp[2]) ? 3'b100 : 3'b101;
							assign node2489 = (inp[3]) ? node2523 : node2490;
								assign node2490 = (inp[0]) ? node2504 : node2491;
									assign node2491 = (inp[11]) ? node2499 : node2492;
										assign node2492 = (inp[7]) ? node2496 : node2493;
											assign node2493 = (inp[9]) ? 3'b100 : 3'b101;
											assign node2496 = (inp[9]) ? 3'b101 : 3'b100;
										assign node2499 = (inp[9]) ? 3'b101 : node2500;
											assign node2500 = (inp[7]) ? 3'b100 : 3'b101;
									assign node2504 = (inp[11]) ? node2516 : node2505;
										assign node2505 = (inp[9]) ? node2511 : node2506;
											assign node2506 = (inp[7]) ? 3'b101 : node2507;
												assign node2507 = (inp[2]) ? 3'b100 : 3'b101;
											assign node2511 = (inp[7]) ? 3'b100 : node2512;
												assign node2512 = (inp[2]) ? 3'b101 : 3'b100;
										assign node2516 = (inp[2]) ? 3'b100 : node2517;
											assign node2517 = (inp[9]) ? node2519 : 3'b100;
												assign node2519 = (inp[7]) ? 3'b101 : 3'b100;
								assign node2523 = (inp[11]) ? node2543 : node2524;
									assign node2524 = (inp[0]) ? node2536 : node2525;
										assign node2525 = (inp[2]) ? node2531 : node2526;
											assign node2526 = (inp[7]) ? node2528 : 3'b111;
												assign node2528 = (inp[9]) ? 3'b111 : 3'b110;
											assign node2531 = (inp[9]) ? 3'b110 : node2532;
												assign node2532 = (inp[7]) ? 3'b111 : 3'b110;
										assign node2536 = (inp[2]) ? node2538 : 3'b110;
											assign node2538 = (inp[9]) ? node2540 : 3'b110;
												assign node2540 = (inp[7]) ? 3'b110 : 3'b111;
									assign node2543 = (inp[2]) ? node2551 : node2544;
										assign node2544 = (inp[9]) ? 3'b111 : node2545;
											assign node2545 = (inp[0]) ? 3'b111 : node2546;
												assign node2546 = (inp[7]) ? 3'b110 : 3'b111;
										assign node2551 = (inp[9]) ? node2555 : node2552;
											assign node2552 = (inp[7]) ? 3'b111 : 3'b110;
											assign node2555 = (inp[7]) ? 3'b110 : 3'b111;
						assign node2558 = (inp[9]) ? node2618 : node2559;
							assign node2559 = (inp[7]) ? node2593 : node2560;
								assign node2560 = (inp[0]) ? node2576 : node2561;
									assign node2561 = (inp[2]) ? node2569 : node2562;
										assign node2562 = (inp[3]) ? node2566 : node2563;
											assign node2563 = (inp[4]) ? 3'b111 : 3'b101;
											assign node2566 = (inp[4]) ? 3'b101 : 3'b111;
										assign node2569 = (inp[4]) ? node2573 : node2570;
											assign node2570 = (inp[3]) ? 3'b110 : 3'b101;
											assign node2573 = (inp[3]) ? 3'b100 : 3'b110;
									assign node2576 = (inp[11]) ? node2584 : node2577;
										assign node2577 = (inp[4]) ? node2581 : node2578;
											assign node2578 = (inp[3]) ? 3'b110 : 3'b100;
											assign node2581 = (inp[3]) ? 3'b100 : 3'b110;
										assign node2584 = (inp[3]) ? node2590 : node2585;
											assign node2585 = (inp[4]) ? 3'b110 : node2586;
												assign node2586 = (inp[2]) ? 3'b100 : 3'b101;
											assign node2590 = (inp[4]) ? 3'b100 : 3'b110;
								assign node2593 = (inp[2]) ? node2609 : node2594;
									assign node2594 = (inp[0]) ? node2604 : node2595;
										assign node2595 = (inp[11]) ? 3'b100 : node2596;
											assign node2596 = (inp[4]) ? node2600 : node2597;
												assign node2597 = (inp[3]) ? 3'b110 : 3'b100;
												assign node2600 = (inp[3]) ? 3'b100 : 3'b110;
										assign node2604 = (inp[3]) ? 3'b111 : node2605;
											assign node2605 = (inp[4]) ? 3'b111 : 3'b100;
									assign node2609 = (inp[4]) ? node2615 : node2610;
										assign node2610 = (inp[3]) ? 3'b111 : node2611;
											assign node2611 = (inp[11]) ? 3'b100 : 3'b101;
										assign node2615 = (inp[3]) ? 3'b101 : 3'b111;
							assign node2618 = (inp[7]) ? node2640 : node2619;
								assign node2619 = (inp[2]) ? node2631 : node2620;
									assign node2620 = (inp[0]) ? node2626 : node2621;
										assign node2621 = (inp[3]) ? node2623 : 3'b100;
											assign node2623 = (inp[4]) ? 3'b100 : 3'b110;
										assign node2626 = (inp[4]) ? 3'b111 : node2627;
											assign node2627 = (inp[3]) ? 3'b111 : 3'b100;
									assign node2631 = (inp[4]) ? node2637 : node2632;
										assign node2632 = (inp[3]) ? 3'b111 : node2633;
											assign node2633 = (inp[11]) ? 3'b100 : 3'b101;
										assign node2637 = (inp[3]) ? 3'b101 : 3'b111;
								assign node2640 = (inp[3]) ? node2648 : node2641;
									assign node2641 = (inp[4]) ? node2643 : 3'b101;
										assign node2643 = (inp[0]) ? 3'b110 : node2644;
											assign node2644 = (inp[2]) ? 3'b110 : 3'b111;
									assign node2648 = (inp[4]) ? 3'b100 : node2649;
										assign node2649 = (inp[2]) ? 3'b110 : node2650;
											assign node2650 = (inp[0]) ? 3'b110 : 3'b111;
					assign node2655 = (inp[11]) ? node2765 : node2656;
						assign node2656 = (inp[9]) ? node2712 : node2657;
							assign node2657 = (inp[7]) ? node2681 : node2658;
								assign node2658 = (inp[0]) ? node2674 : node2659;
									assign node2659 = (inp[2]) ? node2667 : node2660;
										assign node2660 = (inp[4]) ? node2664 : node2661;
											assign node2661 = (inp[8]) ? 3'b111 : 3'b101;
											assign node2664 = (inp[8]) ? 3'b101 : 3'b111;
										assign node2667 = (inp[4]) ? node2671 : node2668;
											assign node2668 = (inp[8]) ? 3'b110 : 3'b101;
											assign node2671 = (inp[8]) ? 3'b100 : 3'b110;
									assign node2674 = (inp[4]) ? node2678 : node2675;
										assign node2675 = (inp[8]) ? 3'b110 : 3'b101;
										assign node2678 = (inp[8]) ? 3'b100 : 3'b110;
								assign node2681 = (inp[0]) ? node2701 : node2682;
									assign node2682 = (inp[2]) ? node2692 : node2683;
										assign node2683 = (inp[3]) ? node2685 : 3'b100;
											assign node2685 = (inp[8]) ? node2689 : node2686;
												assign node2686 = (inp[4]) ? 3'b110 : 3'b100;
												assign node2689 = (inp[4]) ? 3'b100 : 3'b110;
										assign node2692 = (inp[3]) ? 3'b100 : node2693;
											assign node2693 = (inp[8]) ? node2697 : node2694;
												assign node2694 = (inp[4]) ? 3'b111 : 3'b100;
												assign node2697 = (inp[4]) ? 3'b101 : 3'b111;
									assign node2701 = (inp[3]) ? 3'b101 : node2702;
										assign node2702 = (inp[2]) ? node2706 : node2703;
											assign node2703 = (inp[4]) ? 3'b111 : 3'b100;
											assign node2706 = (inp[8]) ? node2708 : 3'b101;
												assign node2708 = (inp[4]) ? 3'b101 : 3'b111;
							assign node2712 = (inp[7]) ? node2740 : node2713;
								assign node2713 = (inp[0]) ? node2725 : node2714;
									assign node2714 = (inp[2]) ? node2720 : node2715;
										assign node2715 = (inp[8]) ? 3'b100 : node2716;
											assign node2716 = (inp[4]) ? 3'b110 : 3'b100;
										assign node2720 = (inp[4]) ? node2722 : 3'b100;
											assign node2722 = (inp[8]) ? 3'b101 : 3'b111;
									assign node2725 = (inp[2]) ? node2733 : node2726;
										assign node2726 = (inp[8]) ? node2730 : node2727;
											assign node2727 = (inp[4]) ? 3'b111 : 3'b100;
											assign node2730 = (inp[4]) ? 3'b101 : 3'b111;
										assign node2733 = (inp[8]) ? node2737 : node2734;
											assign node2734 = (inp[4]) ? 3'b111 : 3'b101;
											assign node2737 = (inp[4]) ? 3'b101 : 3'b111;
								assign node2740 = (inp[0]) ? node2756 : node2741;
									assign node2741 = (inp[2]) ? node2749 : node2742;
										assign node2742 = (inp[4]) ? node2746 : node2743;
											assign node2743 = (inp[8]) ? 3'b111 : 3'b101;
											assign node2746 = (inp[8]) ? 3'b101 : 3'b111;
										assign node2749 = (inp[8]) ? node2753 : node2750;
											assign node2750 = (inp[4]) ? 3'b110 : 3'b101;
											assign node2753 = (inp[4]) ? 3'b100 : 3'b110;
									assign node2756 = (inp[4]) ? node2762 : node2757;
										assign node2757 = (inp[8]) ? 3'b110 : node2758;
											assign node2758 = (inp[2]) ? 3'b100 : 3'b101;
										assign node2762 = (inp[8]) ? 3'b100 : 3'b110;
						assign node2765 = (inp[9]) ? node2817 : node2766;
							assign node2766 = (inp[7]) ? node2794 : node2767;
								assign node2767 = (inp[0]) ? node2785 : node2768;
									assign node2768 = (inp[2]) ? node2778 : node2769;
										assign node2769 = (inp[3]) ? node2773 : node2770;
											assign node2770 = (inp[8]) ? 3'b111 : 3'b101;
											assign node2773 = (inp[4]) ? node2775 : 3'b111;
												assign node2775 = (inp[8]) ? 3'b101 : 3'b111;
										assign node2778 = (inp[8]) ? node2782 : node2779;
											assign node2779 = (inp[4]) ? 3'b110 : 3'b101;
											assign node2782 = (inp[4]) ? 3'b100 : 3'b110;
									assign node2785 = (inp[4]) ? node2791 : node2786;
										assign node2786 = (inp[8]) ? 3'b110 : node2787;
											assign node2787 = (inp[2]) ? 3'b100 : 3'b101;
										assign node2791 = (inp[3]) ? 3'b110 : 3'b100;
								assign node2794 = (inp[0]) ? node2808 : node2795;
									assign node2795 = (inp[2]) ? node2801 : node2796;
										assign node2796 = (inp[4]) ? node2798 : 3'b110;
											assign node2798 = (inp[8]) ? 3'b100 : 3'b110;
										assign node2801 = (inp[8]) ? node2805 : node2802;
											assign node2802 = (inp[4]) ? 3'b111 : 3'b100;
											assign node2805 = (inp[4]) ? 3'b101 : 3'b111;
									assign node2808 = (inp[2]) ? node2810 : 3'b111;
										assign node2810 = (inp[4]) ? node2814 : node2811;
											assign node2811 = (inp[8]) ? 3'b111 : 3'b101;
											assign node2814 = (inp[8]) ? 3'b101 : 3'b111;
							assign node2817 = (inp[3]) ? node2851 : node2818;
								assign node2818 = (inp[7]) ? node2830 : node2819;
									assign node2819 = (inp[8]) ? node2827 : node2820;
										assign node2820 = (inp[4]) ? 3'b111 : node2821;
											assign node2821 = (inp[0]) ? node2823 : 3'b100;
												assign node2823 = (inp[2]) ? 3'b101 : 3'b100;
										assign node2827 = (inp[4]) ? 3'b101 : 3'b111;
									assign node2830 = (inp[0]) ? node2842 : node2831;
										assign node2831 = (inp[2]) ? node2839 : node2832;
											assign node2832 = (inp[8]) ? node2836 : node2833;
												assign node2833 = (inp[4]) ? 3'b111 : 3'b101;
												assign node2836 = (inp[4]) ? 3'b101 : 3'b111;
											assign node2839 = (inp[8]) ? 3'b110 : 3'b101;
										assign node2842 = (inp[2]) ? node2846 : node2843;
											assign node2843 = (inp[4]) ? 3'b100 : 3'b110;
											assign node2846 = (inp[4]) ? node2848 : 3'b100;
												assign node2848 = (inp[8]) ? 3'b100 : 3'b110;
								assign node2851 = (inp[2]) ? node2869 : node2852;
									assign node2852 = (inp[8]) ? node2862 : node2853;
										assign node2853 = (inp[4]) ? node2857 : node2854;
											assign node2854 = (inp[7]) ? 3'b101 : 3'b100;
											assign node2857 = (inp[0]) ? 3'b110 : node2858;
												assign node2858 = (inp[7]) ? 3'b111 : 3'b110;
										assign node2862 = (inp[4]) ? node2864 : 3'b110;
											assign node2864 = (inp[0]) ? node2866 : 3'b101;
												assign node2866 = (inp[7]) ? 3'b100 : 3'b101;
									assign node2869 = (inp[7]) ? node2875 : node2870;
										assign node2870 = (inp[8]) ? node2872 : 3'b100;
											assign node2872 = (inp[4]) ? 3'b101 : 3'b111;
										assign node2875 = (inp[4]) ? 3'b100 : node2876;
											assign node2876 = (inp[8]) ? 3'b110 : 3'b100;
			assign node2880 = (inp[1]) ? node3430 : node2881;
				assign node2881 = (inp[11]) ? node3165 : node2882;
					assign node2882 = (inp[0]) ? node3032 : node2883;
						assign node2883 = (inp[8]) ? node2957 : node2884;
							assign node2884 = (inp[4]) ? node2918 : node2885;
								assign node2885 = (inp[3]) ? node2903 : node2886;
									assign node2886 = (inp[5]) ? node2894 : node2887;
										assign node2887 = (inp[7]) ? node2891 : node2888;
											assign node2888 = (inp[9]) ? 3'b110 : 3'b111;
											assign node2891 = (inp[9]) ? 3'b111 : 3'b110;
										assign node2894 = (inp[2]) ? node2896 : 3'b100;
											assign node2896 = (inp[9]) ? node2900 : node2897;
												assign node2897 = (inp[7]) ? 3'b100 : 3'b101;
												assign node2900 = (inp[7]) ? 3'b101 : 3'b100;
									assign node2903 = (inp[2]) ? node2911 : node2904;
										assign node2904 = (inp[7]) ? node2908 : node2905;
											assign node2905 = (inp[9]) ? 3'b100 : 3'b101;
											assign node2908 = (inp[9]) ? 3'b101 : 3'b100;
										assign node2911 = (inp[7]) ? node2915 : node2912;
											assign node2912 = (inp[9]) ? 3'b100 : 3'b101;
											assign node2915 = (inp[9]) ? 3'b101 : 3'b100;
								assign node2918 = (inp[3]) ? node2938 : node2919;
									assign node2919 = (inp[5]) ? node2929 : node2920;
										assign node2920 = (inp[2]) ? node2922 : 3'b101;
											assign node2922 = (inp[7]) ? node2926 : node2923;
												assign node2923 = (inp[9]) ? 3'b100 : 3'b101;
												assign node2926 = (inp[9]) ? 3'b101 : 3'b100;
										assign node2929 = (inp[9]) ? 3'b110 : node2930;
											assign node2930 = (inp[7]) ? node2934 : node2931;
												assign node2931 = (inp[2]) ? 3'b110 : 3'b111;
												assign node2934 = (inp[2]) ? 3'b111 : 3'b110;
									assign node2938 = (inp[5]) ? node2950 : node2939;
										assign node2939 = (inp[7]) ? node2945 : node2940;
											assign node2940 = (inp[2]) ? 3'b111 : node2941;
												assign node2941 = (inp[9]) ? 3'b110 : 3'b111;
											assign node2945 = (inp[2]) ? 3'b110 : node2946;
												assign node2946 = (inp[9]) ? 3'b111 : 3'b110;
										assign node2950 = (inp[7]) ? 3'b111 : node2951;
											assign node2951 = (inp[2]) ? node2953 : 3'b111;
												assign node2953 = (inp[9]) ? 3'b111 : 3'b110;
							assign node2957 = (inp[4]) ? node2983 : node2958;
								assign node2958 = (inp[3]) ? node2976 : node2959;
									assign node2959 = (inp[5]) ? node2967 : node2960;
										assign node2960 = (inp[9]) ? node2964 : node2961;
											assign node2961 = (inp[7]) ? 3'b100 : 3'b101;
											assign node2964 = (inp[7]) ? 3'b101 : 3'b100;
										assign node2967 = (inp[7]) ? 3'b110 : node2968;
											assign node2968 = (inp[2]) ? node2972 : node2969;
												assign node2969 = (inp[9]) ? 3'b110 : 3'b111;
												assign node2972 = (inp[9]) ? 3'b111 : 3'b110;
									assign node2976 = (inp[2]) ? 3'b110 : node2977;
										assign node2977 = (inp[9]) ? node2979 : 3'b110;
											assign node2979 = (inp[7]) ? 3'b111 : 3'b110;
								assign node2983 = (inp[3]) ? node3011 : node2984;
									assign node2984 = (inp[5]) ? node2998 : node2985;
										assign node2985 = (inp[7]) ? node2993 : node2986;
											assign node2986 = (inp[9]) ? node2990 : node2987;
												assign node2987 = (inp[2]) ? 3'b110 : 3'b111;
												assign node2990 = (inp[2]) ? 3'b111 : 3'b110;
											assign node2993 = (inp[9]) ? node2995 : 3'b110;
												assign node2995 = (inp[2]) ? 3'b110 : 3'b111;
										assign node2998 = (inp[9]) ? node3006 : node2999;
											assign node2999 = (inp[7]) ? node3003 : node3000;
												assign node3000 = (inp[2]) ? 3'b100 : 3'b101;
												assign node3003 = (inp[2]) ? 3'b101 : 3'b100;
											assign node3006 = (inp[7]) ? node3008 : 3'b100;
												assign node3008 = (inp[2]) ? 3'b100 : 3'b101;
									assign node3011 = (inp[7]) ? node3019 : node3012;
										assign node3012 = (inp[9]) ? node3016 : node3013;
											assign node3013 = (inp[2]) ? 3'b100 : 3'b101;
											assign node3016 = (inp[2]) ? 3'b101 : 3'b100;
										assign node3019 = (inp[5]) ? node3027 : node3020;
											assign node3020 = (inp[9]) ? node3024 : node3021;
												assign node3021 = (inp[2]) ? 3'b101 : 3'b100;
												assign node3024 = (inp[2]) ? 3'b100 : 3'b101;
											assign node3027 = (inp[9]) ? node3029 : 3'b101;
												assign node3029 = (inp[2]) ? 3'b100 : 3'b101;
						assign node3032 = (inp[3]) ? node3106 : node3033;
							assign node3033 = (inp[4]) ? node3065 : node3034;
								assign node3034 = (inp[2]) ? node3054 : node3035;
									assign node3035 = (inp[5]) ? node3043 : node3036;
										assign node3036 = (inp[8]) ? 3'b101 : node3037;
											assign node3037 = (inp[7]) ? 3'b111 : node3038;
												assign node3038 = (inp[9]) ? 3'b110 : 3'b111;
										assign node3043 = (inp[8]) ? node3047 : node3044;
											assign node3044 = (inp[7]) ? 3'b100 : 3'b101;
											assign node3047 = (inp[9]) ? node3051 : node3048;
												assign node3048 = (inp[7]) ? 3'b111 : 3'b110;
												assign node3051 = (inp[7]) ? 3'b110 : 3'b111;
									assign node3054 = (inp[8]) ? node3058 : node3055;
										assign node3055 = (inp[5]) ? 3'b101 : 3'b111;
										assign node3058 = (inp[5]) ? 3'b111 : node3059;
											assign node3059 = (inp[7]) ? node3061 : 3'b100;
												assign node3061 = (inp[9]) ? 3'b100 : 3'b101;
								assign node3065 = (inp[2]) ? node3091 : node3066;
									assign node3066 = (inp[7]) ? node3080 : node3067;
										assign node3067 = (inp[9]) ? node3073 : node3068;
											assign node3068 = (inp[8]) ? node3070 : 3'b101;
												assign node3070 = (inp[5]) ? 3'b100 : 3'b110;
											assign node3073 = (inp[8]) ? node3077 : node3074;
												assign node3074 = (inp[5]) ? 3'b111 : 3'b100;
												assign node3077 = (inp[5]) ? 3'b101 : 3'b111;
										assign node3080 = (inp[8]) ? node3088 : node3081;
											assign node3081 = (inp[5]) ? node3085 : node3082;
												assign node3082 = (inp[9]) ? 3'b101 : 3'b100;
												assign node3085 = (inp[9]) ? 3'b110 : 3'b111;
											assign node3088 = (inp[9]) ? 3'b110 : 3'b111;
									assign node3091 = (inp[8]) ? node3101 : node3092;
										assign node3092 = (inp[5]) ? node3094 : 3'b100;
											assign node3094 = (inp[9]) ? node3098 : node3095;
												assign node3095 = (inp[7]) ? 3'b111 : 3'b110;
												assign node3098 = (inp[7]) ? 3'b110 : 3'b111;
										assign node3101 = (inp[7]) ? node3103 : 3'b111;
											assign node3103 = (inp[9]) ? 3'b110 : 3'b111;
							assign node3106 = (inp[2]) ? node3132 : node3107;
								assign node3107 = (inp[7]) ? node3123 : node3108;
									assign node3108 = (inp[9]) ? node3116 : node3109;
										assign node3109 = (inp[4]) ? node3113 : node3110;
											assign node3110 = (inp[8]) ? 3'b110 : 3'b101;
											assign node3113 = (inp[8]) ? 3'b100 : 3'b110;
										assign node3116 = (inp[8]) ? node3120 : node3117;
											assign node3117 = (inp[4]) ? 3'b111 : 3'b100;
											assign node3120 = (inp[4]) ? 3'b101 : 3'b111;
									assign node3123 = (inp[9]) ? node3127 : node3124;
										assign node3124 = (inp[8]) ? 3'b111 : 3'b100;
										assign node3127 = (inp[4]) ? node3129 : 3'b110;
											assign node3129 = (inp[8]) ? 3'b100 : 3'b110;
								assign node3132 = (inp[8]) ? node3148 : node3133;
									assign node3133 = (inp[4]) ? node3141 : node3134;
										assign node3134 = (inp[5]) ? node3136 : 3'b101;
											assign node3136 = (inp[9]) ? 3'b100 : node3137;
												assign node3137 = (inp[7]) ? 3'b101 : 3'b100;
										assign node3141 = (inp[9]) ? node3145 : node3142;
											assign node3142 = (inp[7]) ? 3'b111 : 3'b110;
											assign node3145 = (inp[7]) ? 3'b110 : 3'b111;
									assign node3148 = (inp[4]) ? node3158 : node3149;
										assign node3149 = (inp[5]) ? node3155 : node3150;
											assign node3150 = (inp[7]) ? node3152 : 3'b110;
												assign node3152 = (inp[9]) ? 3'b110 : 3'b111;
											assign node3155 = (inp[9]) ? 3'b111 : 3'b110;
										assign node3158 = (inp[9]) ? node3162 : node3159;
											assign node3159 = (inp[7]) ? 3'b101 : 3'b100;
											assign node3162 = (inp[7]) ? 3'b100 : 3'b101;
					assign node3165 = (inp[2]) ? node3309 : node3166;
						assign node3166 = (inp[8]) ? node3228 : node3167;
							assign node3167 = (inp[4]) ? node3199 : node3168;
								assign node3168 = (inp[5]) ? node3186 : node3169;
									assign node3169 = (inp[3]) ? node3181 : node3170;
										assign node3170 = (inp[0]) ? node3176 : node3171;
											assign node3171 = (inp[7]) ? 3'b011 : node3172;
												assign node3172 = (inp[9]) ? 3'b010 : 3'b011;
											assign node3176 = (inp[9]) ? 3'b010 : node3177;
												assign node3177 = (inp[7]) ? 3'b010 : 3'b011;
										assign node3181 = (inp[9]) ? 3'b000 : node3182;
											assign node3182 = (inp[7]) ? 3'b000 : 3'b001;
									assign node3186 = (inp[0]) ? node3194 : node3187;
										assign node3187 = (inp[7]) ? node3191 : node3188;
											assign node3188 = (inp[9]) ? 3'b000 : 3'b001;
											assign node3191 = (inp[9]) ? 3'b001 : 3'b000;
										assign node3194 = (inp[9]) ? 3'b001 : node3195;
											assign node3195 = (inp[7]) ? 3'b000 : 3'b001;
								assign node3199 = (inp[5]) ? node3215 : node3200;
									assign node3200 = (inp[3]) ? node3206 : node3201;
										assign node3201 = (inp[7]) ? 3'b000 : node3202;
											assign node3202 = (inp[9]) ? 3'b000 : 3'b001;
										assign node3206 = (inp[0]) ? 3'b010 : node3207;
											assign node3207 = (inp[7]) ? node3211 : node3208;
												assign node3208 = (inp[9]) ? 3'b010 : 3'b011;
												assign node3211 = (inp[9]) ? 3'b011 : 3'b010;
									assign node3215 = (inp[9]) ? node3223 : node3216;
										assign node3216 = (inp[7]) ? node3220 : node3217;
											assign node3217 = (inp[0]) ? 3'b010 : 3'b011;
											assign node3220 = (inp[0]) ? 3'b011 : 3'b010;
										assign node3223 = (inp[0]) ? 3'b010 : node3224;
											assign node3224 = (inp[7]) ? 3'b011 : 3'b010;
							assign node3228 = (inp[4]) ? node3266 : node3229;
								assign node3229 = (inp[3]) ? node3247 : node3230;
									assign node3230 = (inp[5]) ? node3238 : node3231;
										assign node3231 = (inp[9]) ? node3235 : node3232;
											assign node3232 = (inp[7]) ? 3'b000 : 3'b001;
											assign node3235 = (inp[7]) ? 3'b001 : 3'b000;
										assign node3238 = (inp[7]) ? node3240 : 3'b011;
											assign node3240 = (inp[9]) ? node3244 : node3241;
												assign node3241 = (inp[0]) ? 3'b011 : 3'b010;
												assign node3244 = (inp[0]) ? 3'b010 : 3'b011;
									assign node3247 = (inp[9]) ? node3261 : node3248;
										assign node3248 = (inp[5]) ? node3254 : node3249;
											assign node3249 = (inp[7]) ? node3251 : 3'b011;
												assign node3251 = (inp[0]) ? 3'b011 : 3'b010;
											assign node3254 = (inp[7]) ? node3258 : node3255;
												assign node3255 = (inp[0]) ? 3'b010 : 3'b011;
												assign node3258 = (inp[0]) ? 3'b011 : 3'b010;
										assign node3261 = (inp[0]) ? 3'b010 : node3262;
											assign node3262 = (inp[7]) ? 3'b011 : 3'b010;
								assign node3266 = (inp[3]) ? node3292 : node3267;
									assign node3267 = (inp[5]) ? node3281 : node3268;
										assign node3268 = (inp[0]) ? node3274 : node3269;
											assign node3269 = (inp[7]) ? 3'b011 : node3270;
												assign node3270 = (inp[9]) ? 3'b010 : 3'b011;
											assign node3274 = (inp[7]) ? node3278 : node3275;
												assign node3275 = (inp[9]) ? 3'b011 : 3'b010;
												assign node3278 = (inp[9]) ? 3'b010 : 3'b011;
										assign node3281 = (inp[9]) ? node3287 : node3282;
											assign node3282 = (inp[0]) ? node3284 : 3'b000;
												assign node3284 = (inp[7]) ? 3'b001 : 3'b000;
											assign node3287 = (inp[0]) ? node3289 : 3'b001;
												assign node3289 = (inp[7]) ? 3'b000 : 3'b001;
									assign node3292 = (inp[7]) ? node3294 : 3'b001;
										assign node3294 = (inp[5]) ? node3302 : node3295;
											assign node3295 = (inp[9]) ? node3299 : node3296;
												assign node3296 = (inp[0]) ? 3'b001 : 3'b000;
												assign node3299 = (inp[0]) ? 3'b000 : 3'b001;
											assign node3302 = (inp[0]) ? node3306 : node3303;
												assign node3303 = (inp[9]) ? 3'b001 : 3'b000;
												assign node3306 = (inp[9]) ? 3'b000 : 3'b001;
						assign node3309 = (inp[5]) ? node3381 : node3310;
							assign node3310 = (inp[0]) ? node3354 : node3311;
								assign node3311 = (inp[7]) ? node3331 : node3312;
									assign node3312 = (inp[3]) ? node3320 : node3313;
										assign node3313 = (inp[9]) ? node3315 : 3'b001;
											assign node3315 = (inp[8]) ? 3'b000 : node3316;
												assign node3316 = (inp[4]) ? 3'b000 : 3'b010;
										assign node3320 = (inp[9]) ? node3326 : node3321;
											assign node3321 = (inp[8]) ? node3323 : 3'b001;
												assign node3323 = (inp[4]) ? 3'b000 : 3'b010;
											assign node3326 = (inp[8]) ? 3'b011 : node3327;
												assign node3327 = (inp[4]) ? 3'b011 : 3'b000;
									assign node3331 = (inp[3]) ? node3339 : node3332;
										assign node3332 = (inp[8]) ? 3'b011 : node3333;
											assign node3333 = (inp[9]) ? 3'b011 : node3334;
												assign node3334 = (inp[4]) ? 3'b000 : 3'b010;
										assign node3339 = (inp[9]) ? node3347 : node3340;
											assign node3340 = (inp[4]) ? node3344 : node3341;
												assign node3341 = (inp[8]) ? 3'b011 : 3'b000;
												assign node3344 = (inp[8]) ? 3'b001 : 3'b011;
											assign node3347 = (inp[8]) ? node3351 : node3348;
												assign node3348 = (inp[4]) ? 3'b010 : 3'b001;
												assign node3351 = (inp[4]) ? 3'b000 : 3'b010;
								assign node3354 = (inp[9]) ? node3364 : node3355;
									assign node3355 = (inp[7]) ? node3361 : node3356;
										assign node3356 = (inp[8]) ? 3'b000 : node3357;
											assign node3357 = (inp[4]) ? 3'b000 : 3'b010;
										assign node3361 = (inp[8]) ? 3'b011 : 3'b001;
									assign node3364 = (inp[7]) ? node3378 : node3365;
										assign node3365 = (inp[8]) ? node3373 : node3366;
											assign node3366 = (inp[3]) ? node3370 : node3367;
												assign node3367 = (inp[4]) ? 3'b001 : 3'b011;
												assign node3370 = (inp[4]) ? 3'b011 : 3'b001;
											assign node3373 = (inp[3]) ? node3375 : 3'b001;
												assign node3375 = (inp[4]) ? 3'b001 : 3'b011;
										assign node3378 = (inp[8]) ? 3'b000 : 3'b010;
							assign node3381 = (inp[4]) ? node3409 : node3382;
								assign node3382 = (inp[8]) ? node3394 : node3383;
									assign node3383 = (inp[3]) ? node3385 : 3'b000;
										assign node3385 = (inp[9]) ? node3387 : 3'b000;
											assign node3387 = (inp[0]) ? node3391 : node3388;
												assign node3388 = (inp[7]) ? 3'b001 : 3'b000;
												assign node3391 = (inp[7]) ? 3'b000 : 3'b001;
									assign node3394 = (inp[0]) ? node3404 : node3395;
										assign node3395 = (inp[3]) ? node3399 : node3396;
											assign node3396 = (inp[7]) ? 3'b011 : 3'b010;
											assign node3399 = (inp[9]) ? node3401 : 3'b010;
												assign node3401 = (inp[7]) ? 3'b010 : 3'b011;
										assign node3404 = (inp[9]) ? node3406 : 3'b010;
											assign node3406 = (inp[7]) ? 3'b010 : 3'b011;
								assign node3409 = (inp[8]) ? node3417 : node3410;
									assign node3410 = (inp[7]) ? node3414 : node3411;
										assign node3411 = (inp[9]) ? 3'b011 : 3'b010;
										assign node3414 = (inp[9]) ? 3'b010 : 3'b011;
									assign node3417 = (inp[3]) ? node3425 : node3418;
										assign node3418 = (inp[9]) ? node3422 : node3419;
											assign node3419 = (inp[7]) ? 3'b001 : 3'b000;
											assign node3422 = (inp[7]) ? 3'b000 : 3'b001;
										assign node3425 = (inp[9]) ? 3'b000 : node3426;
											assign node3426 = (inp[7]) ? 3'b001 : 3'b000;
				assign node3430 = (inp[2]) ? node3642 : node3431;
					assign node3431 = (inp[0]) ? node3545 : node3432;
						assign node3432 = (inp[8]) ? node3478 : node3433;
							assign node3433 = (inp[4]) ? node3457 : node3434;
								assign node3434 = (inp[5]) ? node3448 : node3435;
									assign node3435 = (inp[3]) ? node3443 : node3436;
										assign node3436 = (inp[7]) ? node3440 : node3437;
											assign node3437 = (inp[9]) ? 3'b010 : 3'b011;
											assign node3440 = (inp[9]) ? 3'b011 : 3'b010;
										assign node3443 = (inp[9]) ? node3445 : 3'b001;
											assign node3445 = (inp[7]) ? 3'b001 : 3'b000;
									assign node3448 = (inp[3]) ? 3'b001 : node3449;
										assign node3449 = (inp[9]) ? node3453 : node3450;
											assign node3450 = (inp[7]) ? 3'b000 : 3'b001;
											assign node3453 = (inp[7]) ? 3'b001 : 3'b000;
								assign node3457 = (inp[5]) ? node3471 : node3458;
									assign node3458 = (inp[3]) ? node3466 : node3459;
										assign node3459 = (inp[9]) ? node3463 : node3460;
											assign node3460 = (inp[7]) ? 3'b000 : 3'b001;
											assign node3463 = (inp[7]) ? 3'b001 : 3'b000;
										assign node3466 = (inp[7]) ? node3468 : 3'b011;
											assign node3468 = (inp[9]) ? 3'b011 : 3'b010;
									assign node3471 = (inp[9]) ? node3475 : node3472;
										assign node3472 = (inp[7]) ? 3'b010 : 3'b011;
										assign node3475 = (inp[7]) ? 3'b011 : 3'b010;
							assign node3478 = (inp[4]) ? node3506 : node3479;
								assign node3479 = (inp[3]) ? node3499 : node3480;
									assign node3480 = (inp[5]) ? node3494 : node3481;
										assign node3481 = (inp[11]) ? node3487 : node3482;
											assign node3482 = (inp[7]) ? 3'b000 : node3483;
												assign node3483 = (inp[9]) ? 3'b000 : 3'b001;
											assign node3487 = (inp[9]) ? node3491 : node3488;
												assign node3488 = (inp[7]) ? 3'b000 : 3'b001;
												assign node3491 = (inp[7]) ? 3'b001 : 3'b000;
										assign node3494 = (inp[7]) ? 3'b010 : node3495;
											assign node3495 = (inp[9]) ? 3'b010 : 3'b011;
									assign node3499 = (inp[9]) ? node3503 : node3500;
										assign node3500 = (inp[7]) ? 3'b010 : 3'b011;
										assign node3503 = (inp[7]) ? 3'b011 : 3'b010;
								assign node3506 = (inp[3]) ? node3522 : node3507;
									assign node3507 = (inp[5]) ? node3513 : node3508;
										assign node3508 = (inp[7]) ? 3'b011 : node3509;
											assign node3509 = (inp[9]) ? 3'b010 : 3'b011;
										assign node3513 = (inp[11]) ? node3515 : 3'b001;
											assign node3515 = (inp[7]) ? node3519 : node3516;
												assign node3516 = (inp[9]) ? 3'b000 : 3'b001;
												assign node3519 = (inp[9]) ? 3'b001 : 3'b000;
									assign node3522 = (inp[5]) ? node3530 : node3523;
										assign node3523 = (inp[9]) ? node3527 : node3524;
											assign node3524 = (inp[7]) ? 3'b000 : 3'b001;
											assign node3527 = (inp[7]) ? 3'b001 : 3'b000;
										assign node3530 = (inp[11]) ? node3538 : node3531;
											assign node3531 = (inp[7]) ? node3535 : node3532;
												assign node3532 = (inp[9]) ? 3'b000 : 3'b001;
												assign node3535 = (inp[9]) ? 3'b001 : 3'b000;
											assign node3538 = (inp[9]) ? node3542 : node3539;
												assign node3539 = (inp[7]) ? 3'b000 : 3'b001;
												assign node3542 = (inp[7]) ? 3'b001 : 3'b000;
						assign node3545 = (inp[5]) ? node3611 : node3546;
							assign node3546 = (inp[8]) ? node3584 : node3547;
								assign node3547 = (inp[3]) ? node3561 : node3548;
									assign node3548 = (inp[4]) ? node3554 : node3549;
										assign node3549 = (inp[9]) ? 3'b011 : node3550;
											assign node3550 = (inp[7]) ? 3'b010 : 3'b011;
										assign node3554 = (inp[7]) ? node3558 : node3555;
											assign node3555 = (inp[9]) ? 3'b000 : 3'b001;
											assign node3558 = (inp[9]) ? 3'b001 : 3'b000;
									assign node3561 = (inp[4]) ? node3569 : node3562;
										assign node3562 = (inp[11]) ? node3564 : 3'b001;
											assign node3564 = (inp[7]) ? node3566 : 3'b000;
												assign node3566 = (inp[9]) ? 3'b001 : 3'b000;
										assign node3569 = (inp[11]) ? node3577 : node3570;
											assign node3570 = (inp[7]) ? node3574 : node3571;
												assign node3571 = (inp[9]) ? 3'b011 : 3'b010;
												assign node3574 = (inp[9]) ? 3'b010 : 3'b011;
											assign node3577 = (inp[7]) ? node3581 : node3578;
												assign node3578 = (inp[9]) ? 3'b011 : 3'b010;
												assign node3581 = (inp[9]) ? 3'b010 : 3'b011;
								assign node3584 = (inp[7]) ? node3600 : node3585;
									assign node3585 = (inp[9]) ? node3593 : node3586;
										assign node3586 = (inp[4]) ? node3590 : node3587;
											assign node3587 = (inp[3]) ? 3'b010 : 3'b001;
											assign node3590 = (inp[3]) ? 3'b000 : 3'b010;
										assign node3593 = (inp[3]) ? node3597 : node3594;
											assign node3594 = (inp[4]) ? 3'b011 : 3'b000;
											assign node3597 = (inp[4]) ? 3'b001 : 3'b011;
									assign node3600 = (inp[9]) ? node3606 : node3601;
										assign node3601 = (inp[4]) ? 3'b011 : node3602;
											assign node3602 = (inp[3]) ? 3'b011 : 3'b000;
										assign node3606 = (inp[4]) ? node3608 : 3'b010;
											assign node3608 = (inp[3]) ? 3'b000 : 3'b010;
							assign node3611 = (inp[7]) ? node3627 : node3612;
								assign node3612 = (inp[9]) ? node3620 : node3613;
									assign node3613 = (inp[4]) ? node3617 : node3614;
										assign node3614 = (inp[3]) ? 3'b001 : 3'b010;
										assign node3617 = (inp[8]) ? 3'b000 : 3'b010;
									assign node3620 = (inp[8]) ? node3624 : node3621;
										assign node3621 = (inp[4]) ? 3'b011 : 3'b000;
										assign node3624 = (inp[4]) ? 3'b001 : 3'b011;
								assign node3627 = (inp[9]) ? node3635 : node3628;
									assign node3628 = (inp[8]) ? node3632 : node3629;
										assign node3629 = (inp[4]) ? 3'b011 : 3'b000;
										assign node3632 = (inp[4]) ? 3'b001 : 3'b011;
									assign node3635 = (inp[8]) ? node3639 : node3636;
										assign node3636 = (inp[4]) ? 3'b010 : 3'b001;
										assign node3639 = (inp[4]) ? 3'b000 : 3'b010;
					assign node3642 = (inp[4]) ? node3760 : node3643;
						assign node3643 = (inp[8]) ? node3705 : node3644;
							assign node3644 = (inp[3]) ? node3674 : node3645;
								assign node3645 = (inp[5]) ? node3659 : node3646;
									assign node3646 = (inp[0]) ? node3652 : node3647;
										assign node3647 = (inp[11]) ? node3649 : 3'b010;
											assign node3649 = (inp[7]) ? 3'b011 : 3'b010;
										assign node3652 = (inp[9]) ? node3656 : node3653;
											assign node3653 = (inp[7]) ? 3'b011 : 3'b010;
											assign node3656 = (inp[7]) ? 3'b010 : 3'b011;
									assign node3659 = (inp[11]) ? node3669 : node3660;
										assign node3660 = (inp[0]) ? 3'b000 : node3661;
											assign node3661 = (inp[9]) ? node3665 : node3662;
												assign node3662 = (inp[7]) ? 3'b000 : 3'b001;
												assign node3665 = (inp[7]) ? 3'b001 : 3'b000;
										assign node3669 = (inp[9]) ? 3'b001 : node3670;
											assign node3670 = (inp[0]) ? 3'b001 : 3'b000;
								assign node3674 = (inp[5]) ? node3690 : node3675;
									assign node3675 = (inp[0]) ? node3683 : node3676;
										assign node3676 = (inp[11]) ? 3'b000 : node3677;
											assign node3677 = (inp[7]) ? node3679 : 3'b000;
												assign node3679 = (inp[9]) ? 3'b001 : 3'b000;
										assign node3683 = (inp[7]) ? node3687 : node3684;
											assign node3684 = (inp[9]) ? 3'b001 : 3'b000;
											assign node3687 = (inp[9]) ? 3'b000 : 3'b001;
									assign node3690 = (inp[7]) ? node3698 : node3691;
										assign node3691 = (inp[9]) ? node3695 : node3692;
											assign node3692 = (inp[0]) ? 3'b000 : 3'b001;
											assign node3695 = (inp[0]) ? 3'b001 : 3'b000;
										assign node3698 = (inp[0]) ? node3702 : node3699;
											assign node3699 = (inp[9]) ? 3'b001 : 3'b000;
											assign node3702 = (inp[9]) ? 3'b000 : 3'b001;
							assign node3705 = (inp[5]) ? node3729 : node3706;
								assign node3706 = (inp[3]) ? node3720 : node3707;
									assign node3707 = (inp[0]) ? node3713 : node3708;
										assign node3708 = (inp[7]) ? 3'b000 : node3709;
											assign node3709 = (inp[9]) ? 3'b000 : 3'b001;
										assign node3713 = (inp[9]) ? node3717 : node3714;
											assign node3714 = (inp[7]) ? 3'b001 : 3'b000;
											assign node3717 = (inp[7]) ? 3'b000 : 3'b001;
									assign node3720 = (inp[11]) ? node3726 : node3721;
										assign node3721 = (inp[9]) ? node3723 : 3'b011;
											assign node3723 = (inp[7]) ? 3'b010 : 3'b011;
										assign node3726 = (inp[9]) ? 3'b011 : 3'b010;
								assign node3729 = (inp[3]) ? node3745 : node3730;
									assign node3730 = (inp[0]) ? node3738 : node3731;
										assign node3731 = (inp[9]) ? node3735 : node3732;
											assign node3732 = (inp[7]) ? 3'b011 : 3'b010;
											assign node3735 = (inp[7]) ? 3'b010 : 3'b011;
										assign node3738 = (inp[9]) ? node3742 : node3739;
											assign node3739 = (inp[7]) ? 3'b011 : 3'b010;
											assign node3742 = (inp[7]) ? 3'b010 : 3'b011;
									assign node3745 = (inp[11]) ? node3747 : 3'b010;
										assign node3747 = (inp[0]) ? node3753 : node3748;
											assign node3748 = (inp[7]) ? node3750 : 3'b010;
												assign node3750 = (inp[9]) ? 3'b010 : 3'b011;
											assign node3753 = (inp[9]) ? node3757 : node3754;
												assign node3754 = (inp[7]) ? 3'b011 : 3'b010;
												assign node3757 = (inp[7]) ? 3'b010 : 3'b011;
						assign node3760 = (inp[8]) ? node3820 : node3761;
							assign node3761 = (inp[3]) ? node3783 : node3762;
								assign node3762 = (inp[5]) ? node3770 : node3763;
									assign node3763 = (inp[0]) ? node3765 : 3'b001;
										assign node3765 = (inp[7]) ? node3767 : 3'b000;
											assign node3767 = (inp[9]) ? 3'b000 : 3'b001;
									assign node3770 = (inp[11]) ? node3776 : node3771;
										assign node3771 = (inp[9]) ? 3'b010 : node3772;
											assign node3772 = (inp[7]) ? 3'b011 : 3'b010;
										assign node3776 = (inp[0]) ? 3'b011 : node3777;
											assign node3777 = (inp[7]) ? 3'b010 : node3778;
												assign node3778 = (inp[9]) ? 3'b011 : 3'b010;
								assign node3783 = (inp[11]) ? node3797 : node3784;
									assign node3784 = (inp[5]) ? node3792 : node3785;
										assign node3785 = (inp[7]) ? node3789 : node3786;
											assign node3786 = (inp[9]) ? 3'b011 : 3'b010;
											assign node3789 = (inp[9]) ? 3'b010 : 3'b011;
										assign node3792 = (inp[9]) ? node3794 : 3'b010;
											assign node3794 = (inp[7]) ? 3'b010 : 3'b011;
									assign node3797 = (inp[5]) ? node3811 : node3798;
										assign node3798 = (inp[0]) ? node3806 : node3799;
											assign node3799 = (inp[7]) ? node3803 : node3800;
												assign node3800 = (inp[9]) ? 3'b011 : 3'b010;
												assign node3803 = (inp[9]) ? 3'b010 : 3'b011;
											assign node3806 = (inp[9]) ? node3808 : 3'b010;
												assign node3808 = (inp[7]) ? 3'b010 : 3'b011;
										assign node3811 = (inp[0]) ? node3813 : 3'b011;
											assign node3813 = (inp[9]) ? node3817 : node3814;
												assign node3814 = (inp[7]) ? 3'b011 : 3'b010;
												assign node3817 = (inp[7]) ? 3'b010 : 3'b011;
							assign node3820 = (inp[3]) ? node3836 : node3821;
								assign node3821 = (inp[5]) ? node3829 : node3822;
									assign node3822 = (inp[9]) ? node3826 : node3823;
										assign node3823 = (inp[7]) ? 3'b011 : 3'b010;
										assign node3826 = (inp[7]) ? 3'b010 : 3'b011;
									assign node3829 = (inp[7]) ? node3833 : node3830;
										assign node3830 = (inp[9]) ? 3'b001 : 3'b000;
										assign node3833 = (inp[9]) ? 3'b000 : 3'b001;
								assign node3836 = (inp[7]) ? node3840 : node3837;
									assign node3837 = (inp[9]) ? 3'b001 : 3'b000;
									assign node3840 = (inp[9]) ? 3'b000 : 3'b001;

endmodule