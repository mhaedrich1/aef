module dtc_split25_bm13 (
	input  wire [11-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node5;
	wire [1-1:0] node7;
	wire [1-1:0] node9;
	wire [1-1:0] node10;
	wire [1-1:0] node12;
	wire [1-1:0] node16;
	wire [1-1:0] node17;
	wire [1-1:0] node19;
	wire [1-1:0] node21;
	wire [1-1:0] node22;
	wire [1-1:0] node24;
	wire [1-1:0] node27;
	wire [1-1:0] node28;
	wire [1-1:0] node32;
	wire [1-1:0] node33;
	wire [1-1:0] node35;
	wire [1-1:0] node36;
	wire [1-1:0] node38;
	wire [1-1:0] node42;
	wire [1-1:0] node43;
	wire [1-1:0] node45;
	wire [1-1:0] node46;
	wire [1-1:0] node50;
	wire [1-1:0] node51;
	wire [1-1:0] node52;
	wire [1-1:0] node57;
	wire [1-1:0] node58;
	wire [1-1:0] node59;
	wire [1-1:0] node61;
	wire [1-1:0] node62;
	wire [1-1:0] node64;
	wire [1-1:0] node66;
	wire [1-1:0] node69;
	wire [1-1:0] node72;
	wire [1-1:0] node73;
	wire [1-1:0] node75;
	wire [1-1:0] node76;
	wire [1-1:0] node78;
	wire [1-1:0] node82;
	wire [1-1:0] node83;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node90;
	wire [1-1:0] node91;
	wire [1-1:0] node93;
	wire [1-1:0] node97;
	wire [1-1:0] node98;
	wire [1-1:0] node99;
	wire [1-1:0] node101;
	wire [1-1:0] node104;
	wire [1-1:0] node105;
	wire [1-1:0] node106;
	wire [1-1:0] node108;
	wire [1-1:0] node113;
	wire [1-1:0] node114;
	wire [1-1:0] node115;
	wire [1-1:0] node116;
	wire [1-1:0] node118;
	wire [1-1:0] node124;
	wire [1-1:0] node125;
	wire [1-1:0] node126;
	wire [1-1:0] node127;
	wire [1-1:0] node129;
	wire [1-1:0] node131;
	wire [1-1:0] node132;
	wire [1-1:0] node134;
	wire [1-1:0] node138;
	wire [1-1:0] node139;
	wire [1-1:0] node141;
	wire [1-1:0] node143;
	wire [1-1:0] node146;
	wire [1-1:0] node147;
	wire [1-1:0] node148;
	wire [1-1:0] node150;
	wire [1-1:0] node154;
	wire [1-1:0] node155;
	wire [1-1:0] node159;
	wire [1-1:0] node160;
	wire [1-1:0] node161;
	wire [1-1:0] node163;
	wire [1-1:0] node165;
	wire [1-1:0] node166;
	wire [1-1:0] node170;
	wire [1-1:0] node171;
	wire [1-1:0] node173;
	wire [1-1:0] node174;
	wire [1-1:0] node178;
	wire [1-1:0] node179;
	wire [1-1:0] node180;
	wire [1-1:0] node185;
	wire [1-1:0] node186;
	wire [1-1:0] node187;
	wire [1-1:0] node189;
	wire [1-1:0] node190;
	wire [1-1:0] node196;
	wire [1-1:0] node197;
	wire [1-1:0] node198;
	wire [1-1:0] node200;
	wire [1-1:0] node201;
	wire [1-1:0] node202;
	wire [1-1:0] node204;
	wire [1-1:0] node207;
	wire [1-1:0] node208;
	wire [1-1:0] node212;
	wire [1-1:0] node213;
	wire [1-1:0] node217;
	wire [1-1:0] node218;
	wire [1-1:0] node219;
	wire [1-1:0] node220;
	wire [1-1:0] node222;
	wire [1-1:0] node225;
	wire [1-1:0] node226;
	wire [1-1:0] node230;
	wire [1-1:0] node231;
	wire [1-1:0] node232;
	wire [1-1:0] node238;
	wire [1-1:0] node239;
	wire [1-1:0] node240;
	wire [1-1:0] node241;
	wire [1-1:0] node242;
	wire [1-1:0] node244;

	assign outp = (inp[6]) ? node124 : node1;
		assign node1 = (inp[8]) ? node57 : node2;
			assign node2 = (inp[3]) ? node16 : node3;
				assign node3 = (inp[5]) ? node5 : 1'b1;
					assign node5 = (inp[0]) ? node7 : 1'b1;
						assign node7 = (inp[2]) ? node9 : 1'b1;
							assign node9 = (inp[1]) ? 1'b0 : node10;
								assign node10 = (inp[7]) ? node12 : 1'b1;
									assign node12 = (inp[10]) ? 1'b0 : 1'b1;
				assign node16 = (inp[7]) ? node32 : node17;
					assign node17 = (inp[0]) ? node19 : 1'b1;
						assign node19 = (inp[9]) ? node21 : 1'b1;
							assign node21 = (inp[1]) ? node27 : node22;
								assign node22 = (inp[10]) ? node24 : 1'b1;
									assign node24 = (inp[2]) ? 1'b0 : 1'b1;
								assign node27 = (inp[2]) ? 1'b0 : node28;
									assign node28 = (inp[10]) ? 1'b0 : 1'b1;
					assign node32 = (inp[0]) ? node42 : node33;
						assign node33 = (inp[2]) ? node35 : 1'b1;
							assign node35 = (inp[1]) ? 1'b0 : node36;
								assign node36 = (inp[9]) ? node38 : 1'b1;
									assign node38 = (inp[5]) ? 1'b0 : 1'b1;
						assign node42 = (inp[10]) ? node50 : node43;
							assign node43 = (inp[1]) ? node45 : 1'b1;
								assign node45 = (inp[5]) ? 1'b0 : node46;
									assign node46 = (inp[4]) ? 1'b0 : 1'b1;
							assign node50 = (inp[4]) ? 1'b0 : node51;
								assign node51 = (inp[2]) ? 1'b0 : node52;
									assign node52 = (inp[1]) ? 1'b0 : 1'b0;
			assign node57 = (inp[3]) ? node97 : node58;
				assign node58 = (inp[10]) ? node72 : node59;
					assign node59 = (inp[1]) ? node61 : 1'b1;
						assign node61 = (inp[5]) ? node69 : node62;
							assign node62 = (inp[2]) ? node64 : 1'b1;
								assign node64 = (inp[9]) ? node66 : 1'b1;
									assign node66 = (inp[0]) ? 1'b0 : 1'b1;
							assign node69 = (inp[2]) ? 1'b1 : 1'b0;
					assign node72 = (inp[0]) ? node82 : node73;
						assign node73 = (inp[4]) ? node75 : 1'b1;
							assign node75 = (inp[5]) ? 1'b0 : node76;
								assign node76 = (inp[1]) ? node78 : 1'b1;
									assign node78 = (inp[2]) ? 1'b0 : 1'b1;
						assign node82 = (inp[2]) ? node90 : node83;
							assign node83 = (inp[4]) ? node85 : 1'b1;
								assign node85 = (inp[9]) ? 1'b0 : node86;
									assign node86 = (inp[7]) ? 1'b0 : 1'b1;
							assign node90 = (inp[7]) ? 1'b0 : node91;
								assign node91 = (inp[1]) ? node93 : 1'b0;
									assign node93 = (inp[9]) ? 1'b0 : 1'b1;
				assign node97 = (inp[7]) ? node113 : node98;
					assign node98 = (inp[0]) ? node104 : node99;
						assign node99 = (inp[10]) ? node101 : 1'b1;
							assign node101 = (inp[2]) ? 1'b0 : 1'b1;
						assign node104 = (inp[1]) ? 1'b0 : node105;
							assign node105 = (inp[4]) ? 1'b0 : node106;
								assign node106 = (inp[9]) ? node108 : 1'b1;
									assign node108 = (inp[2]) ? 1'b0 : 1'b1;
					assign node113 = (inp[5]) ? 1'b0 : node114;
						assign node114 = (inp[2]) ? 1'b0 : node115;
							assign node115 = (inp[4]) ? 1'b0 : node116;
								assign node116 = (inp[0]) ? node118 : 1'b1;
									assign node118 = (inp[9]) ? 1'b0 : 1'b1;
		assign node124 = (inp[2]) ? node196 : node125;
			assign node125 = (inp[1]) ? node159 : node126;
				assign node126 = (inp[8]) ? node138 : node127;
					assign node127 = (inp[9]) ? node129 : 1'b1;
						assign node129 = (inp[5]) ? node131 : 1'b1;
							assign node131 = (inp[7]) ? 1'b0 : node132;
								assign node132 = (inp[3]) ? node134 : 1'b1;
									assign node134 = (inp[0]) ? 1'b0 : 1'b0;
					assign node138 = (inp[7]) ? node146 : node139;
						assign node139 = (inp[4]) ? node141 : 1'b1;
							assign node141 = (inp[9]) ? node143 : 1'b1;
								assign node143 = (inp[10]) ? 1'b0 : 1'b1;
						assign node146 = (inp[4]) ? node154 : node147;
							assign node147 = (inp[9]) ? 1'b0 : node148;
								assign node148 = (inp[5]) ? node150 : 1'b1;
									assign node150 = (inp[10]) ? 1'b0 : 1'b1;
							assign node154 = (inp[3]) ? 1'b0 : node155;
								assign node155 = (inp[0]) ? 1'b0 : 1'b1;
				assign node159 = (inp[0]) ? node185 : node160;
					assign node160 = (inp[4]) ? node170 : node161;
						assign node161 = (inp[10]) ? node163 : 1'b1;
							assign node163 = (inp[9]) ? node165 : 1'b1;
								assign node165 = (inp[3]) ? 1'b0 : node166;
									assign node166 = (inp[7]) ? 1'b0 : 1'b1;
						assign node170 = (inp[7]) ? node178 : node171;
							assign node171 = (inp[10]) ? node173 : 1'b1;
								assign node173 = (inp[3]) ? 1'b0 : node174;
									assign node174 = (inp[5]) ? 1'b0 : 1'b1;
							assign node178 = (inp[5]) ? 1'b0 : node179;
								assign node179 = (inp[8]) ? 1'b0 : node180;
									assign node180 = (inp[9]) ? 1'b0 : 1'b1;
					assign node185 = (inp[3]) ? 1'b0 : node186;
						assign node186 = (inp[10]) ? 1'b0 : node187;
							assign node187 = (inp[4]) ? node189 : 1'b1;
								assign node189 = (inp[8]) ? 1'b0 : node190;
									assign node190 = (inp[9]) ? 1'b0 : 1'b1;
			assign node196 = (inp[0]) ? node238 : node197;
				assign node197 = (inp[10]) ? node217 : node198;
					assign node198 = (inp[3]) ? node200 : 1'b1;
						assign node200 = (inp[1]) ? node212 : node201;
							assign node201 = (inp[9]) ? node207 : node202;
								assign node202 = (inp[8]) ? node204 : 1'b1;
									assign node204 = (inp[7]) ? 1'b0 : 1'b1;
								assign node207 = (inp[5]) ? 1'b0 : node208;
									assign node208 = (inp[7]) ? 1'b0 : 1'b1;
							assign node212 = (inp[7]) ? 1'b0 : node213;
								assign node213 = (inp[4]) ? 1'b0 : 1'b1;
					assign node217 = (inp[1]) ? 1'b0 : node218;
						assign node218 = (inp[7]) ? node230 : node219;
							assign node219 = (inp[5]) ? node225 : node220;
								assign node220 = (inp[3]) ? node222 : 1'b1;
									assign node222 = (inp[8]) ? 1'b0 : 1'b1;
								assign node225 = (inp[8]) ? 1'b0 : node226;
									assign node226 = (inp[9]) ? 1'b0 : 1'b1;
							assign node230 = (inp[8]) ? 1'b0 : node231;
								assign node231 = (inp[9]) ? 1'b0 : node232;
									assign node232 = (inp[4]) ? 1'b0 : 1'b1;
				assign node238 = (inp[4]) ? 1'b0 : node239;
					assign node239 = (inp[8]) ? 1'b0 : node240;
						assign node240 = (inp[9]) ? 1'b0 : node241;
							assign node241 = (inp[10]) ? 1'b0 : node242;
								assign node242 = (inp[1]) ? node244 : 1'b1;
									assign node244 = (inp[5]) ? 1'b0 : 1'b1;

endmodule