module dtc_split75_bm49 (
	input  wire [7-1:0] inp,
	output wire [10-1:0] outp
);

	wire [10-1:0] node1;
	wire [10-1:0] node2;
	wire [10-1:0] node3;
	wire [10-1:0] node4;
	wire [10-1:0] node5;
	wire [10-1:0] node6;
	wire [10-1:0] node10;
	wire [10-1:0] node13;
	wire [10-1:0] node14;
	wire [10-1:0] node17;
	wire [10-1:0] node18;
	wire [10-1:0] node21;
	wire [10-1:0] node24;
	wire [10-1:0] node25;
	wire [10-1:0] node26;
	wire [10-1:0] node29;
	wire [10-1:0] node32;
	wire [10-1:0] node33;
	wire [10-1:0] node36;
	wire [10-1:0] node39;
	wire [10-1:0] node40;
	wire [10-1:0] node41;
	wire [10-1:0] node42;
	wire [10-1:0] node43;
	wire [10-1:0] node46;
	wire [10-1:0] node49;
	wire [10-1:0] node50;
	wire [10-1:0] node53;
	wire [10-1:0] node56;
	wire [10-1:0] node57;
	wire [10-1:0] node60;
	wire [10-1:0] node61;
	wire [10-1:0] node64;
	wire [10-1:0] node67;
	wire [10-1:0] node68;
	wire [10-1:0] node69;
	wire [10-1:0] node70;
	wire [10-1:0] node73;
	wire [10-1:0] node76;
	wire [10-1:0] node78;
	wire [10-1:0] node81;
	wire [10-1:0] node82;
	wire [10-1:0] node83;
	wire [10-1:0] node86;
	wire [10-1:0] node89;
	wire [10-1:0] node90;
	wire [10-1:0] node93;
	wire [10-1:0] node96;
	wire [10-1:0] node97;
	wire [10-1:0] node98;
	wire [10-1:0] node99;
	wire [10-1:0] node100;
	wire [10-1:0] node101;
	wire [10-1:0] node105;
	wire [10-1:0] node106;
	wire [10-1:0] node109;
	wire [10-1:0] node112;
	wire [10-1:0] node113;
	wire [10-1:0] node115;
	wire [10-1:0] node118;
	wire [10-1:0] node119;
	wire [10-1:0] node122;
	wire [10-1:0] node125;
	wire [10-1:0] node126;
	wire [10-1:0] node127;
	wire [10-1:0] node128;
	wire [10-1:0] node131;
	wire [10-1:0] node134;
	wire [10-1:0] node135;
	wire [10-1:0] node138;
	wire [10-1:0] node141;
	wire [10-1:0] node142;
	wire [10-1:0] node143;
	wire [10-1:0] node147;
	wire [10-1:0] node149;
	wire [10-1:0] node152;
	wire [10-1:0] node153;
	wire [10-1:0] node154;
	wire [10-1:0] node155;
	wire [10-1:0] node157;
	wire [10-1:0] node160;
	wire [10-1:0] node162;
	wire [10-1:0] node165;
	wire [10-1:0] node166;
	wire [10-1:0] node169;
	wire [10-1:0] node172;
	wire [10-1:0] node173;
	wire [10-1:0] node174;
	wire [10-1:0] node177;
	wire [10-1:0] node178;
	wire [10-1:0] node182;
	wire [10-1:0] node183;
	wire [10-1:0] node185;
	wire [10-1:0] node188;

	assign outp = (inp[3]) ? node96 : node1;
		assign node1 = (inp[1]) ? node39 : node2;
			assign node2 = (inp[0]) ? node24 : node3;
				assign node3 = (inp[4]) ? node13 : node4;
					assign node4 = (inp[6]) ? node10 : node5;
						assign node5 = (inp[5]) ? 10'b1000000110 : node6;
							assign node6 = (inp[2]) ? 10'b1101000010 : 10'b1101010011;
						assign node10 = (inp[2]) ? 10'b1000011110 : 10'b1100001111;
					assign node13 = (inp[2]) ? node17 : node14;
						assign node14 = (inp[5]) ? 10'b1100000001 : 10'b1000001101;
						assign node17 = (inp[6]) ? node21 : node18;
							assign node18 = (inp[5]) ? 10'b1100001000 : 10'b1001000000;
							assign node21 = (inp[5]) ? 10'b1000010000 : 10'b1100010100;
				assign node24 = (inp[5]) ? node32 : node25;
					assign node25 = (inp[2]) ? node29 : node26;
						assign node26 = (inp[6]) ? 10'b0100010111 : 10'b0001000011;
						assign node29 = (inp[6]) ? 10'b0100000110 : 10'b0100011110;
					assign node32 = (inp[4]) ? node36 : node33;
						assign node33 = (inp[6]) ? 10'b0000001001 : 10'b0000000100;
						assign node36 = (inp[6]) ? 10'b0000000010 : 10'b0000011010;
			assign node39 = (inp[0]) ? node67 : node40;
				assign node40 = (inp[2]) ? node56 : node41;
					assign node41 = (inp[6]) ? node49 : node42;
						assign node42 = (inp[4]) ? node46 : node43;
							assign node43 = (inp[5]) ? 10'b0000110110 : 10'b0101110010;
							assign node46 = (inp[5]) ? 10'b0100111000 : 10'b0001110000;
						assign node49 = (inp[4]) ? node53 : node50;
							assign node50 = (inp[5]) ? 10'b0000101010 : 10'b0100101110;
							assign node53 = (inp[5]) ? 10'b0100100000 : 10'b0000101100;
					assign node56 = (inp[4]) ? node60 : node57;
						assign node57 = (inp[5]) ? 10'b0100110001 : 10'b0101100001;
						assign node60 = (inp[6]) ? node64 : node61;
							assign node61 = (inp[5]) ? 10'b0000111011 : 10'b0100111111;
							assign node64 = (inp[5]) ? 10'b0000100011 : 10'b0100100111;
				assign node67 = (inp[2]) ? node81 : node68;
					assign node68 = (inp[6]) ? node76 : node69;
						assign node69 = (inp[4]) ? node73 : node70;
							assign node70 = (inp[5]) ? 10'b1000100111 : 10'b1101100011;
							assign node73 = (inp[5]) ? 10'b1100101001 : 10'b1001100001;
						assign node76 = (inp[5]) ? node78 : 10'b1000111111;
							assign node78 = (inp[4]) ? 10'b1000110001 : 10'b1100110011;
					assign node81 = (inp[6]) ? node89 : node82;
						assign node82 = (inp[4]) ? node86 : node83;
							assign node83 = (inp[5]) ? 10'b1100111010 : 10'b1001110010;
							assign node86 = (inp[5]) ? 10'b1000111000 : 10'b1100111100;
						assign node89 = (inp[5]) ? node93 : node90;
							assign node90 = (inp[4]) ? 10'b1100100100 : 10'b1000101110;
							assign node93 = (inp[4]) ? 10'b1000100000 : 10'b1100100010;
		assign node96 = (inp[1]) ? node152 : node97;
			assign node97 = (inp[2]) ? node125 : node98;
				assign node98 = (inp[0]) ? node112 : node99;
					assign node99 = (inp[6]) ? node105 : node100;
						assign node100 = (inp[5]) ? 10'b1110111000 : node101;
							assign node101 = (inp[4]) ? 10'b1011110000 : 10'b1111110010;
						assign node105 = (inp[5]) ? node109 : node106;
							assign node106 = (inp[4]) ? 10'b1010101100 : 10'b1110101110;
							assign node109 = (inp[4]) ? 10'b1110100000 : 10'b1010101010;
					assign node112 = (inp[4]) ? node118 : node113;
						assign node113 = (inp[6]) ? node115 : 10'b0111110000;
							assign node115 = (inp[5]) ? 10'b0010101000 : 10'b0110101100;
						assign node118 = (inp[6]) ? node122 : node119;
							assign node119 = (inp[5]) ? 10'b0110101010 : 10'b0011100010;
							assign node122 = (inp[5]) ? 10'b0010110010 : 10'b0110110110;
				assign node125 = (inp[0]) ? node141 : node126;
					assign node126 = (inp[4]) ? node134 : node127;
						assign node127 = (inp[6]) ? node131 : node128;
							assign node128 = (inp[5]) ? 10'b1010100101 : 10'b1111100001;
							assign node131 = (inp[5]) ? 10'b1110110001 : 10'b1010111101;
						assign node134 = (inp[6]) ? node138 : node135;
							assign node135 = (inp[5]) ? 10'b1010111011 : 10'b1110111111;
							assign node138 = (inp[5]) ? 10'b1010100011 : 10'b1110100111;
					assign node141 = (inp[6]) ? node147 : node142;
						assign node142 = (inp[4]) ? 10'b0110111101 : node143;
							assign node143 = (inp[5]) ? 10'b0110111011 : 10'b0011110011;
						assign node147 = (inp[5]) ? node149 : 10'b0010101111;
							assign node149 = (inp[4]) ? 10'b0010100001 : 10'b0110100011;
			assign node152 = (inp[2]) ? node172 : node153;
				assign node153 = (inp[6]) ? node165 : node154;
					assign node154 = (inp[5]) ? node160 : node155;
						assign node155 = (inp[0]) ? node157 : 10'b1011000011;
							assign node157 = (inp[4]) ? 10'b0011000001 : 10'b0111000011;
						assign node160 = (inp[4]) ? node162 : 10'b0010000111;
							assign node162 = (inp[0]) ? 10'b0110001001 : 10'b1110001011;
					assign node165 = (inp[4]) ? node169 : node166;
						assign node166 = (inp[0]) ? 10'b0010011111 : 10'b1110001101;
						assign node169 = (inp[5]) ? 10'b1010010011 : 10'b1110010111;
				assign node172 = (inp[0]) ? node182 : node173;
					assign node173 = (inp[5]) ? node177 : node174;
						assign node174 = (inp[6]) ? 10'b1110000110 : 10'b1110011110;
						assign node177 = (inp[4]) ? 10'b1010000010 : node178;
							assign node178 = (inp[6]) ? 10'b1110010000 : 10'b1010000100;
					assign node182 = (inp[4]) ? node188 : node183;
						assign node183 = (inp[6]) ? node185 : 10'b0011010010;
							assign node185 = (inp[5]) ? 10'b0110000010 : 10'b0010001110;
						assign node188 = (inp[6]) ? 10'b0110000100 : 10'b0110011100;

endmodule