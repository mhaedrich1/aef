module dtc_split125_bm79 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node52;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node85;
	wire [3-1:0] node87;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node221;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node297;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node305;
	wire [3-1:0] node306;

	assign outp = (inp[6]) ? node100 : node1;
		assign node1 = (inp[9]) ? node85 : node2;
			assign node2 = (inp[0]) ? node62 : node3;
				assign node3 = (inp[10]) ? node41 : node4;
					assign node4 = (inp[8]) ? node20 : node5;
						assign node5 = (inp[7]) ? node11 : node6;
							assign node6 = (inp[3]) ? 3'b000 : node7;
								assign node7 = (inp[5]) ? 3'b110 : 3'b100;
							assign node11 = (inp[1]) ? node13 : 3'b110;
								assign node13 = (inp[11]) ? node17 : node14;
									assign node14 = (inp[2]) ? 3'b010 : 3'b110;
									assign node17 = (inp[3]) ? 3'b100 : 3'b010;
						assign node20 = (inp[7]) ? node32 : node21;
							assign node21 = (inp[2]) ? node27 : node22;
								assign node22 = (inp[11]) ? 3'b010 : node23;
									assign node23 = (inp[3]) ? 3'b110 : 3'b010;
								assign node27 = (inp[1]) ? 3'b100 : node28;
									assign node28 = (inp[3]) ? 3'b010 : 3'b110;
							assign node32 = (inp[1]) ? node36 : node33;
								assign node33 = (inp[11]) ? 3'b001 : 3'b101;
								assign node36 = (inp[11]) ? node38 : 3'b001;
									assign node38 = (inp[2]) ? 3'b010 : 3'b110;
					assign node41 = (inp[7]) ? node43 : 3'b000;
						assign node43 = (inp[1]) ? node57 : node44;
							assign node44 = (inp[8]) ? node52 : node45;
								assign node45 = (inp[4]) ? node49 : node46;
									assign node46 = (inp[5]) ? 3'b010 : 3'b010;
									assign node49 = (inp[5]) ? 3'b000 : 3'b010;
								assign node52 = (inp[5]) ? node54 : 3'b010;
									assign node54 = (inp[3]) ? 3'b010 : 3'b110;
							assign node57 = (inp[8]) ? 3'b010 : node58;
								assign node58 = (inp[11]) ? 3'b000 : 3'b100;
				assign node62 = (inp[10]) ? 3'b000 : node63;
					assign node63 = (inp[7]) ? node65 : 3'b000;
						assign node65 = (inp[2]) ? node73 : node66;
							assign node66 = (inp[11]) ? 3'b100 : node67;
								assign node67 = (inp[3]) ? 3'b010 : node68;
									assign node68 = (inp[4]) ? 3'b010 : 3'b100;
							assign node73 = (inp[4]) ? node79 : node74;
								assign node74 = (inp[3]) ? 3'b100 : node75;
									assign node75 = (inp[5]) ? 3'b010 : 3'b000;
								assign node79 = (inp[1]) ? 3'b000 : node80;
									assign node80 = (inp[3]) ? 3'b000 : 3'b100;
			assign node85 = (inp[7]) ? node87 : 3'b000;
				assign node87 = (inp[8]) ? node89 : 3'b000;
					assign node89 = (inp[0]) ? 3'b000 : node90;
						assign node90 = (inp[10]) ? 3'b000 : node91;
							assign node91 = (inp[4]) ? 3'b100 : node92;
								assign node92 = (inp[11]) ? 3'b100 : node93;
									assign node93 = (inp[1]) ? 3'b100 : 3'b010;
		assign node100 = (inp[9]) ? node214 : node101;
			assign node101 = (inp[7]) ? node167 : node102;
				assign node102 = (inp[10]) ? node132 : node103;
					assign node103 = (inp[8]) ? node117 : node104;
						assign node104 = (inp[0]) ? node110 : node105;
							assign node105 = (inp[2]) ? node107 : 3'b101;
								assign node107 = (inp[4]) ? 3'b001 : 3'b011;
							assign node110 = (inp[1]) ? node114 : node111;
								assign node111 = (inp[2]) ? 3'b010 : 3'b110;
								assign node114 = (inp[5]) ? 3'b100 : 3'b010;
						assign node117 = (inp[0]) ? node127 : node118;
							assign node118 = (inp[1]) ? node122 : node119;
								assign node119 = (inp[11]) ? 3'b011 : 3'b111;
								assign node122 = (inp[2]) ? node124 : 3'b101;
									assign node124 = (inp[11]) ? 3'b001 : 3'b011;
							assign node127 = (inp[4]) ? node129 : 3'b001;
								assign node129 = (inp[1]) ? 3'b001 : 3'b101;
					assign node132 = (inp[0]) ? node148 : node133;
						assign node133 = (inp[8]) ? node143 : node134;
							assign node134 = (inp[11]) ? node136 : 3'b110;
								assign node136 = (inp[1]) ? node140 : node137;
									assign node137 = (inp[3]) ? 3'b110 : 3'b001;
									assign node140 = (inp[2]) ? 3'b000 : 3'b010;
							assign node143 = (inp[3]) ? node145 : 3'b001;
								assign node145 = (inp[2]) ? 3'b010 : 3'b001;
						assign node148 = (inp[11]) ? node156 : node149;
							assign node149 = (inp[2]) ? node151 : 3'b010;
								assign node151 = (inp[3]) ? node153 : 3'b110;
									assign node153 = (inp[4]) ? 3'b100 : 3'b000;
							assign node156 = (inp[1]) ? node162 : node157;
								assign node157 = (inp[8]) ? node159 : 3'b100;
									assign node159 = (inp[4]) ? 3'b000 : 3'b010;
								assign node162 = (inp[4]) ? 3'b100 : node163;
									assign node163 = (inp[5]) ? 3'b100 : 3'b000;
				assign node167 = (inp[0]) ? node191 : node168;
					assign node168 = (inp[10]) ? node178 : node169;
						assign node169 = (inp[1]) ? node171 : 3'b111;
							assign node171 = (inp[2]) ? node173 : 3'b111;
								assign node173 = (inp[3]) ? 3'b111 : node174;
									assign node174 = (inp[11]) ? 3'b011 : 3'b111;
						assign node178 = (inp[1]) ? node186 : node179;
							assign node179 = (inp[2]) ? node181 : 3'b111;
								assign node181 = (inp[11]) ? node183 : 3'b011;
									assign node183 = (inp[8]) ? 3'b011 : 3'b101;
							assign node186 = (inp[11]) ? node188 : 3'b101;
								assign node188 = (inp[3]) ? 3'b001 : 3'b101;
					assign node191 = (inp[10]) ? node205 : node192;
						assign node192 = (inp[4]) ? node198 : node193;
							assign node193 = (inp[5]) ? 3'b101 : node194;
								assign node194 = (inp[3]) ? 3'b001 : 3'b101;
							assign node198 = (inp[1]) ? 3'b101 : node199;
								assign node199 = (inp[11]) ? 3'b101 : node200;
									assign node200 = (inp[5]) ? 3'b011 : 3'b011;
						assign node205 = (inp[1]) ? node211 : node206;
							assign node206 = (inp[5]) ? 3'b110 : node207;
								assign node207 = (inp[2]) ? 3'b001 : 3'b101;
							assign node211 = (inp[4]) ? 3'b010 : 3'b110;
			assign node214 = (inp[0]) ? node274 : node215;
				assign node215 = (inp[7]) ? node241 : node216;
					assign node216 = (inp[10]) ? node232 : node217;
						assign node217 = (inp[4]) ? node225 : node218;
							assign node218 = (inp[5]) ? 3'b100 : node219;
								assign node219 = (inp[1]) ? node221 : 3'b110;
									assign node221 = (inp[11]) ? 3'b010 : 3'b110;
							assign node225 = (inp[11]) ? 3'b000 : node226;
								assign node226 = (inp[1]) ? 3'b010 : node227;
									assign node227 = (inp[8]) ? 3'b110 : 3'b010;
						assign node232 = (inp[2]) ? 3'b000 : node233;
							assign node233 = (inp[1]) ? node235 : 3'b100;
								assign node235 = (inp[11]) ? 3'b000 : node236;
									assign node236 = (inp[4]) ? 3'b100 : 3'b000;
					assign node241 = (inp[11]) ? node265 : node242;
						assign node242 = (inp[10]) ? node254 : node243;
							assign node243 = (inp[1]) ? node247 : node244;
								assign node244 = (inp[5]) ? 3'b001 : 3'b011;
								assign node247 = (inp[8]) ? node251 : node248;
									assign node248 = (inp[4]) ? 3'b110 : 3'b001;
									assign node251 = (inp[2]) ? 3'b001 : 3'b101;
							assign node254 = (inp[4]) ? node262 : node255;
								assign node255 = (inp[3]) ? node259 : node256;
									assign node256 = (inp[8]) ? 3'b001 : 3'b100;
									assign node259 = (inp[8]) ? 3'b010 : 3'b010;
								assign node262 = (inp[1]) ? 3'b100 : 3'b110;
						assign node265 = (inp[4]) ? node269 : node266;
							assign node266 = (inp[8]) ? 3'b110 : 3'b010;
							assign node269 = (inp[10]) ? node271 : 3'b110;
								assign node271 = (inp[1]) ? 3'b100 : 3'b110;
				assign node274 = (inp[7]) ? node286 : node275;
					assign node275 = (inp[11]) ? 3'b000 : node276;
						assign node276 = (inp[1]) ? 3'b000 : node277;
							assign node277 = (inp[8]) ? node279 : 3'b000;
								assign node279 = (inp[5]) ? 3'b000 : node280;
									assign node280 = (inp[4]) ? 3'b000 : 3'b100;
					assign node286 = (inp[10]) ? node300 : node287;
						assign node287 = (inp[2]) ? node297 : node288;
							assign node288 = (inp[1]) ? node292 : node289;
								assign node289 = (inp[3]) ? 3'b010 : 3'b110;
								assign node292 = (inp[3]) ? 3'b100 : node293;
									assign node293 = (inp[8]) ? 3'b010 : 3'b100;
							assign node297 = (inp[3]) ? 3'b000 : 3'b100;
						assign node300 = (inp[1]) ? 3'b000 : node301;
							assign node301 = (inp[11]) ? node305 : node302;
								assign node302 = (inp[8]) ? 3'b011 : 3'b000;
								assign node305 = (inp[2]) ? 3'b000 : node306;
									assign node306 = (inp[8]) ? 3'b100 : 3'b000;

endmodule