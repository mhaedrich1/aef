module dtc_split33_bm51 (
	input  wire [8-1:0] inp,
	output wire [2-1:0] outp
);

	wire [2-1:0] node1;
	wire [2-1:0] node2;
	wire [2-1:0] node3;
	wire [2-1:0] node4;
	wire [2-1:0] node7;
	wire [2-1:0] node8;
	wire [2-1:0] node10;
	wire [2-1:0] node12;
	wire [2-1:0] node15;
	wire [2-1:0] node16;
	wire [2-1:0] node20;
	wire [2-1:0] node21;
	wire [2-1:0] node22;
	wire [2-1:0] node26;
	wire [2-1:0] node27;
	wire [2-1:0] node30;
	wire [2-1:0] node33;
	wire [2-1:0] node34;
	wire [2-1:0] node35;
	wire [2-1:0] node37;
	wire [2-1:0] node40;
	wire [2-1:0] node43;
	wire [2-1:0] node44;
	wire [2-1:0] node45;
	wire [2-1:0] node50;
	wire [2-1:0] node51;
	wire [2-1:0] node52;
	wire [2-1:0] node53;
	wire [2-1:0] node56;
	wire [2-1:0] node59;
	wire [2-1:0] node60;
	wire [2-1:0] node61;
	wire [2-1:0] node65;
	wire [2-1:0] node68;
	wire [2-1:0] node69;
	wire [2-1:0] node71;
	wire [2-1:0] node72;

	assign outp = (inp[2]) ? node50 : node1;
		assign node1 = (inp[6]) ? node33 : node2;
			assign node2 = (inp[0]) ? node20 : node3;
				assign node3 = (inp[7]) ? node7 : node4;
					assign node4 = (inp[3]) ? 2'b01 : 2'b00;
					assign node7 = (inp[3]) ? node15 : node8;
						assign node8 = (inp[4]) ? node10 : 2'b11;
							assign node10 = (inp[5]) ? node12 : 2'b11;
								assign node12 = (inp[1]) ? 2'b11 : 2'b10;
						assign node15 = (inp[1]) ? 2'b10 : node16;
							assign node16 = (inp[5]) ? 2'b11 : 2'b10;
				assign node20 = (inp[1]) ? node26 : node21;
					assign node21 = (inp[4]) ? 2'b11 : node22;
						assign node22 = (inp[7]) ? 2'b10 : 2'b11;
					assign node26 = (inp[5]) ? node30 : node27;
						assign node27 = (inp[3]) ? 2'b11 : 2'b10;
						assign node30 = (inp[3]) ? 2'b10 : 2'b11;
			assign node33 = (inp[7]) ? node43 : node34;
				assign node34 = (inp[0]) ? node40 : node35;
					assign node35 = (inp[4]) ? node37 : 2'b10;
						assign node37 = (inp[5]) ? 2'b10 : 2'b11;
					assign node40 = (inp[5]) ? 2'b01 : 2'b00;
				assign node43 = (inp[4]) ? 2'b01 : node44;
					assign node44 = (inp[1]) ? 2'b00 : node45;
						assign node45 = (inp[0]) ? 2'b01 : 2'b00;
		assign node50 = (inp[7]) ? node68 : node51;
			assign node51 = (inp[0]) ? node59 : node52;
				assign node52 = (inp[1]) ? node56 : node53;
					assign node53 = (inp[4]) ? 2'b11 : 2'b10;
					assign node56 = (inp[4]) ? 2'b10 : 2'b11;
				assign node59 = (inp[3]) ? node65 : node60;
					assign node60 = (inp[1]) ? 2'b01 : node61;
						assign node61 = (inp[6]) ? 2'b01 : 2'b00;
					assign node65 = (inp[1]) ? 2'b00 : 2'b01;
			assign node68 = (inp[6]) ? 2'b00 : node69;
				assign node69 = (inp[3]) ? node71 : 2'b01;
					assign node71 = (inp[4]) ? 2'b00 : node72;
						assign node72 = (inp[0]) ? 2'b00 : 2'b01;

endmodule