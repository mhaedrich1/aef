module dtc_split33_bm15 (
	input  wire [15-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node7;
	wire [1-1:0] node8;
	wire [1-1:0] node10;
	wire [1-1:0] node12;
	wire [1-1:0] node14;
	wire [1-1:0] node16;
	wire [1-1:0] node19;
	wire [1-1:0] node20;
	wire [1-1:0] node22;
	wire [1-1:0] node24;
	wire [1-1:0] node26;
	wire [1-1:0] node29;
	wire [1-1:0] node31;
	wire [1-1:0] node32;
	wire [1-1:0] node34;
	wire [1-1:0] node37;
	wire [1-1:0] node39;
	wire [1-1:0] node40;
	wire [1-1:0] node44;
	wire [1-1:0] node45;
	wire [1-1:0] node46;
	wire [1-1:0] node48;
	wire [1-1:0] node50;
	wire [1-1:0] node52;
	wire [1-1:0] node54;
	wire [1-1:0] node56;
	wire [1-1:0] node59;
	wire [1-1:0] node60;
	wire [1-1:0] node62;
	wire [1-1:0] node64;
	wire [1-1:0] node66;
	wire [1-1:0] node69;
	wire [1-1:0] node70;
	wire [1-1:0] node71;
	wire [1-1:0] node73;
	wire [1-1:0] node75;
	wire [1-1:0] node79;
	wire [1-1:0] node80;
	wire [1-1:0] node82;
	wire [1-1:0] node83;
	wire [1-1:0] node87;
	wire [1-1:0] node88;
	wire [1-1:0] node90;
	wire [1-1:0] node94;
	wire [1-1:0] node95;
	wire [1-1:0] node96;
	wire [1-1:0] node98;
	wire [1-1:0] node100;
	wire [1-1:0] node102;
	wire [1-1:0] node105;
	wire [1-1:0] node106;
	wire [1-1:0] node108;
	wire [1-1:0] node110;
	wire [1-1:0] node112;
	wire [1-1:0] node115;
	wire [1-1:0] node116;
	wire [1-1:0] node118;
	wire [1-1:0] node120;
	wire [1-1:0] node123;
	wire [1-1:0] node124;
	wire [1-1:0] node126;
	wire [1-1:0] node130;
	wire [1-1:0] node131;
	wire [1-1:0] node132;
	wire [1-1:0] node134;
	wire [1-1:0] node136;
	wire [1-1:0] node139;
	wire [1-1:0] node140;
	wire [1-1:0] node142;
	wire [1-1:0] node144;
	wire [1-1:0] node147;
	wire [1-1:0] node148;
	wire [1-1:0] node149;
	wire [1-1:0] node153;
	wire [1-1:0] node154;
	wire [1-1:0] node158;
	wire [1-1:0] node159;
	wire [1-1:0] node161;
	wire [1-1:0] node162;
	wire [1-1:0] node164;
	wire [1-1:0] node168;
	wire [1-1:0] node169;
	wire [1-1:0] node170;
	wire [1-1:0] node172;
	wire [1-1:0] node175;
	wire [1-1:0] node176;
	wire [1-1:0] node181;
	wire [1-1:0] node182;
	wire [1-1:0] node183;
	wire [1-1:0] node185;
	wire [1-1:0] node186;
	wire [1-1:0] node188;
	wire [1-1:0] node190;
	wire [1-1:0] node192;
	wire [1-1:0] node194;
	wire [1-1:0] node197;
	wire [1-1:0] node198;
	wire [1-1:0] node200;
	wire [1-1:0] node202;
	wire [1-1:0] node205;
	wire [1-1:0] node206;
	wire [1-1:0] node208;
	wire [1-1:0] node209;
	wire [1-1:0] node213;
	wire [1-1:0] node214;
	wire [1-1:0] node216;
	wire [1-1:0] node219;
	wire [1-1:0] node220;
	wire [1-1:0] node224;
	wire [1-1:0] node225;
	wire [1-1:0] node226;
	wire [1-1:0] node228;
	wire [1-1:0] node229;
	wire [1-1:0] node231;
	wire [1-1:0] node233;
	wire [1-1:0] node237;
	wire [1-1:0] node238;
	wire [1-1:0] node240;
	wire [1-1:0] node242;
	wire [1-1:0] node245;
	wire [1-1:0] node246;
	wire [1-1:0] node248;
	wire [1-1:0] node250;
	wire [1-1:0] node253;
	wire [1-1:0] node254;
	wire [1-1:0] node256;
	wire [1-1:0] node260;
	wire [1-1:0] node261;
	wire [1-1:0] node262;
	wire [1-1:0] node264;
	wire [1-1:0] node266;
	wire [1-1:0] node269;
	wire [1-1:0] node270;
	wire [1-1:0] node272;
	wire [1-1:0] node275;
	wire [1-1:0] node276;
	wire [1-1:0] node278;
	wire [1-1:0] node281;
	wire [1-1:0] node282;
	wire [1-1:0] node286;
	wire [1-1:0] node287;
	wire [1-1:0] node288;
	wire [1-1:0] node289;
	wire [1-1:0] node291;
	wire [1-1:0] node294;
	wire [1-1:0] node297;
	wire [1-1:0] node299;
	wire [1-1:0] node300;
	wire [1-1:0] node304;
	wire [1-1:0] node305;
	wire [1-1:0] node307;
	wire [1-1:0] node308;
	wire [1-1:0] node313;
	wire [1-1:0] node314;
	wire [1-1:0] node315;
	wire [1-1:0] node317;
	wire [1-1:0] node319;
	wire [1-1:0] node320;
	wire [1-1:0] node322;
	wire [1-1:0] node323;
	wire [1-1:0] node327;
	wire [1-1:0] node328;
	wire [1-1:0] node331;
	wire [1-1:0] node332;
	wire [1-1:0] node336;
	wire [1-1:0] node337;
	wire [1-1:0] node338;
	wire [1-1:0] node340;
	wire [1-1:0] node342;
	wire [1-1:0] node345;
	wire [1-1:0] node346;
	wire [1-1:0] node348;
	wire [1-1:0] node351;
	wire [1-1:0] node352;
	wire [1-1:0] node355;
	wire [1-1:0] node356;
	wire [1-1:0] node360;
	wire [1-1:0] node361;
	wire [1-1:0] node362;
	wire [1-1:0] node364;
	wire [1-1:0] node367;
	wire [1-1:0] node368;
	wire [1-1:0] node371;
	wire [1-1:0] node372;
	wire [1-1:0] node376;
	wire [1-1:0] node377;
	wire [1-1:0] node378;
	wire [1-1:0] node380;
	wire [1-1:0] node383;
	wire [1-1:0] node387;
	wire [1-1:0] node388;
	wire [1-1:0] node389;
	wire [1-1:0] node391;
	wire [1-1:0] node392;
	wire [1-1:0] node394;
	wire [1-1:0] node397;
	wire [1-1:0] node398;
	wire [1-1:0] node400;
	wire [1-1:0] node403;
	wire [1-1:0] node404;
	wire [1-1:0] node408;
	wire [1-1:0] node409;
	wire [1-1:0] node410;
	wire [1-1:0] node412;
	wire [1-1:0] node415;
	wire [1-1:0] node417;
	wire [1-1:0] node418;
	wire [1-1:0] node422;
	wire [1-1:0] node423;
	wire [1-1:0] node424;
	wire [1-1:0] node426;
	wire [1-1:0] node429;
	wire [1-1:0] node430;
	wire [1-1:0] node435;
	wire [1-1:0] node436;
	wire [1-1:0] node437;
	wire [1-1:0] node439;
	wire [1-1:0] node440;
	wire [1-1:0] node444;
	wire [1-1:0] node445;
	wire [1-1:0] node447;
	wire [1-1:0] node448;
	wire [1-1:0] node452;
	wire [1-1:0] node453;
	wire [1-1:0] node454;
	wire [1-1:0] node459;
	wire [1-1:0] node460;
	wire [1-1:0] node461;
	wire [1-1:0] node462;
	wire [1-1:0] node464;
	wire [1-1:0] node467;
	wire [1-1:0] node470;
	wire [1-1:0] node471;
	wire [1-1:0] node476;
	wire [1-1:0] node477;
	wire [1-1:0] node478;
	wire [1-1:0] node479;
	wire [1-1:0] node480;
	wire [1-1:0] node482;
	wire [1-1:0] node484;
	wire [1-1:0] node486;
	wire [1-1:0] node488;
	wire [1-1:0] node491;
	wire [1-1:0] node492;
	wire [1-1:0] node494;
	wire [1-1:0] node496;
	wire [1-1:0] node498;
	wire [1-1:0] node500;
	wire [1-1:0] node503;
	wire [1-1:0] node504;
	wire [1-1:0] node506;
	wire [1-1:0] node508;
	wire [1-1:0] node511;
	wire [1-1:0] node512;
	wire [1-1:0] node514;
	wire [1-1:0] node516;
	wire [1-1:0] node519;
	wire [1-1:0] node520;
	wire [1-1:0] node523;
	wire [1-1:0] node526;
	wire [1-1:0] node527;
	wire [1-1:0] node529;
	wire [1-1:0] node531;
	wire [1-1:0] node532;
	wire [1-1:0] node534;
	wire [1-1:0] node537;
	wire [1-1:0] node540;
	wire [1-1:0] node541;
	wire [1-1:0] node542;
	wire [1-1:0] node544;
	wire [1-1:0] node545;
	wire [1-1:0] node549;
	wire [1-1:0] node550;
	wire [1-1:0] node552;
	wire [1-1:0] node555;
	wire [1-1:0] node556;
	wire [1-1:0] node560;
	wire [1-1:0] node561;
	wire [1-1:0] node562;
	wire [1-1:0] node564;
	wire [1-1:0] node566;
	wire [1-1:0] node569;
	wire [1-1:0] node572;
	wire [1-1:0] node573;
	wire [1-1:0] node575;
	wire [1-1:0] node576;
	wire [1-1:0] node581;
	wire [1-1:0] node582;
	wire [1-1:0] node583;
	wire [1-1:0] node585;
	wire [1-1:0] node586;
	wire [1-1:0] node588;
	wire [1-1:0] node590;
	wire [1-1:0] node591;
	wire [1-1:0] node595;
	wire [1-1:0] node596;
	wire [1-1:0] node598;
	wire [1-1:0] node600;
	wire [1-1:0] node603;
	wire [1-1:0] node604;
	wire [1-1:0] node606;
	wire [1-1:0] node609;
	wire [1-1:0] node610;
	wire [1-1:0] node614;
	wire [1-1:0] node615;
	wire [1-1:0] node616;
	wire [1-1:0] node618;
	wire [1-1:0] node620;
	wire [1-1:0] node622;
	wire [1-1:0] node625;
	wire [1-1:0] node626;
	wire [1-1:0] node628;
	wire [1-1:0] node630;
	wire [1-1:0] node633;
	wire [1-1:0] node634;
	wire [1-1:0] node638;
	wire [1-1:0] node639;
	wire [1-1:0] node641;
	wire [1-1:0] node643;
	wire [1-1:0] node644;
	wire [1-1:0] node648;
	wire [1-1:0] node649;
	wire [1-1:0] node650;
	wire [1-1:0] node652;
	wire [1-1:0] node657;
	wire [1-1:0] node658;
	wire [1-1:0] node659;
	wire [1-1:0] node660;
	wire [1-1:0] node662;
	wire [1-1:0] node664;
	wire [1-1:0] node666;
	wire [1-1:0] node669;
	wire [1-1:0] node670;
	wire [1-1:0] node672;
	wire [1-1:0] node674;
	wire [1-1:0] node677;
	wire [1-1:0] node678;
	wire [1-1:0] node680;
	wire [1-1:0] node683;
	wire [1-1:0] node684;
	wire [1-1:0] node688;
	wire [1-1:0] node689;
	wire [1-1:0] node690;
	wire [1-1:0] node692;
	wire [1-1:0] node695;
	wire [1-1:0] node696;
	wire [1-1:0] node698;
	wire [1-1:0] node701;
	wire [1-1:0] node702;
	wire [1-1:0] node706;
	wire [1-1:0] node707;
	wire [1-1:0] node708;
	wire [1-1:0] node710;
	wire [1-1:0] node715;
	wire [1-1:0] node716;
	wire [1-1:0] node717;
	wire [1-1:0] node719;
	wire [1-1:0] node720;
	wire [1-1:0] node722;
	wire [1-1:0] node726;
	wire [1-1:0] node727;
	wire [1-1:0] node728;
	wire [1-1:0] node730;
	wire [1-1:0] node735;
	wire [1-1:0] node736;
	wire [1-1:0] node737;
	wire [1-1:0] node739;
	wire [1-1:0] node744;
	wire [1-1:0] node745;
	wire [1-1:0] node746;
	wire [1-1:0] node747;
	wire [1-1:0] node748;
	wire [1-1:0] node750;
	wire [1-1:0] node752;
	wire [1-1:0] node755;
	wire [1-1:0] node756;
	wire [1-1:0] node758;
	wire [1-1:0] node760;
	wire [1-1:0] node762;
	wire [1-1:0] node765;
	wire [1-1:0] node766;
	wire [1-1:0] node768;
	wire [1-1:0] node770;
	wire [1-1:0] node773;
	wire [1-1:0] node774;
	wire [1-1:0] node776;
	wire [1-1:0] node779;
	wire [1-1:0] node780;
	wire [1-1:0] node784;
	wire [1-1:0] node785;
	wire [1-1:0] node786;
	wire [1-1:0] node787;
	wire [1-1:0] node789;
	wire [1-1:0] node793;
	wire [1-1:0] node794;
	wire [1-1:0] node796;
	wire [1-1:0] node798;
	wire [1-1:0] node801;
	wire [1-1:0] node802;
	wire [1-1:0] node803;
	wire [1-1:0] node807;
	wire [1-1:0] node808;
	wire [1-1:0] node812;
	wire [1-1:0] node813;
	wire [1-1:0] node815;
	wire [1-1:0] node816;
	wire [1-1:0] node818;
	wire [1-1:0] node821;
	wire [1-1:0] node822;
	wire [1-1:0] node826;
	wire [1-1:0] node827;
	wire [1-1:0] node828;
	wire [1-1:0] node830;
	wire [1-1:0] node833;
	wire [1-1:0] node834;
	wire [1-1:0] node839;
	wire [1-1:0] node840;
	wire [1-1:0] node841;
	wire [1-1:0] node842;
	wire [1-1:0] node844;
	wire [1-1:0] node846;
	wire [1-1:0] node849;
	wire [1-1:0] node850;
	wire [1-1:0] node852;
	wire [1-1:0] node855;
	wire [1-1:0] node856;
	wire [1-1:0] node858;
	wire [1-1:0] node862;
	wire [1-1:0] node863;
	wire [1-1:0] node864;
	wire [1-1:0] node866;
	wire [1-1:0] node868;
	wire [1-1:0] node871;
	wire [1-1:0] node872;
	wire [1-1:0] node874;
	wire [1-1:0] node878;
	wire [1-1:0] node879;
	wire [1-1:0] node881;
	wire [1-1:0] node882;
	wire [1-1:0] node887;
	wire [1-1:0] node888;
	wire [1-1:0] node889;
	wire [1-1:0] node890;
	wire [1-1:0] node892;
	wire [1-1:0] node894;
	wire [1-1:0] node897;
	wire [1-1:0] node898;
	wire [1-1:0] node900;
	wire [1-1:0] node903;
	wire [1-1:0] node904;
	wire [1-1:0] node908;
	wire [1-1:0] node909;
	wire [1-1:0] node910;
	wire [1-1:0] node912;
	wire [1-1:0] node917;
	wire [1-1:0] node918;
	wire [1-1:0] node919;
	wire [1-1:0] node922;
	wire [1-1:0] node923;
	wire [1-1:0] node924;
	wire [1-1:0] node929;
	wire [1-1:0] node930;
	wire [1-1:0] node931;
	wire [1-1:0] node936;
	wire [1-1:0] node937;
	wire [1-1:0] node938;
	wire [1-1:0] node939;
	wire [1-1:0] node940;
	wire [1-1:0] node942;
	wire [1-1:0] node944;
	wire [1-1:0] node947;
	wire [1-1:0] node948;
	wire [1-1:0] node950;
	wire [1-1:0] node953;
	wire [1-1:0] node954;
	wire [1-1:0] node956;
	wire [1-1:0] node959;
	wire [1-1:0] node960;
	wire [1-1:0] node964;
	wire [1-1:0] node965;
	wire [1-1:0] node966;
	wire [1-1:0] node968;
	wire [1-1:0] node970;
	wire [1-1:0] node973;
	wire [1-1:0] node974;
	wire [1-1:0] node975;
	wire [1-1:0] node979;
	wire [1-1:0] node980;
	wire [1-1:0] node984;
	wire [1-1:0] node985;
	wire [1-1:0] node987;
	wire [1-1:0] node988;
	wire [1-1:0] node993;
	wire [1-1:0] node994;
	wire [1-1:0] node995;
	wire [1-1:0] node997;
	wire [1-1:0] node998;
	wire [1-1:0] node1000;
	wire [1-1:0] node1003;
	wire [1-1:0] node1004;
	wire [1-1:0] node1008;
	wire [1-1:0] node1009;
	wire [1-1:0] node1010;
	wire [1-1:0] node1012;
	wire [1-1:0] node1015;
	wire [1-1:0] node1016;
	wire [1-1:0] node1020;
	wire [1-1:0] node1021;
	wire [1-1:0] node1025;
	wire [1-1:0] node1026;
	wire [1-1:0] node1027;
	wire [1-1:0] node1029;
	wire [1-1:0] node1030;
	wire [1-1:0] node1034;
	wire [1-1:0] node1035;
	wire [1-1:0] node1036;
	wire [1-1:0] node1042;
	wire [1-1:0] node1043;
	wire [1-1:0] node1044;
	wire [1-1:0] node1045;
	wire [1-1:0] node1047;
	wire [1-1:0] node1048;
	wire [1-1:0] node1050;
	wire [1-1:0] node1053;
	wire [1-1:0] node1054;
	wire [1-1:0] node1058;
	wire [1-1:0] node1059;
	wire [1-1:0] node1061;
	wire [1-1:0] node1062;
	wire [1-1:0] node1066;
	wire [1-1:0] node1067;
	wire [1-1:0] node1068;
	wire [1-1:0] node1073;
	wire [1-1:0] node1074;
	wire [1-1:0] node1075;
	wire [1-1:0] node1077;
	wire [1-1:0] node1078;
	wire [1-1:0] node1082;
	wire [1-1:0] node1083;
	wire [1-1:0] node1084;
	wire [1-1:0] node1090;
	wire [1-1:0] node1091;
	wire [1-1:0] node1092;
	wire [1-1:0] node1093;
	wire [1-1:0] node1096;
	wire [1-1:0] node1097;
	wire [1-1:0] node1098;
	wire [1-1:0] node1104;
	wire [1-1:0] node1106;
	wire [1-1:0] node1107;
	wire [1-1:0] node1108;
	wire [1-1:0] node1109;
	wire [1-1:0] node1115;
	wire [1-1:0] node1116;
	wire [1-1:0] node1117;
	wire [1-1:0] node1118;
	wire [1-1:0] node1119;
	wire [1-1:0] node1121;
	wire [1-1:0] node1122;
	wire [1-1:0] node1123;
	wire [1-1:0] node1125;
	wire [1-1:0] node1127;
	wire [1-1:0] node1129;
	wire [1-1:0] node1133;
	wire [1-1:0] node1134;
	wire [1-1:0] node1136;
	wire [1-1:0] node1138;
	wire [1-1:0] node1141;
	wire [1-1:0] node1142;
	wire [1-1:0] node1144;
	wire [1-1:0] node1146;
	wire [1-1:0] node1149;
	wire [1-1:0] node1150;
	wire [1-1:0] node1152;
	wire [1-1:0] node1155;
	wire [1-1:0] node1156;
	wire [1-1:0] node1160;
	wire [1-1:0] node1161;
	wire [1-1:0] node1163;
	wire [1-1:0] node1165;
	wire [1-1:0] node1166;
	wire [1-1:0] node1168;
	wire [1-1:0] node1170;
	wire [1-1:0] node1173;
	wire [1-1:0] node1174;
	wire [1-1:0] node1178;
	wire [1-1:0] node1179;
	wire [1-1:0] node1181;
	wire [1-1:0] node1182;
	wire [1-1:0] node1184;
	wire [1-1:0] node1187;
	wire [1-1:0] node1188;
	wire [1-1:0] node1190;
	wire [1-1:0] node1193;
	wire [1-1:0] node1194;
	wire [1-1:0] node1198;
	wire [1-1:0] node1199;
	wire [1-1:0] node1201;
	wire [1-1:0] node1202;
	wire [1-1:0] node1204;
	wire [1-1:0] node1208;
	wire [1-1:0] node1209;
	wire [1-1:0] node1210;
	wire [1-1:0] node1215;
	wire [1-1:0] node1216;
	wire [1-1:0] node1217;
	wire [1-1:0] node1218;
	wire [1-1:0] node1220;
	wire [1-1:0] node1222;
	wire [1-1:0] node1224;
	wire [1-1:0] node1227;
	wire [1-1:0] node1228;
	wire [1-1:0] node1230;
	wire [1-1:0] node1232;
	wire [1-1:0] node1234;
	wire [1-1:0] node1237;
	wire [1-1:0] node1238;
	wire [1-1:0] node1240;
	wire [1-1:0] node1242;
	wire [1-1:0] node1245;
	wire [1-1:0] node1246;
	wire [1-1:0] node1249;
	wire [1-1:0] node1250;
	wire [1-1:0] node1254;
	wire [1-1:0] node1255;
	wire [1-1:0] node1257;
	wire [1-1:0] node1258;
	wire [1-1:0] node1259;
	wire [1-1:0] node1263;
	wire [1-1:0] node1264;
	wire [1-1:0] node1266;
	wire [1-1:0] node1269;
	wire [1-1:0] node1270;
	wire [1-1:0] node1273;
	wire [1-1:0] node1276;
	wire [1-1:0] node1277;
	wire [1-1:0] node1279;
	wire [1-1:0] node1280;
	wire [1-1:0] node1283;
	wire [1-1:0] node1284;
	wire [1-1:0] node1288;
	wire [1-1:0] node1289;
	wire [1-1:0] node1291;
	wire [1-1:0] node1292;
	wire [1-1:0] node1297;
	wire [1-1:0] node1298;
	wire [1-1:0] node1299;
	wire [1-1:0] node1300;
	wire [1-1:0] node1302;
	wire [1-1:0] node1304;
	wire [1-1:0] node1305;
	wire [1-1:0] node1309;
	wire [1-1:0] node1310;
	wire [1-1:0] node1312;
	wire [1-1:0] node1315;
	wire [1-1:0] node1316;
	wire [1-1:0] node1319;
	wire [1-1:0] node1320;
	wire [1-1:0] node1324;
	wire [1-1:0] node1325;
	wire [1-1:0] node1327;
	wire [1-1:0] node1328;
	wire [1-1:0] node1330;
	wire [1-1:0] node1333;
	wire [1-1:0] node1334;
	wire [1-1:0] node1338;
	wire [1-1:0] node1339;
	wire [1-1:0] node1340;
	wire [1-1:0] node1342;
	wire [1-1:0] node1347;
	wire [1-1:0] node1348;
	wire [1-1:0] node1349;
	wire [1-1:0] node1350;
	wire [1-1:0] node1352;
	wire [1-1:0] node1354;
	wire [1-1:0] node1357;
	wire [1-1:0] node1358;
	wire [1-1:0] node1359;
	wire [1-1:0] node1363;
	wire [1-1:0] node1364;
	wire [1-1:0] node1368;
	wire [1-1:0] node1369;
	wire [1-1:0] node1371;
	wire [1-1:0] node1372;
	wire [1-1:0] node1377;
	wire [1-1:0] node1378;
	wire [1-1:0] node1379;
	wire [1-1:0] node1381;
	wire [1-1:0] node1386;
	wire [1-1:0] node1387;
	wire [1-1:0] node1388;
	wire [1-1:0] node1389;
	wire [1-1:0] node1391;
	wire [1-1:0] node1393;
	wire [1-1:0] node1394;
	wire [1-1:0] node1396;
	wire [1-1:0] node1398;
	wire [1-1:0] node1401;
	wire [1-1:0] node1402;
	wire [1-1:0] node1404;
	wire [1-1:0] node1408;
	wire [1-1:0] node1409;
	wire [1-1:0] node1411;
	wire [1-1:0] node1412;
	wire [1-1:0] node1414;
	wire [1-1:0] node1417;
	wire [1-1:0] node1418;
	wire [1-1:0] node1420;
	wire [1-1:0] node1424;
	wire [1-1:0] node1425;
	wire [1-1:0] node1426;
	wire [1-1:0] node1428;
	wire [1-1:0] node1430;
	wire [1-1:0] node1433;
	wire [1-1:0] node1434;
	wire [1-1:0] node1436;
	wire [1-1:0] node1440;
	wire [1-1:0] node1441;
	wire [1-1:0] node1443;
	wire [1-1:0] node1444;
	wire [1-1:0] node1449;
	wire [1-1:0] node1450;
	wire [1-1:0] node1451;
	wire [1-1:0] node1452;
	wire [1-1:0] node1454;
	wire [1-1:0] node1456;
	wire [1-1:0] node1459;
	wire [1-1:0] node1460;
	wire [1-1:0] node1461;
	wire [1-1:0] node1463;
	wire [1-1:0] node1467;
	wire [1-1:0] node1468;
	wire [1-1:0] node1470;
	wire [1-1:0] node1473;
	wire [1-1:0] node1474;
	wire [1-1:0] node1478;
	wire [1-1:0] node1479;
	wire [1-1:0] node1481;
	wire [1-1:0] node1482;
	wire [1-1:0] node1484;
	wire [1-1:0] node1487;
	wire [1-1:0] node1488;
	wire [1-1:0] node1492;
	wire [1-1:0] node1493;
	wire [1-1:0] node1494;
	wire [1-1:0] node1496;
	wire [1-1:0] node1499;
	wire [1-1:0] node1502;
	wire [1-1:0] node1503;
	wire [1-1:0] node1507;
	wire [1-1:0] node1508;
	wire [1-1:0] node1509;
	wire [1-1:0] node1511;
	wire [1-1:0] node1512;
	wire [1-1:0] node1514;
	wire [1-1:0] node1518;
	wire [1-1:0] node1519;
	wire [1-1:0] node1520;
	wire [1-1:0] node1522;
	wire [1-1:0] node1525;
	wire [1-1:0] node1526;
	wire [1-1:0] node1531;
	wire [1-1:0] node1532;
	wire [1-1:0] node1533;
	wire [1-1:0] node1534;
	wire [1-1:0] node1536;
	wire [1-1:0] node1539;
	wire [1-1:0] node1540;
	wire [1-1:0] node1546;
	wire [1-1:0] node1547;
	wire [1-1:0] node1548;
	wire [1-1:0] node1549;
	wire [1-1:0] node1550;
	wire [1-1:0] node1552;
	wire [1-1:0] node1554;
	wire [1-1:0] node1556;
	wire [1-1:0] node1559;
	wire [1-1:0] node1560;
	wire [1-1:0] node1562;
	wire [1-1:0] node1565;
	wire [1-1:0] node1566;
	wire [1-1:0] node1569;
	wire [1-1:0] node1570;
	wire [1-1:0] node1574;
	wire [1-1:0] node1575;
	wire [1-1:0] node1576;
	wire [1-1:0] node1578;
	wire [1-1:0] node1580;
	wire [1-1:0] node1583;
	wire [1-1:0] node1584;
	wire [1-1:0] node1586;
	wire [1-1:0] node1590;
	wire [1-1:0] node1591;
	wire [1-1:0] node1592;
	wire [1-1:0] node1597;
	wire [1-1:0] node1598;
	wire [1-1:0] node1599;
	wire [1-1:0] node1600;
	wire [1-1:0] node1602;
	wire [1-1:0] node1604;
	wire [1-1:0] node1607;
	wire [1-1:0] node1608;
	wire [1-1:0] node1610;
	wire [1-1:0] node1613;
	wire [1-1:0] node1614;
	wire [1-1:0] node1618;
	wire [1-1:0] node1619;
	wire [1-1:0] node1620;
	wire [1-1:0] node1622;
	wire [1-1:0] node1625;
	wire [1-1:0] node1626;
	wire [1-1:0] node1631;
	wire [1-1:0] node1632;
	wire [1-1:0] node1633;
	wire [1-1:0] node1634;
	wire [1-1:0] node1636;
	wire [1-1:0] node1639;
	wire [1-1:0] node1640;
	wire [1-1:0] node1646;
	wire [1-1:0] node1647;
	wire [1-1:0] node1648;
	wire [1-1:0] node1649;
	wire [1-1:0] node1650;
	wire [1-1:0] node1652;
	wire [1-1:0] node1655;
	wire [1-1:0] node1656;
	wire [1-1:0] node1658;
	wire [1-1:0] node1662;
	wire [1-1:0] node1663;
	wire [1-1:0] node1664;
	wire [1-1:0] node1666;
	wire [1-1:0] node1671;
	wire [1-1:0] node1672;
	wire [1-1:0] node1673;
	wire [1-1:0] node1674;
	wire [1-1:0] node1676;
	wire [1-1:0] node1679;
	wire [1-1:0] node1680;
	wire [1-1:0] node1684;
	wire [1-1:0] node1685;
	wire [1-1:0] node1690;
	wire [1-1:0] node1691;
	wire [1-1:0] node1692;
	wire [1-1:0] node1693;
	wire [1-1:0] node1694;
	wire [1-1:0] node1696;
	wire [1-1:0] node1699;
	wire [1-1:0] node1703;
	wire [1-1:0] node1704;
	wire [1-1:0] node1705;
	wire [1-1:0] node1706;
	wire [1-1:0] node1713;
	wire [1-1:0] node1714;
	wire [1-1:0] node1715;
	wire [1-1:0] node1716;
	wire [1-1:0] node1717;
	wire [1-1:0] node1719;
	wire [1-1:0] node1721;
	wire [1-1:0] node1723;
	wire [1-1:0] node1724;
	wire [1-1:0] node1726;
	wire [1-1:0] node1729;
	wire [1-1:0] node1730;
	wire [1-1:0] node1734;
	wire [1-1:0] node1735;
	wire [1-1:0] node1736;
	wire [1-1:0] node1738;
	wire [1-1:0] node1740;
	wire [1-1:0] node1742;
	wire [1-1:0] node1745;
	wire [1-1:0] node1747;
	wire [1-1:0] node1748;
	wire [1-1:0] node1750;
	wire [1-1:0] node1754;
	wire [1-1:0] node1755;
	wire [1-1:0] node1757;
	wire [1-1:0] node1758;
	wire [1-1:0] node1760;
	wire [1-1:0] node1763;
	wire [1-1:0] node1766;
	wire [1-1:0] node1767;
	wire [1-1:0] node1768;
	wire [1-1:0] node1771;
	wire [1-1:0] node1772;
	wire [1-1:0] node1777;
	wire [1-1:0] node1778;
	wire [1-1:0] node1779;
	wire [1-1:0] node1781;
	wire [1-1:0] node1782;
	wire [1-1:0] node1784;
	wire [1-1:0] node1786;
	wire [1-1:0] node1789;
	wire [1-1:0] node1790;
	wire [1-1:0] node1792;
	wire [1-1:0] node1796;
	wire [1-1:0] node1797;
	wire [1-1:0] node1799;
	wire [1-1:0] node1800;
	wire [1-1:0] node1802;
	wire [1-1:0] node1806;
	wire [1-1:0] node1807;
	wire [1-1:0] node1811;
	wire [1-1:0] node1812;
	wire [1-1:0] node1813;
	wire [1-1:0] node1815;
	wire [1-1:0] node1816;
	wire [1-1:0] node1818;
	wire [1-1:0] node1821;
	wire [1-1:0] node1822;
	wire [1-1:0] node1826;
	wire [1-1:0] node1827;
	wire [1-1:0] node1828;
	wire [1-1:0] node1830;
	wire [1-1:0] node1833;
	wire [1-1:0] node1834;
	wire [1-1:0] node1838;
	wire [1-1:0] node1839;
	wire [1-1:0] node1843;
	wire [1-1:0] node1844;
	wire [1-1:0] node1845;
	wire [1-1:0] node1846;
	wire [1-1:0] node1848;
	wire [1-1:0] node1851;
	wire [1-1:0] node1852;
	wire [1-1:0] node1858;
	wire [1-1:0] node1859;
	wire [1-1:0] node1860;
	wire [1-1:0] node1861;
	wire [1-1:0] node1862;
	wire [1-1:0] node1864;
	wire [1-1:0] node1866;
	wire [1-1:0] node1869;
	wire [1-1:0] node1870;
	wire [1-1:0] node1871;
	wire [1-1:0] node1873;
	wire [1-1:0] node1877;
	wire [1-1:0] node1878;
	wire [1-1:0] node1880;
	wire [1-1:0] node1883;
	wire [1-1:0] node1884;
	wire [1-1:0] node1888;
	wire [1-1:0] node1889;
	wire [1-1:0] node1891;
	wire [1-1:0] node1892;
	wire [1-1:0] node1894;
	wire [1-1:0] node1898;
	wire [1-1:0] node1899;
	wire [1-1:0] node1900;
	wire [1-1:0] node1902;
	wire [1-1:0] node1905;
	wire [1-1:0] node1906;
	wire [1-1:0] node1911;
	wire [1-1:0] node1912;
	wire [1-1:0] node1913;
	wire [1-1:0] node1915;
	wire [1-1:0] node1916;
	wire [1-1:0] node1918;
	wire [1-1:0] node1921;
	wire [1-1:0] node1922;
	wire [1-1:0] node1926;
	wire [1-1:0] node1927;
	wire [1-1:0] node1929;
	wire [1-1:0] node1930;
	wire [1-1:0] node1934;
	wire [1-1:0] node1935;
	wire [1-1:0] node1939;
	wire [1-1:0] node1940;
	wire [1-1:0] node1941;
	wire [1-1:0] node1942;
	wire [1-1:0] node1944;
	wire [1-1:0] node1947;
	wire [1-1:0] node1948;
	wire [1-1:0] node1953;
	wire [1-1:0] node1955;
	wire [1-1:0] node1956;
	wire [1-1:0] node1960;
	wire [1-1:0] node1961;
	wire [1-1:0] node1962;
	wire [1-1:0] node1963;
	wire [1-1:0] node1964;
	wire [1-1:0] node1966;
	wire [1-1:0] node1969;
	wire [1-1:0] node1970;
	wire [1-1:0] node1972;
	wire [1-1:0] node1975;
	wire [1-1:0] node1976;
	wire [1-1:0] node1980;
	wire [1-1:0] node1981;
	wire [1-1:0] node1982;
	wire [1-1:0] node1984;
	wire [1-1:0] node1987;
	wire [1-1:0] node1988;
	wire [1-1:0] node1992;
	wire [1-1:0] node1993;
	wire [1-1:0] node1994;
	wire [1-1:0] node1999;
	wire [1-1:0] node2000;
	wire [1-1:0] node2001;
	wire [1-1:0] node2002;
	wire [1-1:0] node2004;
	wire [1-1:0] node2007;
	wire [1-1:0] node2008;
	wire [1-1:0] node2012;
	wire [1-1:0] node2013;
	wire [1-1:0] node2017;
	wire [1-1:0] node2018;
	wire [1-1:0] node2019;
	wire [1-1:0] node2020;
	wire [1-1:0] node2026;
	wire [1-1:0] node2027;
	wire [1-1:0] node2028;
	wire [1-1:0] node2029;
	wire [1-1:0] node2035;
	wire [1-1:0] node2036;
	wire [1-1:0] node2037;
	wire [1-1:0] node2038;
	wire [1-1:0] node2039;
	wire [1-1:0] node2041;
	wire [1-1:0] node2042;
	wire [1-1:0] node2044;
	wire [1-1:0] node2046;
	wire [1-1:0] node2049;
	wire [1-1:0] node2050;
	wire [1-1:0] node2052;
	wire [1-1:0] node2056;
	wire [1-1:0] node2057;
	wire [1-1:0] node2058;
	wire [1-1:0] node2060;
	wire [1-1:0] node2062;
	wire [1-1:0] node2065;
	wire [1-1:0] node2066;
	wire [1-1:0] node2069;
	wire [1-1:0] node2070;
	wire [1-1:0] node2074;
	wire [1-1:0] node2075;
	wire [1-1:0] node2077;
	wire [1-1:0] node2078;
	wire [1-1:0] node2082;
	wire [1-1:0] node2083;
	wire [1-1:0] node2084;
	wire [1-1:0] node2089;
	wire [1-1:0] node2090;
	wire [1-1:0] node2091;
	wire [1-1:0] node2093;
	wire [1-1:0] node2094;
	wire [1-1:0] node2096;
	wire [1-1:0] node2099;
	wire [1-1:0] node2100;
	wire [1-1:0] node2104;
	wire [1-1:0] node2105;
	wire [1-1:0] node2107;
	wire [1-1:0] node2108;
	wire [1-1:0] node2112;
	wire [1-1:0] node2113;
	wire [1-1:0] node2114;
	wire [1-1:0] node2119;
	wire [1-1:0] node2120;
	wire [1-1:0] node2121;
	wire [1-1:0] node2122;
	wire [1-1:0] node2124;
	wire [1-1:0] node2130;
	wire [1-1:0] node2131;
	wire [1-1:0] node2132;
	wire [1-1:0] node2133;
	wire [1-1:0] node2134;
	wire [1-1:0] node2136;
	wire [1-1:0] node2138;
	wire [1-1:0] node2141;
	wire [1-1:0] node2142;
	wire [1-1:0] node2144;
	wire [1-1:0] node2147;
	wire [1-1:0] node2148;
	wire [1-1:0] node2152;
	wire [1-1:0] node2153;
	wire [1-1:0] node2154;
	wire [1-1:0] node2156;
	wire [1-1:0] node2159;
	wire [1-1:0] node2160;
	wire [1-1:0] node2164;
	wire [1-1:0] node2165;
	wire [1-1:0] node2169;
	wire [1-1:0] node2170;
	wire [1-1:0] node2171;
	wire [1-1:0] node2174;
	wire [1-1:0] node2175;
	wire [1-1:0] node2176;
	wire [1-1:0] node2181;
	wire [1-1:0] node2182;
	wire [1-1:0] node2183;
	wire [1-1:0] node2184;
	wire [1-1:0] node2190;
	wire [1-1:0] node2191;
	wire [1-1:0] node2192;
	wire [1-1:0] node2193;
	wire [1-1:0] node2194;
	wire [1-1:0] node2196;
	wire [1-1:0] node2199;
	wire [1-1:0] node2200;
	wire [1-1:0] node2204;
	wire [1-1:0] node2205;
	wire [1-1:0] node2206;
	wire [1-1:0] node2211;
	wire [1-1:0] node2212;
	wire [1-1:0] node2213;
	wire [1-1:0] node2219;
	wire [1-1:0] node2220;
	wire [1-1:0] node2221;
	wire [1-1:0] node2222;
	wire [1-1:0] node2223;
	wire [1-1:0] node2225;
	wire [1-1:0] node2226;
	wire [1-1:0] node2228;
	wire [1-1:0] node2232;
	wire [1-1:0] node2233;
	wire [1-1:0] node2234;
	wire [1-1:0] node2236;
	wire [1-1:0] node2239;
	wire [1-1:0] node2240;
	wire [1-1:0] node2245;
	wire [1-1:0] node2246;
	wire [1-1:0] node2247;
	wire [1-1:0] node2250;
	wire [1-1:0] node2251;
	wire [1-1:0] node2252;
	wire [1-1:0] node2257;
	wire [1-1:0] node2258;
	wire [1-1:0] node2259;
	wire [1-1:0] node2264;
	wire [1-1:0] node2265;
	wire [1-1:0] node2266;
	wire [1-1:0] node2267;
	wire [1-1:0] node2269;
	wire [1-1:0] node2270;
	wire [1-1:0] node2274;
	wire [1-1:0] node2275;
	wire [1-1:0] node2281;
	wire [1-1:0] node2282;
	wire [1-1:0] node2283;
	wire [1-1:0] node2284;
	wire [1-1:0] node2285;
	wire [1-1:0] node2286;
	wire [1-1:0] node2288;
	wire [1-1:0] node2291;
	wire [1-1:0] node2292;
	wire [1-1:0] node2296;
	wire [1-1:0] node2297;
	wire [1-1:0] node2301;
	wire [1-1:0] node2303;
	wire [1-1:0] node2304;
	wire [1-1:0] node2305;
	wire [1-1:0] node2310;
	wire [1-1:0] node2311;
	wire [1-1:0] node2312;
	wire [1-1:0] node2313;
	wire [1-1:0] node2314;
	wire [1-1:0] node2321;
	wire [1-1:0] node2322;
	wire [1-1:0] node2323;
	wire [1-1:0] node2324;
	wire [1-1:0] node2325;
	wire [1-1:0] node2332;
	wire [1-1:0] node2333;
	wire [1-1:0] node2334;
	wire [1-1:0] node2335;
	wire [1-1:0] node2336;
	wire [1-1:0] node2337;
	wire [1-1:0] node2339;
	wire [1-1:0] node2341;
	wire [1-1:0] node2342;
	wire [1-1:0] node2344;
	wire [1-1:0] node2346;
	wire [1-1:0] node2349;
	wire [1-1:0] node2350;
	wire [1-1:0] node2352;
	wire [1-1:0] node2354;
	wire [1-1:0] node2357;
	wire [1-1:0] node2358;
	wire [1-1:0] node2360;
	wire [1-1:0] node2364;
	wire [1-1:0] node2365;
	wire [1-1:0] node2367;
	wire [1-1:0] node2368;
	wire [1-1:0] node2370;
	wire [1-1:0] node2372;
	wire [1-1:0] node2375;
	wire [1-1:0] node2376;
	wire [1-1:0] node2378;
	wire [1-1:0] node2381;
	wire [1-1:0] node2382;
	wire [1-1:0] node2384;
	wire [1-1:0] node2388;
	wire [1-1:0] node2389;
	wire [1-1:0] node2391;
	wire [1-1:0] node2392;
	wire [1-1:0] node2394;
	wire [1-1:0] node2396;
	wire [1-1:0] node2399;
	wire [1-1:0] node2400;
	wire [1-1:0] node2404;
	wire [1-1:0] node2405;
	wire [1-1:0] node2407;
	wire [1-1:0] node2408;
	wire [1-1:0] node2410;
	wire [1-1:0] node2413;
	wire [1-1:0] node2414;
	wire [1-1:0] node2418;
	wire [1-1:0] node2419;
	wire [1-1:0] node2420;
	wire [1-1:0] node2422;
	wire [1-1:0] node2425;
	wire [1-1:0] node2426;
	wire [1-1:0] node2431;
	wire [1-1:0] node2432;
	wire [1-1:0] node2433;
	wire [1-1:0] node2435;
	wire [1-1:0] node2436;
	wire [1-1:0] node2438;
	wire [1-1:0] node2440;
	wire [1-1:0] node2442;
	wire [1-1:0] node2445;
	wire [1-1:0] node2447;
	wire [1-1:0] node2448;
	wire [1-1:0] node2450;
	wire [1-1:0] node2453;
	wire [1-1:0] node2454;
	wire [1-1:0] node2458;
	wire [1-1:0] node2459;
	wire [1-1:0] node2461;
	wire [1-1:0] node2462;
	wire [1-1:0] node2464;
	wire [1-1:0] node2466;
	wire [1-1:0] node2469;
	wire [1-1:0] node2470;
	wire [1-1:0] node2472;
	wire [1-1:0] node2475;
	wire [1-1:0] node2476;
	wire [1-1:0] node2480;
	wire [1-1:0] node2481;
	wire [1-1:0] node2483;
	wire [1-1:0] node2484;
	wire [1-1:0] node2486;
	wire [1-1:0] node2490;
	wire [1-1:0] node2491;
	wire [1-1:0] node2492;
	wire [1-1:0] node2494;
	wire [1-1:0] node2499;
	wire [1-1:0] node2500;
	wire [1-1:0] node2501;
	wire [1-1:0] node2502;
	wire [1-1:0] node2504;
	wire [1-1:0] node2506;
	wire [1-1:0] node2509;
	wire [1-1:0] node2510;
	wire [1-1:0] node2512;
	wire [1-1:0] node2515;
	wire [1-1:0] node2516;
	wire [1-1:0] node2518;
	wire [1-1:0] node2521;
	wire [1-1:0] node2522;
	wire [1-1:0] node2526;
	wire [1-1:0] node2527;
	wire [1-1:0] node2528;
	wire [1-1:0] node2529;
	wire [1-1:0] node2531;
	wire [1-1:0] node2535;
	wire [1-1:0] node2536;
	wire [1-1:0] node2538;
	wire [1-1:0] node2541;
	wire [1-1:0] node2543;
	wire [1-1:0] node2546;
	wire [1-1:0] node2547;
	wire [1-1:0] node2549;
	wire [1-1:0] node2550;
	wire [1-1:0] node2555;
	wire [1-1:0] node2556;
	wire [1-1:0] node2557;
	wire [1-1:0] node2559;
	wire [1-1:0] node2560;
	wire [1-1:0] node2562;
	wire [1-1:0] node2565;
	wire [1-1:0] node2566;
	wire [1-1:0] node2570;
	wire [1-1:0] node2571;
	wire [1-1:0] node2573;
	wire [1-1:0] node2574;
	wire [1-1:0] node2579;
	wire [1-1:0] node2580;
	wire [1-1:0] node2581;
	wire [1-1:0] node2582;
	wire [1-1:0] node2584;
	wire [1-1:0] node2587;
	wire [1-1:0] node2588;
	wire [1-1:0] node2594;
	wire [1-1:0] node2595;
	wire [1-1:0] node2596;
	wire [1-1:0] node2597;
	wire [1-1:0] node2599;
	wire [1-1:0] node2601;
	wire [1-1:0] node2603;
	wire [1-1:0] node2606;
	wire [1-1:0] node2607;
	wire [1-1:0] node2609;
	wire [1-1:0] node2610;
	wire [1-1:0] node2612;
	wire [1-1:0] node2614;
	wire [1-1:0] node2617;
	wire [1-1:0] node2618;
	wire [1-1:0] node2620;
	wire [1-1:0] node2623;
	wire [1-1:0] node2624;
	wire [1-1:0] node2628;
	wire [1-1:0] node2629;
	wire [1-1:0] node2630;
	wire [1-1:0] node2632;
	wire [1-1:0] node2634;
	wire [1-1:0] node2637;
	wire [1-1:0] node2638;
	wire [1-1:0] node2640;
	wire [1-1:0] node2643;
	wire [1-1:0] node2644;
	wire [1-1:0] node2648;
	wire [1-1:0] node2649;
	wire [1-1:0] node2650;
	wire [1-1:0] node2652;
	wire [1-1:0] node2655;
	wire [1-1:0] node2656;
	wire [1-1:0] node2661;
	wire [1-1:0] node2662;
	wire [1-1:0] node2663;
	wire [1-1:0] node2664;
	wire [1-1:0] node2666;
	wire [1-1:0] node2668;
	wire [1-1:0] node2670;
	wire [1-1:0] node2673;
	wire [1-1:0] node2674;
	wire [1-1:0] node2676;
	wire [1-1:0] node2679;
	wire [1-1:0] node2682;
	wire [1-1:0] node2683;
	wire [1-1:0] node2684;
	wire [1-1:0] node2686;
	wire [1-1:0] node2688;
	wire [1-1:0] node2691;
	wire [1-1:0] node2692;
	wire [1-1:0] node2694;
	wire [1-1:0] node2697;
	wire [1-1:0] node2698;
	wire [1-1:0] node2702;
	wire [1-1:0] node2703;
	wire [1-1:0] node2704;
	wire [1-1:0] node2706;
	wire [1-1:0] node2709;
	wire [1-1:0] node2710;
	wire [1-1:0] node2715;
	wire [1-1:0] node2716;
	wire [1-1:0] node2717;
	wire [1-1:0] node2719;
	wire [1-1:0] node2722;
	wire [1-1:0] node2723;
	wire [1-1:0] node2724;
	wire [1-1:0] node2726;
	wire [1-1:0] node2729;
	wire [1-1:0] node2730;
	wire [1-1:0] node2735;
	wire [1-1:0] node2736;
	wire [1-1:0] node2737;
	wire [1-1:0] node2738;
	wire [1-1:0] node2740;
	wire [1-1:0] node2743;
	wire [1-1:0] node2744;
	wire [1-1:0] node2750;
	wire [1-1:0] node2751;
	wire [1-1:0] node2752;
	wire [1-1:0] node2753;
	wire [1-1:0] node2755;
	wire [1-1:0] node2756;
	wire [1-1:0] node2758;
	wire [1-1:0] node2760;
	wire [1-1:0] node2763;
	wire [1-1:0] node2765;
	wire [1-1:0] node2766;
	wire [1-1:0] node2770;
	wire [1-1:0] node2771;
	wire [1-1:0] node2772;
	wire [1-1:0] node2774;
	wire [1-1:0] node2776;
	wire [1-1:0] node2779;
	wire [1-1:0] node2780;
	wire [1-1:0] node2782;
	wire [1-1:0] node2785;
	wire [1-1:0] node2786;
	wire [1-1:0] node2790;
	wire [1-1:0] node2791;
	wire [1-1:0] node2792;
	wire [1-1:0] node2794;
	wire [1-1:0] node2797;
	wire [1-1:0] node2798;
	wire [1-1:0] node2803;
	wire [1-1:0] node2804;
	wire [1-1:0] node2805;
	wire [1-1:0] node2807;
	wire [1-1:0] node2809;
	wire [1-1:0] node2810;
	wire [1-1:0] node2814;
	wire [1-1:0] node2815;
	wire [1-1:0] node2817;
	wire [1-1:0] node2818;
	wire [1-1:0] node2822;
	wire [1-1:0] node2823;
	wire [1-1:0] node2824;
	wire [1-1:0] node2829;
	wire [1-1:0] node2830;
	wire [1-1:0] node2831;
	wire [1-1:0] node2832;
	wire [1-1:0] node2834;
	wire [1-1:0] node2837;
	wire [1-1:0] node2838;
	wire [1-1:0] node2842;
	wire [1-1:0] node2843;
	wire [1-1:0] node2848;
	wire [1-1:0] node2849;
	wire [1-1:0] node2850;
	wire [1-1:0] node2851;
	wire [1-1:0] node2852;
	wire [1-1:0] node2854;
	wire [1-1:0] node2857;
	wire [1-1:0] node2858;
	wire [1-1:0] node2860;
	wire [1-1:0] node2864;
	wire [1-1:0] node2865;
	wire [1-1:0] node2867;
	wire [1-1:0] node2868;
	wire [1-1:0] node2872;
	wire [1-1:0] node2873;
	wire [1-1:0] node2874;
	wire [1-1:0] node2879;
	wire [1-1:0] node2880;
	wire [1-1:0] node2881;
	wire [1-1:0] node2882;
	wire [1-1:0] node2884;
	wire [1-1:0] node2888;
	wire [1-1:0] node2889;
	wire [1-1:0] node2890;
	wire [1-1:0] node2895;
	wire [1-1:0] node2896;
	wire [1-1:0] node2897;
	wire [1-1:0] node2902;
	wire [1-1:0] node2903;
	wire [1-1:0] node2904;
	wire [1-1:0] node2905;
	wire [1-1:0] node2907;
	wire [1-1:0] node2908;
	wire [1-1:0] node2913;
	wire [1-1:0] node2914;
	wire [1-1:0] node2915;
	wire [1-1:0] node2916;
	wire [1-1:0] node2923;
	wire [1-1:0] node2924;
	wire [1-1:0] node2925;
	wire [1-1:0] node2926;
	wire [1-1:0] node2927;
	wire [1-1:0] node2929;
	wire [1-1:0] node2930;
	wire [1-1:0] node2932;
	wire [1-1:0] node2934;
	wire [1-1:0] node2937;
	wire [1-1:0] node2938;
	wire [1-1:0] node2940;
	wire [1-1:0] node2943;
	wire [1-1:0] node2944;
	wire [1-1:0] node2948;
	wire [1-1:0] node2949;
	wire [1-1:0] node2950;
	wire [1-1:0] node2952;
	wire [1-1:0] node2954;
	wire [1-1:0] node2957;
	wire [1-1:0] node2959;
	wire [1-1:0] node2960;
	wire [1-1:0] node2963;
	wire [1-1:0] node2964;
	wire [1-1:0] node2968;
	wire [1-1:0] node2969;
	wire [1-1:0] node2971;
	wire [1-1:0] node2973;
	wire [1-1:0] node2974;
	wire [1-1:0] node2978;
	wire [1-1:0] node2979;
	wire [1-1:0] node2980;
	wire [1-1:0] node2982;
	wire [1-1:0] node2985;
	wire [1-1:0] node2986;
	wire [1-1:0] node2991;
	wire [1-1:0] node2992;
	wire [1-1:0] node2993;
	wire [1-1:0] node2995;
	wire [1-1:0] node2997;
	wire [1-1:0] node2998;
	wire [1-1:0] node3000;
	wire [1-1:0] node3003;
	wire [1-1:0] node3004;
	wire [1-1:0] node3008;
	wire [1-1:0] node3009;
	wire [1-1:0] node3011;
	wire [1-1:0] node3013;
	wire [1-1:0] node3015;
	wire [1-1:0] node3018;
	wire [1-1:0] node3019;
	wire [1-1:0] node3021;
	wire [1-1:0] node3025;
	wire [1-1:0] node3026;
	wire [1-1:0] node3027;
	wire [1-1:0] node3029;
	wire [1-1:0] node3031;
	wire [1-1:0] node3034;
	wire [1-1:0] node3035;
	wire [1-1:0] node3036;
	wire [1-1:0] node3038;
	wire [1-1:0] node3042;
	wire [1-1:0] node3043;
	wire [1-1:0] node3044;
	wire [1-1:0] node3049;
	wire [1-1:0] node3050;
	wire [1-1:0] node3051;
	wire [1-1:0] node3053;
	wire [1-1:0] node3054;
	wire [1-1:0] node3058;
	wire [1-1:0] node3059;
	wire [1-1:0] node3063;
	wire [1-1:0] node3064;
	wire [1-1:0] node3065;
	wire [1-1:0] node3070;
	wire [1-1:0] node3071;
	wire [1-1:0] node3072;
	wire [1-1:0] node3073;
	wire [1-1:0] node3074;
	wire [1-1:0] node3076;
	wire [1-1:0] node3078;
	wire [1-1:0] node3081;
	wire [1-1:0] node3083;
	wire [1-1:0] node3084;
	wire [1-1:0] node3086;
	wire [1-1:0] node3089;
	wire [1-1:0] node3090;
	wire [1-1:0] node3094;
	wire [1-1:0] node3095;
	wire [1-1:0] node3096;
	wire [1-1:0] node3098;
	wire [1-1:0] node3100;
	wire [1-1:0] node3103;
	wire [1-1:0] node3104;
	wire [1-1:0] node3106;
	wire [1-1:0] node3110;
	wire [1-1:0] node3111;
	wire [1-1:0] node3112;
	wire [1-1:0] node3114;
	wire [1-1:0] node3117;
	wire [1-1:0] node3118;
	wire [1-1:0] node3123;
	wire [1-1:0] node3124;
	wire [1-1:0] node3125;
	wire [1-1:0] node3127;
	wire [1-1:0] node3129;
	wire [1-1:0] node3130;
	wire [1-1:0] node3134;
	wire [1-1:0] node3135;
	wire [1-1:0] node3137;
	wire [1-1:0] node3138;
	wire [1-1:0] node3142;
	wire [1-1:0] node3143;
	wire [1-1:0] node3147;
	wire [1-1:0] node3148;
	wire [1-1:0] node3149;
	wire [1-1:0] node3150;
	wire [1-1:0] node3152;
	wire [1-1:0] node3155;
	wire [1-1:0] node3156;
	wire [1-1:0] node3160;
	wire [1-1:0] node3161;
	wire [1-1:0] node3162;
	wire [1-1:0] node3168;
	wire [1-1:0] node3169;
	wire [1-1:0] node3170;
	wire [1-1:0] node3171;
	wire [1-1:0] node3173;
	wire [1-1:0] node3176;
	wire [1-1:0] node3177;
	wire [1-1:0] node3179;
	wire [1-1:0] node3180;
	wire [1-1:0] node3184;
	wire [1-1:0] node3185;
	wire [1-1:0] node3186;
	wire [1-1:0] node3191;
	wire [1-1:0] node3192;
	wire [1-1:0] node3193;
	wire [1-1:0] node3195;
	wire [1-1:0] node3198;
	wire [1-1:0] node3199;
	wire [1-1:0] node3200;
	wire [1-1:0] node3205;
	wire [1-1:0] node3206;
	wire [1-1:0] node3207;
	wire [1-1:0] node3208;
	wire [1-1:0] node3214;
	wire [1-1:0] node3215;
	wire [1-1:0] node3216;
	wire [1-1:0] node3217;
	wire [1-1:0] node3219;
	wire [1-1:0] node3222;
	wire [1-1:0] node3223;
	wire [1-1:0] node3224;
	wire [1-1:0] node3231;
	wire [1-1:0] node3232;
	wire [1-1:0] node3233;
	wire [1-1:0] node3234;
	wire [1-1:0] node3235;
	wire [1-1:0] node3237;
	wire [1-1:0] node3239;
	wire [1-1:0] node3240;
	wire [1-1:0] node3242;
	wire [1-1:0] node3246;
	wire [1-1:0] node3247;
	wire [1-1:0] node3248;
	wire [1-1:0] node3250;
	wire [1-1:0] node3252;
	wire [1-1:0] node3255;
	wire [1-1:0] node3256;
	wire [1-1:0] node3258;
	wire [1-1:0] node3262;
	wire [1-1:0] node3263;
	wire [1-1:0] node3265;
	wire [1-1:0] node3268;
	wire [1-1:0] node3269;
	wire [1-1:0] node3271;
	wire [1-1:0] node3275;
	wire [1-1:0] node3276;
	wire [1-1:0] node3277;
	wire [1-1:0] node3279;
	wire [1-1:0] node3281;
	wire [1-1:0] node3284;
	wire [1-1:0] node3285;
	wire [1-1:0] node3287;
	wire [1-1:0] node3288;
	wire [1-1:0] node3292;
	wire [1-1:0] node3293;
	wire [1-1:0] node3294;
	wire [1-1:0] node3299;
	wire [1-1:0] node3300;
	wire [1-1:0] node3301;
	wire [1-1:0] node3303;
	wire [1-1:0] node3304;
	wire [1-1:0] node3308;
	wire [1-1:0] node3309;
	wire [1-1:0] node3310;
	wire [1-1:0] node3315;
	wire [1-1:0] node3316;
	wire [1-1:0] node3317;
	wire [1-1:0] node3318;
	wire [1-1:0] node3324;
	wire [1-1:0] node3325;
	wire [1-1:0] node3326;
	wire [1-1:0] node3327;
	wire [1-1:0] node3329;
	wire [1-1:0] node3331;
	wire [1-1:0] node3332;
	wire [1-1:0] node3336;
	wire [1-1:0] node3337;
	wire [1-1:0] node3339;
	wire [1-1:0] node3340;
	wire [1-1:0] node3344;
	wire [1-1:0] node3345;
	wire [1-1:0] node3346;
	wire [1-1:0] node3351;
	wire [1-1:0] node3352;
	wire [1-1:0] node3353;
	wire [1-1:0] node3355;
	wire [1-1:0] node3358;
	wire [1-1:0] node3359;
	wire [1-1:0] node3360;
	wire [1-1:0] node3365;
	wire [1-1:0] node3366;
	wire [1-1:0] node3367;
	wire [1-1:0] node3368;
	wire [1-1:0] node3374;
	wire [1-1:0] node3375;
	wire [1-1:0] node3376;
	wire [1-1:0] node3377;
	wire [1-1:0] node3378;
	wire [1-1:0] node3380;
	wire [1-1:0] node3383;
	wire [1-1:0] node3384;
	wire [1-1:0] node3388;
	wire [1-1:0] node3389;
	wire [1-1:0] node3393;
	wire [1-1:0] node3394;
	wire [1-1:0] node3395;
	wire [1-1:0] node3400;
	wire [1-1:0] node3401;
	wire [1-1:0] node3402;
	wire [1-1:0] node3403;
	wire [1-1:0] node3404;
	wire [1-1:0] node3411;
	wire [1-1:0] node3412;
	wire [1-1:0] node3413;
	wire [1-1:0] node3414;
	wire [1-1:0] node3415;
	wire [1-1:0] node3417;
	wire [1-1:0] node3418;
	wire [1-1:0] node3420;
	wire [1-1:0] node3423;
	wire [1-1:0] node3424;
	wire [1-1:0] node3428;
	wire [1-1:0] node3429;
	wire [1-1:0] node3430;
	wire [1-1:0] node3432;
	wire [1-1:0] node3435;
	wire [1-1:0] node3436;
	wire [1-1:0] node3440;
	wire [1-1:0] node3441;
	wire [1-1:0] node3445;
	wire [1-1:0] node3446;
	wire [1-1:0] node3447;
	wire [1-1:0] node3449;
	wire [1-1:0] node3450;
	wire [1-1:0] node3454;
	wire [1-1:0] node3455;
	wire [1-1:0] node3460;
	wire [1-1:0] node3461;
	wire [1-1:0] node3462;
	wire [1-1:0] node3463;
	wire [1-1:0] node3464;
	wire [1-1:0] node3466;
	wire [1-1:0] node3469;
	wire [1-1:0] node3470;
	wire [1-1:0] node3474;
	wire [1-1:0] node3475;
	wire [1-1:0] node3479;
	wire [1-1:0] node3480;
	wire [1-1:0] node3481;
	wire [1-1:0] node3486;
	wire [1-1:0] node3487;
	wire [1-1:0] node3488;
	wire [1-1:0] node3489;
	wire [1-1:0] node3490;
	wire [1-1:0] node3497;
	wire [1-1:0] node3498;
	wire [1-1:0] node3499;
	wire [1-1:0] node3500;
	wire [1-1:0] node3501;
	wire [1-1:0] node3502;
	wire [1-1:0] node3504;
	wire [1-1:0] node3507;
	wire [1-1:0] node3508;
	wire [1-1:0] node3512;
	wire [1-1:0] node3513;
	wire [1-1:0] node3514;
	wire [1-1:0] node3519;
	wire [1-1:0] node3520;
	wire [1-1:0] node3521;
	wire [1-1:0] node3522;
	wire [1-1:0] node3528;
	wire [1-1:0] node3529;
	wire [1-1:0] node3530;
	wire [1-1:0] node3531;
	wire [1-1:0] node3537;
	wire [1-1:0] node3538;
	wire [1-1:0] node3539;
	wire [1-1:0] node3540;
	wire [1-1:0] node3542;
	wire [1-1:0] node3548;
	wire [1-1:0] node3549;
	wire [1-1:0] node3550;
	wire [1-1:0] node3551;
	wire [1-1:0] node3552;
	wire [1-1:0] node3553;
	wire [1-1:0] node3555;
	wire [1-1:0] node3556;
	wire [1-1:0] node3558;
	wire [1-1:0] node3560;
	wire [1-1:0] node3562;
	wire [1-1:0] node3565;
	wire [1-1:0] node3566;
	wire [1-1:0] node3568;
	wire [1-1:0] node3570;
	wire [1-1:0] node3573;
	wire [1-1:0] node3574;
	wire [1-1:0] node3576;
	wire [1-1:0] node3579;
	wire [1-1:0] node3580;
	wire [1-1:0] node3584;
	wire [1-1:0] node3585;
	wire [1-1:0] node3586;
	wire [1-1:0] node3588;
	wire [1-1:0] node3589;
	wire [1-1:0] node3591;
	wire [1-1:0] node3595;
	wire [1-1:0] node3596;
	wire [1-1:0] node3598;
	wire [1-1:0] node3600;
	wire [1-1:0] node3603;
	wire [1-1:0] node3604;
	wire [1-1:0] node3606;
	wire [1-1:0] node3609;
	wire [1-1:0] node3610;
	wire [1-1:0] node3614;
	wire [1-1:0] node3615;
	wire [1-1:0] node3616;
	wire [1-1:0] node3618;
	wire [1-1:0] node3620;
	wire [1-1:0] node3623;
	wire [1-1:0] node3624;
	wire [1-1:0] node3626;
	wire [1-1:0] node3630;
	wire [1-1:0] node3631;
	wire [1-1:0] node3632;
	wire [1-1:0] node3634;
	wire [1-1:0] node3637;
	wire [1-1:0] node3638;
	wire [1-1:0] node3643;
	wire [1-1:0] node3644;
	wire [1-1:0] node3645;
	wire [1-1:0] node3647;
	wire [1-1:0] node3648;
	wire [1-1:0] node3650;
	wire [1-1:0] node3652;
	wire [1-1:0] node3655;
	wire [1-1:0] node3656;
	wire [1-1:0] node3658;
	wire [1-1:0] node3661;
	wire [1-1:0] node3664;
	wire [1-1:0] node3665;
	wire [1-1:0] node3667;
	wire [1-1:0] node3668;
	wire [1-1:0] node3671;
	wire [1-1:0] node3672;
	wire [1-1:0] node3676;
	wire [1-1:0] node3677;
	wire [1-1:0] node3681;
	wire [1-1:0] node3682;
	wire [1-1:0] node3683;
	wire [1-1:0] node3685;
	wire [1-1:0] node3686;
	wire [1-1:0] node3690;
	wire [1-1:0] node3691;
	wire [1-1:0] node3693;
	wire [1-1:0] node3694;
	wire [1-1:0] node3698;
	wire [1-1:0] node3699;
	wire [1-1:0] node3700;
	wire [1-1:0] node3705;
	wire [1-1:0] node3706;
	wire [1-1:0] node3707;
	wire [1-1:0] node3709;
	wire [1-1:0] node3710;
	wire [1-1:0] node3714;
	wire [1-1:0] node3715;
	wire [1-1:0] node3719;
	wire [1-1:0] node3720;
	wire [1-1:0] node3721;
	wire [1-1:0] node3722;
	wire [1-1:0] node3728;
	wire [1-1:0] node3729;
	wire [1-1:0] node3730;
	wire [1-1:0] node3731;
	wire [1-1:0] node3732;
	wire [1-1:0] node3734;
	wire [1-1:0] node3736;
	wire [1-1:0] node3737;
	wire [1-1:0] node3741;
	wire [1-1:0] node3742;
	wire [1-1:0] node3744;
	wire [1-1:0] node3746;
	wire [1-1:0] node3749;
	wire [1-1:0] node3750;
	wire [1-1:0] node3752;
	wire [1-1:0] node3756;
	wire [1-1:0] node3757;
	wire [1-1:0] node3759;
	wire [1-1:0] node3760;
	wire [1-1:0] node3762;
	wire [1-1:0] node3765;
	wire [1-1:0] node3767;
	wire [1-1:0] node3770;
	wire [1-1:0] node3771;
	wire [1-1:0] node3772;
	wire [1-1:0] node3774;
	wire [1-1:0] node3777;
	wire [1-1:0] node3778;
	wire [1-1:0] node3783;
	wire [1-1:0] node3784;
	wire [1-1:0] node3785;
	wire [1-1:0] node3787;
	wire [1-1:0] node3788;
	wire [1-1:0] node3790;
	wire [1-1:0] node3794;
	wire [1-1:0] node3795;
	wire [1-1:0] node3796;
	wire [1-1:0] node3798;
	wire [1-1:0] node3803;
	wire [1-1:0] node3804;
	wire [1-1:0] node3805;
	wire [1-1:0] node3806;
	wire [1-1:0] node3808;
	wire [1-1:0] node3811;
	wire [1-1:0] node3812;
	wire [1-1:0] node3816;
	wire [1-1:0] node3817;
	wire [1-1:0] node3818;
	wire [1-1:0] node3823;
	wire [1-1:0] node3824;
	wire [1-1:0] node3825;
	wire [1-1:0] node3826;
	wire [1-1:0] node3832;
	wire [1-1:0] node3833;
	wire [1-1:0] node3834;
	wire [1-1:0] node3835;
	wire [1-1:0] node3836;
	wire [1-1:0] node3838;
	wire [1-1:0] node3840;
	wire [1-1:0] node3843;
	wire [1-1:0] node3844;
	wire [1-1:0] node3847;
	wire [1-1:0] node3848;
	wire [1-1:0] node3852;
	wire [1-1:0] node3853;
	wire [1-1:0] node3856;
	wire [1-1:0] node3857;
	wire [1-1:0] node3861;
	wire [1-1:0] node3862;
	wire [1-1:0] node3863;
	wire [1-1:0] node3865;
	wire [1-1:0] node3866;
	wire [1-1:0] node3871;
	wire [1-1:0] node3872;
	wire [1-1:0] node3873;
	wire [1-1:0] node3874;
	wire [1-1:0] node3880;
	wire [1-1:0] node3881;
	wire [1-1:0] node3882;
	wire [1-1:0] node3883;
	wire [1-1:0] node3885;
	wire [1-1:0] node3886;
	wire [1-1:0] node3890;
	wire [1-1:0] node3891;
	wire [1-1:0] node3892;
	wire [1-1:0] node3897;
	wire [1-1:0] node3898;
	wire [1-1:0] node3899;
	wire [1-1:0] node3904;
	wire [1-1:0] node3905;
	wire [1-1:0] node3906;
	wire [1-1:0] node3907;
	wire [1-1:0] node3908;
	wire [1-1:0] node3915;
	wire [1-1:0] node3916;
	wire [1-1:0] node3917;
	wire [1-1:0] node3918;
	wire [1-1:0] node3919;
	wire [1-1:0] node3921;
	wire [1-1:0] node3922;
	wire [1-1:0] node3924;
	wire [1-1:0] node3926;
	wire [1-1:0] node3929;
	wire [1-1:0] node3930;
	wire [1-1:0] node3932;
	wire [1-1:0] node3936;
	wire [1-1:0] node3937;
	wire [1-1:0] node3939;
	wire [1-1:0] node3941;
	wire [1-1:0] node3942;
	wire [1-1:0] node3946;
	wire [1-1:0] node3947;
	wire [1-1:0] node3948;
	wire [1-1:0] node3950;
	wire [1-1:0] node3953;
	wire [1-1:0] node3954;
	wire [1-1:0] node3958;
	wire [1-1:0] node3959;
	wire [1-1:0] node3963;
	wire [1-1:0] node3964;
	wire [1-1:0] node3965;
	wire [1-1:0] node3967;
	wire [1-1:0] node3968;
	wire [1-1:0] node3970;
	wire [1-1:0] node3973;
	wire [1-1:0] node3974;
	wire [1-1:0] node3978;
	wire [1-1:0] node3979;
	wire [1-1:0] node3980;
	wire [1-1:0] node3982;
	wire [1-1:0] node3985;
	wire [1-1:0] node3986;
	wire [1-1:0] node3990;
	wire [1-1:0] node3992;
	wire [1-1:0] node3993;
	wire [1-1:0] node3997;
	wire [1-1:0] node3998;
	wire [1-1:0] node3999;
	wire [1-1:0] node4000;
	wire [1-1:0] node4002;
	wire [1-1:0] node4005;
	wire [1-1:0] node4006;
	wire [1-1:0] node4011;
	wire [1-1:0] node4012;
	wire [1-1:0] node4013;
	wire [1-1:0] node4018;
	wire [1-1:0] node4019;
	wire [1-1:0] node4020;
	wire [1-1:0] node4021;
	wire [1-1:0] node4023;
	wire [1-1:0] node4024;
	wire [1-1:0] node4026;
	wire [1-1:0] node4029;
	wire [1-1:0] node4030;
	wire [1-1:0] node4034;
	wire [1-1:0] node4035;
	wire [1-1:0] node4036;
	wire [1-1:0] node4038;
	wire [1-1:0] node4041;
	wire [1-1:0] node4042;
	wire [1-1:0] node4046;
	wire [1-1:0] node4047;
	wire [1-1:0] node4051;
	wire [1-1:0] node4052;
	wire [1-1:0] node4053;
	wire [1-1:0] node4055;
	wire [1-1:0] node4058;
	wire [1-1:0] node4059;
	wire [1-1:0] node4064;
	wire [1-1:0] node4065;
	wire [1-1:0] node4066;
	wire [1-1:0] node4067;
	wire [1-1:0] node4069;
	wire [1-1:0] node4070;
	wire [1-1:0] node4074;
	wire [1-1:0] node4075;
	wire [1-1:0] node4077;
	wire [1-1:0] node4082;
	wire [1-1:0] node4083;
	wire [1-1:0] node4084;
	wire [1-1:0] node4085;
	wire [1-1:0] node4086;
	wire [1-1:0] node4093;
	wire [1-1:0] node4094;
	wire [1-1:0] node4095;
	wire [1-1:0] node4096;
	wire [1-1:0] node4097;
	wire [1-1:0] node4099;
	wire [1-1:0] node4100;
	wire [1-1:0] node4102;
	wire [1-1:0] node4105;
	wire [1-1:0] node4106;
	wire [1-1:0] node4110;
	wire [1-1:0] node4111;
	wire [1-1:0] node4112;
	wire [1-1:0] node4114;
	wire [1-1:0] node4117;
	wire [1-1:0] node4118;
	wire [1-1:0] node4122;
	wire [1-1:0] node4123;
	wire [1-1:0] node4124;
	wire [1-1:0] node4129;
	wire [1-1:0] node4130;
	wire [1-1:0] node4131;
	wire [1-1:0] node4132;
	wire [1-1:0] node4134;
	wire [1-1:0] node4137;
	wire [1-1:0] node4138;
	wire [1-1:0] node4142;
	wire [1-1:0] node4143;
	wire [1-1:0] node4148;
	wire [1-1:0] node4149;
	wire [1-1:0] node4150;
	wire [1-1:0] node4151;
	wire [1-1:0] node4152;
	wire [1-1:0] node4154;
	wire [1-1:0] node4157;
	wire [1-1:0] node4158;
	wire [1-1:0] node4162;
	wire [1-1:0] node4163;
	wire [1-1:0] node4164;
	wire [1-1:0] node4169;
	wire [1-1:0] node4170;
	wire [1-1:0] node4171;
	wire [1-1:0] node4177;
	wire [1-1:0] node4178;
	wire [1-1:0] node4179;
	wire [1-1:0] node4180;
	wire [1-1:0] node4181;
	wire [1-1:0] node4183;
	wire [1-1:0] node4184;
	wire [1-1:0] node4188;
	wire [1-1:0] node4189;
	wire [1-1:0] node4190;
	wire [1-1:0] node4195;
	wire [1-1:0] node4196;
	wire [1-1:0] node4197;
	wire [1-1:0] node4198;
	wire [1-1:0] node4204;
	wire [1-1:0] node4205;
	wire [1-1:0] node4206;
	wire [1-1:0] node4212;
	wire [1-1:0] node4213;
	wire [1-1:0] node4214;
	wire [1-1:0] node4215;
	wire [1-1:0] node4216;
	wire [1-1:0] node4217;
	wire [1-1:0] node4219;
	wire [1-1:0] node4221;
	wire [1-1:0] node4222;
	wire [1-1:0] node4224;
	wire [1-1:0] node4227;
	wire [1-1:0] node4230;
	wire [1-1:0] node4231;
	wire [1-1:0] node4233;
	wire [1-1:0] node4236;
	wire [1-1:0] node4237;
	wire [1-1:0] node4238;
	wire [1-1:0] node4240;
	wire [1-1:0] node4243;
	wire [1-1:0] node4244;
	wire [1-1:0] node4249;
	wire [1-1:0] node4250;
	wire [1-1:0] node4251;
	wire [1-1:0] node4253;
	wire [1-1:0] node4255;
	wire [1-1:0] node4258;
	wire [1-1:0] node4259;
	wire [1-1:0] node4261;
	wire [1-1:0] node4263;
	wire [1-1:0] node4266;
	wire [1-1:0] node4269;
	wire [1-1:0] node4270;
	wire [1-1:0] node4271;
	wire [1-1:0] node4273;
	wire [1-1:0] node4276;
	wire [1-1:0] node4277;
	wire [1-1:0] node4278;
	wire [1-1:0] node4284;
	wire [1-1:0] node4285;
	wire [1-1:0] node4286;
	wire [1-1:0] node4287;
	wire [1-1:0] node4288;
	wire [1-1:0] node4290;
	wire [1-1:0] node4292;
	wire [1-1:0] node4295;
	wire [1-1:0] node4296;
	wire [1-1:0] node4298;
	wire [1-1:0] node4302;
	wire [1-1:0] node4303;
	wire [1-1:0] node4305;
	wire [1-1:0] node4306;
	wire [1-1:0] node4310;
	wire [1-1:0] node4311;
	wire [1-1:0] node4312;
	wire [1-1:0] node4317;
	wire [1-1:0] node4318;
	wire [1-1:0] node4319;
	wire [1-1:0] node4320;
	wire [1-1:0] node4322;
	wire [1-1:0] node4325;
	wire [1-1:0] node4328;
	wire [1-1:0] node4329;
	wire [1-1:0] node4334;
	wire [1-1:0] node4335;
	wire [1-1:0] node4336;
	wire [1-1:0] node4337;
	wire [1-1:0] node4338;
	wire [1-1:0] node4340;
	wire [1-1:0] node4343;
	wire [1-1:0] node4344;
	wire [1-1:0] node4348;
	wire [1-1:0] node4349;
	wire [1-1:0] node4355;
	wire [1-1:0] node4356;
	wire [1-1:0] node4357;
	wire [1-1:0] node4358;
	wire [1-1:0] node4359;
	wire [1-1:0] node4361;
	wire [1-1:0] node4362;
	wire [1-1:0] node4364;
	wire [1-1:0] node4367;
	wire [1-1:0] node4368;
	wire [1-1:0] node4372;
	wire [1-1:0] node4373;
	wire [1-1:0] node4375;
	wire [1-1:0] node4376;
	wire [1-1:0] node4381;
	wire [1-1:0] node4382;
	wire [1-1:0] node4383;
	wire [1-1:0] node4384;
	wire [1-1:0] node4386;
	wire [1-1:0] node4389;
	wire [1-1:0] node4390;
	wire [1-1:0] node4394;
	wire [1-1:0] node4395;
	wire [1-1:0] node4397;
	wire [1-1:0] node4402;
	wire [1-1:0] node4403;
	wire [1-1:0] node4404;
	wire [1-1:0] node4405;
	wire [1-1:0] node4407;
	wire [1-1:0] node4408;
	wire [1-1:0] node4412;
	wire [1-1:0] node4413;
	wire [1-1:0] node4414;
	wire [1-1:0] node4419;
	wire [1-1:0] node4420;
	wire [1-1:0] node4421;
	wire [1-1:0] node4427;
	wire [1-1:0] node4428;
	wire [1-1:0] node4429;
	wire [1-1:0] node4430;
	wire [1-1:0] node4431;
	wire [1-1:0] node4433;
	wire [1-1:0] node4434;
	wire [1-1:0] node4438;
	wire [1-1:0] node4439;
	wire [1-1:0] node4440;
	wire [1-1:0] node4445;
	wire [1-1:0] node4446;
	wire [1-1:0] node4447;
	wire [1-1:0] node4454;
	wire [1-1:0] node4455;
	wire [1-1:0] node4456;
	wire [1-1:0] node4457;
	wire [1-1:0] node4458;
	wire [1-1:0] node4459;
	wire [1-1:0] node4461;
	wire [1-1:0] node4463;
	wire [1-1:0] node4466;
	wire [1-1:0] node4467;
	wire [1-1:0] node4469;
	wire [1-1:0] node4472;
	wire [1-1:0] node4473;
	wire [1-1:0] node4474;
	wire [1-1:0] node4479;
	wire [1-1:0] node4480;
	wire [1-1:0] node4481;
	wire [1-1:0] node4483;
	wire [1-1:0] node4486;
	wire [1-1:0] node4487;
	wire [1-1:0] node4491;
	wire [1-1:0] node4492;
	wire [1-1:0] node4493;
	wire [1-1:0] node4498;
	wire [1-1:0] node4499;
	wire [1-1:0] node4500;
	wire [1-1:0] node4501;
	wire [1-1:0] node4502;
	wire [1-1:0] node4504;
	wire [1-1:0] node4507;
	wire [1-1:0] node4508;
	wire [1-1:0] node4512;
	wire [1-1:0] node4513;
	wire [1-1:0] node4514;
	wire [1-1:0] node4519;
	wire [1-1:0] node4520;
	wire [1-1:0] node4521;
	wire [1-1:0] node4522;
	wire [1-1:0] node4528;
	wire [1-1:0] node4529;
	wire [1-1:0] node4530;
	wire [1-1:0] node4531;
	wire [1-1:0] node4537;
	wire [1-1:0] node4538;
	wire [1-1:0] node4539;
	wire [1-1:0] node4540;
	wire [1-1:0] node4541;
	wire [1-1:0] node4543;
	wire [1-1:0] node4546;
	wire [1-1:0] node4547;
	wire [1-1:0] node4548;
	wire [1-1:0] node4553;
	wire [1-1:0] node4554;
	wire [1-1:0] node4555;
	wire [1-1:0] node4560;
	wire [1-1:0] node4561;
	wire [1-1:0] node4562;
	wire [1-1:0] node4563;
	wire [1-1:0] node4570;
	wire [1-1:0] node4571;
	wire [1-1:0] node4572;
	wire [1-1:0] node4573;
	wire [1-1:0] node4574;
	wire [1-1:0] node4575;
	wire [1-1:0] node4577;
	wire [1-1:0] node4578;
	wire [1-1:0] node4583;
	wire [1-1:0] node4584;
	wire [1-1:0] node4585;
	wire [1-1:0] node4590;
	wire [1-1:0] node4591;
	wire [1-1:0] node4592;
	wire [1-1:0] node4593;
	wire [1-1:0] node4599;
	wire [1-1:0] node4600;
	wire [1-1:0] node4602;
	wire [1-1:0] node4603;
	wire [1-1:0] node4604;
	wire [1-1:0] node4610;
	wire [1-1:0] node4611;
	wire [1-1:0] node4612;
	wire [1-1:0] node4613;
	wire [1-1:0] node4614;
	wire [1-1:0] node4615;
	wire [1-1:0] node4616;

	assign outp = (inp[2]) ? node2332 : node1;
		assign node1 = (inp[6]) ? node1115 : node2;
			assign node2 = (inp[9]) ? node476 : node3;
				assign node3 = (inp[12]) ? node181 : node4;
					assign node4 = (inp[3]) ? node44 : node5;
						assign node5 = (inp[10]) ? node7 : 1'b1;
							assign node7 = (inp[0]) ? node19 : node8;
								assign node8 = (inp[8]) ? node10 : 1'b1;
									assign node10 = (inp[4]) ? node12 : 1'b1;
										assign node12 = (inp[7]) ? node14 : 1'b1;
											assign node14 = (inp[11]) ? node16 : 1'b1;
												assign node16 = (inp[5]) ? 1'b0 : 1'b1;
								assign node19 = (inp[7]) ? node29 : node20;
									assign node20 = (inp[1]) ? node22 : 1'b1;
										assign node22 = (inp[13]) ? node24 : 1'b1;
											assign node24 = (inp[14]) ? node26 : 1'b1;
												assign node26 = (inp[8]) ? 1'b0 : 1'b1;
									assign node29 = (inp[13]) ? node31 : 1'b1;
										assign node31 = (inp[5]) ? node37 : node32;
											assign node32 = (inp[14]) ? node34 : 1'b1;
												assign node34 = (inp[4]) ? 1'b0 : 1'b1;
											assign node37 = (inp[8]) ? node39 : 1'b1;
												assign node39 = (inp[11]) ? 1'b0 : node40;
													assign node40 = (inp[1]) ? 1'b0 : 1'b0;
						assign node44 = (inp[4]) ? node94 : node45;
							assign node45 = (inp[1]) ? node59 : node46;
								assign node46 = (inp[7]) ? node48 : 1'b1;
									assign node48 = (inp[0]) ? node50 : 1'b1;
										assign node50 = (inp[13]) ? node52 : 1'b1;
											assign node52 = (inp[5]) ? node54 : 1'b1;
												assign node54 = (inp[10]) ? node56 : 1'b1;
													assign node56 = (inp[14]) ? 1'b0 : 1'b1;
								assign node59 = (inp[14]) ? node69 : node60;
									assign node60 = (inp[7]) ? node62 : 1'b1;
										assign node62 = (inp[5]) ? node64 : 1'b1;
											assign node64 = (inp[11]) ? node66 : 1'b1;
												assign node66 = (inp[10]) ? 1'b0 : 1'b1;
									assign node69 = (inp[8]) ? node79 : node70;
										assign node70 = (inp[7]) ? 1'b1 : node71;
											assign node71 = (inp[11]) ? node73 : 1'b1;
												assign node73 = (inp[13]) ? node75 : 1'b1;
													assign node75 = (inp[0]) ? 1'b0 : 1'b1;
										assign node79 = (inp[7]) ? node87 : node80;
											assign node80 = (inp[10]) ? node82 : 1'b1;
												assign node82 = (inp[11]) ? 1'b0 : node83;
													assign node83 = (inp[13]) ? 1'b1 : 1'b1;
											assign node87 = (inp[0]) ? 1'b0 : node88;
												assign node88 = (inp[5]) ? node90 : 1'b1;
													assign node90 = (inp[11]) ? 1'b0 : 1'b1;
							assign node94 = (inp[14]) ? node130 : node95;
								assign node95 = (inp[5]) ? node105 : node96;
									assign node96 = (inp[1]) ? node98 : 1'b1;
										assign node98 = (inp[10]) ? node100 : 1'b1;
											assign node100 = (inp[11]) ? node102 : 1'b1;
												assign node102 = (inp[13]) ? 1'b0 : 1'b1;
									assign node105 = (inp[8]) ? node115 : node106;
										assign node106 = (inp[0]) ? node108 : 1'b1;
											assign node108 = (inp[1]) ? node110 : 1'b1;
												assign node110 = (inp[11]) ? node112 : 1'b1;
													assign node112 = (inp[10]) ? 1'b0 : 1'b1;
										assign node115 = (inp[10]) ? node123 : node116;
											assign node116 = (inp[1]) ? node118 : 1'b1;
												assign node118 = (inp[11]) ? node120 : 1'b1;
													assign node120 = (inp[7]) ? 1'b0 : 1'b1;
											assign node123 = (inp[13]) ? 1'b0 : node124;
												assign node124 = (inp[11]) ? node126 : 1'b1;
													assign node126 = (inp[1]) ? 1'b0 : 1'b1;
								assign node130 = (inp[1]) ? node158 : node131;
									assign node131 = (inp[0]) ? node139 : node132;
										assign node132 = (inp[10]) ? node134 : 1'b1;
											assign node134 = (inp[5]) ? node136 : 1'b1;
												assign node136 = (inp[11]) ? 1'b0 : 1'b1;
										assign node139 = (inp[13]) ? node147 : node140;
											assign node140 = (inp[5]) ? node142 : 1'b1;
												assign node142 = (inp[7]) ? node144 : 1'b1;
													assign node144 = (inp[8]) ? 1'b0 : 1'b1;
											assign node147 = (inp[7]) ? node153 : node148;
												assign node148 = (inp[8]) ? 1'b0 : node149;
													assign node149 = (inp[11]) ? 1'b1 : 1'b1;
												assign node153 = (inp[11]) ? 1'b0 : node154;
													assign node154 = (inp[10]) ? 1'b0 : 1'b1;
									assign node158 = (inp[10]) ? node168 : node159;
										assign node159 = (inp[0]) ? node161 : 1'b1;
											assign node161 = (inp[13]) ? 1'b0 : node162;
												assign node162 = (inp[7]) ? node164 : 1'b1;
													assign node164 = (inp[5]) ? 1'b0 : 1'b1;
										assign node168 = (inp[11]) ? 1'b0 : node169;
											assign node169 = (inp[5]) ? node175 : node170;
												assign node170 = (inp[0]) ? node172 : 1'b1;
													assign node172 = (inp[13]) ? 1'b0 : 1'b1;
												assign node175 = (inp[7]) ? 1'b0 : node176;
													assign node176 = (inp[8]) ? 1'b0 : 1'b1;
					assign node181 = (inp[14]) ? node313 : node182;
						assign node182 = (inp[10]) ? node224 : node183;
							assign node183 = (inp[7]) ? node185 : 1'b1;
								assign node185 = (inp[3]) ? node197 : node186;
									assign node186 = (inp[4]) ? node188 : 1'b1;
										assign node188 = (inp[8]) ? node190 : 1'b1;
											assign node190 = (inp[0]) ? node192 : 1'b1;
												assign node192 = (inp[11]) ? node194 : 1'b1;
													assign node194 = (inp[13]) ? 1'b0 : 1'b1;
									assign node197 = (inp[0]) ? node205 : node198;
										assign node198 = (inp[4]) ? node200 : 1'b1;
											assign node200 = (inp[8]) ? node202 : 1'b1;
												assign node202 = (inp[1]) ? 1'b0 : 1'b1;
										assign node205 = (inp[1]) ? node213 : node206;
											assign node206 = (inp[13]) ? node208 : 1'b1;
												assign node208 = (inp[8]) ? 1'b0 : node209;
													assign node209 = (inp[5]) ? 1'b0 : 1'b1;
											assign node213 = (inp[8]) ? node219 : node214;
												assign node214 = (inp[5]) ? node216 : 1'b1;
													assign node216 = (inp[13]) ? 1'b0 : 1'b0;
												assign node219 = (inp[4]) ? 1'b0 : node220;
													assign node220 = (inp[5]) ? 1'b0 : 1'b0;
							assign node224 = (inp[4]) ? node260 : node225;
								assign node225 = (inp[1]) ? node237 : node226;
									assign node226 = (inp[13]) ? node228 : 1'b1;
										assign node228 = (inp[3]) ? 1'b1 : node229;
											assign node229 = (inp[11]) ? node231 : 1'b1;
												assign node231 = (inp[0]) ? node233 : 1'b1;
													assign node233 = (inp[8]) ? 1'b0 : 1'b1;
									assign node237 = (inp[7]) ? node245 : node238;
										assign node238 = (inp[0]) ? node240 : 1'b1;
											assign node240 = (inp[11]) ? node242 : 1'b1;
												assign node242 = (inp[13]) ? 1'b0 : 1'b1;
										assign node245 = (inp[3]) ? node253 : node246;
											assign node246 = (inp[8]) ? node248 : 1'b1;
												assign node248 = (inp[13]) ? node250 : 1'b1;
													assign node250 = (inp[11]) ? 1'b0 : 1'b1;
											assign node253 = (inp[5]) ? 1'b0 : node254;
												assign node254 = (inp[8]) ? node256 : 1'b1;
													assign node256 = (inp[0]) ? 1'b0 : 1'b1;
								assign node260 = (inp[8]) ? node286 : node261;
									assign node261 = (inp[13]) ? node269 : node262;
										assign node262 = (inp[11]) ? node264 : 1'b1;
											assign node264 = (inp[0]) ? node266 : 1'b1;
												assign node266 = (inp[1]) ? 1'b0 : 1'b1;
										assign node269 = (inp[1]) ? node275 : node270;
											assign node270 = (inp[5]) ? node272 : 1'b1;
												assign node272 = (inp[3]) ? 1'b0 : 1'b1;
											assign node275 = (inp[5]) ? node281 : node276;
												assign node276 = (inp[11]) ? node278 : 1'b1;
													assign node278 = (inp[7]) ? 1'b0 : 1'b1;
												assign node281 = (inp[3]) ? 1'b0 : node282;
													assign node282 = (inp[11]) ? 1'b0 : 1'b1;
									assign node286 = (inp[11]) ? node304 : node287;
										assign node287 = (inp[7]) ? node297 : node288;
											assign node288 = (inp[1]) ? node294 : node289;
												assign node289 = (inp[5]) ? node291 : 1'b1;
													assign node291 = (inp[0]) ? 1'b1 : 1'b1;
												assign node294 = (inp[5]) ? 1'b0 : 1'b1;
											assign node297 = (inp[3]) ? node299 : 1'b1;
												assign node299 = (inp[13]) ? 1'b0 : node300;
													assign node300 = (inp[5]) ? 1'b0 : 1'b1;
										assign node304 = (inp[5]) ? 1'b0 : node305;
											assign node305 = (inp[13]) ? node307 : 1'b1;
												assign node307 = (inp[3]) ? 1'b0 : node308;
													assign node308 = (inp[7]) ? 1'b0 : 1'b1;
						assign node313 = (inp[5]) ? node387 : node314;
							assign node314 = (inp[8]) ? node336 : node315;
								assign node315 = (inp[7]) ? node317 : 1'b1;
									assign node317 = (inp[3]) ? node319 : 1'b1;
										assign node319 = (inp[4]) ? node327 : node320;
											assign node320 = (inp[13]) ? node322 : 1'b1;
												assign node322 = (inp[10]) ? 1'b0 : node323;
													assign node323 = (inp[0]) ? 1'b0 : 1'b1;
											assign node327 = (inp[11]) ? node331 : node328;
												assign node328 = (inp[0]) ? 1'b0 : 1'b1;
												assign node331 = (inp[13]) ? 1'b0 : node332;
													assign node332 = (inp[1]) ? 1'b0 : 1'b1;
								assign node336 = (inp[1]) ? node360 : node337;
									assign node337 = (inp[11]) ? node345 : node338;
										assign node338 = (inp[0]) ? node340 : 1'b1;
											assign node340 = (inp[3]) ? node342 : 1'b1;
												assign node342 = (inp[10]) ? 1'b0 : 1'b1;
										assign node345 = (inp[13]) ? node351 : node346;
											assign node346 = (inp[7]) ? node348 : 1'b1;
												assign node348 = (inp[3]) ? 1'b1 : 1'b0;
											assign node351 = (inp[4]) ? node355 : node352;
												assign node352 = (inp[7]) ? 1'b0 : 1'b1;
												assign node355 = (inp[10]) ? 1'b0 : node356;
													assign node356 = (inp[3]) ? 1'b0 : 1'b0;
									assign node360 = (inp[4]) ? node376 : node361;
										assign node361 = (inp[10]) ? node367 : node362;
											assign node362 = (inp[3]) ? node364 : 1'b1;
												assign node364 = (inp[13]) ? 1'b0 : 1'b1;
											assign node367 = (inp[7]) ? node371 : node368;
												assign node368 = (inp[11]) ? 1'b0 : 1'b1;
												assign node371 = (inp[13]) ? 1'b0 : node372;
													assign node372 = (inp[0]) ? 1'b0 : 1'b1;
										assign node376 = (inp[3]) ? 1'b0 : node377;
											assign node377 = (inp[13]) ? node383 : node378;
												assign node378 = (inp[10]) ? node380 : 1'b1;
													assign node380 = (inp[0]) ? 1'b0 : 1'b1;
												assign node383 = (inp[11]) ? 1'b0 : 1'b1;
							assign node387 = (inp[11]) ? node435 : node388;
								assign node388 = (inp[7]) ? node408 : node389;
									assign node389 = (inp[4]) ? node391 : 1'b1;
										assign node391 = (inp[13]) ? node397 : node392;
											assign node392 = (inp[1]) ? node394 : 1'b1;
												assign node394 = (inp[0]) ? 1'b0 : 1'b1;
											assign node397 = (inp[10]) ? node403 : node398;
												assign node398 = (inp[0]) ? node400 : 1'b1;
													assign node400 = (inp[3]) ? 1'b0 : 1'b1;
												assign node403 = (inp[3]) ? 1'b0 : node404;
													assign node404 = (inp[8]) ? 1'b0 : 1'b1;
									assign node408 = (inp[1]) ? node422 : node409;
										assign node409 = (inp[8]) ? node415 : node410;
											assign node410 = (inp[4]) ? node412 : 1'b1;
												assign node412 = (inp[13]) ? 1'b0 : 1'b1;
											assign node415 = (inp[3]) ? node417 : 1'b1;
												assign node417 = (inp[10]) ? 1'b0 : node418;
													assign node418 = (inp[13]) ? 1'b0 : 1'b1;
										assign node422 = (inp[8]) ? 1'b0 : node423;
											assign node423 = (inp[0]) ? node429 : node424;
												assign node424 = (inp[10]) ? node426 : 1'b1;
													assign node426 = (inp[13]) ? 1'b0 : 1'b1;
												assign node429 = (inp[3]) ? 1'b0 : node430;
													assign node430 = (inp[4]) ? 1'b0 : 1'b1;
								assign node435 = (inp[4]) ? node459 : node436;
									assign node436 = (inp[0]) ? node444 : node437;
										assign node437 = (inp[3]) ? node439 : 1'b1;
											assign node439 = (inp[1]) ? 1'b0 : node440;
												assign node440 = (inp[10]) ? 1'b0 : 1'b1;
										assign node444 = (inp[10]) ? node452 : node445;
											assign node445 = (inp[3]) ? node447 : 1'b1;
												assign node447 = (inp[1]) ? 1'b0 : node448;
													assign node448 = (inp[8]) ? 1'b0 : 1'b1;
											assign node452 = (inp[13]) ? 1'b0 : node453;
												assign node453 = (inp[7]) ? 1'b0 : node454;
													assign node454 = (inp[8]) ? 1'b0 : 1'b1;
									assign node459 = (inp[8]) ? 1'b0 : node460;
										assign node460 = (inp[13]) ? node470 : node461;
											assign node461 = (inp[7]) ? node467 : node462;
												assign node462 = (inp[10]) ? node464 : 1'b1;
													assign node464 = (inp[1]) ? 1'b0 : 1'b1;
												assign node467 = (inp[0]) ? 1'b0 : 1'b1;
											assign node470 = (inp[0]) ? 1'b0 : node471;
												assign node471 = (inp[3]) ? 1'b0 : 1'b1;
				assign node476 = (inp[7]) ? node744 : node477;
					assign node477 = (inp[1]) ? node581 : node478;
						assign node478 = (inp[14]) ? node526 : node479;
							assign node479 = (inp[5]) ? node491 : node480;
								assign node480 = (inp[3]) ? node482 : 1'b1;
									assign node482 = (inp[12]) ? node484 : 1'b1;
										assign node484 = (inp[0]) ? node486 : 1'b1;
											assign node486 = (inp[4]) ? node488 : 1'b1;
												assign node488 = (inp[10]) ? 1'b0 : 1'b1;
								assign node491 = (inp[10]) ? node503 : node492;
									assign node492 = (inp[4]) ? node494 : 1'b1;
										assign node494 = (inp[3]) ? node496 : 1'b1;
											assign node496 = (inp[12]) ? node498 : 1'b1;
												assign node498 = (inp[0]) ? node500 : 1'b1;
													assign node500 = (inp[13]) ? 1'b0 : 1'b1;
									assign node503 = (inp[12]) ? node511 : node504;
										assign node504 = (inp[3]) ? node506 : 1'b1;
											assign node506 = (inp[13]) ? node508 : 1'b1;
												assign node508 = (inp[0]) ? 1'b0 : 1'b1;
										assign node511 = (inp[11]) ? node519 : node512;
											assign node512 = (inp[13]) ? node514 : 1'b1;
												assign node514 = (inp[8]) ? node516 : 1'b1;
													assign node516 = (inp[3]) ? 1'b0 : 1'b0;
											assign node519 = (inp[3]) ? node523 : node520;
												assign node520 = (inp[13]) ? 1'b0 : 1'b1;
												assign node523 = (inp[4]) ? 1'b0 : 1'b1;
							assign node526 = (inp[12]) ? node540 : node527;
								assign node527 = (inp[11]) ? node529 : 1'b1;
									assign node529 = (inp[8]) ? node531 : 1'b1;
										assign node531 = (inp[4]) ? node537 : node532;
											assign node532 = (inp[3]) ? node534 : 1'b1;
												assign node534 = (inp[13]) ? 1'b0 : 1'b1;
											assign node537 = (inp[0]) ? 1'b0 : 1'b1;
								assign node540 = (inp[4]) ? node560 : node541;
									assign node541 = (inp[8]) ? node549 : node542;
										assign node542 = (inp[0]) ? node544 : 1'b1;
											assign node544 = (inp[10]) ? 1'b1 : node545;
												assign node545 = (inp[13]) ? 1'b0 : 1'b1;
										assign node549 = (inp[13]) ? node555 : node550;
											assign node550 = (inp[3]) ? node552 : 1'b1;
												assign node552 = (inp[10]) ? 1'b1 : 1'b0;
											assign node555 = (inp[10]) ? 1'b0 : node556;
												assign node556 = (inp[3]) ? 1'b0 : 1'b1;
									assign node560 = (inp[11]) ? node572 : node561;
										assign node561 = (inp[8]) ? node569 : node562;
											assign node562 = (inp[13]) ? node564 : 1'b1;
												assign node564 = (inp[5]) ? node566 : 1'b1;
													assign node566 = (inp[0]) ? 1'b0 : 1'b1;
											assign node569 = (inp[10]) ? 1'b0 : 1'b1;
										assign node572 = (inp[13]) ? 1'b0 : node573;
											assign node573 = (inp[5]) ? node575 : 1'b1;
												assign node575 = (inp[3]) ? 1'b0 : node576;
													assign node576 = (inp[10]) ? 1'b0 : 1'b1;
						assign node581 = (inp[10]) ? node657 : node582;
							assign node582 = (inp[13]) ? node614 : node583;
								assign node583 = (inp[5]) ? node585 : 1'b1;
									assign node585 = (inp[8]) ? node595 : node586;
										assign node586 = (inp[0]) ? node588 : 1'b1;
											assign node588 = (inp[4]) ? node590 : 1'b1;
												assign node590 = (inp[11]) ? 1'b0 : node591;
													assign node591 = (inp[14]) ? 1'b1 : 1'b1;
										assign node595 = (inp[11]) ? node603 : node596;
											assign node596 = (inp[12]) ? node598 : 1'b1;
												assign node598 = (inp[4]) ? node600 : 1'b1;
													assign node600 = (inp[14]) ? 1'b0 : 1'b1;
											assign node603 = (inp[0]) ? node609 : node604;
												assign node604 = (inp[3]) ? node606 : 1'b1;
													assign node606 = (inp[14]) ? 1'b0 : 1'b1;
												assign node609 = (inp[3]) ? 1'b0 : node610;
													assign node610 = (inp[4]) ? 1'b0 : 1'b1;
								assign node614 = (inp[3]) ? node638 : node615;
									assign node615 = (inp[5]) ? node625 : node616;
										assign node616 = (inp[4]) ? node618 : 1'b1;
											assign node618 = (inp[11]) ? node620 : 1'b1;
												assign node620 = (inp[12]) ? node622 : 1'b1;
													assign node622 = (inp[14]) ? 1'b1 : 1'b0;
										assign node625 = (inp[12]) ? node633 : node626;
											assign node626 = (inp[11]) ? node628 : 1'b1;
												assign node628 = (inp[0]) ? node630 : 1'b1;
													assign node630 = (inp[4]) ? 1'b0 : 1'b1;
											assign node633 = (inp[8]) ? 1'b0 : node634;
												assign node634 = (inp[0]) ? 1'b0 : 1'b1;
									assign node638 = (inp[0]) ? node648 : node639;
										assign node639 = (inp[14]) ? node641 : 1'b1;
											assign node641 = (inp[8]) ? node643 : 1'b1;
												assign node643 = (inp[12]) ? 1'b0 : node644;
													assign node644 = (inp[5]) ? 1'b0 : 1'b1;
										assign node648 = (inp[11]) ? 1'b0 : node649;
											assign node649 = (inp[8]) ? 1'b0 : node650;
												assign node650 = (inp[4]) ? node652 : 1'b1;
													assign node652 = (inp[12]) ? 1'b0 : 1'b1;
							assign node657 = (inp[4]) ? node715 : node658;
								assign node658 = (inp[14]) ? node688 : node659;
									assign node659 = (inp[3]) ? node669 : node660;
										assign node660 = (inp[8]) ? node662 : 1'b1;
											assign node662 = (inp[13]) ? node664 : 1'b1;
												assign node664 = (inp[5]) ? node666 : 1'b1;
													assign node666 = (inp[0]) ? 1'b0 : 1'b1;
										assign node669 = (inp[11]) ? node677 : node670;
											assign node670 = (inp[13]) ? node672 : 1'b1;
												assign node672 = (inp[0]) ? node674 : 1'b1;
													assign node674 = (inp[5]) ? 1'b0 : 1'b1;
											assign node677 = (inp[8]) ? node683 : node678;
												assign node678 = (inp[13]) ? node680 : 1'b1;
													assign node680 = (inp[0]) ? 1'b0 : 1'b1;
												assign node683 = (inp[5]) ? 1'b0 : node684;
													assign node684 = (inp[12]) ? 1'b0 : 1'b1;
									assign node688 = (inp[8]) ? node706 : node689;
										assign node689 = (inp[13]) ? node695 : node690;
											assign node690 = (inp[12]) ? node692 : 1'b1;
												assign node692 = (inp[3]) ? 1'b0 : 1'b1;
											assign node695 = (inp[3]) ? node701 : node696;
												assign node696 = (inp[0]) ? node698 : 1'b1;
													assign node698 = (inp[12]) ? 1'b0 : 1'b1;
												assign node701 = (inp[12]) ? 1'b0 : node702;
													assign node702 = (inp[11]) ? 1'b0 : 1'b1;
										assign node706 = (inp[12]) ? 1'b0 : node707;
											assign node707 = (inp[3]) ? 1'b0 : node708;
												assign node708 = (inp[13]) ? node710 : 1'b1;
													assign node710 = (inp[5]) ? 1'b0 : 1'b1;
								assign node715 = (inp[14]) ? node735 : node716;
									assign node716 = (inp[11]) ? node726 : node717;
										assign node717 = (inp[8]) ? node719 : 1'b1;
											assign node719 = (inp[12]) ? 1'b0 : node720;
												assign node720 = (inp[5]) ? node722 : 1'b1;
													assign node722 = (inp[13]) ? 1'b0 : 1'b1;
										assign node726 = (inp[0]) ? 1'b0 : node727;
											assign node727 = (inp[5]) ? 1'b0 : node728;
												assign node728 = (inp[8]) ? node730 : 1'b1;
													assign node730 = (inp[3]) ? 1'b0 : 1'b1;
									assign node735 = (inp[8]) ? 1'b0 : node736;
										assign node736 = (inp[11]) ? 1'b0 : node737;
											assign node737 = (inp[3]) ? node739 : 1'b1;
												assign node739 = (inp[12]) ? 1'b0 : 1'b1;
					assign node744 = (inp[8]) ? node936 : node745;
						assign node745 = (inp[11]) ? node839 : node746;
							assign node746 = (inp[5]) ? node784 : node747;
								assign node747 = (inp[4]) ? node755 : node748;
									assign node748 = (inp[0]) ? node750 : 1'b1;
										assign node750 = (inp[14]) ? node752 : 1'b1;
											assign node752 = (inp[13]) ? 1'b0 : 1'b1;
									assign node755 = (inp[10]) ? node765 : node756;
										assign node756 = (inp[14]) ? node758 : 1'b1;
											assign node758 = (inp[12]) ? node760 : 1'b1;
												assign node760 = (inp[13]) ? node762 : 1'b1;
													assign node762 = (inp[1]) ? 1'b0 : 1'b1;
										assign node765 = (inp[13]) ? node773 : node766;
											assign node766 = (inp[0]) ? node768 : 1'b1;
												assign node768 = (inp[14]) ? node770 : 1'b1;
													assign node770 = (inp[3]) ? 1'b0 : 1'b1;
											assign node773 = (inp[12]) ? node779 : node774;
												assign node774 = (inp[1]) ? node776 : 1'b1;
													assign node776 = (inp[14]) ? 1'b0 : 1'b1;
												assign node779 = (inp[0]) ? 1'b0 : node780;
													assign node780 = (inp[14]) ? 1'b0 : 1'b1;
								assign node784 = (inp[3]) ? node812 : node785;
									assign node785 = (inp[12]) ? node793 : node786;
										assign node786 = (inp[13]) ? 1'b1 : node787;
											assign node787 = (inp[14]) ? node789 : 1'b1;
												assign node789 = (inp[0]) ? 1'b0 : 1'b1;
										assign node793 = (inp[13]) ? node801 : node794;
											assign node794 = (inp[0]) ? node796 : 1'b1;
												assign node796 = (inp[14]) ? node798 : 1'b1;
													assign node798 = (inp[10]) ? 1'b0 : 1'b1;
											assign node801 = (inp[4]) ? node807 : node802;
												assign node802 = (inp[14]) ? 1'b1 : node803;
													assign node803 = (inp[0]) ? 1'b0 : 1'b1;
												assign node807 = (inp[1]) ? 1'b0 : node808;
													assign node808 = (inp[10]) ? 1'b0 : 1'b1;
									assign node812 = (inp[1]) ? node826 : node813;
										assign node813 = (inp[10]) ? node815 : 1'b1;
											assign node815 = (inp[14]) ? node821 : node816;
												assign node816 = (inp[13]) ? node818 : 1'b1;
													assign node818 = (inp[4]) ? 1'b0 : 1'b1;
												assign node821 = (inp[13]) ? 1'b0 : node822;
													assign node822 = (inp[4]) ? 1'b0 : 1'b1;
										assign node826 = (inp[12]) ? 1'b0 : node827;
											assign node827 = (inp[0]) ? node833 : node828;
												assign node828 = (inp[13]) ? node830 : 1'b1;
													assign node830 = (inp[14]) ? 1'b0 : 1'b1;
												assign node833 = (inp[14]) ? 1'b0 : node834;
													assign node834 = (inp[10]) ? 1'b0 : 1'b1;
							assign node839 = (inp[12]) ? node887 : node840;
								assign node840 = (inp[14]) ? node862 : node841;
									assign node841 = (inp[1]) ? node849 : node842;
										assign node842 = (inp[13]) ? node844 : 1'b1;
											assign node844 = (inp[4]) ? node846 : 1'b1;
												assign node846 = (inp[5]) ? 1'b0 : 1'b1;
										assign node849 = (inp[0]) ? node855 : node850;
											assign node850 = (inp[4]) ? node852 : 1'b1;
												assign node852 = (inp[3]) ? 1'b0 : 1'b1;
											assign node855 = (inp[3]) ? 1'b0 : node856;
												assign node856 = (inp[10]) ? node858 : 1'b1;
													assign node858 = (inp[5]) ? 1'b0 : 1'b1;
									assign node862 = (inp[0]) ? node878 : node863;
										assign node863 = (inp[13]) ? node871 : node864;
											assign node864 = (inp[5]) ? node866 : 1'b1;
												assign node866 = (inp[4]) ? node868 : 1'b1;
													assign node868 = (inp[1]) ? 1'b0 : 1'b1;
											assign node871 = (inp[5]) ? 1'b0 : node872;
												assign node872 = (inp[1]) ? node874 : 1'b1;
													assign node874 = (inp[3]) ? 1'b0 : 1'b0;
										assign node878 = (inp[1]) ? 1'b0 : node879;
											assign node879 = (inp[13]) ? node881 : 1'b1;
												assign node881 = (inp[10]) ? 1'b0 : node882;
													assign node882 = (inp[5]) ? 1'b0 : 1'b0;
								assign node887 = (inp[10]) ? node917 : node888;
									assign node888 = (inp[4]) ? node908 : node889;
										assign node889 = (inp[1]) ? node897 : node890;
											assign node890 = (inp[3]) ? node892 : 1'b1;
												assign node892 = (inp[5]) ? node894 : 1'b1;
													assign node894 = (inp[0]) ? 1'b0 : 1'b1;
											assign node897 = (inp[14]) ? node903 : node898;
												assign node898 = (inp[3]) ? node900 : 1'b1;
													assign node900 = (inp[5]) ? 1'b0 : 1'b1;
												assign node903 = (inp[0]) ? 1'b0 : node904;
													assign node904 = (inp[5]) ? 1'b0 : 1'b1;
										assign node908 = (inp[5]) ? 1'b0 : node909;
											assign node909 = (inp[0]) ? 1'b0 : node910;
												assign node910 = (inp[13]) ? node912 : 1'b1;
													assign node912 = (inp[1]) ? 1'b0 : 1'b1;
									assign node917 = (inp[3]) ? node929 : node918;
										assign node918 = (inp[1]) ? node922 : node919;
											assign node919 = (inp[5]) ? 1'b0 : 1'b1;
											assign node922 = (inp[0]) ? 1'b0 : node923;
												assign node923 = (inp[4]) ? 1'b0 : node924;
													assign node924 = (inp[14]) ? 1'b0 : 1'b0;
										assign node929 = (inp[5]) ? 1'b0 : node930;
											assign node930 = (inp[0]) ? 1'b0 : node931;
												assign node931 = (inp[14]) ? 1'b0 : 1'b1;
						assign node936 = (inp[10]) ? node1042 : node937;
							assign node937 = (inp[3]) ? node993 : node938;
								assign node938 = (inp[4]) ? node964 : node939;
									assign node939 = (inp[11]) ? node947 : node940;
										assign node940 = (inp[14]) ? node942 : 1'b1;
											assign node942 = (inp[13]) ? node944 : 1'b1;
												assign node944 = (inp[12]) ? 1'b0 : 1'b1;
										assign node947 = (inp[5]) ? node953 : node948;
											assign node948 = (inp[1]) ? node950 : 1'b1;
												assign node950 = (inp[13]) ? 1'b0 : 1'b1;
											assign node953 = (inp[0]) ? node959 : node954;
												assign node954 = (inp[13]) ? node956 : 1'b1;
													assign node956 = (inp[14]) ? 1'b0 : 1'b1;
												assign node959 = (inp[12]) ? 1'b0 : node960;
													assign node960 = (inp[14]) ? 1'b0 : 1'b1;
									assign node964 = (inp[0]) ? node984 : node965;
										assign node965 = (inp[13]) ? node973 : node966;
											assign node966 = (inp[1]) ? node968 : 1'b1;
												assign node968 = (inp[12]) ? node970 : 1'b1;
													assign node970 = (inp[14]) ? 1'b0 : 1'b1;
											assign node973 = (inp[12]) ? node979 : node974;
												assign node974 = (inp[5]) ? 1'b1 : node975;
													assign node975 = (inp[1]) ? 1'b0 : 1'b1;
												assign node979 = (inp[11]) ? 1'b0 : node980;
													assign node980 = (inp[1]) ? 1'b0 : 1'b1;
										assign node984 = (inp[14]) ? 1'b0 : node985;
											assign node985 = (inp[5]) ? node987 : 1'b1;
												assign node987 = (inp[11]) ? 1'b0 : node988;
													assign node988 = (inp[13]) ? 1'b0 : 1'b1;
								assign node993 = (inp[11]) ? node1025 : node994;
									assign node994 = (inp[14]) ? node1008 : node995;
										assign node995 = (inp[5]) ? node997 : 1'b1;
											assign node997 = (inp[0]) ? node1003 : node998;
												assign node998 = (inp[13]) ? node1000 : 1'b1;
													assign node1000 = (inp[4]) ? 1'b0 : 1'b1;
												assign node1003 = (inp[13]) ? 1'b0 : node1004;
													assign node1004 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1008 = (inp[1]) ? node1020 : node1009;
											assign node1009 = (inp[0]) ? node1015 : node1010;
												assign node1010 = (inp[5]) ? node1012 : 1'b1;
													assign node1012 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1015 = (inp[12]) ? 1'b0 : node1016;
													assign node1016 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1020 = (inp[13]) ? 1'b0 : node1021;
												assign node1021 = (inp[12]) ? 1'b0 : 1'b1;
									assign node1025 = (inp[1]) ? 1'b0 : node1026;
										assign node1026 = (inp[0]) ? node1034 : node1027;
											assign node1027 = (inp[12]) ? node1029 : 1'b1;
												assign node1029 = (inp[13]) ? 1'b0 : node1030;
													assign node1030 = (inp[5]) ? 1'b0 : 1'b1;
											assign node1034 = (inp[14]) ? 1'b0 : node1035;
												assign node1035 = (inp[13]) ? 1'b0 : node1036;
													assign node1036 = (inp[5]) ? 1'b0 : 1'b1;
							assign node1042 = (inp[0]) ? node1090 : node1043;
								assign node1043 = (inp[13]) ? node1073 : node1044;
									assign node1044 = (inp[1]) ? node1058 : node1045;
										assign node1045 = (inp[14]) ? node1047 : 1'b1;
											assign node1047 = (inp[4]) ? node1053 : node1048;
												assign node1048 = (inp[3]) ? node1050 : 1'b1;
													assign node1050 = (inp[5]) ? 1'b0 : 1'b1;
												assign node1053 = (inp[11]) ? 1'b0 : node1054;
													assign node1054 = (inp[5]) ? 1'b0 : 1'b1;
										assign node1058 = (inp[12]) ? node1066 : node1059;
											assign node1059 = (inp[3]) ? node1061 : 1'b1;
												assign node1061 = (inp[5]) ? 1'b0 : node1062;
													assign node1062 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1066 = (inp[11]) ? 1'b0 : node1067;
												assign node1067 = (inp[4]) ? 1'b0 : node1068;
													assign node1068 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1073 = (inp[3]) ? 1'b0 : node1074;
										assign node1074 = (inp[1]) ? node1082 : node1075;
											assign node1075 = (inp[14]) ? node1077 : 1'b1;
												assign node1077 = (inp[4]) ? 1'b0 : node1078;
													assign node1078 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1082 = (inp[12]) ? 1'b0 : node1083;
												assign node1083 = (inp[4]) ? 1'b0 : node1084;
													assign node1084 = (inp[5]) ? 1'b0 : 1'b1;
								assign node1090 = (inp[14]) ? node1104 : node1091;
									assign node1091 = (inp[1]) ? 1'b0 : node1092;
										assign node1092 = (inp[3]) ? node1096 : node1093;
											assign node1093 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1096 = (inp[13]) ? 1'b0 : node1097;
												assign node1097 = (inp[12]) ? 1'b0 : node1098;
													assign node1098 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1104 = (inp[1]) ? node1106 : 1'b0;
										assign node1106 = (inp[11]) ? 1'b0 : node1107;
											assign node1107 = (inp[3]) ? 1'b0 : node1108;
												assign node1108 = (inp[5]) ? 1'b0 : node1109;
													assign node1109 = (inp[4]) ? 1'b0 : 1'b0;
			assign node1115 = (inp[0]) ? node1713 : node1116;
				assign node1116 = (inp[5]) ? node1386 : node1117;
					assign node1117 = (inp[10]) ? node1215 : node1118;
						assign node1118 = (inp[4]) ? node1160 : node1119;
							assign node1119 = (inp[12]) ? node1121 : 1'b1;
								assign node1121 = (inp[13]) ? node1133 : node1122;
									assign node1122 = (inp[11]) ? 1'b1 : node1123;
										assign node1123 = (inp[7]) ? node1125 : 1'b1;
											assign node1125 = (inp[1]) ? node1127 : 1'b1;
												assign node1127 = (inp[14]) ? node1129 : 1'b1;
													assign node1129 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1133 = (inp[7]) ? node1141 : node1134;
										assign node1134 = (inp[3]) ? node1136 : 1'b1;
											assign node1136 = (inp[8]) ? node1138 : 1'b1;
												assign node1138 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1141 = (inp[14]) ? node1149 : node1142;
											assign node1142 = (inp[3]) ? node1144 : 1'b1;
												assign node1144 = (inp[9]) ? node1146 : 1'b1;
													assign node1146 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1149 = (inp[1]) ? node1155 : node1150;
												assign node1150 = (inp[11]) ? node1152 : 1'b1;
													assign node1152 = (inp[8]) ? 1'b0 : 1'b1;
												assign node1155 = (inp[3]) ? 1'b0 : node1156;
													assign node1156 = (inp[8]) ? 1'b0 : 1'b1;
							assign node1160 = (inp[11]) ? node1178 : node1161;
								assign node1161 = (inp[7]) ? node1163 : 1'b1;
									assign node1163 = (inp[1]) ? node1165 : 1'b1;
										assign node1165 = (inp[8]) ? node1173 : node1166;
											assign node1166 = (inp[9]) ? node1168 : 1'b1;
												assign node1168 = (inp[13]) ? node1170 : 1'b1;
													assign node1170 = (inp[14]) ? 1'b0 : 1'b0;
											assign node1173 = (inp[12]) ? 1'b0 : node1174;
												assign node1174 = (inp[13]) ? 1'b0 : 1'b1;
								assign node1178 = (inp[1]) ? node1198 : node1179;
									assign node1179 = (inp[8]) ? node1181 : 1'b1;
										assign node1181 = (inp[12]) ? node1187 : node1182;
											assign node1182 = (inp[3]) ? node1184 : 1'b1;
												assign node1184 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1187 = (inp[7]) ? node1193 : node1188;
												assign node1188 = (inp[3]) ? node1190 : 1'b1;
													assign node1190 = (inp[14]) ? 1'b0 : 1'b1;
												assign node1193 = (inp[13]) ? 1'b0 : node1194;
													assign node1194 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1198 = (inp[14]) ? node1208 : node1199;
										assign node1199 = (inp[7]) ? node1201 : 1'b1;
											assign node1201 = (inp[9]) ? 1'b0 : node1202;
												assign node1202 = (inp[13]) ? node1204 : 1'b1;
													assign node1204 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1208 = (inp[8]) ? 1'b0 : node1209;
											assign node1209 = (inp[9]) ? 1'b0 : node1210;
												assign node1210 = (inp[3]) ? 1'b0 : 1'b1;
						assign node1215 = (inp[12]) ? node1297 : node1216;
							assign node1216 = (inp[3]) ? node1254 : node1217;
								assign node1217 = (inp[1]) ? node1227 : node1218;
									assign node1218 = (inp[8]) ? node1220 : 1'b1;
										assign node1220 = (inp[13]) ? node1222 : 1'b1;
											assign node1222 = (inp[4]) ? node1224 : 1'b1;
												assign node1224 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1227 = (inp[4]) ? node1237 : node1228;
										assign node1228 = (inp[14]) ? node1230 : 1'b1;
											assign node1230 = (inp[11]) ? node1232 : 1'b1;
												assign node1232 = (inp[7]) ? node1234 : 1'b1;
													assign node1234 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1237 = (inp[11]) ? node1245 : node1238;
											assign node1238 = (inp[8]) ? node1240 : 1'b1;
												assign node1240 = (inp[9]) ? node1242 : 1'b1;
													assign node1242 = (inp[13]) ? 1'b0 : 1'b1;
											assign node1245 = (inp[13]) ? node1249 : node1246;
												assign node1246 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1249 = (inp[7]) ? 1'b0 : node1250;
													assign node1250 = (inp[8]) ? 1'b0 : 1'b1;
								assign node1254 = (inp[13]) ? node1276 : node1255;
									assign node1255 = (inp[11]) ? node1257 : 1'b1;
										assign node1257 = (inp[9]) ? node1263 : node1258;
											assign node1258 = (inp[4]) ? 1'b1 : node1259;
												assign node1259 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1263 = (inp[4]) ? node1269 : node1264;
												assign node1264 = (inp[7]) ? node1266 : 1'b1;
													assign node1266 = (inp[14]) ? 1'b0 : 1'b1;
												assign node1269 = (inp[1]) ? node1273 : node1270;
													assign node1270 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1273 = (inp[7]) ? 1'b0 : 1'b0;
									assign node1276 = (inp[8]) ? node1288 : node1277;
										assign node1277 = (inp[11]) ? node1279 : 1'b1;
											assign node1279 = (inp[4]) ? node1283 : node1280;
												assign node1280 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1283 = (inp[1]) ? 1'b0 : node1284;
													assign node1284 = (inp[14]) ? 1'b0 : 1'b0;
										assign node1288 = (inp[14]) ? 1'b0 : node1289;
											assign node1289 = (inp[4]) ? node1291 : 1'b1;
												assign node1291 = (inp[1]) ? 1'b0 : node1292;
													assign node1292 = (inp[9]) ? 1'b0 : 1'b1;
							assign node1297 = (inp[14]) ? node1347 : node1298;
								assign node1298 = (inp[9]) ? node1324 : node1299;
									assign node1299 = (inp[4]) ? node1309 : node1300;
										assign node1300 = (inp[13]) ? node1302 : 1'b1;
											assign node1302 = (inp[1]) ? node1304 : 1'b1;
												assign node1304 = (inp[7]) ? 1'b0 : node1305;
													assign node1305 = (inp[3]) ? 1'b1 : 1'b1;
										assign node1309 = (inp[11]) ? node1315 : node1310;
											assign node1310 = (inp[3]) ? node1312 : 1'b1;
												assign node1312 = (inp[13]) ? 1'b0 : 1'b1;
											assign node1315 = (inp[8]) ? node1319 : node1316;
												assign node1316 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1319 = (inp[7]) ? 1'b0 : node1320;
													assign node1320 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1324 = (inp[7]) ? node1338 : node1325;
										assign node1325 = (inp[8]) ? node1327 : 1'b1;
											assign node1327 = (inp[3]) ? node1333 : node1328;
												assign node1328 = (inp[4]) ? node1330 : 1'b1;
													assign node1330 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1333 = (inp[11]) ? 1'b0 : node1334;
													assign node1334 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1338 = (inp[1]) ? 1'b0 : node1339;
											assign node1339 = (inp[13]) ? 1'b0 : node1340;
												assign node1340 = (inp[11]) ? node1342 : 1'b1;
													assign node1342 = (inp[3]) ? 1'b0 : 1'b1;
								assign node1347 = (inp[3]) ? node1377 : node1348;
									assign node1348 = (inp[1]) ? node1368 : node1349;
										assign node1349 = (inp[9]) ? node1357 : node1350;
											assign node1350 = (inp[7]) ? node1352 : 1'b1;
												assign node1352 = (inp[13]) ? node1354 : 1'b1;
													assign node1354 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1357 = (inp[8]) ? node1363 : node1358;
												assign node1358 = (inp[13]) ? 1'b0 : node1359;
													assign node1359 = (inp[11]) ? 1'b1 : 1'b1;
												assign node1363 = (inp[11]) ? 1'b0 : node1364;
													assign node1364 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1368 = (inp[7]) ? 1'b0 : node1369;
											assign node1369 = (inp[9]) ? node1371 : 1'b1;
												assign node1371 = (inp[4]) ? 1'b0 : node1372;
													assign node1372 = (inp[13]) ? 1'b0 : 1'b1;
									assign node1377 = (inp[7]) ? 1'b0 : node1378;
										assign node1378 = (inp[11]) ? 1'b0 : node1379;
											assign node1379 = (inp[1]) ? node1381 : 1'b1;
												assign node1381 = (inp[4]) ? 1'b0 : 1'b1;
					assign node1386 = (inp[11]) ? node1546 : node1387;
						assign node1387 = (inp[8]) ? node1449 : node1388;
							assign node1388 = (inp[10]) ? node1408 : node1389;
								assign node1389 = (inp[12]) ? node1391 : 1'b1;
									assign node1391 = (inp[13]) ? node1393 : 1'b1;
										assign node1393 = (inp[9]) ? node1401 : node1394;
											assign node1394 = (inp[4]) ? node1396 : 1'b1;
												assign node1396 = (inp[1]) ? node1398 : 1'b1;
													assign node1398 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1401 = (inp[7]) ? 1'b0 : node1402;
												assign node1402 = (inp[14]) ? node1404 : 1'b1;
													assign node1404 = (inp[4]) ? 1'b0 : 1'b1;
								assign node1408 = (inp[7]) ? node1424 : node1409;
									assign node1409 = (inp[3]) ? node1411 : 1'b1;
										assign node1411 = (inp[1]) ? node1417 : node1412;
											assign node1412 = (inp[4]) ? node1414 : 1'b1;
												assign node1414 = (inp[9]) ? 1'b0 : 1'b1;
											assign node1417 = (inp[13]) ? 1'b0 : node1418;
												assign node1418 = (inp[12]) ? node1420 : 1'b1;
													assign node1420 = (inp[4]) ? 1'b0 : 1'b1;
									assign node1424 = (inp[4]) ? node1440 : node1425;
										assign node1425 = (inp[13]) ? node1433 : node1426;
											assign node1426 = (inp[9]) ? node1428 : 1'b1;
												assign node1428 = (inp[1]) ? node1430 : 1'b1;
													assign node1430 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1433 = (inp[9]) ? 1'b0 : node1434;
												assign node1434 = (inp[1]) ? node1436 : 1'b1;
													assign node1436 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1440 = (inp[14]) ? 1'b0 : node1441;
											assign node1441 = (inp[12]) ? node1443 : 1'b1;
												assign node1443 = (inp[1]) ? 1'b0 : node1444;
													assign node1444 = (inp[9]) ? 1'b0 : 1'b1;
							assign node1449 = (inp[4]) ? node1507 : node1450;
								assign node1450 = (inp[7]) ? node1478 : node1451;
									assign node1451 = (inp[3]) ? node1459 : node1452;
										assign node1452 = (inp[12]) ? node1454 : 1'b1;
											assign node1454 = (inp[9]) ? node1456 : 1'b1;
												assign node1456 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1459 = (inp[14]) ? node1467 : node1460;
											assign node1460 = (inp[12]) ? 1'b1 : node1461;
												assign node1461 = (inp[1]) ? node1463 : 1'b1;
													assign node1463 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1467 = (inp[1]) ? node1473 : node1468;
												assign node1468 = (inp[9]) ? node1470 : 1'b1;
													assign node1470 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1473 = (inp[12]) ? 1'b0 : node1474;
													assign node1474 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1478 = (inp[13]) ? node1492 : node1479;
										assign node1479 = (inp[10]) ? node1481 : 1'b1;
											assign node1481 = (inp[14]) ? node1487 : node1482;
												assign node1482 = (inp[3]) ? node1484 : 1'b1;
													assign node1484 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1487 = (inp[1]) ? 1'b0 : node1488;
													assign node1488 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1492 = (inp[9]) ? node1502 : node1493;
											assign node1493 = (inp[14]) ? node1499 : node1494;
												assign node1494 = (inp[1]) ? node1496 : 1'b1;
													assign node1496 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1499 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1502 = (inp[10]) ? 1'b0 : node1503;
												assign node1503 = (inp[3]) ? 1'b0 : 1'b1;
								assign node1507 = (inp[1]) ? node1531 : node1508;
									assign node1508 = (inp[12]) ? node1518 : node1509;
										assign node1509 = (inp[7]) ? node1511 : 1'b1;
											assign node1511 = (inp[9]) ? 1'b0 : node1512;
												assign node1512 = (inp[13]) ? node1514 : 1'b1;
													assign node1514 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1518 = (inp[9]) ? 1'b0 : node1519;
											assign node1519 = (inp[10]) ? node1525 : node1520;
												assign node1520 = (inp[3]) ? node1522 : 1'b1;
													assign node1522 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1525 = (inp[7]) ? 1'b0 : node1526;
													assign node1526 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1531 = (inp[10]) ? 1'b0 : node1532;
										assign node1532 = (inp[13]) ? 1'b0 : node1533;
											assign node1533 = (inp[9]) ? node1539 : node1534;
												assign node1534 = (inp[3]) ? node1536 : 1'b1;
													assign node1536 = (inp[12]) ? 1'b0 : 1'b1;
												assign node1539 = (inp[12]) ? 1'b0 : node1540;
													assign node1540 = (inp[7]) ? 1'b0 : 1'b1;
						assign node1546 = (inp[1]) ? node1646 : node1547;
							assign node1547 = (inp[12]) ? node1597 : node1548;
								assign node1548 = (inp[14]) ? node1574 : node1549;
									assign node1549 = (inp[10]) ? node1559 : node1550;
										assign node1550 = (inp[13]) ? node1552 : 1'b1;
											assign node1552 = (inp[4]) ? node1554 : 1'b1;
												assign node1554 = (inp[8]) ? node1556 : 1'b1;
													assign node1556 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1559 = (inp[13]) ? node1565 : node1560;
											assign node1560 = (inp[9]) ? node1562 : 1'b1;
												assign node1562 = (inp[8]) ? 1'b0 : 1'b1;
											assign node1565 = (inp[7]) ? node1569 : node1566;
												assign node1566 = (inp[8]) ? 1'b0 : 1'b1;
												assign node1569 = (inp[9]) ? 1'b0 : node1570;
													assign node1570 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1574 = (inp[3]) ? node1590 : node1575;
										assign node1575 = (inp[4]) ? node1583 : node1576;
											assign node1576 = (inp[9]) ? node1578 : 1'b1;
												assign node1578 = (inp[13]) ? node1580 : 1'b1;
													assign node1580 = (inp[8]) ? 1'b0 : 1'b1;
											assign node1583 = (inp[7]) ? 1'b0 : node1584;
												assign node1584 = (inp[13]) ? node1586 : 1'b1;
													assign node1586 = (inp[8]) ? 1'b1 : 1'b0;
										assign node1590 = (inp[8]) ? 1'b0 : node1591;
											assign node1591 = (inp[10]) ? 1'b0 : node1592;
												assign node1592 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1597 = (inp[8]) ? node1631 : node1598;
									assign node1598 = (inp[13]) ? node1618 : node1599;
										assign node1599 = (inp[10]) ? node1607 : node1600;
											assign node1600 = (inp[3]) ? node1602 : 1'b1;
												assign node1602 = (inp[7]) ? node1604 : 1'b1;
													assign node1604 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1607 = (inp[4]) ? node1613 : node1608;
												assign node1608 = (inp[9]) ? node1610 : 1'b1;
													assign node1610 = (inp[14]) ? 1'b0 : 1'b1;
												assign node1613 = (inp[14]) ? 1'b0 : node1614;
													assign node1614 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1618 = (inp[4]) ? 1'b0 : node1619;
											assign node1619 = (inp[3]) ? node1625 : node1620;
												assign node1620 = (inp[9]) ? node1622 : 1'b1;
													assign node1622 = (inp[14]) ? 1'b0 : 1'b1;
												assign node1625 = (inp[7]) ? 1'b0 : node1626;
													assign node1626 = (inp[14]) ? 1'b0 : 1'b1;
									assign node1631 = (inp[10]) ? 1'b0 : node1632;
										assign node1632 = (inp[3]) ? 1'b0 : node1633;
											assign node1633 = (inp[4]) ? node1639 : node1634;
												assign node1634 = (inp[13]) ? node1636 : 1'b1;
													assign node1636 = (inp[14]) ? 1'b0 : 1'b1;
												assign node1639 = (inp[7]) ? 1'b0 : node1640;
													assign node1640 = (inp[14]) ? 1'b1 : 1'b0;
							assign node1646 = (inp[13]) ? node1690 : node1647;
								assign node1647 = (inp[10]) ? node1671 : node1648;
									assign node1648 = (inp[8]) ? node1662 : node1649;
										assign node1649 = (inp[3]) ? node1655 : node1650;
											assign node1650 = (inp[7]) ? node1652 : 1'b1;
												assign node1652 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1655 = (inp[12]) ? 1'b0 : node1656;
												assign node1656 = (inp[14]) ? node1658 : 1'b1;
													assign node1658 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1662 = (inp[14]) ? 1'b0 : node1663;
											assign node1663 = (inp[9]) ? 1'b0 : node1664;
												assign node1664 = (inp[3]) ? node1666 : 1'b1;
													assign node1666 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1671 = (inp[14]) ? 1'b0 : node1672;
										assign node1672 = (inp[12]) ? node1684 : node1673;
											assign node1673 = (inp[3]) ? node1679 : node1674;
												assign node1674 = (inp[8]) ? node1676 : 1'b1;
													assign node1676 = (inp[4]) ? 1'b0 : 1'b1;
												assign node1679 = (inp[7]) ? 1'b0 : node1680;
													assign node1680 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1684 = (inp[8]) ? 1'b0 : node1685;
												assign node1685 = (inp[3]) ? 1'b0 : 1'b1;
								assign node1690 = (inp[12]) ? 1'b0 : node1691;
									assign node1691 = (inp[14]) ? node1703 : node1692;
										assign node1692 = (inp[4]) ? 1'b0 : node1693;
											assign node1693 = (inp[9]) ? node1699 : node1694;
												assign node1694 = (inp[10]) ? node1696 : 1'b1;
													assign node1696 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1699 = (inp[10]) ? 1'b1 : 1'b0;
										assign node1703 = (inp[3]) ? 1'b0 : node1704;
											assign node1704 = (inp[8]) ? 1'b0 : node1705;
												assign node1705 = (inp[10]) ? 1'b0 : node1706;
													assign node1706 = (inp[9]) ? 1'b0 : 1'b1;
				assign node1713 = (inp[1]) ? node2035 : node1714;
					assign node1714 = (inp[8]) ? node1858 : node1715;
						assign node1715 = (inp[7]) ? node1777 : node1716;
							assign node1716 = (inp[9]) ? node1734 : node1717;
								assign node1717 = (inp[14]) ? node1719 : 1'b1;
									assign node1719 = (inp[3]) ? node1721 : 1'b1;
										assign node1721 = (inp[5]) ? node1723 : 1'b1;
											assign node1723 = (inp[13]) ? node1729 : node1724;
												assign node1724 = (inp[11]) ? node1726 : 1'b1;
													assign node1726 = (inp[12]) ? 1'b0 : 1'b1;
												assign node1729 = (inp[4]) ? 1'b0 : node1730;
													assign node1730 = (inp[10]) ? 1'b0 : 1'b1;
								assign node1734 = (inp[12]) ? node1754 : node1735;
									assign node1735 = (inp[11]) ? node1745 : node1736;
										assign node1736 = (inp[14]) ? node1738 : 1'b1;
											assign node1738 = (inp[4]) ? node1740 : 1'b1;
												assign node1740 = (inp[5]) ? node1742 : 1'b1;
													assign node1742 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1745 = (inp[13]) ? node1747 : 1'b1;
											assign node1747 = (inp[5]) ? 1'b0 : node1748;
												assign node1748 = (inp[14]) ? node1750 : 1'b1;
													assign node1750 = (inp[4]) ? 1'b0 : 1'b1;
									assign node1754 = (inp[3]) ? node1766 : node1755;
										assign node1755 = (inp[5]) ? node1757 : 1'b1;
											assign node1757 = (inp[11]) ? node1763 : node1758;
												assign node1758 = (inp[4]) ? node1760 : 1'b1;
													assign node1760 = (inp[14]) ? 1'b0 : 1'b1;
												assign node1763 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1766 = (inp[10]) ? 1'b0 : node1767;
											assign node1767 = (inp[11]) ? node1771 : node1768;
												assign node1768 = (inp[14]) ? 1'b0 : 1'b1;
												assign node1771 = (inp[13]) ? 1'b0 : node1772;
													assign node1772 = (inp[4]) ? 1'b0 : 1'b1;
							assign node1777 = (inp[14]) ? node1811 : node1778;
								assign node1778 = (inp[10]) ? node1796 : node1779;
									assign node1779 = (inp[12]) ? node1781 : 1'b1;
										assign node1781 = (inp[13]) ? node1789 : node1782;
											assign node1782 = (inp[3]) ? node1784 : 1'b1;
												assign node1784 = (inp[9]) ? node1786 : 1'b1;
													assign node1786 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1789 = (inp[4]) ? 1'b0 : node1790;
												assign node1790 = (inp[3]) ? node1792 : 1'b1;
													assign node1792 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1796 = (inp[5]) ? node1806 : node1797;
										assign node1797 = (inp[13]) ? node1799 : 1'b1;
											assign node1799 = (inp[3]) ? 1'b0 : node1800;
												assign node1800 = (inp[9]) ? node1802 : 1'b1;
													assign node1802 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1806 = (inp[9]) ? 1'b0 : node1807;
											assign node1807 = (inp[13]) ? 1'b0 : 1'b1;
								assign node1811 = (inp[4]) ? node1843 : node1812;
									assign node1812 = (inp[9]) ? node1826 : node1813;
										assign node1813 = (inp[11]) ? node1815 : 1'b1;
											assign node1815 = (inp[10]) ? node1821 : node1816;
												assign node1816 = (inp[13]) ? node1818 : 1'b1;
													assign node1818 = (inp[5]) ? 1'b0 : 1'b1;
												assign node1821 = (inp[13]) ? 1'b0 : node1822;
													assign node1822 = (inp[12]) ? 1'b0 : 1'b0;
										assign node1826 = (inp[12]) ? node1838 : node1827;
											assign node1827 = (inp[13]) ? node1833 : node1828;
												assign node1828 = (inp[10]) ? node1830 : 1'b1;
													assign node1830 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1833 = (inp[10]) ? 1'b0 : node1834;
													assign node1834 = (inp[5]) ? 1'b0 : 1'b1;
											assign node1838 = (inp[11]) ? 1'b0 : node1839;
												assign node1839 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1843 = (inp[9]) ? 1'b0 : node1844;
										assign node1844 = (inp[5]) ? 1'b0 : node1845;
											assign node1845 = (inp[13]) ? node1851 : node1846;
												assign node1846 = (inp[3]) ? node1848 : 1'b1;
													assign node1848 = (inp[10]) ? 1'b0 : 1'b1;
												assign node1851 = (inp[12]) ? 1'b0 : node1852;
													assign node1852 = (inp[11]) ? 1'b0 : 1'b1;
						assign node1858 = (inp[10]) ? node1960 : node1859;
							assign node1859 = (inp[4]) ? node1911 : node1860;
								assign node1860 = (inp[9]) ? node1888 : node1861;
									assign node1861 = (inp[7]) ? node1869 : node1862;
										assign node1862 = (inp[12]) ? node1864 : 1'b1;
											assign node1864 = (inp[13]) ? node1866 : 1'b1;
												assign node1866 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1869 = (inp[11]) ? node1877 : node1870;
											assign node1870 = (inp[13]) ? 1'b1 : node1871;
												assign node1871 = (inp[3]) ? node1873 : 1'b1;
													assign node1873 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1877 = (inp[13]) ? node1883 : node1878;
												assign node1878 = (inp[14]) ? node1880 : 1'b1;
													assign node1880 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1883 = (inp[5]) ? 1'b0 : node1884;
													assign node1884 = (inp[12]) ? 1'b0 : 1'b1;
									assign node1888 = (inp[5]) ? node1898 : node1889;
										assign node1889 = (inp[12]) ? node1891 : 1'b1;
											assign node1891 = (inp[7]) ? 1'b0 : node1892;
												assign node1892 = (inp[11]) ? node1894 : 1'b1;
													assign node1894 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1898 = (inp[14]) ? 1'b0 : node1899;
											assign node1899 = (inp[13]) ? node1905 : node1900;
												assign node1900 = (inp[7]) ? node1902 : 1'b1;
													assign node1902 = (inp[12]) ? 1'b0 : 1'b1;
												assign node1905 = (inp[11]) ? 1'b0 : node1906;
													assign node1906 = (inp[12]) ? 1'b0 : 1'b1;
								assign node1911 = (inp[13]) ? node1939 : node1912;
									assign node1912 = (inp[7]) ? node1926 : node1913;
										assign node1913 = (inp[14]) ? node1915 : 1'b1;
											assign node1915 = (inp[11]) ? node1921 : node1916;
												assign node1916 = (inp[3]) ? node1918 : 1'b1;
													assign node1918 = (inp[12]) ? 1'b0 : 1'b1;
												assign node1921 = (inp[9]) ? 1'b0 : node1922;
													assign node1922 = (inp[5]) ? 1'b0 : 1'b1;
										assign node1926 = (inp[11]) ? node1934 : node1927;
											assign node1927 = (inp[12]) ? node1929 : 1'b1;
												assign node1929 = (inp[9]) ? 1'b0 : node1930;
													assign node1930 = (inp[5]) ? 1'b0 : 1'b1;
											assign node1934 = (inp[3]) ? 1'b0 : node1935;
												assign node1935 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1939 = (inp[11]) ? node1953 : node1940;
										assign node1940 = (inp[14]) ? 1'b0 : node1941;
											assign node1941 = (inp[12]) ? node1947 : node1942;
												assign node1942 = (inp[3]) ? node1944 : 1'b1;
													assign node1944 = (inp[5]) ? 1'b0 : 1'b1;
												assign node1947 = (inp[7]) ? 1'b0 : node1948;
													assign node1948 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1953 = (inp[14]) ? node1955 : 1'b0;
											assign node1955 = (inp[5]) ? 1'b0 : node1956;
												assign node1956 = (inp[7]) ? 1'b0 : 1'b1;
							assign node1960 = (inp[4]) ? node2026 : node1961;
								assign node1961 = (inp[12]) ? node1999 : node1962;
									assign node1962 = (inp[5]) ? node1980 : node1963;
										assign node1963 = (inp[3]) ? node1969 : node1964;
											assign node1964 = (inp[9]) ? node1966 : 1'b1;
												assign node1966 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1969 = (inp[11]) ? node1975 : node1970;
												assign node1970 = (inp[14]) ? node1972 : 1'b1;
													assign node1972 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1975 = (inp[13]) ? 1'b0 : node1976;
													assign node1976 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1980 = (inp[14]) ? node1992 : node1981;
											assign node1981 = (inp[13]) ? node1987 : node1982;
												assign node1982 = (inp[3]) ? node1984 : 1'b1;
													assign node1984 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1987 = (inp[9]) ? 1'b0 : node1988;
													assign node1988 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1992 = (inp[9]) ? 1'b0 : node1993;
												assign node1993 = (inp[7]) ? 1'b0 : node1994;
													assign node1994 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1999 = (inp[3]) ? node2017 : node2000;
										assign node2000 = (inp[14]) ? node2012 : node2001;
											assign node2001 = (inp[5]) ? node2007 : node2002;
												assign node2002 = (inp[9]) ? node2004 : 1'b1;
													assign node2004 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2007 = (inp[13]) ? 1'b0 : node2008;
													assign node2008 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2012 = (inp[13]) ? 1'b0 : node2013;
												assign node2013 = (inp[9]) ? 1'b0 : 1'b1;
										assign node2017 = (inp[13]) ? 1'b0 : node2018;
											assign node2018 = (inp[9]) ? 1'b0 : node2019;
												assign node2019 = (inp[7]) ? 1'b0 : node2020;
													assign node2020 = (inp[11]) ? 1'b0 : 1'b1;
								assign node2026 = (inp[3]) ? 1'b0 : node2027;
									assign node2027 = (inp[5]) ? 1'b0 : node2028;
										assign node2028 = (inp[7]) ? 1'b0 : node2029;
											assign node2029 = (inp[12]) ? 1'b0 : 1'b1;
					assign node2035 = (inp[12]) ? node2219 : node2036;
						assign node2036 = (inp[3]) ? node2130 : node2037;
							assign node2037 = (inp[5]) ? node2089 : node2038;
								assign node2038 = (inp[9]) ? node2056 : node2039;
									assign node2039 = (inp[7]) ? node2041 : 1'b1;
										assign node2041 = (inp[4]) ? node2049 : node2042;
											assign node2042 = (inp[10]) ? node2044 : 1'b1;
												assign node2044 = (inp[11]) ? node2046 : 1'b1;
													assign node2046 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2049 = (inp[13]) ? 1'b0 : node2050;
												assign node2050 = (inp[11]) ? node2052 : 1'b1;
													assign node2052 = (inp[14]) ? 1'b0 : 1'b1;
									assign node2056 = (inp[10]) ? node2074 : node2057;
										assign node2057 = (inp[4]) ? node2065 : node2058;
											assign node2058 = (inp[14]) ? node2060 : 1'b1;
												assign node2060 = (inp[13]) ? node2062 : 1'b1;
													assign node2062 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2065 = (inp[13]) ? node2069 : node2066;
												assign node2066 = (inp[8]) ? 1'b0 : 1'b1;
												assign node2069 = (inp[14]) ? 1'b0 : node2070;
													assign node2070 = (inp[8]) ? 1'b1 : 1'b0;
										assign node2074 = (inp[14]) ? node2082 : node2075;
											assign node2075 = (inp[8]) ? node2077 : 1'b1;
												assign node2077 = (inp[7]) ? 1'b0 : node2078;
													assign node2078 = (inp[4]) ? 1'b0 : 1'b1;
											assign node2082 = (inp[11]) ? 1'b0 : node2083;
												assign node2083 = (inp[7]) ? 1'b0 : node2084;
													assign node2084 = (inp[13]) ? 1'b0 : 1'b1;
								assign node2089 = (inp[11]) ? node2119 : node2090;
									assign node2090 = (inp[14]) ? node2104 : node2091;
										assign node2091 = (inp[4]) ? node2093 : 1'b1;
											assign node2093 = (inp[7]) ? node2099 : node2094;
												assign node2094 = (inp[8]) ? node2096 : 1'b1;
													assign node2096 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2099 = (inp[9]) ? 1'b0 : node2100;
													assign node2100 = (inp[8]) ? 1'b0 : 1'b1;
										assign node2104 = (inp[4]) ? node2112 : node2105;
											assign node2105 = (inp[13]) ? node2107 : 1'b1;
												assign node2107 = (inp[9]) ? 1'b0 : node2108;
													assign node2108 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2112 = (inp[10]) ? 1'b0 : node2113;
												assign node2113 = (inp[8]) ? 1'b0 : node2114;
													assign node2114 = (inp[7]) ? 1'b0 : 1'b1;
									assign node2119 = (inp[10]) ? 1'b0 : node2120;
										assign node2120 = (inp[13]) ? 1'b0 : node2121;
											assign node2121 = (inp[9]) ? 1'b0 : node2122;
												assign node2122 = (inp[4]) ? node2124 : 1'b1;
													assign node2124 = (inp[8]) ? 1'b0 : 1'b1;
							assign node2130 = (inp[8]) ? node2190 : node2131;
								assign node2131 = (inp[14]) ? node2169 : node2132;
									assign node2132 = (inp[9]) ? node2152 : node2133;
										assign node2133 = (inp[5]) ? node2141 : node2134;
											assign node2134 = (inp[7]) ? node2136 : 1'b1;
												assign node2136 = (inp[11]) ? node2138 : 1'b1;
													assign node2138 = (inp[4]) ? 1'b0 : 1'b1;
											assign node2141 = (inp[13]) ? node2147 : node2142;
												assign node2142 = (inp[10]) ? node2144 : 1'b1;
													assign node2144 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2147 = (inp[7]) ? 1'b0 : node2148;
													assign node2148 = (inp[4]) ? 1'b0 : 1'b1;
										assign node2152 = (inp[4]) ? node2164 : node2153;
											assign node2153 = (inp[5]) ? node2159 : node2154;
												assign node2154 = (inp[10]) ? node2156 : 1'b1;
													assign node2156 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2159 = (inp[7]) ? 1'b0 : node2160;
													assign node2160 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2164 = (inp[7]) ? 1'b0 : node2165;
												assign node2165 = (inp[13]) ? 1'b0 : 1'b1;
									assign node2169 = (inp[10]) ? node2181 : node2170;
										assign node2170 = (inp[13]) ? node2174 : node2171;
											assign node2171 = (inp[4]) ? 1'b0 : 1'b1;
											assign node2174 = (inp[5]) ? 1'b0 : node2175;
												assign node2175 = (inp[9]) ? 1'b0 : node2176;
													assign node2176 = (inp[7]) ? 1'b0 : 1'b1;
										assign node2181 = (inp[11]) ? 1'b0 : node2182;
											assign node2182 = (inp[7]) ? 1'b0 : node2183;
												assign node2183 = (inp[5]) ? 1'b0 : node2184;
													assign node2184 = (inp[13]) ? 1'b0 : 1'b1;
								assign node2190 = (inp[10]) ? 1'b0 : node2191;
									assign node2191 = (inp[7]) ? node2211 : node2192;
										assign node2192 = (inp[4]) ? node2204 : node2193;
											assign node2193 = (inp[11]) ? node2199 : node2194;
												assign node2194 = (inp[9]) ? node2196 : 1'b1;
													assign node2196 = (inp[14]) ? 1'b0 : 1'b1;
												assign node2199 = (inp[14]) ? 1'b0 : node2200;
													assign node2200 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2204 = (inp[13]) ? 1'b0 : node2205;
												assign node2205 = (inp[9]) ? 1'b0 : node2206;
													assign node2206 = (inp[5]) ? 1'b0 : 1'b1;
										assign node2211 = (inp[11]) ? 1'b0 : node2212;
											assign node2212 = (inp[4]) ? 1'b0 : node2213;
												assign node2213 = (inp[5]) ? 1'b0 : 1'b1;
						assign node2219 = (inp[10]) ? node2281 : node2220;
							assign node2220 = (inp[8]) ? node2264 : node2221;
								assign node2221 = (inp[9]) ? node2245 : node2222;
									assign node2222 = (inp[5]) ? node2232 : node2223;
										assign node2223 = (inp[14]) ? node2225 : 1'b1;
											assign node2225 = (inp[3]) ? 1'b0 : node2226;
												assign node2226 = (inp[4]) ? node2228 : 1'b1;
													assign node2228 = (inp[7]) ? 1'b0 : 1'b1;
										assign node2232 = (inp[7]) ? 1'b0 : node2233;
											assign node2233 = (inp[11]) ? node2239 : node2234;
												assign node2234 = (inp[4]) ? node2236 : 1'b1;
													assign node2236 = (inp[14]) ? 1'b0 : 1'b0;
												assign node2239 = (inp[13]) ? 1'b0 : node2240;
													assign node2240 = (inp[14]) ? 1'b0 : 1'b1;
									assign node2245 = (inp[7]) ? node2257 : node2246;
										assign node2246 = (inp[3]) ? node2250 : node2247;
											assign node2247 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2250 = (inp[5]) ? 1'b0 : node2251;
												assign node2251 = (inp[14]) ? 1'b0 : node2252;
													assign node2252 = (inp[13]) ? 1'b0 : 1'b1;
										assign node2257 = (inp[14]) ? 1'b0 : node2258;
											assign node2258 = (inp[13]) ? 1'b0 : node2259;
												assign node2259 = (inp[11]) ? 1'b0 : 1'b1;
								assign node2264 = (inp[11]) ? 1'b0 : node2265;
									assign node2265 = (inp[7]) ? 1'b0 : node2266;
										assign node2266 = (inp[3]) ? node2274 : node2267;
											assign node2267 = (inp[13]) ? node2269 : 1'b1;
												assign node2269 = (inp[5]) ? 1'b0 : node2270;
													assign node2270 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2274 = (inp[5]) ? 1'b0 : node2275;
												assign node2275 = (inp[14]) ? 1'b0 : 1'b1;
							assign node2281 = (inp[9]) ? node2321 : node2282;
								assign node2282 = (inp[11]) ? node2310 : node2283;
									assign node2283 = (inp[5]) ? node2301 : node2284;
										assign node2284 = (inp[4]) ? node2296 : node2285;
											assign node2285 = (inp[7]) ? node2291 : node2286;
												assign node2286 = (inp[13]) ? node2288 : 1'b1;
													assign node2288 = (inp[8]) ? 1'b0 : 1'b1;
												assign node2291 = (inp[14]) ? 1'b0 : node2292;
													assign node2292 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2296 = (inp[8]) ? 1'b0 : node2297;
												assign node2297 = (inp[13]) ? 1'b0 : 1'b1;
										assign node2301 = (inp[13]) ? node2303 : 1'b0;
											assign node2303 = (inp[3]) ? 1'b0 : node2304;
												assign node2304 = (inp[14]) ? 1'b0 : node2305;
													assign node2305 = (inp[4]) ? 1'b0 : 1'b1;
									assign node2310 = (inp[3]) ? 1'b0 : node2311;
										assign node2311 = (inp[13]) ? 1'b0 : node2312;
											assign node2312 = (inp[7]) ? 1'b0 : node2313;
												assign node2313 = (inp[14]) ? 1'b0 : node2314;
													assign node2314 = (inp[4]) ? 1'b0 : 1'b1;
								assign node2321 = (inp[13]) ? 1'b0 : node2322;
									assign node2322 = (inp[14]) ? 1'b0 : node2323;
										assign node2323 = (inp[4]) ? 1'b0 : node2324;
											assign node2324 = (inp[3]) ? 1'b0 : node2325;
												assign node2325 = (inp[5]) ? 1'b0 : 1'b1;
		assign node2332 = (inp[4]) ? node3548 : node2333;
			assign node2333 = (inp[1]) ? node2923 : node2334;
				assign node2334 = (inp[5]) ? node2594 : node2335;
					assign node2335 = (inp[11]) ? node2431 : node2336;
						assign node2336 = (inp[8]) ? node2364 : node2337;
							assign node2337 = (inp[10]) ? node2339 : 1'b1;
								assign node2339 = (inp[6]) ? node2341 : 1'b1;
									assign node2341 = (inp[12]) ? node2349 : node2342;
										assign node2342 = (inp[9]) ? node2344 : 1'b1;
											assign node2344 = (inp[13]) ? node2346 : 1'b1;
												assign node2346 = (inp[0]) ? 1'b0 : 1'b1;
										assign node2349 = (inp[14]) ? node2357 : node2350;
											assign node2350 = (inp[3]) ? node2352 : 1'b1;
												assign node2352 = (inp[0]) ? node2354 : 1'b1;
													assign node2354 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2357 = (inp[0]) ? 1'b0 : node2358;
												assign node2358 = (inp[3]) ? node2360 : 1'b1;
													assign node2360 = (inp[9]) ? 1'b0 : 1'b1;
							assign node2364 = (inp[6]) ? node2388 : node2365;
								assign node2365 = (inp[12]) ? node2367 : 1'b1;
									assign node2367 = (inp[13]) ? node2375 : node2368;
										assign node2368 = (inp[3]) ? node2370 : 1'b1;
											assign node2370 = (inp[14]) ? node2372 : 1'b1;
												assign node2372 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2375 = (inp[9]) ? node2381 : node2376;
											assign node2376 = (inp[14]) ? node2378 : 1'b1;
												assign node2378 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2381 = (inp[10]) ? 1'b0 : node2382;
												assign node2382 = (inp[7]) ? node2384 : 1'b1;
													assign node2384 = (inp[0]) ? 1'b0 : 1'b1;
								assign node2388 = (inp[10]) ? node2404 : node2389;
									assign node2389 = (inp[13]) ? node2391 : 1'b1;
										assign node2391 = (inp[9]) ? node2399 : node2392;
											assign node2392 = (inp[3]) ? node2394 : 1'b1;
												assign node2394 = (inp[0]) ? node2396 : 1'b1;
													assign node2396 = (inp[7]) ? 1'b0 : 1'b0;
											assign node2399 = (inp[7]) ? 1'b0 : node2400;
												assign node2400 = (inp[0]) ? 1'b0 : 1'b1;
									assign node2404 = (inp[0]) ? node2418 : node2405;
										assign node2405 = (inp[14]) ? node2407 : 1'b1;
											assign node2407 = (inp[9]) ? node2413 : node2408;
												assign node2408 = (inp[12]) ? node2410 : 1'b1;
													assign node2410 = (inp[3]) ? 1'b0 : 1'b1;
												assign node2413 = (inp[13]) ? 1'b0 : node2414;
													assign node2414 = (inp[7]) ? 1'b0 : 1'b1;
										assign node2418 = (inp[3]) ? 1'b0 : node2419;
											assign node2419 = (inp[12]) ? node2425 : node2420;
												assign node2420 = (inp[14]) ? node2422 : 1'b1;
													assign node2422 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2425 = (inp[14]) ? 1'b0 : node2426;
													assign node2426 = (inp[13]) ? 1'b0 : 1'b1;
						assign node2431 = (inp[12]) ? node2499 : node2432;
							assign node2432 = (inp[10]) ? node2458 : node2433;
								assign node2433 = (inp[9]) ? node2435 : 1'b1;
									assign node2435 = (inp[14]) ? node2445 : node2436;
										assign node2436 = (inp[13]) ? node2438 : 1'b1;
											assign node2438 = (inp[8]) ? node2440 : 1'b1;
												assign node2440 = (inp[7]) ? node2442 : 1'b1;
													assign node2442 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2445 = (inp[6]) ? node2447 : 1'b1;
											assign node2447 = (inp[13]) ? node2453 : node2448;
												assign node2448 = (inp[8]) ? node2450 : 1'b1;
													assign node2450 = (inp[3]) ? 1'b0 : 1'b1;
												assign node2453 = (inp[3]) ? 1'b0 : node2454;
													assign node2454 = (inp[0]) ? 1'b0 : 1'b1;
								assign node2458 = (inp[3]) ? node2480 : node2459;
									assign node2459 = (inp[9]) ? node2461 : 1'b1;
										assign node2461 = (inp[6]) ? node2469 : node2462;
											assign node2462 = (inp[13]) ? node2464 : 1'b1;
												assign node2464 = (inp[7]) ? node2466 : 1'b1;
													assign node2466 = (inp[0]) ? 1'b0 : 1'b1;
											assign node2469 = (inp[13]) ? node2475 : node2470;
												assign node2470 = (inp[0]) ? node2472 : 1'b1;
													assign node2472 = (inp[14]) ? 1'b0 : 1'b1;
												assign node2475 = (inp[8]) ? 1'b0 : node2476;
													assign node2476 = (inp[7]) ? 1'b0 : 1'b1;
									assign node2480 = (inp[7]) ? node2490 : node2481;
										assign node2481 = (inp[6]) ? node2483 : 1'b1;
											assign node2483 = (inp[0]) ? 1'b0 : node2484;
												assign node2484 = (inp[13]) ? node2486 : 1'b1;
													assign node2486 = (inp[8]) ? 1'b0 : 1'b1;
										assign node2490 = (inp[13]) ? 1'b0 : node2491;
											assign node2491 = (inp[6]) ? 1'b0 : node2492;
												assign node2492 = (inp[8]) ? node2494 : 1'b1;
													assign node2494 = (inp[0]) ? 1'b0 : 1'b0;
							assign node2499 = (inp[14]) ? node2555 : node2500;
								assign node2500 = (inp[3]) ? node2526 : node2501;
									assign node2501 = (inp[10]) ? node2509 : node2502;
										assign node2502 = (inp[9]) ? node2504 : 1'b1;
											assign node2504 = (inp[6]) ? node2506 : 1'b1;
												assign node2506 = (inp[0]) ? 1'b0 : 1'b1;
										assign node2509 = (inp[7]) ? node2515 : node2510;
											assign node2510 = (inp[6]) ? node2512 : 1'b1;
												assign node2512 = (inp[8]) ? 1'b1 : 1'b0;
											assign node2515 = (inp[8]) ? node2521 : node2516;
												assign node2516 = (inp[6]) ? node2518 : 1'b1;
													assign node2518 = (inp[9]) ? 1'b0 : 1'b1;
												assign node2521 = (inp[0]) ? 1'b0 : node2522;
													assign node2522 = (inp[9]) ? 1'b0 : 1'b1;
									assign node2526 = (inp[0]) ? node2546 : node2527;
										assign node2527 = (inp[7]) ? node2535 : node2528;
											assign node2528 = (inp[13]) ? 1'b1 : node2529;
												assign node2529 = (inp[6]) ? node2531 : 1'b1;
													assign node2531 = (inp[9]) ? 1'b1 : 1'b1;
											assign node2535 = (inp[8]) ? node2541 : node2536;
												assign node2536 = (inp[6]) ? node2538 : 1'b1;
													assign node2538 = (inp[9]) ? 1'b0 : 1'b1;
												assign node2541 = (inp[10]) ? node2543 : 1'b0;
													assign node2543 = (inp[13]) ? 1'b0 : 1'b1;
										assign node2546 = (inp[13]) ? 1'b0 : node2547;
											assign node2547 = (inp[10]) ? node2549 : 1'b1;
												assign node2549 = (inp[8]) ? 1'b0 : node2550;
													assign node2550 = (inp[6]) ? 1'b0 : 1'b1;
								assign node2555 = (inp[7]) ? node2579 : node2556;
									assign node2556 = (inp[13]) ? node2570 : node2557;
										assign node2557 = (inp[6]) ? node2559 : 1'b1;
											assign node2559 = (inp[9]) ? node2565 : node2560;
												assign node2560 = (inp[3]) ? node2562 : 1'b1;
													assign node2562 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2565 = (inp[10]) ? 1'b0 : node2566;
													assign node2566 = (inp[8]) ? 1'b0 : 1'b1;
										assign node2570 = (inp[0]) ? 1'b0 : node2571;
											assign node2571 = (inp[6]) ? node2573 : 1'b1;
												assign node2573 = (inp[8]) ? 1'b0 : node2574;
													assign node2574 = (inp[3]) ? 1'b0 : 1'b1;
									assign node2579 = (inp[6]) ? 1'b0 : node2580;
										assign node2580 = (inp[0]) ? 1'b0 : node2581;
											assign node2581 = (inp[13]) ? node2587 : node2582;
												assign node2582 = (inp[9]) ? node2584 : 1'b1;
													assign node2584 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2587 = (inp[8]) ? 1'b0 : node2588;
													assign node2588 = (inp[9]) ? 1'b0 : 1'b1;
					assign node2594 = (inp[9]) ? node2750 : node2595;
						assign node2595 = (inp[13]) ? node2661 : node2596;
							assign node2596 = (inp[12]) ? node2606 : node2597;
								assign node2597 = (inp[14]) ? node2599 : 1'b1;
									assign node2599 = (inp[11]) ? node2601 : 1'b1;
										assign node2601 = (inp[7]) ? node2603 : 1'b1;
											assign node2603 = (inp[8]) ? 1'b0 : 1'b1;
								assign node2606 = (inp[14]) ? node2628 : node2607;
									assign node2607 = (inp[0]) ? node2609 : 1'b1;
										assign node2609 = (inp[11]) ? node2617 : node2610;
											assign node2610 = (inp[10]) ? node2612 : 1'b1;
												assign node2612 = (inp[3]) ? node2614 : 1'b1;
													assign node2614 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2617 = (inp[7]) ? node2623 : node2618;
												assign node2618 = (inp[10]) ? node2620 : 1'b1;
													assign node2620 = (inp[3]) ? 1'b0 : 1'b1;
												assign node2623 = (inp[3]) ? 1'b0 : node2624;
													assign node2624 = (inp[10]) ? 1'b0 : 1'b1;
									assign node2628 = (inp[8]) ? node2648 : node2629;
										assign node2629 = (inp[10]) ? node2637 : node2630;
											assign node2630 = (inp[11]) ? node2632 : 1'b1;
												assign node2632 = (inp[7]) ? node2634 : 1'b1;
													assign node2634 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2637 = (inp[6]) ? node2643 : node2638;
												assign node2638 = (inp[11]) ? node2640 : 1'b1;
													assign node2640 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2643 = (inp[11]) ? 1'b0 : node2644;
													assign node2644 = (inp[7]) ? 1'b0 : 1'b1;
										assign node2648 = (inp[11]) ? 1'b0 : node2649;
											assign node2649 = (inp[3]) ? node2655 : node2650;
												assign node2650 = (inp[10]) ? node2652 : 1'b1;
													assign node2652 = (inp[0]) ? 1'b0 : 1'b1;
												assign node2655 = (inp[6]) ? 1'b0 : node2656;
													assign node2656 = (inp[0]) ? 1'b0 : 1'b1;
							assign node2661 = (inp[0]) ? node2715 : node2662;
								assign node2662 = (inp[6]) ? node2682 : node2663;
									assign node2663 = (inp[8]) ? node2673 : node2664;
										assign node2664 = (inp[11]) ? node2666 : 1'b1;
											assign node2666 = (inp[14]) ? node2668 : 1'b1;
												assign node2668 = (inp[12]) ? node2670 : 1'b1;
													assign node2670 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2673 = (inp[10]) ? node2679 : node2674;
											assign node2674 = (inp[12]) ? node2676 : 1'b1;
												assign node2676 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2679 = (inp[3]) ? 1'b0 : 1'b1;
									assign node2682 = (inp[14]) ? node2702 : node2683;
										assign node2683 = (inp[11]) ? node2691 : node2684;
											assign node2684 = (inp[7]) ? node2686 : 1'b1;
												assign node2686 = (inp[10]) ? node2688 : 1'b1;
													assign node2688 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2691 = (inp[3]) ? node2697 : node2692;
												assign node2692 = (inp[7]) ? node2694 : 1'b1;
													assign node2694 = (inp[8]) ? 1'b0 : 1'b1;
												assign node2697 = (inp[8]) ? 1'b0 : node2698;
													assign node2698 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2702 = (inp[7]) ? 1'b0 : node2703;
											assign node2703 = (inp[3]) ? node2709 : node2704;
												assign node2704 = (inp[8]) ? node2706 : 1'b1;
													assign node2706 = (inp[12]) ? 1'b0 : 1'b1;
												assign node2709 = (inp[8]) ? 1'b0 : node2710;
													assign node2710 = (inp[10]) ? 1'b0 : 1'b1;
								assign node2715 = (inp[3]) ? node2735 : node2716;
									assign node2716 = (inp[14]) ? node2722 : node2717;
										assign node2717 = (inp[11]) ? node2719 : 1'b1;
											assign node2719 = (inp[12]) ? 1'b0 : 1'b1;
										assign node2722 = (inp[8]) ? 1'b0 : node2723;
											assign node2723 = (inp[10]) ? node2729 : node2724;
												assign node2724 = (inp[6]) ? node2726 : 1'b1;
													assign node2726 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2729 = (inp[6]) ? 1'b0 : node2730;
													assign node2730 = (inp[7]) ? 1'b0 : 1'b1;
									assign node2735 = (inp[10]) ? 1'b0 : node2736;
										assign node2736 = (inp[14]) ? 1'b0 : node2737;
											assign node2737 = (inp[11]) ? node2743 : node2738;
												assign node2738 = (inp[6]) ? node2740 : 1'b1;
													assign node2740 = (inp[8]) ? 1'b0 : 1'b1;
												assign node2743 = (inp[12]) ? 1'b0 : node2744;
													assign node2744 = (inp[8]) ? 1'b0 : 1'b1;
						assign node2750 = (inp[0]) ? node2848 : node2751;
							assign node2751 = (inp[3]) ? node2803 : node2752;
								assign node2752 = (inp[13]) ? node2770 : node2753;
									assign node2753 = (inp[7]) ? node2755 : 1'b1;
										assign node2755 = (inp[11]) ? node2763 : node2756;
											assign node2756 = (inp[10]) ? node2758 : 1'b1;
												assign node2758 = (inp[8]) ? node2760 : 1'b1;
													assign node2760 = (inp[12]) ? 1'b0 : 1'b1;
											assign node2763 = (inp[14]) ? node2765 : 1'b1;
												assign node2765 = (inp[8]) ? 1'b0 : node2766;
													assign node2766 = (inp[6]) ? 1'b0 : 1'b1;
									assign node2770 = (inp[6]) ? node2790 : node2771;
										assign node2771 = (inp[8]) ? node2779 : node2772;
											assign node2772 = (inp[14]) ? node2774 : 1'b1;
												assign node2774 = (inp[12]) ? node2776 : 1'b1;
													assign node2776 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2779 = (inp[12]) ? node2785 : node2780;
												assign node2780 = (inp[7]) ? node2782 : 1'b1;
													assign node2782 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2785 = (inp[7]) ? 1'b0 : node2786;
													assign node2786 = (inp[14]) ? 1'b0 : 1'b1;
										assign node2790 = (inp[12]) ? 1'b0 : node2791;
											assign node2791 = (inp[14]) ? node2797 : node2792;
												assign node2792 = (inp[8]) ? node2794 : 1'b1;
													assign node2794 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2797 = (inp[7]) ? 1'b0 : node2798;
													assign node2798 = (inp[8]) ? 1'b0 : 1'b1;
								assign node2803 = (inp[14]) ? node2829 : node2804;
									assign node2804 = (inp[6]) ? node2814 : node2805;
										assign node2805 = (inp[11]) ? node2807 : 1'b1;
											assign node2807 = (inp[8]) ? node2809 : 1'b1;
												assign node2809 = (inp[13]) ? 1'b0 : node2810;
													assign node2810 = (inp[7]) ? 1'b0 : 1'b1;
										assign node2814 = (inp[7]) ? node2822 : node2815;
											assign node2815 = (inp[11]) ? node2817 : 1'b1;
												assign node2817 = (inp[12]) ? 1'b0 : node2818;
													assign node2818 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2822 = (inp[8]) ? 1'b0 : node2823;
												assign node2823 = (inp[12]) ? 1'b0 : node2824;
													assign node2824 = (inp[13]) ? 1'b0 : 1'b1;
									assign node2829 = (inp[7]) ? 1'b0 : node2830;
										assign node2830 = (inp[6]) ? node2842 : node2831;
											assign node2831 = (inp[12]) ? node2837 : node2832;
												assign node2832 = (inp[8]) ? node2834 : 1'b1;
													assign node2834 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2837 = (inp[10]) ? 1'b0 : node2838;
													assign node2838 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2842 = (inp[10]) ? 1'b0 : node2843;
												assign node2843 = (inp[11]) ? 1'b0 : 1'b1;
							assign node2848 = (inp[10]) ? node2902 : node2849;
								assign node2849 = (inp[12]) ? node2879 : node2850;
									assign node2850 = (inp[7]) ? node2864 : node2851;
										assign node2851 = (inp[11]) ? node2857 : node2852;
											assign node2852 = (inp[3]) ? node2854 : 1'b1;
												assign node2854 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2857 = (inp[6]) ? 1'b0 : node2858;
												assign node2858 = (inp[13]) ? node2860 : 1'b1;
													assign node2860 = (inp[14]) ? 1'b0 : 1'b1;
										assign node2864 = (inp[14]) ? node2872 : node2865;
											assign node2865 = (inp[3]) ? node2867 : 1'b1;
												assign node2867 = (inp[11]) ? 1'b0 : node2868;
													assign node2868 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2872 = (inp[6]) ? 1'b0 : node2873;
												assign node2873 = (inp[3]) ? 1'b0 : node2874;
													assign node2874 = (inp[13]) ? 1'b0 : 1'b1;
									assign node2879 = (inp[8]) ? node2895 : node2880;
										assign node2880 = (inp[14]) ? node2888 : node2881;
											assign node2881 = (inp[6]) ? 1'b0 : node2882;
												assign node2882 = (inp[13]) ? node2884 : 1'b1;
													assign node2884 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2888 = (inp[3]) ? 1'b0 : node2889;
												assign node2889 = (inp[11]) ? 1'b0 : node2890;
													assign node2890 = (inp[7]) ? 1'b0 : 1'b1;
										assign node2895 = (inp[13]) ? 1'b0 : node2896;
											assign node2896 = (inp[3]) ? 1'b0 : node2897;
												assign node2897 = (inp[6]) ? 1'b0 : 1'b1;
								assign node2902 = (inp[3]) ? 1'b0 : node2903;
									assign node2903 = (inp[13]) ? node2913 : node2904;
										assign node2904 = (inp[6]) ? 1'b0 : node2905;
											assign node2905 = (inp[8]) ? node2907 : 1'b1;
												assign node2907 = (inp[7]) ? 1'b0 : node2908;
													assign node2908 = (inp[14]) ? 1'b0 : 1'b0;
										assign node2913 = (inp[11]) ? 1'b0 : node2914;
											assign node2914 = (inp[12]) ? 1'b0 : node2915;
												assign node2915 = (inp[7]) ? 1'b0 : node2916;
													assign node2916 = (inp[8]) ? 1'b0 : 1'b1;
				assign node2923 = (inp[6]) ? node3231 : node2924;
					assign node2924 = (inp[10]) ? node3070 : node2925;
						assign node2925 = (inp[11]) ? node2991 : node2926;
							assign node2926 = (inp[3]) ? node2948 : node2927;
								assign node2927 = (inp[8]) ? node2929 : 1'b1;
									assign node2929 = (inp[9]) ? node2937 : node2930;
										assign node2930 = (inp[13]) ? node2932 : 1'b1;
											assign node2932 = (inp[0]) ? node2934 : 1'b1;
												assign node2934 = (inp[7]) ? 1'b0 : 1'b1;
										assign node2937 = (inp[7]) ? node2943 : node2938;
											assign node2938 = (inp[14]) ? node2940 : 1'b1;
												assign node2940 = (inp[12]) ? 1'b0 : 1'b1;
											assign node2943 = (inp[14]) ? 1'b0 : node2944;
												assign node2944 = (inp[5]) ? 1'b0 : 1'b1;
								assign node2948 = (inp[13]) ? node2968 : node2949;
									assign node2949 = (inp[8]) ? node2957 : node2950;
										assign node2950 = (inp[0]) ? node2952 : 1'b1;
											assign node2952 = (inp[9]) ? node2954 : 1'b1;
												assign node2954 = (inp[5]) ? 1'b0 : 1'b1;
										assign node2957 = (inp[7]) ? node2959 : 1'b1;
											assign node2959 = (inp[9]) ? node2963 : node2960;
												assign node2960 = (inp[0]) ? 1'b0 : 1'b1;
												assign node2963 = (inp[12]) ? 1'b0 : node2964;
													assign node2964 = (inp[5]) ? 1'b0 : 1'b1;
									assign node2968 = (inp[14]) ? node2978 : node2969;
										assign node2969 = (inp[0]) ? node2971 : 1'b1;
											assign node2971 = (inp[8]) ? node2973 : 1'b1;
												assign node2973 = (inp[9]) ? 1'b0 : node2974;
													assign node2974 = (inp[5]) ? 1'b0 : 1'b1;
										assign node2978 = (inp[12]) ? 1'b0 : node2979;
											assign node2979 = (inp[0]) ? node2985 : node2980;
												assign node2980 = (inp[8]) ? node2982 : 1'b1;
													assign node2982 = (inp[5]) ? 1'b0 : 1'b1;
												assign node2985 = (inp[9]) ? 1'b0 : node2986;
													assign node2986 = (inp[7]) ? 1'b0 : 1'b1;
							assign node2991 = (inp[8]) ? node3025 : node2992;
								assign node2992 = (inp[5]) ? node3008 : node2993;
									assign node2993 = (inp[13]) ? node2995 : 1'b1;
										assign node2995 = (inp[3]) ? node2997 : 1'b1;
											assign node2997 = (inp[14]) ? node3003 : node2998;
												assign node2998 = (inp[7]) ? node3000 : 1'b1;
													assign node3000 = (inp[0]) ? 1'b0 : 1'b1;
												assign node3003 = (inp[7]) ? 1'b0 : node3004;
													assign node3004 = (inp[0]) ? 1'b0 : 1'b1;
									assign node3008 = (inp[7]) ? node3018 : node3009;
										assign node3009 = (inp[3]) ? node3011 : 1'b1;
											assign node3011 = (inp[0]) ? node3013 : 1'b1;
												assign node3013 = (inp[13]) ? node3015 : 1'b0;
													assign node3015 = (inp[9]) ? 1'b0 : 1'b0;
										assign node3018 = (inp[13]) ? 1'b0 : node3019;
											assign node3019 = (inp[3]) ? node3021 : 1'b1;
												assign node3021 = (inp[0]) ? 1'b0 : 1'b1;
								assign node3025 = (inp[9]) ? node3049 : node3026;
									assign node3026 = (inp[13]) ? node3034 : node3027;
										assign node3027 = (inp[12]) ? node3029 : 1'b1;
											assign node3029 = (inp[5]) ? node3031 : 1'b1;
												assign node3031 = (inp[3]) ? 1'b0 : 1'b1;
										assign node3034 = (inp[3]) ? node3042 : node3035;
											assign node3035 = (inp[0]) ? 1'b0 : node3036;
												assign node3036 = (inp[5]) ? node3038 : 1'b1;
													assign node3038 = (inp[7]) ? 1'b0 : 1'b1;
											assign node3042 = (inp[14]) ? 1'b0 : node3043;
												assign node3043 = (inp[7]) ? 1'b0 : node3044;
													assign node3044 = (inp[12]) ? 1'b0 : 1'b1;
									assign node3049 = (inp[7]) ? node3063 : node3050;
										assign node3050 = (inp[14]) ? node3058 : node3051;
											assign node3051 = (inp[5]) ? node3053 : 1'b1;
												assign node3053 = (inp[13]) ? 1'b0 : node3054;
													assign node3054 = (inp[0]) ? 1'b0 : 1'b1;
											assign node3058 = (inp[0]) ? 1'b0 : node3059;
												assign node3059 = (inp[3]) ? 1'b0 : 1'b1;
										assign node3063 = (inp[3]) ? 1'b0 : node3064;
											assign node3064 = (inp[14]) ? 1'b0 : node3065;
												assign node3065 = (inp[12]) ? 1'b0 : 1'b1;
						assign node3070 = (inp[14]) ? node3168 : node3071;
							assign node3071 = (inp[0]) ? node3123 : node3072;
								assign node3072 = (inp[8]) ? node3094 : node3073;
									assign node3073 = (inp[9]) ? node3081 : node3074;
										assign node3074 = (inp[7]) ? node3076 : 1'b1;
											assign node3076 = (inp[13]) ? node3078 : 1'b1;
												assign node3078 = (inp[5]) ? 1'b0 : 1'b1;
										assign node3081 = (inp[3]) ? node3083 : 1'b1;
											assign node3083 = (inp[5]) ? node3089 : node3084;
												assign node3084 = (inp[7]) ? node3086 : 1'b1;
													assign node3086 = (inp[13]) ? 1'b0 : 1'b1;
												assign node3089 = (inp[7]) ? 1'b0 : node3090;
													assign node3090 = (inp[11]) ? 1'b0 : 1'b1;
									assign node3094 = (inp[3]) ? node3110 : node3095;
										assign node3095 = (inp[12]) ? node3103 : node3096;
											assign node3096 = (inp[7]) ? node3098 : 1'b1;
												assign node3098 = (inp[11]) ? node3100 : 1'b1;
													assign node3100 = (inp[5]) ? 1'b0 : 1'b1;
											assign node3103 = (inp[5]) ? 1'b0 : node3104;
												assign node3104 = (inp[9]) ? node3106 : 1'b1;
													assign node3106 = (inp[13]) ? 1'b0 : 1'b1;
										assign node3110 = (inp[5]) ? 1'b0 : node3111;
											assign node3111 = (inp[7]) ? node3117 : node3112;
												assign node3112 = (inp[9]) ? node3114 : 1'b1;
													assign node3114 = (inp[11]) ? 1'b0 : 1'b1;
												assign node3117 = (inp[13]) ? 1'b0 : node3118;
													assign node3118 = (inp[9]) ? 1'b0 : 1'b1;
								assign node3123 = (inp[13]) ? node3147 : node3124;
									assign node3124 = (inp[11]) ? node3134 : node3125;
										assign node3125 = (inp[7]) ? node3127 : 1'b1;
											assign node3127 = (inp[8]) ? node3129 : 1'b1;
												assign node3129 = (inp[3]) ? 1'b0 : node3130;
													assign node3130 = (inp[5]) ? 1'b0 : 1'b1;
										assign node3134 = (inp[3]) ? node3142 : node3135;
											assign node3135 = (inp[12]) ? node3137 : 1'b1;
												assign node3137 = (inp[5]) ? 1'b0 : node3138;
													assign node3138 = (inp[7]) ? 1'b0 : 1'b1;
											assign node3142 = (inp[9]) ? 1'b0 : node3143;
												assign node3143 = (inp[5]) ? 1'b0 : 1'b1;
									assign node3147 = (inp[12]) ? 1'b0 : node3148;
										assign node3148 = (inp[9]) ? node3160 : node3149;
											assign node3149 = (inp[8]) ? node3155 : node3150;
												assign node3150 = (inp[3]) ? node3152 : 1'b1;
													assign node3152 = (inp[11]) ? 1'b0 : 1'b1;
												assign node3155 = (inp[11]) ? 1'b0 : node3156;
													assign node3156 = (inp[5]) ? 1'b0 : 1'b1;
											assign node3160 = (inp[11]) ? 1'b0 : node3161;
												assign node3161 = (inp[8]) ? 1'b0 : node3162;
													assign node3162 = (inp[3]) ? 1'b0 : 1'b0;
							assign node3168 = (inp[0]) ? node3214 : node3169;
								assign node3169 = (inp[12]) ? node3191 : node3170;
									assign node3170 = (inp[8]) ? node3176 : node3171;
										assign node3171 = (inp[13]) ? node3173 : 1'b1;
											assign node3173 = (inp[3]) ? 1'b0 : 1'b1;
										assign node3176 = (inp[5]) ? node3184 : node3177;
											assign node3177 = (inp[11]) ? node3179 : 1'b1;
												assign node3179 = (inp[9]) ? 1'b0 : node3180;
													assign node3180 = (inp[3]) ? 1'b0 : 1'b1;
											assign node3184 = (inp[7]) ? 1'b0 : node3185;
												assign node3185 = (inp[13]) ? 1'b0 : node3186;
													assign node3186 = (inp[9]) ? 1'b0 : 1'b1;
									assign node3191 = (inp[3]) ? node3205 : node3192;
										assign node3192 = (inp[9]) ? node3198 : node3193;
											assign node3193 = (inp[11]) ? node3195 : 1'b1;
												assign node3195 = (inp[13]) ? 1'b0 : 1'b1;
											assign node3198 = (inp[7]) ? 1'b0 : node3199;
												assign node3199 = (inp[13]) ? 1'b0 : node3200;
													assign node3200 = (inp[8]) ? 1'b0 : 1'b1;
										assign node3205 = (inp[5]) ? 1'b0 : node3206;
											assign node3206 = (inp[8]) ? 1'b0 : node3207;
												assign node3207 = (inp[11]) ? 1'b0 : node3208;
													assign node3208 = (inp[9]) ? 1'b0 : 1'b1;
								assign node3214 = (inp[8]) ? 1'b0 : node3215;
									assign node3215 = (inp[3]) ? 1'b0 : node3216;
										assign node3216 = (inp[7]) ? node3222 : node3217;
											assign node3217 = (inp[13]) ? node3219 : 1'b1;
												assign node3219 = (inp[5]) ? 1'b0 : 1'b1;
											assign node3222 = (inp[9]) ? 1'b0 : node3223;
												assign node3223 = (inp[11]) ? 1'b0 : node3224;
													assign node3224 = (inp[12]) ? 1'b0 : 1'b1;
					assign node3231 = (inp[12]) ? node3411 : node3232;
						assign node3232 = (inp[7]) ? node3324 : node3233;
							assign node3233 = (inp[3]) ? node3275 : node3234;
								assign node3234 = (inp[10]) ? node3246 : node3235;
									assign node3235 = (inp[5]) ? node3237 : 1'b1;
										assign node3237 = (inp[8]) ? node3239 : 1'b1;
											assign node3239 = (inp[9]) ? 1'b0 : node3240;
												assign node3240 = (inp[11]) ? node3242 : 1'b1;
													assign node3242 = (inp[0]) ? 1'b0 : 1'b0;
									assign node3246 = (inp[13]) ? node3262 : node3247;
										assign node3247 = (inp[8]) ? node3255 : node3248;
											assign node3248 = (inp[11]) ? node3250 : 1'b1;
												assign node3250 = (inp[9]) ? node3252 : 1'b1;
													assign node3252 = (inp[5]) ? 1'b0 : 1'b1;
											assign node3255 = (inp[9]) ? 1'b0 : node3256;
												assign node3256 = (inp[14]) ? node3258 : 1'b1;
													assign node3258 = (inp[11]) ? 1'b0 : 1'b1;
										assign node3262 = (inp[5]) ? node3268 : node3263;
											assign node3263 = (inp[9]) ? node3265 : 1'b1;
												assign node3265 = (inp[14]) ? 1'b0 : 1'b1;
											assign node3268 = (inp[9]) ? 1'b0 : node3269;
												assign node3269 = (inp[11]) ? node3271 : 1'b1;
													assign node3271 = (inp[14]) ? 1'b0 : 1'b0;
								assign node3275 = (inp[14]) ? node3299 : node3276;
									assign node3276 = (inp[8]) ? node3284 : node3277;
										assign node3277 = (inp[0]) ? node3279 : 1'b1;
											assign node3279 = (inp[10]) ? node3281 : 1'b1;
												assign node3281 = (inp[5]) ? 1'b0 : 1'b1;
										assign node3284 = (inp[13]) ? node3292 : node3285;
											assign node3285 = (inp[5]) ? node3287 : 1'b1;
												assign node3287 = (inp[9]) ? 1'b0 : node3288;
													assign node3288 = (inp[10]) ? 1'b0 : 1'b1;
											assign node3292 = (inp[11]) ? 1'b0 : node3293;
												assign node3293 = (inp[0]) ? 1'b0 : node3294;
													assign node3294 = (inp[9]) ? 1'b0 : 1'b1;
									assign node3299 = (inp[9]) ? node3315 : node3300;
										assign node3300 = (inp[0]) ? node3308 : node3301;
											assign node3301 = (inp[11]) ? node3303 : 1'b1;
												assign node3303 = (inp[8]) ? 1'b0 : node3304;
													assign node3304 = (inp[10]) ? 1'b0 : 1'b1;
											assign node3308 = (inp[13]) ? 1'b0 : node3309;
												assign node3309 = (inp[11]) ? 1'b0 : node3310;
													assign node3310 = (inp[5]) ? 1'b0 : 1'b1;
										assign node3315 = (inp[8]) ? 1'b0 : node3316;
											assign node3316 = (inp[11]) ? 1'b0 : node3317;
												assign node3317 = (inp[13]) ? 1'b0 : node3318;
													assign node3318 = (inp[10]) ? 1'b0 : 1'b1;
							assign node3324 = (inp[8]) ? node3374 : node3325;
								assign node3325 = (inp[3]) ? node3351 : node3326;
									assign node3326 = (inp[9]) ? node3336 : node3327;
										assign node3327 = (inp[0]) ? node3329 : 1'b1;
											assign node3329 = (inp[14]) ? node3331 : 1'b1;
												assign node3331 = (inp[5]) ? 1'b0 : node3332;
													assign node3332 = (inp[10]) ? 1'b0 : 1'b1;
										assign node3336 = (inp[13]) ? node3344 : node3337;
											assign node3337 = (inp[14]) ? node3339 : 1'b1;
												assign node3339 = (inp[5]) ? 1'b0 : node3340;
													assign node3340 = (inp[10]) ? 1'b0 : 1'b1;
											assign node3344 = (inp[10]) ? 1'b0 : node3345;
												assign node3345 = (inp[14]) ? 1'b0 : node3346;
													assign node3346 = (inp[5]) ? 1'b0 : 1'b1;
									assign node3351 = (inp[10]) ? node3365 : node3352;
										assign node3352 = (inp[5]) ? node3358 : node3353;
											assign node3353 = (inp[0]) ? node3355 : 1'b1;
												assign node3355 = (inp[14]) ? 1'b0 : 1'b1;
											assign node3358 = (inp[14]) ? 1'b0 : node3359;
												assign node3359 = (inp[11]) ? 1'b0 : node3360;
													assign node3360 = (inp[9]) ? 1'b0 : 1'b1;
										assign node3365 = (inp[9]) ? 1'b0 : node3366;
											assign node3366 = (inp[13]) ? 1'b0 : node3367;
												assign node3367 = (inp[14]) ? 1'b0 : node3368;
													assign node3368 = (inp[0]) ? 1'b0 : 1'b1;
								assign node3374 = (inp[13]) ? node3400 : node3375;
									assign node3375 = (inp[14]) ? node3393 : node3376;
										assign node3376 = (inp[0]) ? node3388 : node3377;
											assign node3377 = (inp[5]) ? node3383 : node3378;
												assign node3378 = (inp[3]) ? node3380 : 1'b1;
													assign node3380 = (inp[10]) ? 1'b0 : 1'b1;
												assign node3383 = (inp[11]) ? 1'b0 : node3384;
													assign node3384 = (inp[10]) ? 1'b1 : 1'b0;
											assign node3388 = (inp[10]) ? 1'b0 : node3389;
												assign node3389 = (inp[11]) ? 1'b0 : 1'b1;
										assign node3393 = (inp[10]) ? 1'b0 : node3394;
											assign node3394 = (inp[9]) ? 1'b0 : node3395;
												assign node3395 = (inp[5]) ? 1'b0 : 1'b1;
									assign node3400 = (inp[9]) ? 1'b0 : node3401;
										assign node3401 = (inp[14]) ? 1'b0 : node3402;
											assign node3402 = (inp[11]) ? 1'b0 : node3403;
												assign node3403 = (inp[0]) ? 1'b0 : node3404;
													assign node3404 = (inp[3]) ? 1'b0 : 1'b1;
						assign node3411 = (inp[7]) ? node3497 : node3412;
							assign node3412 = (inp[5]) ? node3460 : node3413;
								assign node3413 = (inp[9]) ? node3445 : node3414;
									assign node3414 = (inp[11]) ? node3428 : node3415;
										assign node3415 = (inp[10]) ? node3417 : 1'b1;
											assign node3417 = (inp[0]) ? node3423 : node3418;
												assign node3418 = (inp[14]) ? node3420 : 1'b1;
													assign node3420 = (inp[8]) ? 1'b0 : 1'b1;
												assign node3423 = (inp[8]) ? 1'b0 : node3424;
													assign node3424 = (inp[14]) ? 1'b0 : 1'b1;
										assign node3428 = (inp[13]) ? node3440 : node3429;
											assign node3429 = (inp[8]) ? node3435 : node3430;
												assign node3430 = (inp[0]) ? node3432 : 1'b1;
													assign node3432 = (inp[14]) ? 1'b1 : 1'b0;
												assign node3435 = (inp[10]) ? 1'b0 : node3436;
													assign node3436 = (inp[14]) ? 1'b0 : 1'b1;
											assign node3440 = (inp[3]) ? 1'b0 : node3441;
												assign node3441 = (inp[0]) ? 1'b0 : 1'b1;
									assign node3445 = (inp[10]) ? 1'b0 : node3446;
										assign node3446 = (inp[13]) ? node3454 : node3447;
											assign node3447 = (inp[0]) ? node3449 : 1'b1;
												assign node3449 = (inp[14]) ? 1'b0 : node3450;
													assign node3450 = (inp[8]) ? 1'b0 : 1'b1;
											assign node3454 = (inp[8]) ? 1'b0 : node3455;
												assign node3455 = (inp[11]) ? 1'b0 : 1'b1;
								assign node3460 = (inp[11]) ? node3486 : node3461;
									assign node3461 = (inp[10]) ? node3479 : node3462;
										assign node3462 = (inp[8]) ? node3474 : node3463;
											assign node3463 = (inp[3]) ? node3469 : node3464;
												assign node3464 = (inp[13]) ? node3466 : 1'b1;
													assign node3466 = (inp[14]) ? 1'b0 : 1'b1;
												assign node3469 = (inp[13]) ? 1'b0 : node3470;
													assign node3470 = (inp[9]) ? 1'b0 : 1'b1;
											assign node3474 = (inp[14]) ? 1'b0 : node3475;
												assign node3475 = (inp[13]) ? 1'b0 : 1'b1;
										assign node3479 = (inp[9]) ? 1'b0 : node3480;
											assign node3480 = (inp[8]) ? 1'b0 : node3481;
												assign node3481 = (inp[14]) ? 1'b0 : 1'b1;
									assign node3486 = (inp[8]) ? 1'b0 : node3487;
										assign node3487 = (inp[0]) ? 1'b0 : node3488;
											assign node3488 = (inp[14]) ? 1'b0 : node3489;
												assign node3489 = (inp[10]) ? 1'b0 : node3490;
													assign node3490 = (inp[9]) ? 1'b0 : 1'b1;
							assign node3497 = (inp[5]) ? node3537 : node3498;
								assign node3498 = (inp[9]) ? node3528 : node3499;
									assign node3499 = (inp[10]) ? node3519 : node3500;
										assign node3500 = (inp[0]) ? node3512 : node3501;
											assign node3501 = (inp[8]) ? node3507 : node3502;
												assign node3502 = (inp[3]) ? node3504 : 1'b1;
													assign node3504 = (inp[14]) ? 1'b0 : 1'b1;
												assign node3507 = (inp[11]) ? 1'b0 : node3508;
													assign node3508 = (inp[14]) ? 1'b0 : 1'b1;
											assign node3512 = (inp[11]) ? 1'b0 : node3513;
												assign node3513 = (inp[3]) ? 1'b0 : node3514;
													assign node3514 = (inp[14]) ? 1'b0 : 1'b1;
										assign node3519 = (inp[13]) ? 1'b0 : node3520;
											assign node3520 = (inp[11]) ? 1'b0 : node3521;
												assign node3521 = (inp[8]) ? 1'b0 : node3522;
													assign node3522 = (inp[14]) ? 1'b0 : 1'b1;
									assign node3528 = (inp[13]) ? 1'b0 : node3529;
										assign node3529 = (inp[14]) ? 1'b0 : node3530;
											assign node3530 = (inp[3]) ? 1'b0 : node3531;
												assign node3531 = (inp[11]) ? 1'b0 : 1'b1;
								assign node3537 = (inp[13]) ? 1'b0 : node3538;
									assign node3538 = (inp[3]) ? 1'b0 : node3539;
										assign node3539 = (inp[8]) ? 1'b0 : node3540;
											assign node3540 = (inp[9]) ? node3542 : 1'b0;
												assign node3542 = (inp[14]) ? 1'b0 : 1'b1;
			assign node3548 = (inp[13]) ? node4212 : node3549;
				assign node3549 = (inp[0]) ? node3915 : node3550;
					assign node3550 = (inp[12]) ? node3728 : node3551;
						assign node3551 = (inp[1]) ? node3643 : node3552;
							assign node3552 = (inp[7]) ? node3584 : node3553;
								assign node3553 = (inp[3]) ? node3555 : 1'b1;
									assign node3555 = (inp[5]) ? node3565 : node3556;
										assign node3556 = (inp[8]) ? node3558 : 1'b1;
											assign node3558 = (inp[10]) ? node3560 : 1'b1;
												assign node3560 = (inp[14]) ? node3562 : 1'b1;
													assign node3562 = (inp[6]) ? 1'b0 : 1'b1;
										assign node3565 = (inp[11]) ? node3573 : node3566;
											assign node3566 = (inp[9]) ? node3568 : 1'b1;
												assign node3568 = (inp[6]) ? node3570 : 1'b1;
													assign node3570 = (inp[8]) ? 1'b0 : 1'b1;
											assign node3573 = (inp[6]) ? node3579 : node3574;
												assign node3574 = (inp[8]) ? node3576 : 1'b1;
													assign node3576 = (inp[10]) ? 1'b0 : 1'b1;
												assign node3579 = (inp[8]) ? 1'b0 : node3580;
													assign node3580 = (inp[14]) ? 1'b0 : 1'b1;
								assign node3584 = (inp[11]) ? node3614 : node3585;
									assign node3585 = (inp[3]) ? node3595 : node3586;
										assign node3586 = (inp[8]) ? node3588 : 1'b1;
											assign node3588 = (inp[9]) ? 1'b1 : node3589;
												assign node3589 = (inp[10]) ? node3591 : 1'b1;
													assign node3591 = (inp[5]) ? 1'b0 : 1'b1;
										assign node3595 = (inp[9]) ? node3603 : node3596;
											assign node3596 = (inp[14]) ? node3598 : 1'b1;
												assign node3598 = (inp[5]) ? node3600 : 1'b1;
													assign node3600 = (inp[10]) ? 1'b0 : 1'b1;
											assign node3603 = (inp[5]) ? node3609 : node3604;
												assign node3604 = (inp[8]) ? node3606 : 1'b1;
													assign node3606 = (inp[14]) ? 1'b0 : 1'b1;
												assign node3609 = (inp[6]) ? 1'b0 : node3610;
													assign node3610 = (inp[14]) ? 1'b0 : 1'b1;
									assign node3614 = (inp[14]) ? node3630 : node3615;
										assign node3615 = (inp[6]) ? node3623 : node3616;
											assign node3616 = (inp[10]) ? node3618 : 1'b1;
												assign node3618 = (inp[5]) ? node3620 : 1'b1;
													assign node3620 = (inp[8]) ? 1'b0 : 1'b1;
											assign node3623 = (inp[5]) ? 1'b0 : node3624;
												assign node3624 = (inp[3]) ? node3626 : 1'b1;
													assign node3626 = (inp[10]) ? 1'b0 : 1'b1;
										assign node3630 = (inp[3]) ? 1'b0 : node3631;
											assign node3631 = (inp[9]) ? node3637 : node3632;
												assign node3632 = (inp[6]) ? node3634 : 1'b1;
													assign node3634 = (inp[8]) ? 1'b0 : 1'b1;
												assign node3637 = (inp[10]) ? 1'b0 : node3638;
													assign node3638 = (inp[6]) ? 1'b0 : 1'b1;
							assign node3643 = (inp[5]) ? node3681 : node3644;
								assign node3644 = (inp[3]) ? node3664 : node3645;
									assign node3645 = (inp[9]) ? node3647 : 1'b1;
										assign node3647 = (inp[6]) ? node3655 : node3648;
											assign node3648 = (inp[8]) ? node3650 : 1'b1;
												assign node3650 = (inp[11]) ? node3652 : 1'b1;
													assign node3652 = (inp[7]) ? 1'b0 : 1'b1;
											assign node3655 = (inp[7]) ? node3661 : node3656;
												assign node3656 = (inp[8]) ? node3658 : 1'b1;
													assign node3658 = (inp[10]) ? 1'b0 : 1'b1;
												assign node3661 = (inp[11]) ? 1'b0 : 1'b1;
									assign node3664 = (inp[8]) ? node3676 : node3665;
										assign node3665 = (inp[11]) ? node3667 : 1'b1;
											assign node3667 = (inp[10]) ? node3671 : node3668;
												assign node3668 = (inp[14]) ? 1'b0 : 1'b1;
												assign node3671 = (inp[9]) ? 1'b0 : node3672;
													assign node3672 = (inp[14]) ? 1'b0 : 1'b1;
										assign node3676 = (inp[6]) ? 1'b0 : node3677;
											assign node3677 = (inp[10]) ? 1'b0 : 1'b1;
								assign node3681 = (inp[7]) ? node3705 : node3682;
									assign node3682 = (inp[9]) ? node3690 : node3683;
										assign node3683 = (inp[11]) ? node3685 : 1'b1;
											assign node3685 = (inp[10]) ? 1'b0 : node3686;
												assign node3686 = (inp[3]) ? 1'b0 : 1'b1;
										assign node3690 = (inp[14]) ? node3698 : node3691;
											assign node3691 = (inp[8]) ? node3693 : 1'b1;
												assign node3693 = (inp[10]) ? 1'b0 : node3694;
													assign node3694 = (inp[3]) ? 1'b0 : 1'b1;
											assign node3698 = (inp[11]) ? 1'b0 : node3699;
												assign node3699 = (inp[3]) ? 1'b0 : node3700;
													assign node3700 = (inp[8]) ? 1'b0 : 1'b1;
									assign node3705 = (inp[10]) ? node3719 : node3706;
										assign node3706 = (inp[8]) ? node3714 : node3707;
											assign node3707 = (inp[6]) ? node3709 : 1'b1;
												assign node3709 = (inp[9]) ? 1'b0 : node3710;
													assign node3710 = (inp[11]) ? 1'b0 : 1'b1;
											assign node3714 = (inp[3]) ? 1'b0 : node3715;
												assign node3715 = (inp[9]) ? 1'b0 : 1'b1;
										assign node3719 = (inp[3]) ? 1'b0 : node3720;
											assign node3720 = (inp[9]) ? 1'b0 : node3721;
												assign node3721 = (inp[14]) ? 1'b0 : node3722;
													assign node3722 = (inp[11]) ? 1'b0 : 1'b1;
						assign node3728 = (inp[3]) ? node3832 : node3729;
							assign node3729 = (inp[7]) ? node3783 : node3730;
								assign node3730 = (inp[1]) ? node3756 : node3731;
									assign node3731 = (inp[14]) ? node3741 : node3732;
										assign node3732 = (inp[11]) ? node3734 : 1'b1;
											assign node3734 = (inp[6]) ? node3736 : 1'b1;
												assign node3736 = (inp[9]) ? 1'b1 : node3737;
													assign node3737 = (inp[8]) ? 1'b0 : 1'b1;
										assign node3741 = (inp[5]) ? node3749 : node3742;
											assign node3742 = (inp[9]) ? node3744 : 1'b1;
												assign node3744 = (inp[8]) ? node3746 : 1'b1;
													assign node3746 = (inp[10]) ? 1'b0 : 1'b1;
											assign node3749 = (inp[11]) ? 1'b0 : node3750;
												assign node3750 = (inp[8]) ? node3752 : 1'b1;
													assign node3752 = (inp[6]) ? 1'b0 : 1'b1;
									assign node3756 = (inp[11]) ? node3770 : node3757;
										assign node3757 = (inp[14]) ? node3759 : 1'b1;
											assign node3759 = (inp[5]) ? node3765 : node3760;
												assign node3760 = (inp[9]) ? node3762 : 1'b1;
													assign node3762 = (inp[6]) ? 1'b0 : 1'b1;
												assign node3765 = (inp[10]) ? node3767 : 1'b0;
													assign node3767 = (inp[8]) ? 1'b0 : 1'b1;
										assign node3770 = (inp[10]) ? 1'b0 : node3771;
											assign node3771 = (inp[6]) ? node3777 : node3772;
												assign node3772 = (inp[5]) ? node3774 : 1'b1;
													assign node3774 = (inp[8]) ? 1'b0 : 1'b1;
												assign node3777 = (inp[8]) ? 1'b0 : node3778;
													assign node3778 = (inp[14]) ? 1'b0 : 1'b1;
								assign node3783 = (inp[14]) ? node3803 : node3784;
									assign node3784 = (inp[11]) ? node3794 : node3785;
										assign node3785 = (inp[10]) ? node3787 : 1'b1;
											assign node3787 = (inp[6]) ? 1'b0 : node3788;
												assign node3788 = (inp[8]) ? node3790 : 1'b1;
													assign node3790 = (inp[5]) ? 1'b0 : 1'b1;
										assign node3794 = (inp[9]) ? 1'b0 : node3795;
											assign node3795 = (inp[1]) ? 1'b0 : node3796;
												assign node3796 = (inp[10]) ? node3798 : 1'b1;
													assign node3798 = (inp[8]) ? 1'b0 : 1'b1;
									assign node3803 = (inp[8]) ? node3823 : node3804;
										assign node3804 = (inp[5]) ? node3816 : node3805;
											assign node3805 = (inp[11]) ? node3811 : node3806;
												assign node3806 = (inp[1]) ? node3808 : 1'b1;
													assign node3808 = (inp[6]) ? 1'b0 : 1'b1;
												assign node3811 = (inp[9]) ? 1'b0 : node3812;
													assign node3812 = (inp[1]) ? 1'b0 : 1'b1;
											assign node3816 = (inp[10]) ? 1'b0 : node3817;
												assign node3817 = (inp[11]) ? 1'b0 : node3818;
													assign node3818 = (inp[9]) ? 1'b0 : 1'b1;
										assign node3823 = (inp[10]) ? 1'b0 : node3824;
											assign node3824 = (inp[6]) ? 1'b0 : node3825;
												assign node3825 = (inp[1]) ? 1'b0 : node3826;
													assign node3826 = (inp[9]) ? 1'b0 : 1'b1;
							assign node3832 = (inp[6]) ? node3880 : node3833;
								assign node3833 = (inp[1]) ? node3861 : node3834;
									assign node3834 = (inp[8]) ? node3852 : node3835;
										assign node3835 = (inp[9]) ? node3843 : node3836;
											assign node3836 = (inp[5]) ? node3838 : 1'b1;
												assign node3838 = (inp[11]) ? node3840 : 1'b1;
													assign node3840 = (inp[10]) ? 1'b0 : 1'b1;
											assign node3843 = (inp[14]) ? node3847 : node3844;
												assign node3844 = (inp[11]) ? 1'b0 : 1'b1;
												assign node3847 = (inp[5]) ? 1'b0 : node3848;
													assign node3848 = (inp[7]) ? 1'b0 : 1'b1;
										assign node3852 = (inp[11]) ? node3856 : node3853;
											assign node3853 = (inp[7]) ? 1'b0 : 1'b1;
											assign node3856 = (inp[5]) ? 1'b0 : node3857;
												assign node3857 = (inp[9]) ? 1'b0 : 1'b1;
									assign node3861 = (inp[14]) ? node3871 : node3862;
										assign node3862 = (inp[7]) ? 1'b0 : node3863;
											assign node3863 = (inp[10]) ? node3865 : 1'b1;
												assign node3865 = (inp[9]) ? 1'b0 : node3866;
													assign node3866 = (inp[11]) ? 1'b0 : 1'b1;
										assign node3871 = (inp[10]) ? 1'b0 : node3872;
											assign node3872 = (inp[8]) ? 1'b0 : node3873;
												assign node3873 = (inp[5]) ? 1'b0 : node3874;
													assign node3874 = (inp[9]) ? 1'b0 : 1'b1;
								assign node3880 = (inp[11]) ? node3904 : node3881;
									assign node3881 = (inp[1]) ? node3897 : node3882;
										assign node3882 = (inp[9]) ? node3890 : node3883;
											assign node3883 = (inp[8]) ? node3885 : 1'b1;
												assign node3885 = (inp[14]) ? 1'b0 : node3886;
													assign node3886 = (inp[5]) ? 1'b0 : 1'b1;
											assign node3890 = (inp[5]) ? 1'b0 : node3891;
												assign node3891 = (inp[7]) ? 1'b0 : node3892;
													assign node3892 = (inp[10]) ? 1'b0 : 1'b1;
										assign node3897 = (inp[10]) ? 1'b0 : node3898;
											assign node3898 = (inp[8]) ? 1'b0 : node3899;
												assign node3899 = (inp[5]) ? 1'b0 : 1'b1;
									assign node3904 = (inp[14]) ? 1'b0 : node3905;
										assign node3905 = (inp[5]) ? 1'b0 : node3906;
											assign node3906 = (inp[7]) ? 1'b0 : node3907;
												assign node3907 = (inp[10]) ? 1'b0 : node3908;
													assign node3908 = (inp[8]) ? 1'b0 : 1'b1;
					assign node3915 = (inp[11]) ? node4093 : node3916;
						assign node3916 = (inp[14]) ? node4018 : node3917;
							assign node3917 = (inp[6]) ? node3963 : node3918;
								assign node3918 = (inp[1]) ? node3936 : node3919;
									assign node3919 = (inp[10]) ? node3921 : 1'b1;
										assign node3921 = (inp[5]) ? node3929 : node3922;
											assign node3922 = (inp[7]) ? node3924 : 1'b1;
												assign node3924 = (inp[3]) ? node3926 : 1'b1;
													assign node3926 = (inp[8]) ? 1'b0 : 1'b1;
											assign node3929 = (inp[8]) ? 1'b0 : node3930;
												assign node3930 = (inp[7]) ? node3932 : 1'b1;
													assign node3932 = (inp[12]) ? 1'b0 : 1'b1;
									assign node3936 = (inp[7]) ? node3946 : node3937;
										assign node3937 = (inp[12]) ? node3939 : 1'b1;
											assign node3939 = (inp[3]) ? node3941 : 1'b1;
												assign node3941 = (inp[8]) ? 1'b0 : node3942;
													assign node3942 = (inp[10]) ? 1'b0 : 1'b1;
										assign node3946 = (inp[3]) ? node3958 : node3947;
											assign node3947 = (inp[12]) ? node3953 : node3948;
												assign node3948 = (inp[9]) ? node3950 : 1'b1;
													assign node3950 = (inp[10]) ? 1'b0 : 1'b1;
												assign node3953 = (inp[10]) ? 1'b0 : node3954;
													assign node3954 = (inp[8]) ? 1'b0 : 1'b1;
											assign node3958 = (inp[5]) ? 1'b0 : node3959;
												assign node3959 = (inp[10]) ? 1'b0 : 1'b1;
								assign node3963 = (inp[10]) ? node3997 : node3964;
									assign node3964 = (inp[3]) ? node3978 : node3965;
										assign node3965 = (inp[7]) ? node3967 : 1'b1;
											assign node3967 = (inp[8]) ? node3973 : node3968;
												assign node3968 = (inp[12]) ? node3970 : 1'b1;
													assign node3970 = (inp[5]) ? 1'b0 : 1'b1;
												assign node3973 = (inp[9]) ? 1'b0 : node3974;
													assign node3974 = (inp[12]) ? 1'b0 : 1'b1;
										assign node3978 = (inp[12]) ? node3990 : node3979;
											assign node3979 = (inp[1]) ? node3985 : node3980;
												assign node3980 = (inp[8]) ? node3982 : 1'b1;
													assign node3982 = (inp[7]) ? 1'b0 : 1'b1;
												assign node3985 = (inp[9]) ? 1'b0 : node3986;
													assign node3986 = (inp[8]) ? 1'b0 : 1'b0;
											assign node3990 = (inp[5]) ? node3992 : 1'b0;
												assign node3992 = (inp[9]) ? 1'b0 : node3993;
													assign node3993 = (inp[7]) ? 1'b0 : 1'b0;
									assign node3997 = (inp[5]) ? node4011 : node3998;
										assign node3998 = (inp[7]) ? 1'b0 : node3999;
											assign node3999 = (inp[1]) ? node4005 : node4000;
												assign node4000 = (inp[12]) ? node4002 : 1'b1;
													assign node4002 = (inp[8]) ? 1'b0 : 1'b1;
												assign node4005 = (inp[9]) ? 1'b0 : node4006;
													assign node4006 = (inp[12]) ? 1'b0 : 1'b1;
										assign node4011 = (inp[12]) ? 1'b0 : node4012;
											assign node4012 = (inp[1]) ? 1'b0 : node4013;
												assign node4013 = (inp[8]) ? 1'b0 : 1'b1;
							assign node4018 = (inp[7]) ? node4064 : node4019;
								assign node4019 = (inp[3]) ? node4051 : node4020;
									assign node4020 = (inp[1]) ? node4034 : node4021;
										assign node4021 = (inp[5]) ? node4023 : 1'b1;
											assign node4023 = (inp[8]) ? node4029 : node4024;
												assign node4024 = (inp[12]) ? node4026 : 1'b1;
													assign node4026 = (inp[9]) ? 1'b0 : 1'b1;
												assign node4029 = (inp[9]) ? 1'b0 : node4030;
													assign node4030 = (inp[12]) ? 1'b0 : 1'b1;
										assign node4034 = (inp[12]) ? node4046 : node4035;
											assign node4035 = (inp[10]) ? node4041 : node4036;
												assign node4036 = (inp[8]) ? node4038 : 1'b1;
													assign node4038 = (inp[9]) ? 1'b0 : 1'b1;
												assign node4041 = (inp[6]) ? 1'b0 : node4042;
													assign node4042 = (inp[5]) ? 1'b0 : 1'b1;
											assign node4046 = (inp[10]) ? 1'b0 : node4047;
												assign node4047 = (inp[9]) ? 1'b0 : 1'b1;
									assign node4051 = (inp[10]) ? 1'b0 : node4052;
										assign node4052 = (inp[9]) ? node4058 : node4053;
											assign node4053 = (inp[5]) ? node4055 : 1'b1;
												assign node4055 = (inp[1]) ? 1'b0 : 1'b1;
											assign node4058 = (inp[12]) ? 1'b0 : node4059;
												assign node4059 = (inp[6]) ? 1'b0 : 1'b1;
								assign node4064 = (inp[10]) ? node4082 : node4065;
									assign node4065 = (inp[5]) ? 1'b0 : node4066;
										assign node4066 = (inp[1]) ? node4074 : node4067;
											assign node4067 = (inp[8]) ? node4069 : 1'b1;
												assign node4069 = (inp[9]) ? 1'b0 : node4070;
													assign node4070 = (inp[6]) ? 1'b0 : 1'b1;
											assign node4074 = (inp[12]) ? 1'b0 : node4075;
												assign node4075 = (inp[8]) ? node4077 : 1'b0;
													assign node4077 = (inp[3]) ? 1'b0 : 1'b1;
									assign node4082 = (inp[8]) ? 1'b0 : node4083;
										assign node4083 = (inp[3]) ? 1'b0 : node4084;
											assign node4084 = (inp[12]) ? 1'b0 : node4085;
												assign node4085 = (inp[6]) ? 1'b0 : node4086;
													assign node4086 = (inp[1]) ? 1'b0 : 1'b1;
						assign node4093 = (inp[9]) ? node4177 : node4094;
							assign node4094 = (inp[8]) ? node4148 : node4095;
								assign node4095 = (inp[12]) ? node4129 : node4096;
									assign node4096 = (inp[3]) ? node4110 : node4097;
										assign node4097 = (inp[1]) ? node4099 : 1'b1;
											assign node4099 = (inp[7]) ? node4105 : node4100;
												assign node4100 = (inp[6]) ? node4102 : 1'b1;
													assign node4102 = (inp[10]) ? 1'b0 : 1'b1;
												assign node4105 = (inp[14]) ? 1'b0 : node4106;
													assign node4106 = (inp[6]) ? 1'b0 : 1'b1;
										assign node4110 = (inp[10]) ? node4122 : node4111;
											assign node4111 = (inp[5]) ? node4117 : node4112;
												assign node4112 = (inp[14]) ? node4114 : 1'b1;
													assign node4114 = (inp[6]) ? 1'b0 : 1'b1;
												assign node4117 = (inp[14]) ? 1'b0 : node4118;
													assign node4118 = (inp[7]) ? 1'b0 : 1'b1;
											assign node4122 = (inp[1]) ? 1'b0 : node4123;
												assign node4123 = (inp[7]) ? 1'b0 : node4124;
													assign node4124 = (inp[6]) ? 1'b0 : 1'b1;
									assign node4129 = (inp[5]) ? 1'b0 : node4130;
										assign node4130 = (inp[10]) ? node4142 : node4131;
											assign node4131 = (inp[14]) ? node4137 : node4132;
												assign node4132 = (inp[6]) ? node4134 : 1'b1;
													assign node4134 = (inp[3]) ? 1'b0 : 1'b1;
												assign node4137 = (inp[7]) ? 1'b0 : node4138;
													assign node4138 = (inp[6]) ? 1'b0 : 1'b1;
											assign node4142 = (inp[3]) ? 1'b0 : node4143;
												assign node4143 = (inp[7]) ? 1'b0 : 1'b1;
								assign node4148 = (inp[7]) ? 1'b0 : node4149;
									assign node4149 = (inp[6]) ? node4169 : node4150;
										assign node4150 = (inp[10]) ? node4162 : node4151;
											assign node4151 = (inp[14]) ? node4157 : node4152;
												assign node4152 = (inp[3]) ? node4154 : 1'b1;
													assign node4154 = (inp[5]) ? 1'b0 : 1'b1;
												assign node4157 = (inp[1]) ? 1'b0 : node4158;
													assign node4158 = (inp[3]) ? 1'b0 : 1'b1;
											assign node4162 = (inp[1]) ? 1'b0 : node4163;
												assign node4163 = (inp[5]) ? 1'b0 : node4164;
													assign node4164 = (inp[12]) ? 1'b0 : 1'b1;
										assign node4169 = (inp[10]) ? 1'b0 : node4170;
											assign node4170 = (inp[3]) ? 1'b0 : node4171;
												assign node4171 = (inp[12]) ? 1'b0 : 1'b1;
							assign node4177 = (inp[1]) ? 1'b0 : node4178;
								assign node4178 = (inp[5]) ? node4204 : node4179;
									assign node4179 = (inp[12]) ? node4195 : node4180;
										assign node4180 = (inp[10]) ? node4188 : node4181;
											assign node4181 = (inp[6]) ? node4183 : 1'b1;
												assign node4183 = (inp[7]) ? 1'b0 : node4184;
													assign node4184 = (inp[14]) ? 1'b0 : 1'b1;
											assign node4188 = (inp[14]) ? 1'b0 : node4189;
												assign node4189 = (inp[3]) ? 1'b0 : node4190;
													assign node4190 = (inp[7]) ? 1'b1 : 1'b0;
										assign node4195 = (inp[6]) ? 1'b0 : node4196;
											assign node4196 = (inp[7]) ? 1'b0 : node4197;
												assign node4197 = (inp[14]) ? 1'b0 : node4198;
													assign node4198 = (inp[3]) ? 1'b0 : 1'b1;
									assign node4204 = (inp[3]) ? 1'b0 : node4205;
										assign node4205 = (inp[12]) ? 1'b0 : node4206;
											assign node4206 = (inp[14]) ? 1'b0 : 1'b1;
				assign node4212 = (inp[10]) ? node4454 : node4213;
					assign node4213 = (inp[0]) ? node4355 : node4214;
						assign node4214 = (inp[7]) ? node4284 : node4215;
							assign node4215 = (inp[12]) ? node4249 : node4216;
								assign node4216 = (inp[14]) ? node4230 : node4217;
									assign node4217 = (inp[6]) ? node4219 : 1'b1;
										assign node4219 = (inp[9]) ? node4221 : 1'b1;
											assign node4221 = (inp[8]) ? node4227 : node4222;
												assign node4222 = (inp[1]) ? node4224 : 1'b1;
													assign node4224 = (inp[5]) ? 1'b0 : 1'b1;
												assign node4227 = (inp[5]) ? 1'b0 : 1'b1;
									assign node4230 = (inp[5]) ? node4236 : node4231;
										assign node4231 = (inp[8]) ? node4233 : 1'b1;
											assign node4233 = (inp[9]) ? 1'b0 : 1'b1;
										assign node4236 = (inp[3]) ? 1'b0 : node4237;
											assign node4237 = (inp[11]) ? node4243 : node4238;
												assign node4238 = (inp[1]) ? node4240 : 1'b1;
													assign node4240 = (inp[8]) ? 1'b0 : 1'b1;
												assign node4243 = (inp[6]) ? 1'b0 : node4244;
													assign node4244 = (inp[1]) ? 1'b0 : 1'b1;
								assign node4249 = (inp[8]) ? node4269 : node4250;
									assign node4250 = (inp[3]) ? node4258 : node4251;
										assign node4251 = (inp[6]) ? node4253 : 1'b1;
											assign node4253 = (inp[5]) ? node4255 : 1'b1;
												assign node4255 = (inp[11]) ? 1'b0 : 1'b1;
										assign node4258 = (inp[14]) ? node4266 : node4259;
											assign node4259 = (inp[9]) ? node4261 : 1'b1;
												assign node4261 = (inp[6]) ? node4263 : 1'b1;
													assign node4263 = (inp[5]) ? 1'b0 : 1'b0;
											assign node4266 = (inp[1]) ? 1'b0 : 1'b1;
									assign node4269 = (inp[11]) ? 1'b0 : node4270;
										assign node4270 = (inp[9]) ? node4276 : node4271;
											assign node4271 = (inp[6]) ? node4273 : 1'b1;
												assign node4273 = (inp[3]) ? 1'b0 : 1'b1;
											assign node4276 = (inp[5]) ? 1'b0 : node4277;
												assign node4277 = (inp[6]) ? 1'b0 : node4278;
													assign node4278 = (inp[1]) ? 1'b0 : 1'b1;
							assign node4284 = (inp[6]) ? node4334 : node4285;
								assign node4285 = (inp[11]) ? node4317 : node4286;
									assign node4286 = (inp[9]) ? node4302 : node4287;
										assign node4287 = (inp[5]) ? node4295 : node4288;
											assign node4288 = (inp[1]) ? node4290 : 1'b1;
												assign node4290 = (inp[8]) ? node4292 : 1'b1;
													assign node4292 = (inp[14]) ? 1'b0 : 1'b1;
											assign node4295 = (inp[8]) ? 1'b0 : node4296;
												assign node4296 = (inp[3]) ? node4298 : 1'b1;
													assign node4298 = (inp[14]) ? 1'b0 : 1'b1;
										assign node4302 = (inp[12]) ? node4310 : node4303;
											assign node4303 = (inp[14]) ? node4305 : 1'b1;
												assign node4305 = (inp[1]) ? 1'b0 : node4306;
													assign node4306 = (inp[8]) ? 1'b0 : 1'b1;
											assign node4310 = (inp[3]) ? 1'b0 : node4311;
												assign node4311 = (inp[8]) ? 1'b0 : node4312;
													assign node4312 = (inp[14]) ? 1'b0 : 1'b1;
									assign node4317 = (inp[8]) ? 1'b0 : node4318;
										assign node4318 = (inp[3]) ? node4328 : node4319;
											assign node4319 = (inp[12]) ? node4325 : node4320;
												assign node4320 = (inp[1]) ? node4322 : 1'b1;
													assign node4322 = (inp[14]) ? 1'b0 : 1'b1;
												assign node4325 = (inp[9]) ? 1'b0 : 1'b1;
											assign node4328 = (inp[1]) ? 1'b0 : node4329;
												assign node4329 = (inp[9]) ? 1'b1 : 1'b0;
								assign node4334 = (inp[1]) ? 1'b0 : node4335;
									assign node4335 = (inp[9]) ? 1'b0 : node4336;
										assign node4336 = (inp[8]) ? node4348 : node4337;
											assign node4337 = (inp[12]) ? node4343 : node4338;
												assign node4338 = (inp[14]) ? node4340 : 1'b1;
													assign node4340 = (inp[3]) ? 1'b0 : 1'b1;
												assign node4343 = (inp[3]) ? 1'b0 : node4344;
													assign node4344 = (inp[14]) ? 1'b0 : 1'b1;
											assign node4348 = (inp[3]) ? 1'b0 : node4349;
												assign node4349 = (inp[11]) ? 1'b0 : 1'b1;
						assign node4355 = (inp[1]) ? node4427 : node4356;
							assign node4356 = (inp[11]) ? node4402 : node4357;
								assign node4357 = (inp[5]) ? node4381 : node4358;
									assign node4358 = (inp[12]) ? node4372 : node4359;
										assign node4359 = (inp[8]) ? node4361 : 1'b1;
											assign node4361 = (inp[9]) ? node4367 : node4362;
												assign node4362 = (inp[3]) ? node4364 : 1'b1;
													assign node4364 = (inp[7]) ? 1'b0 : 1'b1;
												assign node4367 = (inp[7]) ? 1'b0 : node4368;
													assign node4368 = (inp[3]) ? 1'b0 : 1'b1;
										assign node4372 = (inp[3]) ? 1'b0 : node4373;
											assign node4373 = (inp[7]) ? node4375 : 1'b1;
												assign node4375 = (inp[6]) ? 1'b0 : node4376;
													assign node4376 = (inp[8]) ? 1'b0 : 1'b1;
									assign node4381 = (inp[14]) ? 1'b0 : node4382;
										assign node4382 = (inp[8]) ? node4394 : node4383;
											assign node4383 = (inp[9]) ? node4389 : node4384;
												assign node4384 = (inp[7]) ? node4386 : 1'b1;
													assign node4386 = (inp[6]) ? 1'b0 : 1'b1;
												assign node4389 = (inp[12]) ? 1'b0 : node4390;
													assign node4390 = (inp[6]) ? 1'b0 : 1'b1;
											assign node4394 = (inp[6]) ? 1'b0 : node4395;
												assign node4395 = (inp[9]) ? node4397 : 1'b0;
													assign node4397 = (inp[7]) ? 1'b0 : 1'b1;
								assign node4402 = (inp[12]) ? 1'b0 : node4403;
									assign node4403 = (inp[8]) ? node4419 : node4404;
										assign node4404 = (inp[5]) ? node4412 : node4405;
											assign node4405 = (inp[9]) ? node4407 : 1'b1;
												assign node4407 = (inp[6]) ? 1'b0 : node4408;
													assign node4408 = (inp[7]) ? 1'b0 : 1'b1;
											assign node4412 = (inp[7]) ? 1'b0 : node4413;
												assign node4413 = (inp[6]) ? 1'b0 : node4414;
													assign node4414 = (inp[9]) ? 1'b0 : 1'b1;
										assign node4419 = (inp[7]) ? 1'b0 : node4420;
											assign node4420 = (inp[14]) ? 1'b0 : node4421;
												assign node4421 = (inp[5]) ? 1'b0 : 1'b1;
							assign node4427 = (inp[14]) ? 1'b0 : node4428;
								assign node4428 = (inp[7]) ? 1'b0 : node4429;
									assign node4429 = (inp[9]) ? node4445 : node4430;
										assign node4430 = (inp[5]) ? node4438 : node4431;
											assign node4431 = (inp[6]) ? node4433 : 1'b1;
												assign node4433 = (inp[8]) ? 1'b0 : node4434;
													assign node4434 = (inp[3]) ? 1'b0 : 1'b1;
											assign node4438 = (inp[12]) ? 1'b0 : node4439;
												assign node4439 = (inp[8]) ? 1'b0 : node4440;
													assign node4440 = (inp[11]) ? 1'b0 : 1'b1;
										assign node4445 = (inp[12]) ? 1'b0 : node4446;
											assign node4446 = (inp[5]) ? 1'b0 : node4447;
												assign node4447 = (inp[8]) ? 1'b0 : 1'b1;
					assign node4454 = (inp[3]) ? node4570 : node4455;
						assign node4455 = (inp[9]) ? node4537 : node4456;
							assign node4456 = (inp[7]) ? node4498 : node4457;
								assign node4457 = (inp[11]) ? node4479 : node4458;
									assign node4458 = (inp[0]) ? node4466 : node4459;
										assign node4459 = (inp[5]) ? node4461 : 1'b1;
											assign node4461 = (inp[14]) ? node4463 : 1'b1;
												assign node4463 = (inp[1]) ? 1'b0 : 1'b1;
										assign node4466 = (inp[6]) ? node4472 : node4467;
											assign node4467 = (inp[1]) ? node4469 : 1'b1;
												assign node4469 = (inp[8]) ? 1'b0 : 1'b1;
											assign node4472 = (inp[5]) ? 1'b0 : node4473;
												assign node4473 = (inp[1]) ? 1'b0 : node4474;
													assign node4474 = (inp[14]) ? 1'b0 : 1'b1;
									assign node4479 = (inp[8]) ? node4491 : node4480;
										assign node4480 = (inp[6]) ? node4486 : node4481;
											assign node4481 = (inp[14]) ? node4483 : 1'b1;
												assign node4483 = (inp[12]) ? 1'b0 : 1'b1;
											assign node4486 = (inp[5]) ? 1'b0 : node4487;
												assign node4487 = (inp[0]) ? 1'b0 : 1'b1;
										assign node4491 = (inp[1]) ? 1'b0 : node4492;
											assign node4492 = (inp[12]) ? 1'b0 : node4493;
												assign node4493 = (inp[5]) ? 1'b0 : 1'b1;
								assign node4498 = (inp[8]) ? node4528 : node4499;
									assign node4499 = (inp[12]) ? node4519 : node4500;
										assign node4500 = (inp[5]) ? node4512 : node4501;
											assign node4501 = (inp[14]) ? node4507 : node4502;
												assign node4502 = (inp[1]) ? node4504 : 1'b1;
													assign node4504 = (inp[0]) ? 1'b0 : 1'b1;
												assign node4507 = (inp[6]) ? 1'b0 : node4508;
													assign node4508 = (inp[1]) ? 1'b0 : 1'b1;
											assign node4512 = (inp[14]) ? 1'b0 : node4513;
												assign node4513 = (inp[11]) ? 1'b0 : node4514;
													assign node4514 = (inp[1]) ? 1'b0 : 1'b1;
										assign node4519 = (inp[6]) ? 1'b0 : node4520;
											assign node4520 = (inp[0]) ? 1'b0 : node4521;
												assign node4521 = (inp[11]) ? 1'b0 : node4522;
													assign node4522 = (inp[5]) ? 1'b0 : 1'b1;
									assign node4528 = (inp[0]) ? 1'b0 : node4529;
										assign node4529 = (inp[1]) ? 1'b0 : node4530;
											assign node4530 = (inp[14]) ? 1'b0 : node4531;
												assign node4531 = (inp[11]) ? 1'b0 : 1'b1;
							assign node4537 = (inp[5]) ? 1'b0 : node4538;
								assign node4538 = (inp[12]) ? node4560 : node4539;
									assign node4539 = (inp[8]) ? node4553 : node4540;
										assign node4540 = (inp[6]) ? node4546 : node4541;
											assign node4541 = (inp[11]) ? node4543 : 1'b1;
												assign node4543 = (inp[7]) ? 1'b0 : 1'b1;
											assign node4546 = (inp[14]) ? 1'b0 : node4547;
												assign node4547 = (inp[1]) ? 1'b0 : node4548;
													assign node4548 = (inp[11]) ? 1'b0 : 1'b1;
										assign node4553 = (inp[7]) ? 1'b0 : node4554;
											assign node4554 = (inp[6]) ? 1'b0 : node4555;
												assign node4555 = (inp[0]) ? 1'b0 : 1'b1;
									assign node4560 = (inp[11]) ? 1'b0 : node4561;
										assign node4561 = (inp[1]) ? 1'b0 : node4562;
											assign node4562 = (inp[8]) ? 1'b0 : node4563;
												assign node4563 = (inp[6]) ? 1'b0 : 1'b1;
						assign node4570 = (inp[12]) ? node4610 : node4571;
							assign node4571 = (inp[9]) ? node4599 : node4572;
								assign node4572 = (inp[11]) ? node4590 : node4573;
									assign node4573 = (inp[5]) ? node4583 : node4574;
										assign node4574 = (inp[8]) ? 1'b0 : node4575;
											assign node4575 = (inp[6]) ? node4577 : 1'b1;
												assign node4577 = (inp[1]) ? 1'b0 : node4578;
													assign node4578 = (inp[0]) ? 1'b0 : 1'b1;
										assign node4583 = (inp[6]) ? 1'b0 : node4584;
											assign node4584 = (inp[14]) ? 1'b0 : node4585;
												assign node4585 = (inp[8]) ? 1'b1 : 1'b0;
									assign node4590 = (inp[0]) ? 1'b0 : node4591;
										assign node4591 = (inp[7]) ? 1'b0 : node4592;
											assign node4592 = (inp[1]) ? 1'b0 : node4593;
												assign node4593 = (inp[6]) ? 1'b0 : 1'b1;
								assign node4599 = (inp[0]) ? 1'b0 : node4600;
									assign node4600 = (inp[7]) ? node4602 : 1'b0;
										assign node4602 = (inp[8]) ? 1'b0 : node4603;
											assign node4603 = (inp[5]) ? 1'b0 : node4604;
												assign node4604 = (inp[6]) ? 1'b0 : 1'b1;
							assign node4610 = (inp[1]) ? 1'b0 : node4611;
								assign node4611 = (inp[11]) ? 1'b0 : node4612;
									assign node4612 = (inp[6]) ? 1'b0 : node4613;
										assign node4613 = (inp[14]) ? 1'b0 : node4614;
											assign node4614 = (inp[0]) ? 1'b0 : node4615;
												assign node4615 = (inp[7]) ? 1'b0 : node4616;
													assign node4616 = (inp[9]) ? 1'b0 : 1'b1;

endmodule