module dtc_split66_bm58 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node61;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node204;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node265;
	wire [3-1:0] node268;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node284;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node292;
	wire [3-1:0] node296;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node316;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node322;
	wire [3-1:0] node325;
	wire [3-1:0] node326;

	assign outp = (inp[6]) ? node2 : 3'b000;
		assign node2 = (inp[0]) ? node208 : node3;
			assign node3 = (inp[4]) ? node87 : node4;
				assign node4 = (inp[9]) ? node34 : node5;
					assign node5 = (inp[1]) ? 3'b000 : node6;
						assign node6 = (inp[8]) ? node22 : node7;
							assign node7 = (inp[11]) ? 3'b000 : node8;
								assign node8 = (inp[10]) ? node14 : node9;
									assign node9 = (inp[2]) ? node11 : 3'b000;
										assign node11 = (inp[3]) ? 3'b000 : 3'b100;
									assign node14 = (inp[7]) ? node16 : 3'b100;
										assign node16 = (inp[2]) ? 3'b100 : node17;
											assign node17 = (inp[3]) ? 3'b000 : 3'b100;
							assign node22 = (inp[11]) ? node24 : 3'b100;
								assign node24 = (inp[3]) ? node26 : 3'b100;
									assign node26 = (inp[10]) ? node28 : 3'b000;
										assign node28 = (inp[7]) ? node30 : 3'b100;
											assign node30 = (inp[2]) ? 3'b100 : 3'b000;
					assign node34 = (inp[1]) ? node70 : node35;
						assign node35 = (inp[10]) ? node53 : node36;
							assign node36 = (inp[8]) ? node44 : node37;
								assign node37 = (inp[11]) ? 3'b100 : node38;
									assign node38 = (inp[3]) ? node40 : 3'b000;
										assign node40 = (inp[2]) ? 3'b000 : 3'b100;
								assign node44 = (inp[2]) ? node46 : 3'b000;
									assign node46 = (inp[5]) ? 3'b000 : node47;
										assign node47 = (inp[3]) ? 3'b000 : node48;
											assign node48 = (inp[11]) ? 3'b000 : 3'b100;
							assign node53 = (inp[8]) ? node61 : node54;
								assign node54 = (inp[3]) ? node56 : 3'b000;
									assign node56 = (inp[2]) ? 3'b000 : node57;
										assign node57 = (inp[11]) ? 3'b100 : 3'b000;
								assign node61 = (inp[11]) ? node63 : 3'b100;
									assign node63 = (inp[2]) ? 3'b100 : node64;
										assign node64 = (inp[7]) ? 3'b000 : node65;
											assign node65 = (inp[3]) ? 3'b000 : 3'b100;
						assign node70 = (inp[8]) ? node72 : 3'b100;
							assign node72 = (inp[10]) ? node80 : node73;
								assign node73 = (inp[11]) ? 3'b100 : node74;
									assign node74 = (inp[2]) ? 3'b000 : node75;
										assign node75 = (inp[3]) ? 3'b100 : 3'b000;
								assign node80 = (inp[2]) ? 3'b000 : node81;
									assign node81 = (inp[11]) ? node83 : 3'b000;
										assign node83 = (inp[3]) ? 3'b100 : 3'b000;
				assign node87 = (inp[9]) ? node123 : node88;
					assign node88 = (inp[1]) ? node90 : 3'b100;
						assign node90 = (inp[8]) ? node106 : node91;
							assign node91 = (inp[11]) ? 3'b000 : node92;
								assign node92 = (inp[3]) ? node100 : node93;
									assign node93 = (inp[7]) ? node95 : 3'b100;
										assign node95 = (inp[2]) ? 3'b100 : node96;
											assign node96 = (inp[10]) ? 3'b100 : 3'b000;
									assign node100 = (inp[10]) ? node102 : 3'b000;
										assign node102 = (inp[2]) ? 3'b100 : 3'b000;
							assign node106 = (inp[11]) ? node108 : 3'b100;
								assign node108 = (inp[10]) ? node116 : node109;
									assign node109 = (inp[3]) ? 3'b000 : node110;
										assign node110 = (inp[2]) ? 3'b100 : node111;
											assign node111 = (inp[7]) ? 3'b000 : 3'b100;
									assign node116 = (inp[2]) ? 3'b100 : node117;
										assign node117 = (inp[7]) ? node119 : 3'b100;
											assign node119 = (inp[3]) ? 3'b000 : 3'b100;
					assign node123 = (inp[8]) ? node169 : node124;
						assign node124 = (inp[1]) ? node148 : node125;
							assign node125 = (inp[10]) ? node135 : node126;
								assign node126 = (inp[3]) ? 3'b001 : node127;
									assign node127 = (inp[11]) ? node131 : node128;
										assign node128 = (inp[2]) ? 3'b101 : 3'b001;
										assign node131 = (inp[2]) ? 3'b001 : 3'b100;
								assign node135 = (inp[11]) ? node141 : node136;
									assign node136 = (inp[3]) ? 3'b101 : node137;
										assign node137 = (inp[2]) ? 3'b101 : 3'b001;
									assign node141 = (inp[2]) ? 3'b001 : node142;
										assign node142 = (inp[3]) ? node144 : 3'b101;
											assign node144 = (inp[7]) ? 3'b001 : 3'b101;
							assign node148 = (inp[10]) ? node162 : node149;
								assign node149 = (inp[11]) ? node157 : node150;
									assign node150 = (inp[7]) ? node152 : 3'b100;
										assign node152 = (inp[2]) ? 3'b100 : node153;
											assign node153 = (inp[3]) ? 3'b000 : 3'b100;
									assign node157 = (inp[3]) ? 3'b000 : node158;
										assign node158 = (inp[2]) ? 3'b100 : 3'b000;
								assign node162 = (inp[11]) ? node166 : node163;
									assign node163 = (inp[2]) ? 3'b101 : 3'b001;
									assign node166 = (inp[2]) ? 3'b001 : 3'b100;
						assign node169 = (inp[2]) ? node199 : node170;
							assign node170 = (inp[10]) ? node192 : node171;
								assign node171 = (inp[1]) ? node181 : node172;
									assign node172 = (inp[11]) ? node176 : node173;
										assign node173 = (inp[3]) ? 3'b100 : 3'b000;
										assign node176 = (inp[7]) ? 3'b000 : node177;
											assign node177 = (inp[3]) ? 3'b000 : 3'b100;
									assign node181 = (inp[5]) ? node183 : 3'b001;
										assign node183 = (inp[7]) ? node189 : node184;
											assign node184 = (inp[3]) ? 3'b101 : node185;
												assign node185 = (inp[11]) ? 3'b001 : 3'b101;
											assign node189 = (inp[11]) ? 3'b101 : 3'b001;
								assign node192 = (inp[11]) ? node196 : node193;
									assign node193 = (inp[7]) ? 3'b011 : 3'b111;
									assign node196 = (inp[7]) ? 3'b010 : 3'b110;
							assign node199 = (inp[10]) ? 3'b000 : node200;
								assign node200 = (inp[1]) ? node204 : node201;
									assign node201 = (inp[3]) ? 3'b001 : 3'b101;
									assign node204 = (inp[3]) ? 3'b000 : 3'b100;
			assign node208 = (inp[9]) ? node210 : 3'b000;
				assign node210 = (inp[1]) ? node284 : node211;
					assign node211 = (inp[4]) ? node235 : node212;
						assign node212 = (inp[8]) ? node224 : node213;
							assign node213 = (inp[11]) ? 3'b000 : node214;
								assign node214 = (inp[10]) ? 3'b100 : node215;
									assign node215 = (inp[3]) ? 3'b000 : node216;
										assign node216 = (inp[2]) ? 3'b100 : node217;
											assign node217 = (inp[7]) ? 3'b000 : 3'b100;
							assign node224 = (inp[3]) ? node226 : 3'b100;
								assign node226 = (inp[11]) ? node228 : 3'b100;
									assign node228 = (inp[10]) ? node230 : 3'b000;
										assign node230 = (inp[7]) ? node232 : 3'b100;
											assign node232 = (inp[2]) ? 3'b100 : 3'b000;
						assign node235 = (inp[8]) ? node257 : node236;
							assign node236 = (inp[10]) ? node244 : node237;
								assign node237 = (inp[11]) ? 3'b100 : node238;
									assign node238 = (inp[2]) ? 3'b000 : node239;
										assign node239 = (inp[3]) ? 3'b100 : 3'b000;
								assign node244 = (inp[11]) ? node252 : node245;
									assign node245 = (inp[2]) ? 3'b100 : node246;
										assign node246 = (inp[3]) ? 3'b000 : node247;
											assign node247 = (inp[7]) ? 3'b000 : 3'b100;
									assign node252 = (inp[2]) ? 3'b000 : node253;
										assign node253 = (inp[3]) ? 3'b100 : 3'b000;
							assign node257 = (inp[10]) ? node275 : node258;
								assign node258 = (inp[3]) ? node268 : node259;
									assign node259 = (inp[11]) ? node265 : node260;
										assign node260 = (inp[2]) ? 3'b101 : node261;
											assign node261 = (inp[7]) ? 3'b001 : 3'b101;
										assign node265 = (inp[2]) ? 3'b101 : 3'b100;
									assign node268 = (inp[7]) ? node270 : 3'b001;
										assign node270 = (inp[11]) ? node272 : 3'b001;
											assign node272 = (inp[2]) ? 3'b001 : 3'b000;
								assign node275 = (inp[2]) ? 3'b000 : node276;
									assign node276 = (inp[11]) ? node280 : node277;
										assign node277 = (inp[7]) ? 3'b001 : 3'b101;
										assign node280 = (inp[7]) ? 3'b000 : 3'b100;
					assign node284 = (inp[4]) ? node286 : 3'b000;
						assign node286 = (inp[11]) ? node316 : node287;
							assign node287 = (inp[8]) ? node303 : node288;
								assign node288 = (inp[10]) ? node296 : node289;
									assign node289 = (inp[3]) ? 3'b000 : node290;
										assign node290 = (inp[7]) ? node292 : 3'b100;
											assign node292 = (inp[2]) ? 3'b100 : 3'b000;
									assign node296 = (inp[7]) ? node298 : 3'b100;
										assign node298 = (inp[2]) ? 3'b100 : node299;
											assign node299 = (inp[3]) ? 3'b000 : 3'b100;
								assign node303 = (inp[2]) ? node311 : node304;
									assign node304 = (inp[10]) ? node308 : node305;
										assign node305 = (inp[3]) ? 3'b100 : 3'b000;
										assign node308 = (inp[7]) ? 3'b001 : 3'b101;
									assign node311 = (inp[3]) ? 3'b000 : node312;
										assign node312 = (inp[10]) ? 3'b000 : 3'b100;
							assign node316 = (inp[8]) ? node318 : 3'b000;
								assign node318 = (inp[7]) ? 3'b000 : node319;
									assign node319 = (inp[2]) ? node325 : node320;
										assign node320 = (inp[3]) ? node322 : 3'b100;
											assign node322 = (inp[10]) ? 3'b100 : 3'b000;
										assign node325 = (inp[3]) ? 3'b000 : node326;
											assign node326 = (inp[10]) ? 3'b000 : 3'b100;

endmodule