module dtc_split66_bm61 (
	input  wire [12-1:0] inp,
	output wire [11-1:0] outp
);

	wire [11-1:0] node1;
	wire [11-1:0] node2;
	wire [11-1:0] node3;
	wire [11-1:0] node4;
	wire [11-1:0] node5;
	wire [11-1:0] node6;
	wire [11-1:0] node7;
	wire [11-1:0] node8;
	wire [11-1:0] node9;
	wire [11-1:0] node10;
	wire [11-1:0] node14;
	wire [11-1:0] node15;
	wire [11-1:0] node16;
	wire [11-1:0] node19;
	wire [11-1:0] node22;
	wire [11-1:0] node25;
	wire [11-1:0] node26;
	wire [11-1:0] node27;
	wire [11-1:0] node28;
	wire [11-1:0] node31;
	wire [11-1:0] node34;
	wire [11-1:0] node37;
	wire [11-1:0] node38;
	wire [11-1:0] node39;
	wire [11-1:0] node42;
	wire [11-1:0] node45;
	wire [11-1:0] node47;
	wire [11-1:0] node50;
	wire [11-1:0] node51;
	wire [11-1:0] node52;
	wire [11-1:0] node53;
	wire [11-1:0] node54;
	wire [11-1:0] node57;
	wire [11-1:0] node60;
	wire [11-1:0] node63;
	wire [11-1:0] node64;
	wire [11-1:0] node66;
	wire [11-1:0] node69;
	wire [11-1:0] node71;
	wire [11-1:0] node74;
	wire [11-1:0] node75;
	wire [11-1:0] node76;
	wire [11-1:0] node77;
	wire [11-1:0] node82;
	wire [11-1:0] node83;
	wire [11-1:0] node85;
	wire [11-1:0] node88;
	wire [11-1:0] node89;
	wire [11-1:0] node93;
	wire [11-1:0] node94;
	wire [11-1:0] node95;
	wire [11-1:0] node96;
	wire [11-1:0] node97;
	wire [11-1:0] node99;
	wire [11-1:0] node102;
	wire [11-1:0] node103;
	wire [11-1:0] node106;
	wire [11-1:0] node109;
	wire [11-1:0] node110;
	wire [11-1:0] node113;
	wire [11-1:0] node116;
	wire [11-1:0] node117;
	wire [11-1:0] node118;
	wire [11-1:0] node121;
	wire [11-1:0] node123;
	wire [11-1:0] node126;
	wire [11-1:0] node127;
	wire [11-1:0] node128;
	wire [11-1:0] node131;
	wire [11-1:0] node134;
	wire [11-1:0] node135;
	wire [11-1:0] node139;
	wire [11-1:0] node140;
	wire [11-1:0] node141;
	wire [11-1:0] node142;
	wire [11-1:0] node143;
	wire [11-1:0] node146;
	wire [11-1:0] node149;
	wire [11-1:0] node152;
	wire [11-1:0] node153;
	wire [11-1:0] node156;
	wire [11-1:0] node157;
	wire [11-1:0] node161;
	wire [11-1:0] node162;
	wire [11-1:0] node163;
	wire [11-1:0] node164;
	wire [11-1:0] node167;
	wire [11-1:0] node170;
	wire [11-1:0] node172;
	wire [11-1:0] node175;
	wire [11-1:0] node177;
	wire [11-1:0] node180;
	wire [11-1:0] node181;
	wire [11-1:0] node182;
	wire [11-1:0] node183;
	wire [11-1:0] node184;
	wire [11-1:0] node185;
	wire [11-1:0] node187;
	wire [11-1:0] node190;
	wire [11-1:0] node193;
	wire [11-1:0] node194;
	wire [11-1:0] node196;
	wire [11-1:0] node199;
	wire [11-1:0] node202;
	wire [11-1:0] node203;
	wire [11-1:0] node204;
	wire [11-1:0] node205;
	wire [11-1:0] node208;
	wire [11-1:0] node211;
	wire [11-1:0] node214;
	wire [11-1:0] node215;
	wire [11-1:0] node216;
	wire [11-1:0] node219;
	wire [11-1:0] node223;
	wire [11-1:0] node224;
	wire [11-1:0] node225;
	wire [11-1:0] node226;
	wire [11-1:0] node227;
	wire [11-1:0] node231;
	wire [11-1:0] node234;
	wire [11-1:0] node235;
	wire [11-1:0] node236;
	wire [11-1:0] node240;
	wire [11-1:0] node241;
	wire [11-1:0] node245;
	wire [11-1:0] node246;
	wire [11-1:0] node247;
	wire [11-1:0] node250;
	wire [11-1:0] node251;
	wire [11-1:0] node255;
	wire [11-1:0] node258;
	wire [11-1:0] node259;
	wire [11-1:0] node260;
	wire [11-1:0] node261;
	wire [11-1:0] node263;
	wire [11-1:0] node264;
	wire [11-1:0] node268;
	wire [11-1:0] node270;
	wire [11-1:0] node271;
	wire [11-1:0] node275;
	wire [11-1:0] node276;
	wire [11-1:0] node278;
	wire [11-1:0] node281;
	wire [11-1:0] node282;
	wire [11-1:0] node284;
	wire [11-1:0] node287;
	wire [11-1:0] node290;
	wire [11-1:0] node291;
	wire [11-1:0] node292;
	wire [11-1:0] node293;
	wire [11-1:0] node296;
	wire [11-1:0] node299;
	wire [11-1:0] node300;
	wire [11-1:0] node301;
	wire [11-1:0] node304;
	wire [11-1:0] node307;
	wire [11-1:0] node310;
	wire [11-1:0] node311;
	wire [11-1:0] node313;
	wire [11-1:0] node314;
	wire [11-1:0] node318;
	wire [11-1:0] node320;
	wire [11-1:0] node323;
	wire [11-1:0] node324;
	wire [11-1:0] node325;
	wire [11-1:0] node326;
	wire [11-1:0] node327;
	wire [11-1:0] node328;
	wire [11-1:0] node329;
	wire [11-1:0] node330;
	wire [11-1:0] node334;
	wire [11-1:0] node335;
	wire [11-1:0] node338;
	wire [11-1:0] node341;
	wire [11-1:0] node342;
	wire [11-1:0] node345;
	wire [11-1:0] node348;
	wire [11-1:0] node349;
	wire [11-1:0] node350;
	wire [11-1:0] node351;
	wire [11-1:0] node355;
	wire [11-1:0] node356;
	wire [11-1:0] node359;
	wire [11-1:0] node362;
	wire [11-1:0] node363;
	wire [11-1:0] node366;
	wire [11-1:0] node368;
	wire [11-1:0] node371;
	wire [11-1:0] node372;
	wire [11-1:0] node373;
	wire [11-1:0] node374;
	wire [11-1:0] node377;
	wire [11-1:0] node378;
	wire [11-1:0] node382;
	wire [11-1:0] node383;
	wire [11-1:0] node385;
	wire [11-1:0] node388;
	wire [11-1:0] node391;
	wire [11-1:0] node392;
	wire [11-1:0] node393;
	wire [11-1:0] node395;
	wire [11-1:0] node398;
	wire [11-1:0] node401;
	wire [11-1:0] node402;
	wire [11-1:0] node403;
	wire [11-1:0] node406;
	wire [11-1:0] node409;
	wire [11-1:0] node410;
	wire [11-1:0] node414;
	wire [11-1:0] node415;
	wire [11-1:0] node416;
	wire [11-1:0] node417;
	wire [11-1:0] node418;
	wire [11-1:0] node421;
	wire [11-1:0] node422;
	wire [11-1:0] node425;
	wire [11-1:0] node428;
	wire [11-1:0] node429;
	wire [11-1:0] node431;
	wire [11-1:0] node435;
	wire [11-1:0] node436;
	wire [11-1:0] node437;
	wire [11-1:0] node438;
	wire [11-1:0] node441;
	wire [11-1:0] node444;
	wire [11-1:0] node446;
	wire [11-1:0] node449;
	wire [11-1:0] node450;
	wire [11-1:0] node452;
	wire [11-1:0] node455;
	wire [11-1:0] node458;
	wire [11-1:0] node459;
	wire [11-1:0] node460;
	wire [11-1:0] node461;
	wire [11-1:0] node463;
	wire [11-1:0] node466;
	wire [11-1:0] node469;
	wire [11-1:0] node470;
	wire [11-1:0] node471;
	wire [11-1:0] node475;
	wire [11-1:0] node476;
	wire [11-1:0] node479;
	wire [11-1:0] node482;
	wire [11-1:0] node483;
	wire [11-1:0] node484;
	wire [11-1:0] node486;
	wire [11-1:0] node489;
	wire [11-1:0] node492;
	wire [11-1:0] node493;
	wire [11-1:0] node496;
	wire [11-1:0] node498;
	wire [11-1:0] node501;
	wire [11-1:0] node502;
	wire [11-1:0] node503;
	wire [11-1:0] node504;
	wire [11-1:0] node505;
	wire [11-1:0] node506;
	wire [11-1:0] node510;
	wire [11-1:0] node511;
	wire [11-1:0] node512;
	wire [11-1:0] node516;
	wire [11-1:0] node517;
	wire [11-1:0] node521;
	wire [11-1:0] node522;
	wire [11-1:0] node523;
	wire [11-1:0] node524;
	wire [11-1:0] node528;
	wire [11-1:0] node529;
	wire [11-1:0] node532;
	wire [11-1:0] node535;
	wire [11-1:0] node536;
	wire [11-1:0] node537;
	wire [11-1:0] node541;
	wire [11-1:0] node544;
	wire [11-1:0] node545;
	wire [11-1:0] node546;
	wire [11-1:0] node547;
	wire [11-1:0] node548;
	wire [11-1:0] node552;
	wire [11-1:0] node555;
	wire [11-1:0] node557;
	wire [11-1:0] node559;
	wire [11-1:0] node562;
	wire [11-1:0] node563;
	wire [11-1:0] node564;
	wire [11-1:0] node567;
	wire [11-1:0] node570;
	wire [11-1:0] node571;
	wire [11-1:0] node572;
	wire [11-1:0] node576;
	wire [11-1:0] node578;
	wire [11-1:0] node581;
	wire [11-1:0] node582;
	wire [11-1:0] node583;
	wire [11-1:0] node584;
	wire [11-1:0] node586;
	wire [11-1:0] node589;
	wire [11-1:0] node590;
	wire [11-1:0] node592;
	wire [11-1:0] node595;
	wire [11-1:0] node596;
	wire [11-1:0] node599;
	wire [11-1:0] node602;
	wire [11-1:0] node603;
	wire [11-1:0] node604;
	wire [11-1:0] node605;
	wire [11-1:0] node608;
	wire [11-1:0] node611;
	wire [11-1:0] node613;
	wire [11-1:0] node616;
	wire [11-1:0] node617;
	wire [11-1:0] node619;
	wire [11-1:0] node622;
	wire [11-1:0] node623;
	wire [11-1:0] node627;
	wire [11-1:0] node628;
	wire [11-1:0] node629;
	wire [11-1:0] node630;
	wire [11-1:0] node633;
	wire [11-1:0] node635;
	wire [11-1:0] node638;
	wire [11-1:0] node639;
	wire [11-1:0] node640;
	wire [11-1:0] node643;
	wire [11-1:0] node646;
	wire [11-1:0] node647;
	wire [11-1:0] node651;
	wire [11-1:0] node652;
	wire [11-1:0] node653;
	wire [11-1:0] node654;
	wire [11-1:0] node658;
	wire [11-1:0] node659;
	wire [11-1:0] node662;
	wire [11-1:0] node665;
	wire [11-1:0] node666;
	wire [11-1:0] node668;
	wire [11-1:0] node671;
	wire [11-1:0] node673;
	wire [11-1:0] node676;
	wire [11-1:0] node677;
	wire [11-1:0] node678;
	wire [11-1:0] node679;
	wire [11-1:0] node680;
	wire [11-1:0] node681;
	wire [11-1:0] node682;
	wire [11-1:0] node683;
	wire [11-1:0] node687;
	wire [11-1:0] node688;
	wire [11-1:0] node691;
	wire [11-1:0] node692;
	wire [11-1:0] node695;
	wire [11-1:0] node698;
	wire [11-1:0] node699;
	wire [11-1:0] node700;
	wire [11-1:0] node701;
	wire [11-1:0] node705;
	wire [11-1:0] node707;
	wire [11-1:0] node710;
	wire [11-1:0] node711;
	wire [11-1:0] node713;
	wire [11-1:0] node716;
	wire [11-1:0] node717;
	wire [11-1:0] node720;
	wire [11-1:0] node723;
	wire [11-1:0] node724;
	wire [11-1:0] node725;
	wire [11-1:0] node726;
	wire [11-1:0] node727;
	wire [11-1:0] node732;
	wire [11-1:0] node733;
	wire [11-1:0] node735;
	wire [11-1:0] node738;
	wire [11-1:0] node741;
	wire [11-1:0] node742;
	wire [11-1:0] node743;
	wire [11-1:0] node744;
	wire [11-1:0] node747;
	wire [11-1:0] node750;
	wire [11-1:0] node751;
	wire [11-1:0] node755;
	wire [11-1:0] node756;
	wire [11-1:0] node757;
	wire [11-1:0] node760;
	wire [11-1:0] node763;
	wire [11-1:0] node765;
	wire [11-1:0] node768;
	wire [11-1:0] node769;
	wire [11-1:0] node770;
	wire [11-1:0] node771;
	wire [11-1:0] node772;
	wire [11-1:0] node774;
	wire [11-1:0] node777;
	wire [11-1:0] node780;
	wire [11-1:0] node781;
	wire [11-1:0] node782;
	wire [11-1:0] node785;
	wire [11-1:0] node788;
	wire [11-1:0] node791;
	wire [11-1:0] node792;
	wire [11-1:0] node794;
	wire [11-1:0] node796;
	wire [11-1:0] node799;
	wire [11-1:0] node801;
	wire [11-1:0] node802;
	wire [11-1:0] node805;
	wire [11-1:0] node808;
	wire [11-1:0] node809;
	wire [11-1:0] node810;
	wire [11-1:0] node811;
	wire [11-1:0] node814;
	wire [11-1:0] node816;
	wire [11-1:0] node819;
	wire [11-1:0] node820;
	wire [11-1:0] node823;
	wire [11-1:0] node824;
	wire [11-1:0] node828;
	wire [11-1:0] node829;
	wire [11-1:0] node830;
	wire [11-1:0] node831;
	wire [11-1:0] node835;
	wire [11-1:0] node838;
	wire [11-1:0] node839;
	wire [11-1:0] node840;
	wire [11-1:0] node843;
	wire [11-1:0] node846;
	wire [11-1:0] node849;
	wire [11-1:0] node850;
	wire [11-1:0] node851;
	wire [11-1:0] node852;
	wire [11-1:0] node853;
	wire [11-1:0] node854;
	wire [11-1:0] node855;
	wire [11-1:0] node858;
	wire [11-1:0] node861;
	wire [11-1:0] node864;
	wire [11-1:0] node865;
	wire [11-1:0] node866;
	wire [11-1:0] node870;
	wire [11-1:0] node873;
	wire [11-1:0] node874;
	wire [11-1:0] node875;
	wire [11-1:0] node878;
	wire [11-1:0] node880;
	wire [11-1:0] node883;
	wire [11-1:0] node884;
	wire [11-1:0] node885;
	wire [11-1:0] node889;
	wire [11-1:0] node890;
	wire [11-1:0] node893;
	wire [11-1:0] node896;
	wire [11-1:0] node897;
	wire [11-1:0] node898;
	wire [11-1:0] node899;
	wire [11-1:0] node902;
	wire [11-1:0] node905;
	wire [11-1:0] node906;
	wire [11-1:0] node907;
	wire [11-1:0] node911;
	wire [11-1:0] node914;
	wire [11-1:0] node915;
	wire [11-1:0] node916;
	wire [11-1:0] node919;
	wire [11-1:0] node920;
	wire [11-1:0] node923;
	wire [11-1:0] node926;
	wire [11-1:0] node927;
	wire [11-1:0] node930;
	wire [11-1:0] node933;
	wire [11-1:0] node934;
	wire [11-1:0] node935;
	wire [11-1:0] node936;
	wire [11-1:0] node937;
	wire [11-1:0] node939;
	wire [11-1:0] node942;
	wire [11-1:0] node943;
	wire [11-1:0] node946;
	wire [11-1:0] node949;
	wire [11-1:0] node950;
	wire [11-1:0] node952;
	wire [11-1:0] node955;
	wire [11-1:0] node956;
	wire [11-1:0] node959;
	wire [11-1:0] node962;
	wire [11-1:0] node963;
	wire [11-1:0] node965;
	wire [11-1:0] node966;
	wire [11-1:0] node970;
	wire [11-1:0] node972;
	wire [11-1:0] node973;
	wire [11-1:0] node976;
	wire [11-1:0] node979;
	wire [11-1:0] node980;
	wire [11-1:0] node981;
	wire [11-1:0] node982;
	wire [11-1:0] node985;
	wire [11-1:0] node988;
	wire [11-1:0] node989;
	wire [11-1:0] node992;
	wire [11-1:0] node995;
	wire [11-1:0] node996;
	wire [11-1:0] node997;
	wire [11-1:0] node1000;
	wire [11-1:0] node1003;
	wire [11-1:0] node1004;
	wire [11-1:0] node1006;
	wire [11-1:0] node1009;
	wire [11-1:0] node1010;
	wire [11-1:0] node1014;
	wire [11-1:0] node1015;
	wire [11-1:0] node1016;
	wire [11-1:0] node1017;
	wire [11-1:0] node1018;
	wire [11-1:0] node1019;
	wire [11-1:0] node1020;
	wire [11-1:0] node1023;
	wire [11-1:0] node1024;
	wire [11-1:0] node1028;
	wire [11-1:0] node1029;
	wire [11-1:0] node1030;
	wire [11-1:0] node1034;
	wire [11-1:0] node1035;
	wire [11-1:0] node1038;
	wire [11-1:0] node1041;
	wire [11-1:0] node1042;
	wire [11-1:0] node1043;
	wire [11-1:0] node1044;
	wire [11-1:0] node1047;
	wire [11-1:0] node1050;
	wire [11-1:0] node1051;
	wire [11-1:0] node1055;
	wire [11-1:0] node1056;
	wire [11-1:0] node1059;
	wire [11-1:0] node1060;
	wire [11-1:0] node1063;
	wire [11-1:0] node1066;
	wire [11-1:0] node1067;
	wire [11-1:0] node1068;
	wire [11-1:0] node1069;
	wire [11-1:0] node1070;
	wire [11-1:0] node1074;
	wire [11-1:0] node1075;
	wire [11-1:0] node1079;
	wire [11-1:0] node1080;
	wire [11-1:0] node1083;
	wire [11-1:0] node1084;
	wire [11-1:0] node1087;
	wire [11-1:0] node1090;
	wire [11-1:0] node1091;
	wire [11-1:0] node1092;
	wire [11-1:0] node1094;
	wire [11-1:0] node1097;
	wire [11-1:0] node1098;
	wire [11-1:0] node1102;
	wire [11-1:0] node1103;
	wire [11-1:0] node1106;
	wire [11-1:0] node1108;
	wire [11-1:0] node1111;
	wire [11-1:0] node1112;
	wire [11-1:0] node1113;
	wire [11-1:0] node1114;
	wire [11-1:0] node1115;
	wire [11-1:0] node1118;
	wire [11-1:0] node1121;
	wire [11-1:0] node1122;
	wire [11-1:0] node1123;
	wire [11-1:0] node1126;
	wire [11-1:0] node1129;
	wire [11-1:0] node1130;
	wire [11-1:0] node1134;
	wire [11-1:0] node1135;
	wire [11-1:0] node1136;
	wire [11-1:0] node1137;
	wire [11-1:0] node1141;
	wire [11-1:0] node1143;
	wire [11-1:0] node1146;
	wire [11-1:0] node1147;
	wire [11-1:0] node1148;
	wire [11-1:0] node1152;
	wire [11-1:0] node1155;
	wire [11-1:0] node1156;
	wire [11-1:0] node1157;
	wire [11-1:0] node1158;
	wire [11-1:0] node1159;
	wire [11-1:0] node1163;
	wire [11-1:0] node1164;
	wire [11-1:0] node1167;
	wire [11-1:0] node1170;
	wire [11-1:0] node1171;
	wire [11-1:0] node1172;
	wire [11-1:0] node1176;
	wire [11-1:0] node1179;
	wire [11-1:0] node1180;
	wire [11-1:0] node1181;
	wire [11-1:0] node1182;
	wire [11-1:0] node1185;
	wire [11-1:0] node1188;
	wire [11-1:0] node1189;
	wire [11-1:0] node1192;
	wire [11-1:0] node1195;
	wire [11-1:0] node1196;
	wire [11-1:0] node1198;
	wire [11-1:0] node1201;
	wire [11-1:0] node1204;
	wire [11-1:0] node1205;
	wire [11-1:0] node1206;
	wire [11-1:0] node1207;
	wire [11-1:0] node1208;
	wire [11-1:0] node1209;
	wire [11-1:0] node1210;
	wire [11-1:0] node1213;
	wire [11-1:0] node1216;
	wire [11-1:0] node1219;
	wire [11-1:0] node1222;
	wire [11-1:0] node1223;
	wire [11-1:0] node1225;
	wire [11-1:0] node1227;
	wire [11-1:0] node1230;
	wire [11-1:0] node1231;
	wire [11-1:0] node1232;
	wire [11-1:0] node1236;
	wire [11-1:0] node1238;
	wire [11-1:0] node1241;
	wire [11-1:0] node1242;
	wire [11-1:0] node1243;
	wire [11-1:0] node1244;
	wire [11-1:0] node1245;
	wire [11-1:0] node1249;
	wire [11-1:0] node1252;
	wire [11-1:0] node1253;
	wire [11-1:0] node1254;
	wire [11-1:0] node1257;
	wire [11-1:0] node1260;
	wire [11-1:0] node1261;
	wire [11-1:0] node1265;
	wire [11-1:0] node1266;
	wire [11-1:0] node1267;
	wire [11-1:0] node1268;
	wire [11-1:0] node1271;
	wire [11-1:0] node1274;
	wire [11-1:0] node1275;
	wire [11-1:0] node1278;
	wire [11-1:0] node1281;
	wire [11-1:0] node1282;
	wire [11-1:0] node1284;
	wire [11-1:0] node1287;
	wire [11-1:0] node1289;
	wire [11-1:0] node1292;
	wire [11-1:0] node1293;
	wire [11-1:0] node1294;
	wire [11-1:0] node1295;
	wire [11-1:0] node1296;
	wire [11-1:0] node1299;
	wire [11-1:0] node1301;
	wire [11-1:0] node1304;
	wire [11-1:0] node1305;
	wire [11-1:0] node1306;
	wire [11-1:0] node1310;
	wire [11-1:0] node1313;
	wire [11-1:0] node1314;
	wire [11-1:0] node1315;
	wire [11-1:0] node1316;
	wire [11-1:0] node1320;
	wire [11-1:0] node1323;
	wire [11-1:0] node1324;
	wire [11-1:0] node1328;
	wire [11-1:0] node1329;
	wire [11-1:0] node1330;
	wire [11-1:0] node1331;
	wire [11-1:0] node1332;
	wire [11-1:0] node1336;
	wire [11-1:0] node1337;
	wire [11-1:0] node1340;
	wire [11-1:0] node1343;
	wire [11-1:0] node1344;
	wire [11-1:0] node1347;
	wire [11-1:0] node1350;
	wire [11-1:0] node1351;
	wire [11-1:0] node1352;
	wire [11-1:0] node1353;
	wire [11-1:0] node1357;
	wire [11-1:0] node1360;
	wire [11-1:0] node1361;
	wire [11-1:0] node1364;
	wire [11-1:0] node1365;
	wire [11-1:0] node1368;
	wire [11-1:0] node1371;
	wire [11-1:0] node1372;
	wire [11-1:0] node1373;
	wire [11-1:0] node1374;
	wire [11-1:0] node1375;
	wire [11-1:0] node1376;
	wire [11-1:0] node1377;
	wire [11-1:0] node1378;
	wire [11-1:0] node1379;
	wire [11-1:0] node1380;
	wire [11-1:0] node1384;
	wire [11-1:0] node1385;
	wire [11-1:0] node1389;
	wire [11-1:0] node1390;
	wire [11-1:0] node1393;
	wire [11-1:0] node1394;
	wire [11-1:0] node1398;
	wire [11-1:0] node1399;
	wire [11-1:0] node1400;
	wire [11-1:0] node1401;
	wire [11-1:0] node1404;
	wire [11-1:0] node1407;
	wire [11-1:0] node1410;
	wire [11-1:0] node1411;
	wire [11-1:0] node1413;
	wire [11-1:0] node1416;
	wire [11-1:0] node1417;
	wire [11-1:0] node1421;
	wire [11-1:0] node1422;
	wire [11-1:0] node1423;
	wire [11-1:0] node1425;
	wire [11-1:0] node1427;
	wire [11-1:0] node1430;
	wire [11-1:0] node1431;
	wire [11-1:0] node1432;
	wire [11-1:0] node1436;
	wire [11-1:0] node1437;
	wire [11-1:0] node1440;
	wire [11-1:0] node1443;
	wire [11-1:0] node1444;
	wire [11-1:0] node1445;
	wire [11-1:0] node1446;
	wire [11-1:0] node1450;
	wire [11-1:0] node1452;
	wire [11-1:0] node1455;
	wire [11-1:0] node1456;
	wire [11-1:0] node1457;
	wire [11-1:0] node1460;
	wire [11-1:0] node1463;
	wire [11-1:0] node1464;
	wire [11-1:0] node1468;
	wire [11-1:0] node1469;
	wire [11-1:0] node1470;
	wire [11-1:0] node1471;
	wire [11-1:0] node1472;
	wire [11-1:0] node1473;
	wire [11-1:0] node1477;
	wire [11-1:0] node1480;
	wire [11-1:0] node1481;
	wire [11-1:0] node1482;
	wire [11-1:0] node1486;
	wire [11-1:0] node1487;
	wire [11-1:0] node1491;
	wire [11-1:0] node1492;
	wire [11-1:0] node1493;
	wire [11-1:0] node1496;
	wire [11-1:0] node1498;
	wire [11-1:0] node1501;
	wire [11-1:0] node1502;
	wire [11-1:0] node1503;
	wire [11-1:0] node1507;
	wire [11-1:0] node1510;
	wire [11-1:0] node1511;
	wire [11-1:0] node1512;
	wire [11-1:0] node1513;
	wire [11-1:0] node1516;
	wire [11-1:0] node1519;
	wire [11-1:0] node1520;
	wire [11-1:0] node1521;
	wire [11-1:0] node1524;
	wire [11-1:0] node1527;
	wire [11-1:0] node1530;
	wire [11-1:0] node1531;
	wire [11-1:0] node1532;
	wire [11-1:0] node1533;
	wire [11-1:0] node1536;
	wire [11-1:0] node1539;
	wire [11-1:0] node1542;
	wire [11-1:0] node1543;
	wire [11-1:0] node1546;
	wire [11-1:0] node1547;
	wire [11-1:0] node1550;
	wire [11-1:0] node1553;
	wire [11-1:0] node1554;
	wire [11-1:0] node1555;
	wire [11-1:0] node1556;
	wire [11-1:0] node1557;
	wire [11-1:0] node1558;
	wire [11-1:0] node1559;
	wire [11-1:0] node1562;
	wire [11-1:0] node1565;
	wire [11-1:0] node1568;
	wire [11-1:0] node1569;
	wire [11-1:0] node1571;
	wire [11-1:0] node1574;
	wire [11-1:0] node1576;
	wire [11-1:0] node1579;
	wire [11-1:0] node1580;
	wire [11-1:0] node1581;
	wire [11-1:0] node1584;
	wire [11-1:0] node1585;
	wire [11-1:0] node1588;
	wire [11-1:0] node1591;
	wire [11-1:0] node1592;
	wire [11-1:0] node1593;
	wire [11-1:0] node1597;
	wire [11-1:0] node1600;
	wire [11-1:0] node1601;
	wire [11-1:0] node1602;
	wire [11-1:0] node1603;
	wire [11-1:0] node1606;
	wire [11-1:0] node1609;
	wire [11-1:0] node1611;
	wire [11-1:0] node1614;
	wire [11-1:0] node1615;
	wire [11-1:0] node1616;
	wire [11-1:0] node1619;
	wire [11-1:0] node1622;
	wire [11-1:0] node1624;
	wire [11-1:0] node1625;
	wire [11-1:0] node1629;
	wire [11-1:0] node1630;
	wire [11-1:0] node1631;
	wire [11-1:0] node1632;
	wire [11-1:0] node1633;
	wire [11-1:0] node1634;
	wire [11-1:0] node1637;
	wire [11-1:0] node1640;
	wire [11-1:0] node1643;
	wire [11-1:0] node1644;
	wire [11-1:0] node1645;
	wire [11-1:0] node1648;
	wire [11-1:0] node1652;
	wire [11-1:0] node1653;
	wire [11-1:0] node1654;
	wire [11-1:0] node1657;
	wire [11-1:0] node1660;
	wire [11-1:0] node1661;
	wire [11-1:0] node1662;
	wire [11-1:0] node1666;
	wire [11-1:0] node1667;
	wire [11-1:0] node1670;
	wire [11-1:0] node1673;
	wire [11-1:0] node1674;
	wire [11-1:0] node1675;
	wire [11-1:0] node1676;
	wire [11-1:0] node1679;
	wire [11-1:0] node1681;
	wire [11-1:0] node1684;
	wire [11-1:0] node1685;
	wire [11-1:0] node1688;
	wire [11-1:0] node1691;
	wire [11-1:0] node1692;
	wire [11-1:0] node1693;
	wire [11-1:0] node1696;
	wire [11-1:0] node1697;
	wire [11-1:0] node1701;
	wire [11-1:0] node1702;
	wire [11-1:0] node1704;
	wire [11-1:0] node1707;
	wire [11-1:0] node1710;
	wire [11-1:0] node1711;
	wire [11-1:0] node1712;
	wire [11-1:0] node1713;
	wire [11-1:0] node1714;
	wire [11-1:0] node1715;
	wire [11-1:0] node1716;
	wire [11-1:0] node1719;
	wire [11-1:0] node1722;
	wire [11-1:0] node1723;
	wire [11-1:0] node1724;
	wire [11-1:0] node1728;
	wire [11-1:0] node1731;
	wire [11-1:0] node1732;
	wire [11-1:0] node1734;
	wire [11-1:0] node1735;
	wire [11-1:0] node1739;
	wire [11-1:0] node1740;
	wire [11-1:0] node1741;
	wire [11-1:0] node1744;
	wire [11-1:0] node1747;
	wire [11-1:0] node1748;
	wire [11-1:0] node1751;
	wire [11-1:0] node1754;
	wire [11-1:0] node1755;
	wire [11-1:0] node1756;
	wire [11-1:0] node1757;
	wire [11-1:0] node1759;
	wire [11-1:0] node1762;
	wire [11-1:0] node1764;
	wire [11-1:0] node1767;
	wire [11-1:0] node1768;
	wire [11-1:0] node1771;
	wire [11-1:0] node1772;
	wire [11-1:0] node1776;
	wire [11-1:0] node1777;
	wire [11-1:0] node1778;
	wire [11-1:0] node1779;
	wire [11-1:0] node1783;
	wire [11-1:0] node1785;
	wire [11-1:0] node1788;
	wire [11-1:0] node1789;
	wire [11-1:0] node1792;
	wire [11-1:0] node1794;
	wire [11-1:0] node1797;
	wire [11-1:0] node1798;
	wire [11-1:0] node1799;
	wire [11-1:0] node1800;
	wire [11-1:0] node1801;
	wire [11-1:0] node1802;
	wire [11-1:0] node1806;
	wire [11-1:0] node1807;
	wire [11-1:0] node1811;
	wire [11-1:0] node1812;
	wire [11-1:0] node1814;
	wire [11-1:0] node1817;
	wire [11-1:0] node1820;
	wire [11-1:0] node1821;
	wire [11-1:0] node1823;
	wire [11-1:0] node1825;
	wire [11-1:0] node1828;
	wire [11-1:0] node1829;
	wire [11-1:0] node1832;
	wire [11-1:0] node1834;
	wire [11-1:0] node1837;
	wire [11-1:0] node1838;
	wire [11-1:0] node1839;
	wire [11-1:0] node1840;
	wire [11-1:0] node1843;
	wire [11-1:0] node1844;
	wire [11-1:0] node1848;
	wire [11-1:0] node1849;
	wire [11-1:0] node1850;
	wire [11-1:0] node1855;
	wire [11-1:0] node1856;
	wire [11-1:0] node1857;
	wire [11-1:0] node1860;
	wire [11-1:0] node1862;
	wire [11-1:0] node1865;
	wire [11-1:0] node1866;
	wire [11-1:0] node1867;
	wire [11-1:0] node1870;
	wire [11-1:0] node1873;
	wire [11-1:0] node1876;
	wire [11-1:0] node1877;
	wire [11-1:0] node1878;
	wire [11-1:0] node1879;
	wire [11-1:0] node1880;
	wire [11-1:0] node1881;
	wire [11-1:0] node1882;
	wire [11-1:0] node1886;
	wire [11-1:0] node1889;
	wire [11-1:0] node1891;
	wire [11-1:0] node1893;
	wire [11-1:0] node1896;
	wire [11-1:0] node1897;
	wire [11-1:0] node1898;
	wire [11-1:0] node1899;
	wire [11-1:0] node1903;
	wire [11-1:0] node1906;
	wire [11-1:0] node1908;
	wire [11-1:0] node1911;
	wire [11-1:0] node1912;
	wire [11-1:0] node1913;
	wire [11-1:0] node1914;
	wire [11-1:0] node1916;
	wire [11-1:0] node1919;
	wire [11-1:0] node1921;
	wire [11-1:0] node1924;
	wire [11-1:0] node1925;
	wire [11-1:0] node1927;
	wire [11-1:0] node1930;
	wire [11-1:0] node1933;
	wire [11-1:0] node1934;
	wire [11-1:0] node1935;
	wire [11-1:0] node1936;
	wire [11-1:0] node1939;
	wire [11-1:0] node1942;
	wire [11-1:0] node1943;
	wire [11-1:0] node1947;
	wire [11-1:0] node1948;
	wire [11-1:0] node1951;
	wire [11-1:0] node1954;
	wire [11-1:0] node1955;
	wire [11-1:0] node1956;
	wire [11-1:0] node1957;
	wire [11-1:0] node1958;
	wire [11-1:0] node1961;
	wire [11-1:0] node1962;
	wire [11-1:0] node1965;
	wire [11-1:0] node1968;
	wire [11-1:0] node1971;
	wire [11-1:0] node1972;
	wire [11-1:0] node1974;
	wire [11-1:0] node1975;
	wire [11-1:0] node1979;
	wire [11-1:0] node1980;
	wire [11-1:0] node1983;
	wire [11-1:0] node1984;
	wire [11-1:0] node1988;
	wire [11-1:0] node1989;
	wire [11-1:0] node1990;
	wire [11-1:0] node1992;
	wire [11-1:0] node1993;
	wire [11-1:0] node1996;
	wire [11-1:0] node1999;
	wire [11-1:0] node2000;
	wire [11-1:0] node2001;
	wire [11-1:0] node2004;
	wire [11-1:0] node2008;
	wire [11-1:0] node2009;
	wire [11-1:0] node2010;
	wire [11-1:0] node2011;
	wire [11-1:0] node2015;
	wire [11-1:0] node2018;
	wire [11-1:0] node2019;
	wire [11-1:0] node2020;
	wire [11-1:0] node2025;
	wire [11-1:0] node2026;
	wire [11-1:0] node2027;
	wire [11-1:0] node2028;
	wire [11-1:0] node2029;
	wire [11-1:0] node2030;
	wire [11-1:0] node2031;
	wire [11-1:0] node2032;
	wire [11-1:0] node2035;
	wire [11-1:0] node2038;
	wire [11-1:0] node2039;
	wire [11-1:0] node2040;
	wire [11-1:0] node2043;
	wire [11-1:0] node2046;
	wire [11-1:0] node2048;
	wire [11-1:0] node2051;
	wire [11-1:0] node2052;
	wire [11-1:0] node2053;
	wire [11-1:0] node2055;
	wire [11-1:0] node2058;
	wire [11-1:0] node2061;
	wire [11-1:0] node2062;
	wire [11-1:0] node2065;
	wire [11-1:0] node2067;
	wire [11-1:0] node2070;
	wire [11-1:0] node2071;
	wire [11-1:0] node2072;
	wire [11-1:0] node2074;
	wire [11-1:0] node2077;
	wire [11-1:0] node2078;
	wire [11-1:0] node2079;
	wire [11-1:0] node2082;
	wire [11-1:0] node2085;
	wire [11-1:0] node2086;
	wire [11-1:0] node2090;
	wire [11-1:0] node2091;
	wire [11-1:0] node2092;
	wire [11-1:0] node2095;
	wire [11-1:0] node2098;
	wire [11-1:0] node2100;
	wire [11-1:0] node2103;
	wire [11-1:0] node2104;
	wire [11-1:0] node2105;
	wire [11-1:0] node2106;
	wire [11-1:0] node2107;
	wire [11-1:0] node2109;
	wire [11-1:0] node2112;
	wire [11-1:0] node2115;
	wire [11-1:0] node2116;
	wire [11-1:0] node2117;
	wire [11-1:0] node2122;
	wire [11-1:0] node2123;
	wire [11-1:0] node2124;
	wire [11-1:0] node2125;
	wire [11-1:0] node2129;
	wire [11-1:0] node2132;
	wire [11-1:0] node2133;
	wire [11-1:0] node2135;
	wire [11-1:0] node2138;
	wire [11-1:0] node2139;
	wire [11-1:0] node2143;
	wire [11-1:0] node2144;
	wire [11-1:0] node2145;
	wire [11-1:0] node2147;
	wire [11-1:0] node2148;
	wire [11-1:0] node2151;
	wire [11-1:0] node2154;
	wire [11-1:0] node2155;
	wire [11-1:0] node2158;
	wire [11-1:0] node2161;
	wire [11-1:0] node2162;
	wire [11-1:0] node2163;
	wire [11-1:0] node2166;
	wire [11-1:0] node2168;
	wire [11-1:0] node2171;
	wire [11-1:0] node2172;
	wire [11-1:0] node2175;
	wire [11-1:0] node2176;
	wire [11-1:0] node2179;
	wire [11-1:0] node2182;
	wire [11-1:0] node2183;
	wire [11-1:0] node2184;
	wire [11-1:0] node2185;
	wire [11-1:0] node2186;
	wire [11-1:0] node2187;
	wire [11-1:0] node2188;
	wire [11-1:0] node2191;
	wire [11-1:0] node2194;
	wire [11-1:0] node2195;
	wire [11-1:0] node2198;
	wire [11-1:0] node2201;
	wire [11-1:0] node2203;
	wire [11-1:0] node2205;
	wire [11-1:0] node2208;
	wire [11-1:0] node2209;
	wire [11-1:0] node2210;
	wire [11-1:0] node2212;
	wire [11-1:0] node2215;
	wire [11-1:0] node2216;
	wire [11-1:0] node2219;
	wire [11-1:0] node2222;
	wire [11-1:0] node2223;
	wire [11-1:0] node2224;
	wire [11-1:0] node2227;
	wire [11-1:0] node2230;
	wire [11-1:0] node2231;
	wire [11-1:0] node2234;
	wire [11-1:0] node2237;
	wire [11-1:0] node2238;
	wire [11-1:0] node2239;
	wire [11-1:0] node2240;
	wire [11-1:0] node2241;
	wire [11-1:0] node2245;
	wire [11-1:0] node2248;
	wire [11-1:0] node2250;
	wire [11-1:0] node2251;
	wire [11-1:0] node2255;
	wire [11-1:0] node2256;
	wire [11-1:0] node2257;
	wire [11-1:0] node2260;
	wire [11-1:0] node2262;
	wire [11-1:0] node2265;
	wire [11-1:0] node2266;
	wire [11-1:0] node2269;
	wire [11-1:0] node2270;
	wire [11-1:0] node2274;
	wire [11-1:0] node2275;
	wire [11-1:0] node2276;
	wire [11-1:0] node2277;
	wire [11-1:0] node2278;
	wire [11-1:0] node2280;
	wire [11-1:0] node2284;
	wire [11-1:0] node2285;
	wire [11-1:0] node2287;
	wire [11-1:0] node2290;
	wire [11-1:0] node2293;
	wire [11-1:0] node2294;
	wire [11-1:0] node2295;
	wire [11-1:0] node2296;
	wire [11-1:0] node2299;
	wire [11-1:0] node2302;
	wire [11-1:0] node2303;
	wire [11-1:0] node2307;
	wire [11-1:0] node2308;
	wire [11-1:0] node2311;
	wire [11-1:0] node2312;
	wire [11-1:0] node2316;
	wire [11-1:0] node2317;
	wire [11-1:0] node2318;
	wire [11-1:0] node2319;
	wire [11-1:0] node2321;
	wire [11-1:0] node2324;
	wire [11-1:0] node2326;
	wire [11-1:0] node2329;
	wire [11-1:0] node2330;
	wire [11-1:0] node2331;
	wire [11-1:0] node2334;
	wire [11-1:0] node2337;
	wire [11-1:0] node2338;
	wire [11-1:0] node2342;
	wire [11-1:0] node2343;
	wire [11-1:0] node2344;
	wire [11-1:0] node2345;
	wire [11-1:0] node2348;
	wire [11-1:0] node2351;
	wire [11-1:0] node2354;
	wire [11-1:0] node2355;
	wire [11-1:0] node2356;
	wire [11-1:0] node2361;
	wire [11-1:0] node2362;
	wire [11-1:0] node2363;
	wire [11-1:0] node2364;
	wire [11-1:0] node2365;
	wire [11-1:0] node2366;
	wire [11-1:0] node2367;
	wire [11-1:0] node2368;
	wire [11-1:0] node2372;
	wire [11-1:0] node2375;
	wire [11-1:0] node2376;
	wire [11-1:0] node2378;
	wire [11-1:0] node2381;
	wire [11-1:0] node2384;
	wire [11-1:0] node2385;
	wire [11-1:0] node2386;
	wire [11-1:0] node2387;
	wire [11-1:0] node2390;
	wire [11-1:0] node2393;
	wire [11-1:0] node2394;
	wire [11-1:0] node2397;
	wire [11-1:0] node2400;
	wire [11-1:0] node2401;
	wire [11-1:0] node2402;
	wire [11-1:0] node2405;
	wire [11-1:0] node2408;
	wire [11-1:0] node2411;
	wire [11-1:0] node2412;
	wire [11-1:0] node2413;
	wire [11-1:0] node2414;
	wire [11-1:0] node2415;
	wire [11-1:0] node2419;
	wire [11-1:0] node2422;
	wire [11-1:0] node2423;
	wire [11-1:0] node2425;
	wire [11-1:0] node2428;
	wire [11-1:0] node2431;
	wire [11-1:0] node2432;
	wire [11-1:0] node2433;
	wire [11-1:0] node2437;
	wire [11-1:0] node2438;
	wire [11-1:0] node2439;
	wire [11-1:0] node2443;
	wire [11-1:0] node2444;
	wire [11-1:0] node2448;
	wire [11-1:0] node2449;
	wire [11-1:0] node2450;
	wire [11-1:0] node2451;
	wire [11-1:0] node2452;
	wire [11-1:0] node2455;
	wire [11-1:0] node2456;
	wire [11-1:0] node2460;
	wire [11-1:0] node2463;
	wire [11-1:0] node2464;
	wire [11-1:0] node2465;
	wire [11-1:0] node2468;
	wire [11-1:0] node2470;
	wire [11-1:0] node2473;
	wire [11-1:0] node2474;
	wire [11-1:0] node2476;
	wire [11-1:0] node2479;
	wire [11-1:0] node2482;
	wire [11-1:0] node2483;
	wire [11-1:0] node2484;
	wire [11-1:0] node2485;
	wire [11-1:0] node2487;
	wire [11-1:0] node2490;
	wire [11-1:0] node2491;
	wire [11-1:0] node2495;
	wire [11-1:0] node2496;
	wire [11-1:0] node2499;
	wire [11-1:0] node2502;
	wire [11-1:0] node2503;
	wire [11-1:0] node2506;
	wire [11-1:0] node2508;
	wire [11-1:0] node2510;
	wire [11-1:0] node2513;
	wire [11-1:0] node2514;
	wire [11-1:0] node2515;
	wire [11-1:0] node2516;
	wire [11-1:0] node2517;
	wire [11-1:0] node2518;
	wire [11-1:0] node2521;
	wire [11-1:0] node2522;
	wire [11-1:0] node2526;
	wire [11-1:0] node2527;
	wire [11-1:0] node2528;
	wire [11-1:0] node2533;
	wire [11-1:0] node2534;
	wire [11-1:0] node2535;
	wire [11-1:0] node2538;
	wire [11-1:0] node2541;
	wire [11-1:0] node2542;
	wire [11-1:0] node2543;
	wire [11-1:0] node2547;
	wire [11-1:0] node2548;
	wire [11-1:0] node2552;
	wire [11-1:0] node2553;
	wire [11-1:0] node2554;
	wire [11-1:0] node2555;
	wire [11-1:0] node2556;
	wire [11-1:0] node2559;
	wire [11-1:0] node2562;
	wire [11-1:0] node2565;
	wire [11-1:0] node2566;
	wire [11-1:0] node2567;
	wire [11-1:0] node2571;
	wire [11-1:0] node2574;
	wire [11-1:0] node2575;
	wire [11-1:0] node2576;
	wire [11-1:0] node2577;
	wire [11-1:0] node2582;
	wire [11-1:0] node2583;
	wire [11-1:0] node2586;
	wire [11-1:0] node2587;
	wire [11-1:0] node2591;
	wire [11-1:0] node2592;
	wire [11-1:0] node2593;
	wire [11-1:0] node2594;
	wire [11-1:0] node2595;
	wire [11-1:0] node2597;
	wire [11-1:0] node2600;
	wire [11-1:0] node2602;
	wire [11-1:0] node2605;
	wire [11-1:0] node2606;
	wire [11-1:0] node2607;
	wire [11-1:0] node2611;
	wire [11-1:0] node2614;
	wire [11-1:0] node2615;
	wire [11-1:0] node2616;
	wire [11-1:0] node2620;
	wire [11-1:0] node2621;
	wire [11-1:0] node2623;
	wire [11-1:0] node2626;
	wire [11-1:0] node2627;
	wire [11-1:0] node2631;
	wire [11-1:0] node2632;
	wire [11-1:0] node2633;
	wire [11-1:0] node2635;
	wire [11-1:0] node2636;
	wire [11-1:0] node2639;
	wire [11-1:0] node2642;
	wire [11-1:0] node2643;
	wire [11-1:0] node2645;
	wire [11-1:0] node2648;
	wire [11-1:0] node2650;
	wire [11-1:0] node2653;
	wire [11-1:0] node2654;
	wire [11-1:0] node2655;
	wire [11-1:0] node2656;
	wire [11-1:0] node2659;
	wire [11-1:0] node2662;
	wire [11-1:0] node2663;
	wire [11-1:0] node2666;
	wire [11-1:0] node2669;
	wire [11-1:0] node2670;
	wire [11-1:0] node2671;
	wire [11-1:0] node2676;
	wire [11-1:0] node2677;
	wire [11-1:0] node2678;
	wire [11-1:0] node2679;
	wire [11-1:0] node2680;
	wire [11-1:0] node2681;
	wire [11-1:0] node2682;
	wire [11-1:0] node2683;
	wire [11-1:0] node2684;
	wire [11-1:0] node2685;
	wire [11-1:0] node2686;
	wire [11-1:0] node2690;
	wire [11-1:0] node2691;
	wire [11-1:0] node2694;
	wire [11-1:0] node2697;
	wire [11-1:0] node2698;
	wire [11-1:0] node2701;
	wire [11-1:0] node2703;
	wire [11-1:0] node2706;
	wire [11-1:0] node2707;
	wire [11-1:0] node2708;
	wire [11-1:0] node2711;
	wire [11-1:0] node2714;
	wire [11-1:0] node2715;
	wire [11-1:0] node2716;
	wire [11-1:0] node2721;
	wire [11-1:0] node2722;
	wire [11-1:0] node2723;
	wire [11-1:0] node2724;
	wire [11-1:0] node2727;
	wire [11-1:0] node2728;
	wire [11-1:0] node2732;
	wire [11-1:0] node2733;
	wire [11-1:0] node2734;
	wire [11-1:0] node2737;
	wire [11-1:0] node2740;
	wire [11-1:0] node2741;
	wire [11-1:0] node2745;
	wire [11-1:0] node2746;
	wire [11-1:0] node2747;
	wire [11-1:0] node2748;
	wire [11-1:0] node2752;
	wire [11-1:0] node2754;
	wire [11-1:0] node2757;
	wire [11-1:0] node2758;
	wire [11-1:0] node2761;
	wire [11-1:0] node2762;
	wire [11-1:0] node2766;
	wire [11-1:0] node2767;
	wire [11-1:0] node2768;
	wire [11-1:0] node2769;
	wire [11-1:0] node2770;
	wire [11-1:0] node2773;
	wire [11-1:0] node2776;
	wire [11-1:0] node2777;
	wire [11-1:0] node2779;
	wire [11-1:0] node2782;
	wire [11-1:0] node2785;
	wire [11-1:0] node2786;
	wire [11-1:0] node2787;
	wire [11-1:0] node2790;
	wire [11-1:0] node2791;
	wire [11-1:0] node2794;
	wire [11-1:0] node2797;
	wire [11-1:0] node2798;
	wire [11-1:0] node2800;
	wire [11-1:0] node2803;
	wire [11-1:0] node2805;
	wire [11-1:0] node2808;
	wire [11-1:0] node2809;
	wire [11-1:0] node2810;
	wire [11-1:0] node2811;
	wire [11-1:0] node2814;
	wire [11-1:0] node2817;
	wire [11-1:0] node2818;
	wire [11-1:0] node2819;
	wire [11-1:0] node2823;
	wire [11-1:0] node2824;
	wire [11-1:0] node2828;
	wire [11-1:0] node2829;
	wire [11-1:0] node2831;
	wire [11-1:0] node2833;
	wire [11-1:0] node2836;
	wire [11-1:0] node2837;
	wire [11-1:0] node2840;
	wire [11-1:0] node2842;
	wire [11-1:0] node2845;
	wire [11-1:0] node2846;
	wire [11-1:0] node2847;
	wire [11-1:0] node2848;
	wire [11-1:0] node2849;
	wire [11-1:0] node2851;
	wire [11-1:0] node2852;
	wire [11-1:0] node2855;
	wire [11-1:0] node2858;
	wire [11-1:0] node2859;
	wire [11-1:0] node2860;
	wire [11-1:0] node2865;
	wire [11-1:0] node2866;
	wire [11-1:0] node2867;
	wire [11-1:0] node2869;
	wire [11-1:0] node2872;
	wire [11-1:0] node2875;
	wire [11-1:0] node2877;
	wire [11-1:0] node2880;
	wire [11-1:0] node2881;
	wire [11-1:0] node2882;
	wire [11-1:0] node2883;
	wire [11-1:0] node2886;
	wire [11-1:0] node2888;
	wire [11-1:0] node2891;
	wire [11-1:0] node2892;
	wire [11-1:0] node2893;
	wire [11-1:0] node2896;
	wire [11-1:0] node2899;
	wire [11-1:0] node2902;
	wire [11-1:0] node2903;
	wire [11-1:0] node2904;
	wire [11-1:0] node2906;
	wire [11-1:0] node2909;
	wire [11-1:0] node2912;
	wire [11-1:0] node2914;
	wire [11-1:0] node2917;
	wire [11-1:0] node2918;
	wire [11-1:0] node2919;
	wire [11-1:0] node2920;
	wire [11-1:0] node2922;
	wire [11-1:0] node2923;
	wire [11-1:0] node2926;
	wire [11-1:0] node2929;
	wire [11-1:0] node2930;
	wire [11-1:0] node2933;
	wire [11-1:0] node2936;
	wire [11-1:0] node2937;
	wire [11-1:0] node2938;
	wire [11-1:0] node2939;
	wire [11-1:0] node2943;
	wire [11-1:0] node2945;
	wire [11-1:0] node2948;
	wire [11-1:0] node2949;
	wire [11-1:0] node2951;
	wire [11-1:0] node2954;
	wire [11-1:0] node2956;
	wire [11-1:0] node2959;
	wire [11-1:0] node2960;
	wire [11-1:0] node2961;
	wire [11-1:0] node2962;
	wire [11-1:0] node2965;
	wire [11-1:0] node2967;
	wire [11-1:0] node2970;
	wire [11-1:0] node2971;
	wire [11-1:0] node2975;
	wire [11-1:0] node2976;
	wire [11-1:0] node2977;
	wire [11-1:0] node2980;
	wire [11-1:0] node2983;
	wire [11-1:0] node2984;
	wire [11-1:0] node2986;
	wire [11-1:0] node2989;
	wire [11-1:0] node2992;
	wire [11-1:0] node2993;
	wire [11-1:0] node2994;
	wire [11-1:0] node2995;
	wire [11-1:0] node2996;
	wire [11-1:0] node2997;
	wire [11-1:0] node2998;
	wire [11-1:0] node3002;
	wire [11-1:0] node3003;
	wire [11-1:0] node3006;
	wire [11-1:0] node3007;
	wire [11-1:0] node3010;
	wire [11-1:0] node3013;
	wire [11-1:0] node3014;
	wire [11-1:0] node3015;
	wire [11-1:0] node3016;
	wire [11-1:0] node3019;
	wire [11-1:0] node3022;
	wire [11-1:0] node3025;
	wire [11-1:0] node3026;
	wire [11-1:0] node3027;
	wire [11-1:0] node3030;
	wire [11-1:0] node3033;
	wire [11-1:0] node3036;
	wire [11-1:0] node3037;
	wire [11-1:0] node3038;
	wire [11-1:0] node3039;
	wire [11-1:0] node3042;
	wire [11-1:0] node3043;
	wire [11-1:0] node3046;
	wire [11-1:0] node3049;
	wire [11-1:0] node3050;
	wire [11-1:0] node3051;
	wire [11-1:0] node3054;
	wire [11-1:0] node3057;
	wire [11-1:0] node3060;
	wire [11-1:0] node3061;
	wire [11-1:0] node3062;
	wire [11-1:0] node3065;
	wire [11-1:0] node3066;
	wire [11-1:0] node3069;
	wire [11-1:0] node3072;
	wire [11-1:0] node3073;
	wire [11-1:0] node3075;
	wire [11-1:0] node3078;
	wire [11-1:0] node3080;
	wire [11-1:0] node3083;
	wire [11-1:0] node3084;
	wire [11-1:0] node3085;
	wire [11-1:0] node3086;
	wire [11-1:0] node3087;
	wire [11-1:0] node3088;
	wire [11-1:0] node3092;
	wire [11-1:0] node3093;
	wire [11-1:0] node3096;
	wire [11-1:0] node3099;
	wire [11-1:0] node3100;
	wire [11-1:0] node3103;
	wire [11-1:0] node3105;
	wire [11-1:0] node3108;
	wire [11-1:0] node3109;
	wire [11-1:0] node3110;
	wire [11-1:0] node3111;
	wire [11-1:0] node3115;
	wire [11-1:0] node3118;
	wire [11-1:0] node3119;
	wire [11-1:0] node3122;
	wire [11-1:0] node3123;
	wire [11-1:0] node3126;
	wire [11-1:0] node3129;
	wire [11-1:0] node3130;
	wire [11-1:0] node3131;
	wire [11-1:0] node3132;
	wire [11-1:0] node3133;
	wire [11-1:0] node3137;
	wire [11-1:0] node3139;
	wire [11-1:0] node3142;
	wire [11-1:0] node3143;
	wire [11-1:0] node3145;
	wire [11-1:0] node3148;
	wire [11-1:0] node3149;
	wire [11-1:0] node3152;
	wire [11-1:0] node3155;
	wire [11-1:0] node3156;
	wire [11-1:0] node3158;
	wire [11-1:0] node3161;
	wire [11-1:0] node3162;
	wire [11-1:0] node3164;
	wire [11-1:0] node3167;
	wire [11-1:0] node3168;
	wire [11-1:0] node3171;
	wire [11-1:0] node3174;
	wire [11-1:0] node3175;
	wire [11-1:0] node3176;
	wire [11-1:0] node3177;
	wire [11-1:0] node3178;
	wire [11-1:0] node3179;
	wire [11-1:0] node3180;
	wire [11-1:0] node3183;
	wire [11-1:0] node3186;
	wire [11-1:0] node3188;
	wire [11-1:0] node3191;
	wire [11-1:0] node3192;
	wire [11-1:0] node3193;
	wire [11-1:0] node3197;
	wire [11-1:0] node3198;
	wire [11-1:0] node3202;
	wire [11-1:0] node3203;
	wire [11-1:0] node3204;
	wire [11-1:0] node3207;
	wire [11-1:0] node3210;
	wire [11-1:0] node3211;
	wire [11-1:0] node3212;
	wire [11-1:0] node3216;
	wire [11-1:0] node3218;
	wire [11-1:0] node3221;
	wire [11-1:0] node3222;
	wire [11-1:0] node3223;
	wire [11-1:0] node3224;
	wire [11-1:0] node3226;
	wire [11-1:0] node3230;
	wire [11-1:0] node3232;
	wire [11-1:0] node3233;
	wire [11-1:0] node3236;
	wire [11-1:0] node3239;
	wire [11-1:0] node3240;
	wire [11-1:0] node3241;
	wire [11-1:0] node3242;
	wire [11-1:0] node3246;
	wire [11-1:0] node3249;
	wire [11-1:0] node3250;
	wire [11-1:0] node3251;
	wire [11-1:0] node3255;
	wire [11-1:0] node3256;
	wire [11-1:0] node3260;
	wire [11-1:0] node3261;
	wire [11-1:0] node3262;
	wire [11-1:0] node3263;
	wire [11-1:0] node3264;
	wire [11-1:0] node3265;
	wire [11-1:0] node3269;
	wire [11-1:0] node3270;
	wire [11-1:0] node3274;
	wire [11-1:0] node3275;
	wire [11-1:0] node3276;
	wire [11-1:0] node3279;
	wire [11-1:0] node3282;
	wire [11-1:0] node3285;
	wire [11-1:0] node3286;
	wire [11-1:0] node3287;
	wire [11-1:0] node3289;
	wire [11-1:0] node3293;
	wire [11-1:0] node3294;
	wire [11-1:0] node3296;
	wire [11-1:0] node3299;
	wire [11-1:0] node3300;
	wire [11-1:0] node3304;
	wire [11-1:0] node3305;
	wire [11-1:0] node3306;
	wire [11-1:0] node3307;
	wire [11-1:0] node3308;
	wire [11-1:0] node3311;
	wire [11-1:0] node3314;
	wire [11-1:0] node3316;
	wire [11-1:0] node3319;
	wire [11-1:0] node3320;
	wire [11-1:0] node3323;
	wire [11-1:0] node3325;
	wire [11-1:0] node3328;
	wire [11-1:0] node3329;
	wire [11-1:0] node3330;
	wire [11-1:0] node3332;
	wire [11-1:0] node3335;
	wire [11-1:0] node3338;
	wire [11-1:0] node3339;
	wire [11-1:0] node3341;
	wire [11-1:0] node3344;
	wire [11-1:0] node3347;
	wire [11-1:0] node3348;
	wire [11-1:0] node3349;
	wire [11-1:0] node3350;
	wire [11-1:0] node3351;
	wire [11-1:0] node3352;
	wire [11-1:0] node3353;
	wire [11-1:0] node3354;
	wire [11-1:0] node3355;
	wire [11-1:0] node3359;
	wire [11-1:0] node3360;
	wire [11-1:0] node3364;
	wire [11-1:0] node3365;
	wire [11-1:0] node3366;
	wire [11-1:0] node3369;
	wire [11-1:0] node3373;
	wire [11-1:0] node3374;
	wire [11-1:0] node3375;
	wire [11-1:0] node3378;
	wire [11-1:0] node3381;
	wire [11-1:0] node3382;
	wire [11-1:0] node3385;
	wire [11-1:0] node3386;
	wire [11-1:0] node3389;
	wire [11-1:0] node3392;
	wire [11-1:0] node3393;
	wire [11-1:0] node3394;
	wire [11-1:0] node3395;
	wire [11-1:0] node3397;
	wire [11-1:0] node3401;
	wire [11-1:0] node3402;
	wire [11-1:0] node3406;
	wire [11-1:0] node3407;
	wire [11-1:0] node3408;
	wire [11-1:0] node3409;
	wire [11-1:0] node3413;
	wire [11-1:0] node3414;
	wire [11-1:0] node3417;
	wire [11-1:0] node3420;
	wire [11-1:0] node3421;
	wire [11-1:0] node3422;
	wire [11-1:0] node3425;
	wire [11-1:0] node3428;
	wire [11-1:0] node3430;
	wire [11-1:0] node3433;
	wire [11-1:0] node3434;
	wire [11-1:0] node3435;
	wire [11-1:0] node3436;
	wire [11-1:0] node3438;
	wire [11-1:0] node3441;
	wire [11-1:0] node3442;
	wire [11-1:0] node3445;
	wire [11-1:0] node3446;
	wire [11-1:0] node3450;
	wire [11-1:0] node3451;
	wire [11-1:0] node3452;
	wire [11-1:0] node3453;
	wire [11-1:0] node3456;
	wire [11-1:0] node3460;
	wire [11-1:0] node3461;
	wire [11-1:0] node3464;
	wire [11-1:0] node3466;
	wire [11-1:0] node3469;
	wire [11-1:0] node3470;
	wire [11-1:0] node3471;
	wire [11-1:0] node3473;
	wire [11-1:0] node3474;
	wire [11-1:0] node3477;
	wire [11-1:0] node3480;
	wire [11-1:0] node3481;
	wire [11-1:0] node3482;
	wire [11-1:0] node3486;
	wire [11-1:0] node3487;
	wire [11-1:0] node3490;
	wire [11-1:0] node3493;
	wire [11-1:0] node3494;
	wire [11-1:0] node3495;
	wire [11-1:0] node3496;
	wire [11-1:0] node3500;
	wire [11-1:0] node3503;
	wire [11-1:0] node3504;
	wire [11-1:0] node3506;
	wire [11-1:0] node3509;
	wire [11-1:0] node3510;
	wire [11-1:0] node3513;
	wire [11-1:0] node3516;
	wire [11-1:0] node3517;
	wire [11-1:0] node3518;
	wire [11-1:0] node3519;
	wire [11-1:0] node3520;
	wire [11-1:0] node3521;
	wire [11-1:0] node3523;
	wire [11-1:0] node3526;
	wire [11-1:0] node3529;
	wire [11-1:0] node3530;
	wire [11-1:0] node3532;
	wire [11-1:0] node3535;
	wire [11-1:0] node3536;
	wire [11-1:0] node3540;
	wire [11-1:0] node3541;
	wire [11-1:0] node3542;
	wire [11-1:0] node3544;
	wire [11-1:0] node3547;
	wire [11-1:0] node3548;
	wire [11-1:0] node3551;
	wire [11-1:0] node3554;
	wire [11-1:0] node3555;
	wire [11-1:0] node3558;
	wire [11-1:0] node3561;
	wire [11-1:0] node3562;
	wire [11-1:0] node3563;
	wire [11-1:0] node3564;
	wire [11-1:0] node3565;
	wire [11-1:0] node3568;
	wire [11-1:0] node3572;
	wire [11-1:0] node3573;
	wire [11-1:0] node3575;
	wire [11-1:0] node3578;
	wire [11-1:0] node3581;
	wire [11-1:0] node3582;
	wire [11-1:0] node3583;
	wire [11-1:0] node3584;
	wire [11-1:0] node3587;
	wire [11-1:0] node3590;
	wire [11-1:0] node3593;
	wire [11-1:0] node3594;
	wire [11-1:0] node3597;
	wire [11-1:0] node3600;
	wire [11-1:0] node3601;
	wire [11-1:0] node3602;
	wire [11-1:0] node3603;
	wire [11-1:0] node3604;
	wire [11-1:0] node3605;
	wire [11-1:0] node3609;
	wire [11-1:0] node3610;
	wire [11-1:0] node3614;
	wire [11-1:0] node3615;
	wire [11-1:0] node3618;
	wire [11-1:0] node3621;
	wire [11-1:0] node3622;
	wire [11-1:0] node3623;
	wire [11-1:0] node3624;
	wire [11-1:0] node3627;
	wire [11-1:0] node3630;
	wire [11-1:0] node3631;
	wire [11-1:0] node3635;
	wire [11-1:0] node3636;
	wire [11-1:0] node3637;
	wire [11-1:0] node3641;
	wire [11-1:0] node3642;
	wire [11-1:0] node3645;
	wire [11-1:0] node3648;
	wire [11-1:0] node3649;
	wire [11-1:0] node3650;
	wire [11-1:0] node3651;
	wire [11-1:0] node3654;
	wire [11-1:0] node3655;
	wire [11-1:0] node3658;
	wire [11-1:0] node3661;
	wire [11-1:0] node3662;
	wire [11-1:0] node3663;
	wire [11-1:0] node3666;
	wire [11-1:0] node3669;
	wire [11-1:0] node3670;
	wire [11-1:0] node3673;
	wire [11-1:0] node3676;
	wire [11-1:0] node3677;
	wire [11-1:0] node3678;
	wire [11-1:0] node3679;
	wire [11-1:0] node3682;
	wire [11-1:0] node3685;
	wire [11-1:0] node3686;
	wire [11-1:0] node3690;
	wire [11-1:0] node3691;
	wire [11-1:0] node3693;
	wire [11-1:0] node3696;
	wire [11-1:0] node3699;
	wire [11-1:0] node3700;
	wire [11-1:0] node3701;
	wire [11-1:0] node3702;
	wire [11-1:0] node3703;
	wire [11-1:0] node3704;
	wire [11-1:0] node3705;
	wire [11-1:0] node3707;
	wire [11-1:0] node3710;
	wire [11-1:0] node3713;
	wire [11-1:0] node3714;
	wire [11-1:0] node3717;
	wire [11-1:0] node3718;
	wire [11-1:0] node3721;
	wire [11-1:0] node3724;
	wire [11-1:0] node3725;
	wire [11-1:0] node3727;
	wire [11-1:0] node3730;
	wire [11-1:0] node3731;
	wire [11-1:0] node3734;
	wire [11-1:0] node3737;
	wire [11-1:0] node3738;
	wire [11-1:0] node3739;
	wire [11-1:0] node3740;
	wire [11-1:0] node3741;
	wire [11-1:0] node3745;
	wire [11-1:0] node3748;
	wire [11-1:0] node3749;
	wire [11-1:0] node3753;
	wire [11-1:0] node3754;
	wire [11-1:0] node3755;
	wire [11-1:0] node3757;
	wire [11-1:0] node3760;
	wire [11-1:0] node3763;
	wire [11-1:0] node3766;
	wire [11-1:0] node3767;
	wire [11-1:0] node3768;
	wire [11-1:0] node3769;
	wire [11-1:0] node3770;
	wire [11-1:0] node3771;
	wire [11-1:0] node3775;
	wire [11-1:0] node3778;
	wire [11-1:0] node3779;
	wire [11-1:0] node3780;
	wire [11-1:0] node3783;
	wire [11-1:0] node3786;
	wire [11-1:0] node3789;
	wire [11-1:0] node3790;
	wire [11-1:0] node3791;
	wire [11-1:0] node3792;
	wire [11-1:0] node3795;
	wire [11-1:0] node3798;
	wire [11-1:0] node3799;
	wire [11-1:0] node3802;
	wire [11-1:0] node3805;
	wire [11-1:0] node3806;
	wire [11-1:0] node3808;
	wire [11-1:0] node3811;
	wire [11-1:0] node3813;
	wire [11-1:0] node3816;
	wire [11-1:0] node3817;
	wire [11-1:0] node3818;
	wire [11-1:0] node3819;
	wire [11-1:0] node3821;
	wire [11-1:0] node3824;
	wire [11-1:0] node3825;
	wire [11-1:0] node3829;
	wire [11-1:0] node3830;
	wire [11-1:0] node3832;
	wire [11-1:0] node3835;
	wire [11-1:0] node3838;
	wire [11-1:0] node3839;
	wire [11-1:0] node3840;
	wire [11-1:0] node3843;
	wire [11-1:0] node3845;
	wire [11-1:0] node3848;
	wire [11-1:0] node3849;
	wire [11-1:0] node3852;
	wire [11-1:0] node3853;
	wire [11-1:0] node3857;
	wire [11-1:0] node3858;
	wire [11-1:0] node3859;
	wire [11-1:0] node3860;
	wire [11-1:0] node3861;
	wire [11-1:0] node3863;
	wire [11-1:0] node3866;
	wire [11-1:0] node3868;
	wire [11-1:0] node3871;
	wire [11-1:0] node3872;
	wire [11-1:0] node3874;
	wire [11-1:0] node3877;
	wire [11-1:0] node3879;
	wire [11-1:0] node3880;
	wire [11-1:0] node3884;
	wire [11-1:0] node3885;
	wire [11-1:0] node3886;
	wire [11-1:0] node3887;
	wire [11-1:0] node3888;
	wire [11-1:0] node3891;
	wire [11-1:0] node3894;
	wire [11-1:0] node3897;
	wire [11-1:0] node3898;
	wire [11-1:0] node3899;
	wire [11-1:0] node3903;
	wire [11-1:0] node3904;
	wire [11-1:0] node3908;
	wire [11-1:0] node3909;
	wire [11-1:0] node3910;
	wire [11-1:0] node3911;
	wire [11-1:0] node3914;
	wire [11-1:0] node3917;
	wire [11-1:0] node3918;
	wire [11-1:0] node3922;
	wire [11-1:0] node3924;
	wire [11-1:0] node3927;
	wire [11-1:0] node3928;
	wire [11-1:0] node3929;
	wire [11-1:0] node3930;
	wire [11-1:0] node3931;
	wire [11-1:0] node3932;
	wire [11-1:0] node3936;
	wire [11-1:0] node3937;
	wire [11-1:0] node3941;
	wire [11-1:0] node3942;
	wire [11-1:0] node3945;
	wire [11-1:0] node3947;
	wire [11-1:0] node3950;
	wire [11-1:0] node3951;
	wire [11-1:0] node3953;
	wire [11-1:0] node3955;
	wire [11-1:0] node3958;
	wire [11-1:0] node3959;
	wire [11-1:0] node3961;
	wire [11-1:0] node3964;
	wire [11-1:0] node3965;
	wire [11-1:0] node3969;
	wire [11-1:0] node3970;
	wire [11-1:0] node3971;
	wire [11-1:0] node3972;
	wire [11-1:0] node3974;
	wire [11-1:0] node3977;
	wire [11-1:0] node3979;
	wire [11-1:0] node3982;
	wire [11-1:0] node3983;
	wire [11-1:0] node3986;
	wire [11-1:0] node3987;
	wire [11-1:0] node3991;
	wire [11-1:0] node3992;
	wire [11-1:0] node3993;
	wire [11-1:0] node3995;
	wire [11-1:0] node3998;
	wire [11-1:0] node3999;
	wire [11-1:0] node4003;
	wire [11-1:0] node4004;
	wire [11-1:0] node4005;
	wire [11-1:0] node4009;
	wire [11-1:0] node4012;
	wire [11-1:0] node4013;
	wire [11-1:0] node4014;
	wire [11-1:0] node4015;
	wire [11-1:0] node4016;
	wire [11-1:0] node4017;
	wire [11-1:0] node4018;
	wire [11-1:0] node4019;
	wire [11-1:0] node4020;
	wire [11-1:0] node4023;
	wire [11-1:0] node4026;
	wire [11-1:0] node4027;
	wire [11-1:0] node4028;
	wire [11-1:0] node4032;
	wire [11-1:0] node4033;
	wire [11-1:0] node4036;
	wire [11-1:0] node4039;
	wire [11-1:0] node4040;
	wire [11-1:0] node4041;
	wire [11-1:0] node4044;
	wire [11-1:0] node4046;
	wire [11-1:0] node4049;
	wire [11-1:0] node4051;
	wire [11-1:0] node4053;
	wire [11-1:0] node4056;
	wire [11-1:0] node4057;
	wire [11-1:0] node4058;
	wire [11-1:0] node4059;
	wire [11-1:0] node4063;
	wire [11-1:0] node4065;
	wire [11-1:0] node4068;
	wire [11-1:0] node4069;
	wire [11-1:0] node4070;
	wire [11-1:0] node4073;
	wire [11-1:0] node4076;
	wire [11-1:0] node4077;
	wire [11-1:0] node4080;
	wire [11-1:0] node4083;
	wire [11-1:0] node4084;
	wire [11-1:0] node4085;
	wire [11-1:0] node4086;
	wire [11-1:0] node4087;
	wire [11-1:0] node4090;
	wire [11-1:0] node4091;
	wire [11-1:0] node4094;
	wire [11-1:0] node4097;
	wire [11-1:0] node4098;
	wire [11-1:0] node4101;
	wire [11-1:0] node4104;
	wire [11-1:0] node4105;
	wire [11-1:0] node4106;
	wire [11-1:0] node4107;
	wire [11-1:0] node4111;
	wire [11-1:0] node4112;
	wire [11-1:0] node4116;
	wire [11-1:0] node4117;
	wire [11-1:0] node4118;
	wire [11-1:0] node4123;
	wire [11-1:0] node4124;
	wire [11-1:0] node4125;
	wire [11-1:0] node4126;
	wire [11-1:0] node4129;
	wire [11-1:0] node4130;
	wire [11-1:0] node4133;
	wire [11-1:0] node4136;
	wire [11-1:0] node4137;
	wire [11-1:0] node4140;
	wire [11-1:0] node4143;
	wire [11-1:0] node4144;
	wire [11-1:0] node4145;
	wire [11-1:0] node4148;
	wire [11-1:0] node4151;
	wire [11-1:0] node4152;
	wire [11-1:0] node4155;
	wire [11-1:0] node4158;
	wire [11-1:0] node4159;
	wire [11-1:0] node4160;
	wire [11-1:0] node4161;
	wire [11-1:0] node4162;
	wire [11-1:0] node4163;
	wire [11-1:0] node4164;
	wire [11-1:0] node4167;
	wire [11-1:0] node4171;
	wire [11-1:0] node4172;
	wire [11-1:0] node4174;
	wire [11-1:0] node4177;
	wire [11-1:0] node4178;
	wire [11-1:0] node4182;
	wire [11-1:0] node4183;
	wire [11-1:0] node4184;
	wire [11-1:0] node4185;
	wire [11-1:0] node4189;
	wire [11-1:0] node4192;
	wire [11-1:0] node4193;
	wire [11-1:0] node4195;
	wire [11-1:0] node4198;
	wire [11-1:0] node4199;
	wire [11-1:0] node4202;
	wire [11-1:0] node4205;
	wire [11-1:0] node4206;
	wire [11-1:0] node4207;
	wire [11-1:0] node4208;
	wire [11-1:0] node4211;
	wire [11-1:0] node4214;
	wire [11-1:0] node4215;
	wire [11-1:0] node4216;
	wire [11-1:0] node4219;
	wire [11-1:0] node4222;
	wire [11-1:0] node4223;
	wire [11-1:0] node4226;
	wire [11-1:0] node4229;
	wire [11-1:0] node4230;
	wire [11-1:0] node4231;
	wire [11-1:0] node4233;
	wire [11-1:0] node4237;
	wire [11-1:0] node4238;
	wire [11-1:0] node4241;
	wire [11-1:0] node4244;
	wire [11-1:0] node4245;
	wire [11-1:0] node4246;
	wire [11-1:0] node4247;
	wire [11-1:0] node4248;
	wire [11-1:0] node4249;
	wire [11-1:0] node4252;
	wire [11-1:0] node4255;
	wire [11-1:0] node4257;
	wire [11-1:0] node4260;
	wire [11-1:0] node4261;
	wire [11-1:0] node4263;
	wire [11-1:0] node4266;
	wire [11-1:0] node4267;
	wire [11-1:0] node4271;
	wire [11-1:0] node4272;
	wire [11-1:0] node4273;
	wire [11-1:0] node4276;
	wire [11-1:0] node4277;
	wire [11-1:0] node4280;
	wire [11-1:0] node4283;
	wire [11-1:0] node4284;
	wire [11-1:0] node4285;
	wire [11-1:0] node4289;
	wire [11-1:0] node4292;
	wire [11-1:0] node4293;
	wire [11-1:0] node4294;
	wire [11-1:0] node4295;
	wire [11-1:0] node4296;
	wire [11-1:0] node4300;
	wire [11-1:0] node4303;
	wire [11-1:0] node4304;
	wire [11-1:0] node4307;
	wire [11-1:0] node4310;
	wire [11-1:0] node4311;
	wire [11-1:0] node4313;
	wire [11-1:0] node4314;
	wire [11-1:0] node4318;
	wire [11-1:0] node4319;
	wire [11-1:0] node4321;
	wire [11-1:0] node4324;
	wire [11-1:0] node4325;
	wire [11-1:0] node4329;
	wire [11-1:0] node4330;
	wire [11-1:0] node4331;
	wire [11-1:0] node4332;
	wire [11-1:0] node4333;
	wire [11-1:0] node4334;
	wire [11-1:0] node4335;
	wire [11-1:0] node4336;
	wire [11-1:0] node4340;
	wire [11-1:0] node4342;
	wire [11-1:0] node4345;
	wire [11-1:0] node4346;
	wire [11-1:0] node4347;
	wire [11-1:0] node4352;
	wire [11-1:0] node4353;
	wire [11-1:0] node4354;
	wire [11-1:0] node4357;
	wire [11-1:0] node4360;
	wire [11-1:0] node4361;
	wire [11-1:0] node4362;
	wire [11-1:0] node4365;
	wire [11-1:0] node4368;
	wire [11-1:0] node4371;
	wire [11-1:0] node4372;
	wire [11-1:0] node4373;
	wire [11-1:0] node4374;
	wire [11-1:0] node4375;
	wire [11-1:0] node4378;
	wire [11-1:0] node4381;
	wire [11-1:0] node4384;
	wire [11-1:0] node4385;
	wire [11-1:0] node4386;
	wire [11-1:0] node4389;
	wire [11-1:0] node4392;
	wire [11-1:0] node4393;
	wire [11-1:0] node4396;
	wire [11-1:0] node4399;
	wire [11-1:0] node4400;
	wire [11-1:0] node4401;
	wire [11-1:0] node4404;
	wire [11-1:0] node4405;
	wire [11-1:0] node4409;
	wire [11-1:0] node4410;
	wire [11-1:0] node4411;
	wire [11-1:0] node4414;
	wire [11-1:0] node4417;
	wire [11-1:0] node4420;
	wire [11-1:0] node4421;
	wire [11-1:0] node4422;
	wire [11-1:0] node4423;
	wire [11-1:0] node4425;
	wire [11-1:0] node4427;
	wire [11-1:0] node4430;
	wire [11-1:0] node4431;
	wire [11-1:0] node4434;
	wire [11-1:0] node4437;
	wire [11-1:0] node4438;
	wire [11-1:0] node4439;
	wire [11-1:0] node4442;
	wire [11-1:0] node4443;
	wire [11-1:0] node4446;
	wire [11-1:0] node4449;
	wire [11-1:0] node4450;
	wire [11-1:0] node4451;
	wire [11-1:0] node4455;
	wire [11-1:0] node4456;
	wire [11-1:0] node4459;
	wire [11-1:0] node4462;
	wire [11-1:0] node4463;
	wire [11-1:0] node4464;
	wire [11-1:0] node4465;
	wire [11-1:0] node4469;
	wire [11-1:0] node4470;
	wire [11-1:0] node4472;
	wire [11-1:0] node4475;
	wire [11-1:0] node4476;
	wire [11-1:0] node4480;
	wire [11-1:0] node4481;
	wire [11-1:0] node4482;
	wire [11-1:0] node4485;
	wire [11-1:0] node4487;
	wire [11-1:0] node4490;
	wire [11-1:0] node4491;
	wire [11-1:0] node4494;
	wire [11-1:0] node4497;
	wire [11-1:0] node4498;
	wire [11-1:0] node4499;
	wire [11-1:0] node4500;
	wire [11-1:0] node4501;
	wire [11-1:0] node4502;
	wire [11-1:0] node4503;
	wire [11-1:0] node4506;
	wire [11-1:0] node4509;
	wire [11-1:0] node4510;
	wire [11-1:0] node4514;
	wire [11-1:0] node4515;
	wire [11-1:0] node4516;
	wire [11-1:0] node4520;
	wire [11-1:0] node4523;
	wire [11-1:0] node4524;
	wire [11-1:0] node4525;
	wire [11-1:0] node4526;
	wire [11-1:0] node4530;
	wire [11-1:0] node4531;
	wire [11-1:0] node4534;
	wire [11-1:0] node4537;
	wire [11-1:0] node4538;
	wire [11-1:0] node4539;
	wire [11-1:0] node4544;
	wire [11-1:0] node4545;
	wire [11-1:0] node4546;
	wire [11-1:0] node4547;
	wire [11-1:0] node4548;
	wire [11-1:0] node4551;
	wire [11-1:0] node4554;
	wire [11-1:0] node4555;
	wire [11-1:0] node4558;
	wire [11-1:0] node4561;
	wire [11-1:0] node4562;
	wire [11-1:0] node4565;
	wire [11-1:0] node4567;
	wire [11-1:0] node4570;
	wire [11-1:0] node4571;
	wire [11-1:0] node4572;
	wire [11-1:0] node4573;
	wire [11-1:0] node4577;
	wire [11-1:0] node4580;
	wire [11-1:0] node4581;
	wire [11-1:0] node4582;
	wire [11-1:0] node4586;
	wire [11-1:0] node4589;
	wire [11-1:0] node4590;
	wire [11-1:0] node4591;
	wire [11-1:0] node4592;
	wire [11-1:0] node4594;
	wire [11-1:0] node4596;
	wire [11-1:0] node4599;
	wire [11-1:0] node4600;
	wire [11-1:0] node4601;
	wire [11-1:0] node4604;
	wire [11-1:0] node4607;
	wire [11-1:0] node4610;
	wire [11-1:0] node4611;
	wire [11-1:0] node4612;
	wire [11-1:0] node4613;
	wire [11-1:0] node4616;
	wire [11-1:0] node4619;
	wire [11-1:0] node4620;
	wire [11-1:0] node4624;
	wire [11-1:0] node4625;
	wire [11-1:0] node4628;
	wire [11-1:0] node4631;
	wire [11-1:0] node4632;
	wire [11-1:0] node4633;
	wire [11-1:0] node4635;
	wire [11-1:0] node4637;
	wire [11-1:0] node4640;
	wire [11-1:0] node4641;
	wire [11-1:0] node4644;
	wire [11-1:0] node4645;
	wire [11-1:0] node4649;
	wire [11-1:0] node4650;
	wire [11-1:0] node4651;
	wire [11-1:0] node4652;
	wire [11-1:0] node4655;
	wire [11-1:0] node4658;
	wire [11-1:0] node4659;
	wire [11-1:0] node4662;
	wire [11-1:0] node4665;
	wire [11-1:0] node4666;
	wire [11-1:0] node4670;
	wire [11-1:0] node4671;
	wire [11-1:0] node4672;
	wire [11-1:0] node4673;
	wire [11-1:0] node4674;
	wire [11-1:0] node4675;
	wire [11-1:0] node4676;
	wire [11-1:0] node4677;
	wire [11-1:0] node4679;
	wire [11-1:0] node4682;
	wire [11-1:0] node4685;
	wire [11-1:0] node4686;
	wire [11-1:0] node4687;
	wire [11-1:0] node4690;
	wire [11-1:0] node4694;
	wire [11-1:0] node4695;
	wire [11-1:0] node4696;
	wire [11-1:0] node4697;
	wire [11-1:0] node4701;
	wire [11-1:0] node4704;
	wire [11-1:0] node4705;
	wire [11-1:0] node4708;
	wire [11-1:0] node4709;
	wire [11-1:0] node4713;
	wire [11-1:0] node4714;
	wire [11-1:0] node4715;
	wire [11-1:0] node4716;
	wire [11-1:0] node4720;
	wire [11-1:0] node4721;
	wire [11-1:0] node4724;
	wire [11-1:0] node4725;
	wire [11-1:0] node4728;
	wire [11-1:0] node4731;
	wire [11-1:0] node4732;
	wire [11-1:0] node4734;
	wire [11-1:0] node4737;
	wire [11-1:0] node4738;
	wire [11-1:0] node4741;
	wire [11-1:0] node4742;
	wire [11-1:0] node4746;
	wire [11-1:0] node4747;
	wire [11-1:0] node4748;
	wire [11-1:0] node4749;
	wire [11-1:0] node4750;
	wire [11-1:0] node4751;
	wire [11-1:0] node4754;
	wire [11-1:0] node4757;
	wire [11-1:0] node4758;
	wire [11-1:0] node4762;
	wire [11-1:0] node4763;
	wire [11-1:0] node4765;
	wire [11-1:0] node4768;
	wire [11-1:0] node4771;
	wire [11-1:0] node4772;
	wire [11-1:0] node4773;
	wire [11-1:0] node4776;
	wire [11-1:0] node4777;
	wire [11-1:0] node4781;
	wire [11-1:0] node4782;
	wire [11-1:0] node4784;
	wire [11-1:0] node4787;
	wire [11-1:0] node4789;
	wire [11-1:0] node4792;
	wire [11-1:0] node4793;
	wire [11-1:0] node4794;
	wire [11-1:0] node4796;
	wire [11-1:0] node4797;
	wire [11-1:0] node4801;
	wire [11-1:0] node4802;
	wire [11-1:0] node4804;
	wire [11-1:0] node4808;
	wire [11-1:0] node4809;
	wire [11-1:0] node4810;
	wire [11-1:0] node4811;
	wire [11-1:0] node4814;
	wire [11-1:0] node4817;
	wire [11-1:0] node4819;
	wire [11-1:0] node4822;
	wire [11-1:0] node4823;
	wire [11-1:0] node4824;
	wire [11-1:0] node4828;
	wire [11-1:0] node4829;
	wire [11-1:0] node4833;
	wire [11-1:0] node4834;
	wire [11-1:0] node4835;
	wire [11-1:0] node4836;
	wire [11-1:0] node4837;
	wire [11-1:0] node4838;
	wire [11-1:0] node4839;
	wire [11-1:0] node4842;
	wire [11-1:0] node4845;
	wire [11-1:0] node4848;
	wire [11-1:0] node4849;
	wire [11-1:0] node4850;
	wire [11-1:0] node4854;
	wire [11-1:0] node4855;
	wire [11-1:0] node4859;
	wire [11-1:0] node4860;
	wire [11-1:0] node4861;
	wire [11-1:0] node4864;
	wire [11-1:0] node4866;
	wire [11-1:0] node4869;
	wire [11-1:0] node4870;
	wire [11-1:0] node4871;
	wire [11-1:0] node4874;
	wire [11-1:0] node4877;
	wire [11-1:0] node4880;
	wire [11-1:0] node4881;
	wire [11-1:0] node4882;
	wire [11-1:0] node4883;
	wire [11-1:0] node4886;
	wire [11-1:0] node4889;
	wire [11-1:0] node4890;
	wire [11-1:0] node4892;
	wire [11-1:0] node4895;
	wire [11-1:0] node4896;
	wire [11-1:0] node4900;
	wire [11-1:0] node4901;
	wire [11-1:0] node4902;
	wire [11-1:0] node4904;
	wire [11-1:0] node4907;
	wire [11-1:0] node4910;
	wire [11-1:0] node4911;
	wire [11-1:0] node4914;
	wire [11-1:0] node4917;
	wire [11-1:0] node4918;
	wire [11-1:0] node4919;
	wire [11-1:0] node4920;
	wire [11-1:0] node4921;
	wire [11-1:0] node4924;
	wire [11-1:0] node4925;
	wire [11-1:0] node4929;
	wire [11-1:0] node4932;
	wire [11-1:0] node4933;
	wire [11-1:0] node4935;
	wire [11-1:0] node4937;
	wire [11-1:0] node4940;
	wire [11-1:0] node4941;
	wire [11-1:0] node4944;
	wire [11-1:0] node4946;
	wire [11-1:0] node4949;
	wire [11-1:0] node4950;
	wire [11-1:0] node4951;
	wire [11-1:0] node4952;
	wire [11-1:0] node4955;
	wire [11-1:0] node4956;
	wire [11-1:0] node4960;
	wire [11-1:0] node4961;
	wire [11-1:0] node4964;
	wire [11-1:0] node4967;
	wire [11-1:0] node4968;
	wire [11-1:0] node4969;
	wire [11-1:0] node4970;
	wire [11-1:0] node4973;
	wire [11-1:0] node4977;
	wire [11-1:0] node4978;
	wire [11-1:0] node4982;
	wire [11-1:0] node4983;
	wire [11-1:0] node4984;
	wire [11-1:0] node4985;
	wire [11-1:0] node4986;
	wire [11-1:0] node4987;
	wire [11-1:0] node4988;
	wire [11-1:0] node4990;
	wire [11-1:0] node4994;
	wire [11-1:0] node4995;
	wire [11-1:0] node4996;
	wire [11-1:0] node4999;
	wire [11-1:0] node5002;
	wire [11-1:0] node5004;
	wire [11-1:0] node5007;
	wire [11-1:0] node5008;
	wire [11-1:0] node5010;
	wire [11-1:0] node5011;
	wire [11-1:0] node5015;
	wire [11-1:0] node5016;
	wire [11-1:0] node5019;
	wire [11-1:0] node5021;
	wire [11-1:0] node5024;
	wire [11-1:0] node5025;
	wire [11-1:0] node5026;
	wire [11-1:0] node5027;
	wire [11-1:0] node5030;
	wire [11-1:0] node5033;
	wire [11-1:0] node5034;
	wire [11-1:0] node5037;
	wire [11-1:0] node5040;
	wire [11-1:0] node5041;
	wire [11-1:0] node5043;
	wire [11-1:0] node5044;
	wire [11-1:0] node5048;
	wire [11-1:0] node5049;
	wire [11-1:0] node5050;
	wire [11-1:0] node5054;
	wire [11-1:0] node5055;
	wire [11-1:0] node5059;
	wire [11-1:0] node5060;
	wire [11-1:0] node5061;
	wire [11-1:0] node5062;
	wire [11-1:0] node5063;
	wire [11-1:0] node5064;
	wire [11-1:0] node5068;
	wire [11-1:0] node5070;
	wire [11-1:0] node5073;
	wire [11-1:0] node5074;
	wire [11-1:0] node5077;
	wire [11-1:0] node5080;
	wire [11-1:0] node5081;
	wire [11-1:0] node5082;
	wire [11-1:0] node5084;
	wire [11-1:0] node5087;
	wire [11-1:0] node5088;
	wire [11-1:0] node5091;
	wire [11-1:0] node5094;
	wire [11-1:0] node5095;
	wire [11-1:0] node5097;
	wire [11-1:0] node5101;
	wire [11-1:0] node5102;
	wire [11-1:0] node5103;
	wire [11-1:0] node5105;
	wire [11-1:0] node5106;
	wire [11-1:0] node5109;
	wire [11-1:0] node5112;
	wire [11-1:0] node5113;
	wire [11-1:0] node5115;
	wire [11-1:0] node5118;
	wire [11-1:0] node5121;
	wire [11-1:0] node5122;
	wire [11-1:0] node5123;
	wire [11-1:0] node5124;
	wire [11-1:0] node5127;
	wire [11-1:0] node5130;
	wire [11-1:0] node5132;
	wire [11-1:0] node5135;
	wire [11-1:0] node5136;
	wire [11-1:0] node5139;
	wire [11-1:0] node5142;
	wire [11-1:0] node5143;
	wire [11-1:0] node5144;
	wire [11-1:0] node5145;
	wire [11-1:0] node5146;
	wire [11-1:0] node5147;
	wire [11-1:0] node5150;
	wire [11-1:0] node5152;
	wire [11-1:0] node5155;
	wire [11-1:0] node5157;
	wire [11-1:0] node5159;
	wire [11-1:0] node5162;
	wire [11-1:0] node5163;
	wire [11-1:0] node5164;
	wire [11-1:0] node5167;
	wire [11-1:0] node5169;
	wire [11-1:0] node5172;
	wire [11-1:0] node5174;
	wire [11-1:0] node5177;
	wire [11-1:0] node5178;
	wire [11-1:0] node5179;
	wire [11-1:0] node5180;
	wire [11-1:0] node5181;
	wire [11-1:0] node5185;
	wire [11-1:0] node5187;
	wire [11-1:0] node5190;
	wire [11-1:0] node5191;
	wire [11-1:0] node5195;
	wire [11-1:0] node5196;
	wire [11-1:0] node5198;
	wire [11-1:0] node5199;
	wire [11-1:0] node5203;
	wire [11-1:0] node5204;
	wire [11-1:0] node5207;
	wire [11-1:0] node5210;
	wire [11-1:0] node5211;
	wire [11-1:0] node5212;
	wire [11-1:0] node5213;
	wire [11-1:0] node5214;
	wire [11-1:0] node5215;
	wire [11-1:0] node5219;
	wire [11-1:0] node5220;
	wire [11-1:0] node5223;
	wire [11-1:0] node5226;
	wire [11-1:0] node5227;
	wire [11-1:0] node5230;
	wire [11-1:0] node5231;
	wire [11-1:0] node5235;
	wire [11-1:0] node5236;
	wire [11-1:0] node5237;
	wire [11-1:0] node5238;
	wire [11-1:0] node5241;
	wire [11-1:0] node5244;
	wire [11-1:0] node5247;
	wire [11-1:0] node5249;
	wire [11-1:0] node5250;
	wire [11-1:0] node5254;
	wire [11-1:0] node5255;
	wire [11-1:0] node5256;
	wire [11-1:0] node5257;
	wire [11-1:0] node5260;
	wire [11-1:0] node5263;
	wire [11-1:0] node5265;
	wire [11-1:0] node5268;
	wire [11-1:0] node5269;
	wire [11-1:0] node5270;
	wire [11-1:0] node5271;
	wire [11-1:0] node5274;
	wire [11-1:0] node5277;
	wire [11-1:0] node5280;
	wire [11-1:0] node5282;

	assign outp = (inp[1]) ? node2676 : node1;
		assign node1 = (inp[7]) ? node1371 : node2;
			assign node2 = (inp[2]) ? node676 : node3;
				assign node3 = (inp[0]) ? node323 : node4;
					assign node4 = (inp[4]) ? node180 : node5;
						assign node5 = (inp[10]) ? node93 : node6;
							assign node6 = (inp[3]) ? node50 : node7;
								assign node7 = (inp[9]) ? node25 : node8;
									assign node8 = (inp[5]) ? node14 : node9;
										assign node9 = (inp[11]) ? 11'b01010000010 : node10;
											assign node10 = (inp[8]) ? 11'b01000101010 : 11'b01001100010;
										assign node14 = (inp[11]) ? node22 : node15;
											assign node15 = (inp[8]) ? node19 : node16;
												assign node16 = (inp[6]) ? 11'b01001011011 : 11'b01001111010;
												assign node19 = (inp[6]) ? 11'b01000111011 : 11'b01000011011;
											assign node22 = (inp[8]) ? 11'b01001011010 : 11'b01000011000;
									assign node25 = (inp[11]) ? node37 : node26;
										assign node26 = (inp[5]) ? node34 : node27;
											assign node27 = (inp[6]) ? node31 : node28;
												assign node28 = (inp[8]) ? 11'b01010101011 : 11'b01001101011;
												assign node31 = (inp[8]) ? 11'b01010001000 : 11'b01000100000;
											assign node34 = (inp[6]) ? 11'b01001111011 : 11'b01010111010;
										assign node37 = (inp[5]) ? node45 : node38;
											assign node38 = (inp[6]) ? node42 : node39;
												assign node39 = (inp[8]) ? 11'b01110111001 : 11'b01101111011;
												assign node42 = (inp[8]) ? 11'b01101011010 : 11'b01111111001;
											assign node45 = (inp[6]) ? node47 : 11'b01001101010;
												assign node47 = (inp[8]) ? 11'b01010101001 : 11'b01111001011;
								assign node50 = (inp[9]) ? node74 : node51;
									assign node51 = (inp[11]) ? node63 : node52;
										assign node52 = (inp[8]) ? node60 : node53;
											assign node53 = (inp[6]) ? node57 : node54;
												assign node54 = (inp[5]) ? 11'b11001111010 : 11'b11001101011;
												assign node57 = (inp[5]) ? 11'b11011011011 : 11'b11011100010;
											assign node60 = (inp[6]) ? 11'b11000111001 : 11'b11000011011;
										assign node63 = (inp[5]) ? node69 : node64;
											assign node64 = (inp[8]) ? node66 : 11'b11000010010;
												assign node66 = (inp[6]) ? 11'b11101111000 : 11'b11100011001;
											assign node69 = (inp[6]) ? node71 : 11'b11010001010;
												assign node71 = (inp[8]) ? 11'b11001101011 : 11'b11100001001;
									assign node74 = (inp[5]) ? node82 : node75;
										assign node75 = (inp[6]) ? 11'b11111001110 : node76;
											assign node76 = (inp[8]) ? 11'b11100101101 : node77;
												assign node77 = (inp[11]) ? 11'b11101101111 : 11'b11001101111;
										assign node82 = (inp[6]) ? node88 : node83;
											assign node83 = (inp[8]) ? node85 : 11'b11011111100;
												assign node85 = (inp[11]) ? 11'b11100111110 : 11'b11000111100;
											assign node88 = (inp[11]) ? 11'b11010011111 : node89;
												assign node89 = (inp[8]) ? 11'b11010111111 : 11'b11001111111;
							assign node93 = (inp[3]) ? node139 : node94;
								assign node94 = (inp[9]) ? node116 : node95;
									assign node95 = (inp[5]) ? node109 : node96;
										assign node96 = (inp[11]) ? node102 : node97;
											assign node97 = (inp[8]) ? node99 : 11'b11000100010;
												assign node99 = (inp[6]) ? 11'b11011001010 : 11'b11001101011;
											assign node102 = (inp[8]) ? node106 : node103;
												assign node103 = (inp[6]) ? 11'b11011101011 : 11'b11000101011;
												assign node106 = (inp[6]) ? 11'b11110101000 : 11'b11111101001;
										assign node109 = (inp[6]) ? node113 : node110;
											assign node110 = (inp[11]) ? 11'b11010011010 : 11'b11100111010;
											assign node113 = (inp[11]) ? 11'b11110011001 : 11'b11110111001;
									assign node116 = (inp[5]) ? node126 : node117;
										assign node117 = (inp[8]) ? node121 : node118;
											assign node118 = (inp[6]) ? 11'b11110111101 : 11'b11100111111;
											assign node121 = (inp[6]) ? node123 : 11'b11001111101;
												assign node123 = (inp[11]) ? 11'b11011011100 : 11'b11001011110;
										assign node126 = (inp[6]) ? node134 : node127;
											assign node127 = (inp[11]) ? node131 : node128;
												assign node128 = (inp[8]) ? 11'b11000101100 : 11'b11100101110;
												assign node131 = (inp[8]) ? 11'b11110101110 : 11'b11111101100;
											assign node134 = (inp[11]) ? 11'b11100001101 : node135;
												assign node135 = (inp[8]) ? 11'b11010101111 : 11'b11111101111;
								assign node139 = (inp[8]) ? node161 : node140;
									assign node140 = (inp[6]) ? node152 : node141;
										assign node141 = (inp[5]) ? node149 : node142;
											assign node142 = (inp[9]) ? node146 : node143;
												assign node143 = (inp[11]) ? 11'b01000111111 : 11'b01000101111;
												assign node146 = (inp[11]) ? 11'b01010111111 : 11'b01000111111;
											assign node149 = (inp[9]) ? 11'b01000101100 : 11'b01100111110;
										assign node152 = (inp[11]) ? node156 : node153;
											assign node153 = (inp[5]) ? 11'b01110011101 : 11'b01010100110;
											assign node156 = (inp[9]) ? 11'b01010001101 : node157;
												assign node157 = (inp[5]) ? 11'b01001001111 : 11'b01001111101;
									assign node161 = (inp[5]) ? node175 : node162;
										assign node162 = (inp[6]) ? node170 : node163;
											assign node163 = (inp[11]) ? node167 : node164;
												assign node164 = (inp[9]) ? 11'b01110111111 : 11'b01100101111;
												assign node167 = (inp[9]) ? 11'b01101111101 : 11'b01011111101;
											assign node170 = (inp[9]) ? node172 : 11'b01010111110;
												assign node172 = (inp[11]) ? 11'b01100011100 : 11'b01111011110;
										assign node175 = (inp[6]) ? node177 : 11'b01111111110;
											assign node177 = (inp[9]) ? 11'b01111101111 : 11'b01011101101;
						assign node180 = (inp[3]) ? node258 : node181;
							assign node181 = (inp[10]) ? node223 : node182;
								assign node182 = (inp[11]) ? node202 : node183;
									assign node183 = (inp[5]) ? node193 : node184;
										assign node184 = (inp[6]) ? node190 : node185;
											assign node185 = (inp[8]) ? node187 : 11'b01101001111;
												assign node187 = (inp[9]) ? 11'b01110001111 : 11'b01100101111;
											assign node190 = (inp[9]) ? 11'b01111101100 : 11'b01100001110;
										assign node193 = (inp[6]) ? node199 : node194;
											assign node194 = (inp[8]) ? node196 : 11'b01111011110;
												assign node196 = (inp[9]) ? 11'b01101011100 : 11'b01111111100;
											assign node199 = (inp[9]) ? 11'b01100111111 : 11'b01010111111;
									assign node202 = (inp[5]) ? node214 : node203;
										assign node203 = (inp[8]) ? node211 : node204;
											assign node204 = (inp[9]) ? node208 : node205;
												assign node205 = (inp[6]) ? 11'b01011101111 : 11'b01011001111;
												assign node208 = (inp[6]) ? 11'b01001011101 : 11'b01011011111;
											assign node211 = (inp[6]) ? 11'b01010011100 : 11'b01110101101;
										assign node214 = (inp[8]) ? 11'b01101001111 : node215;
											assign node215 = (inp[9]) ? node219 : node216;
												assign node216 = (inp[6]) ? 11'b01001111100 : 11'b01000111100;
												assign node219 = (inp[6]) ? 11'b01011101110 : 11'b01010001100;
								assign node223 = (inp[5]) ? node245 : node224;
									assign node224 = (inp[11]) ? node234 : node225;
										assign node225 = (inp[9]) ? node231 : node226;
											assign node226 = (inp[8]) ? 11'b11110011100 : node227;
												assign node227 = (inp[6]) ? 11'b11001010110 : 11'b11000011111;
											assign node231 = (inp[6]) ? 11'b11000101010 : 11'b11001001001;
										assign node234 = (inp[8]) ? node240 : node235;
											assign node235 = (inp[9]) ? 11'b11100011011 : node236;
												assign node236 = (inp[6]) ? 11'b11110111111 : 11'b11110011111;
											assign node240 = (inp[6]) ? 11'b11111111001 : node241;
												assign node241 = (inp[9]) ? 11'b11111011011 : 11'b11111011101;
									assign node245 = (inp[9]) ? node255 : node246;
										assign node246 = (inp[11]) ? node250 : node247;
											assign node247 = (inp[6]) ? 11'b11000001111 : 11'b11010001110;
											assign node250 = (inp[8]) ? 11'b11110101100 : node251;
												assign node251 = (inp[6]) ? 11'b11010101110 : 11'b11001001100;
										assign node255 = (inp[6]) ? 11'b11001101000 : 11'b11011001000;
							assign node258 = (inp[10]) ? node290 : node259;
								assign node259 = (inp[9]) ? node275 : node260;
									assign node260 = (inp[5]) ? node268 : node261;
										assign node261 = (inp[8]) ? node263 : 11'b11111001111;
											assign node263 = (inp[11]) ? 11'b11010101101 : node264;
												assign node264 = (inp[6]) ? 11'b11000001100 : 11'b11001001111;
										assign node268 = (inp[11]) ? node270 : 11'b11111011110;
											assign node270 = (inp[6]) ? 11'b11100111101 : node271;
												assign node271 = (inp[8]) ? 11'b11101111100 : 11'b11101011100;
									assign node275 = (inp[5]) ? node281 : node276;
										assign node276 = (inp[6]) ? node278 : 11'b11011011011;
											assign node278 = (inp[8]) ? 11'b11000011000 : 11'b11011011001;
										assign node281 = (inp[6]) ? node287 : node282;
											assign node282 = (inp[11]) ? node284 : 11'b11110001000;
												assign node284 = (inp[8]) ? 11'b11101001000 : 11'b11111001000;
											assign node287 = (inp[8]) ? 11'b11101001001 : 11'b11101101000;
								assign node290 = (inp[5]) ? node310 : node291;
									assign node291 = (inp[9]) ? node299 : node292;
										assign node292 = (inp[6]) ? node296 : node293;
											assign node293 = (inp[8]) ? 11'b01010001011 : 11'b01100001011;
											assign node296 = (inp[8]) ? 11'b01001101000 : 11'b01110000010;
										assign node299 = (inp[11]) ? node307 : node300;
											assign node300 = (inp[6]) ? node304 : node301;
												assign node301 = (inp[8]) ? 11'b01101011001 : 11'b01100011011;
												assign node304 = (inp[8]) ? 11'b01111111010 : 11'b01111010000;
											assign node307 = (inp[8]) ? 11'b01111011011 : 11'b01110011011;
									assign node310 = (inp[6]) ? node318 : node311;
										assign node311 = (inp[9]) ? node313 : 11'b01001011000;
											assign node313 = (inp[11]) ? 11'b01110001000 : node314;
												assign node314 = (inp[8]) ? 11'b01101001010 : 11'b01100001000;
										assign node318 = (inp[8]) ? node320 : 11'b01111001011;
											assign node320 = (inp[9]) ? 11'b01110001001 : 11'b01111001011;
					assign node323 = (inp[3]) ? node501 : node324;
						assign node324 = (inp[4]) ? node414 : node325;
							assign node325 = (inp[11]) ? node371 : node326;
								assign node326 = (inp[6]) ? node348 : node327;
									assign node327 = (inp[5]) ? node341 : node328;
										assign node328 = (inp[8]) ? node334 : node329;
											assign node329 = (inp[10]) ? 11'b01000101101 : node330;
												assign node330 = (inp[9]) ? 11'b01001101101 : 11'b01001101001;
											assign node334 = (inp[9]) ? node338 : node335;
												assign node335 = (inp[10]) ? 11'b01101101101 : 11'b01100001000;
												assign node338 = (inp[10]) ? 11'b01111111001 : 11'b01110101101;
										assign node341 = (inp[10]) ? node345 : node342;
											assign node342 = (inp[8]) ? 11'b01110101100 : 11'b01001101100;
											assign node345 = (inp[9]) ? 11'b01100111000 : 11'b01100101100;
									assign node348 = (inp[5]) ? node362 : node349;
										assign node349 = (inp[8]) ? node355 : node350;
											assign node350 = (inp[9]) ? 11'b01010110010 : node351;
												assign node351 = (inp[10]) ? 11'b01010100100 : 11'b01011100000;
											assign node355 = (inp[10]) ? node359 : node356;
												assign node356 = (inp[9]) ? 11'b01100001110 : 11'b01110101000;
												assign node359 = (inp[9]) ? 11'b01101011000 : 11'b01111001100;
										assign node362 = (inp[9]) ? node366 : node363;
											assign node363 = (inp[8]) ? 11'b01001101111 : 11'b01110001111;
											assign node366 = (inp[10]) ? node368 : 11'b01101101101;
												assign node368 = (inp[8]) ? 11'b01010111001 : 11'b01111111001;
								assign node371 = (inp[9]) ? node391 : node372;
									assign node372 = (inp[8]) ? node382 : node373;
										assign node373 = (inp[10]) ? node377 : node374;
											assign node374 = (inp[5]) ? 11'b01001111010 : 11'b01001111001;
											assign node377 = (inp[5]) ? 11'b01000011101 : node378;
												assign node378 = (inp[6]) ? 11'b01011111101 : 11'b01000111101;
										assign node382 = (inp[5]) ? node388 : node383;
											assign node383 = (inp[6]) ? node385 : 11'b01111111111;
												assign node385 = (inp[10]) ? 11'b01100111100 : 11'b01111111010;
											assign node388 = (inp[10]) ? 11'b01110011100 : 11'b01110011001;
									assign node391 = (inp[10]) ? node401 : node392;
										assign node392 = (inp[6]) ? node398 : node393;
											assign node393 = (inp[8]) ? node395 : 11'b01101111101;
												assign node395 = (inp[5]) ? 11'b01001111100 : 11'b01000111111;
											assign node398 = (inp[8]) ? 11'b01010111111 : 11'b01110111111;
										assign node401 = (inp[6]) ? node409 : node402;
											assign node402 = (inp[5]) ? node406 : node403;
												assign node403 = (inp[8]) ? 11'b01101101011 : 11'b01010101001;
												assign node406 = (inp[8]) ? 11'b01010101000 : 11'b01110101010;
											assign node409 = (inp[8]) ? 11'b01110001010 : node410;
												assign node410 = (inp[5]) ? 11'b01100001011 : 11'b01000101001;
							assign node414 = (inp[11]) ? node458 : node415;
								assign node415 = (inp[6]) ? node435 : node416;
									assign node416 = (inp[5]) ? node428 : node417;
										assign node417 = (inp[9]) ? node421 : node418;
											assign node418 = (inp[8]) ? 11'b01100101001 : 11'b01000011101;
											assign node421 = (inp[8]) ? node425 : node422;
												assign node422 = (inp[10]) ? 11'b01100011001 : 11'b01101011101;
												assign node425 = (inp[10]) ? 11'b01001011011 : 11'b01010011101;
										assign node428 = (inp[8]) ? 11'b01010011110 : node429;
											assign node429 = (inp[10]) ? node431 : 11'b01111011100;
												assign node431 = (inp[9]) ? 11'b01100011010 : 11'b01010011100;
									assign node435 = (inp[5]) ? node449 : node436;
										assign node436 = (inp[8]) ? node444 : node437;
											assign node437 = (inp[9]) ? node441 : node438;
												assign node438 = (inp[10]) ? 11'b01011010100 : 11'b01010100000;
												assign node441 = (inp[10]) ? 11'b01111010010 : 11'b01110010110;
											assign node444 = (inp[9]) ? node446 : 11'b01111111110;
												assign node446 = (inp[10]) ? 11'b01010111000 : 11'b01001111100;
										assign node449 = (inp[10]) ? node455 : node450;
											assign node450 = (inp[8]) ? node452 : 11'b01100101011;
												assign node452 = (inp[9]) ? 11'b01001011111 : 11'b01001001011;
											assign node455 = (inp[9]) ? 11'b01111011001 : 11'b01110011101;
								assign node458 = (inp[5]) ? node482 : node459;
									assign node459 = (inp[6]) ? node469 : node460;
										assign node460 = (inp[9]) ? node466 : node461;
											assign node461 = (inp[10]) ? node463 : 11'b01110111011;
												assign node463 = (inp[8]) ? 11'b01001001101 : 11'b01110001101;
											assign node466 = (inp[10]) ? 11'b01011001001 : 11'b01011001101;
										assign node469 = (inp[8]) ? node475 : node470;
											assign node470 = (inp[10]) ? 11'b01100101111 : node471;
												assign node471 = (inp[9]) ? 11'b01001001111 : 11'b01001111001;
											assign node475 = (inp[10]) ? node479 : node476;
												assign node476 = (inp[9]) ? 11'b01110001110 : 11'b01100011000;
												assign node479 = (inp[9]) ? 11'b01001101001 : 11'b01011001100;
									assign node482 = (inp[8]) ? node492 : node483;
										assign node483 = (inp[6]) ? node489 : node484;
											assign node484 = (inp[9]) ? node486 : 11'b01100001110;
												assign node486 = (inp[10]) ? 11'b01110001010 : 11'b01111001110;
											assign node489 = (inp[10]) ? 11'b01110101100 : 11'b01111111010;
										assign node492 = (inp[9]) ? node496 : node493;
											assign node493 = (inp[10]) ? 11'b01010101110 : 11'b01010111011;
											assign node496 = (inp[10]) ? node498 : 11'b01001001110;
												assign node498 = (inp[6]) ? 11'b01000001011 : 11'b01010001010;
						assign node501 = (inp[10]) ? node581 : node502;
							assign node502 = (inp[8]) ? node544 : node503;
								assign node503 = (inp[4]) ? node521 : node504;
									assign node504 = (inp[9]) ? node510 : node505;
										assign node505 = (inp[5]) ? 11'b01101001011 : node506;
											assign node506 = (inp[6]) ? 11'b01001100000 : 11'b01001101001;
										assign node510 = (inp[5]) ? node516 : node511;
											assign node511 = (inp[6]) ? 11'b01001110010 : node512;
												assign node512 = (inp[11]) ? 11'b01101111001 : 11'b01001111001;
											assign node516 = (inp[11]) ? 11'b01011111010 : node517;
												assign node517 = (inp[6]) ? 11'b01101111001 : 11'b01101111000;
									assign node521 = (inp[9]) ? node535 : node522;
										assign node522 = (inp[6]) ? node528 : node523;
											assign node523 = (inp[5]) ? 11'b01111011000 : node524;
												assign node524 = (inp[11]) ? 11'b01111011001 : 11'b01001011001;
											assign node528 = (inp[11]) ? node532 : node529;
												assign node529 = (inp[5]) ? 11'b01111111011 : 11'b01001010000;
												assign node532 = (inp[5]) ? 11'b01001111000 : 11'b01110111001;
										assign node535 = (inp[5]) ? node541 : node536;
											assign node536 = (inp[11]) ? 11'b01110001011 : node537;
												assign node537 = (inp[6]) ? 11'b01101000010 : 11'b01101001001;
											assign node541 = (inp[6]) ? 11'b01011101010 : 11'b01011001010;
								assign node544 = (inp[5]) ? node562 : node545;
									assign node545 = (inp[4]) ? node555 : node546;
										assign node546 = (inp[9]) ? node552 : node547;
											assign node547 = (inp[6]) ? 11'b01010101010 : node548;
												assign node548 = (inp[11]) ? 11'b01011101011 : 11'b01001101001;
											assign node552 = (inp[6]) ? 11'b01101011010 : 11'b01101111011;
										assign node555 = (inp[9]) ? node557 : 11'b01111011000;
											assign node557 = (inp[11]) ? node559 : 11'b01110101000;
												assign node559 = (inp[6]) ? 11'b01111101011 : 11'b01110001001;
									assign node562 = (inp[4]) ? node570 : node563;
										assign node563 = (inp[9]) ? node567 : node564;
											assign node564 = (inp[11]) ? 11'b01110001000 : 11'b01100001001;
											assign node567 = (inp[6]) ? 11'b01010111001 : 11'b01100111010;
										assign node570 = (inp[9]) ? node576 : node571;
											assign node571 = (inp[6]) ? 11'b01110011011 : node572;
												assign node572 = (inp[11]) ? 11'b01010111010 : 11'b01110111010;
											assign node576 = (inp[6]) ? node578 : 11'b01010001010;
												assign node578 = (inp[11]) ? 11'b01010001011 : 11'b01011001011;
							assign node581 = (inp[4]) ? node627 : node582;
								assign node582 = (inp[5]) ? node602 : node583;
									assign node583 = (inp[11]) ? node589 : node584;
										assign node584 = (inp[6]) ? node586 : 11'b01000101001;
											assign node586 = (inp[9]) ? 11'b01000100000 : 11'b01000100010;
										assign node589 = (inp[9]) ? node595 : node590;
											assign node590 = (inp[8]) ? node592 : 11'b01100101001;
												assign node592 = (inp[6]) ? 11'b01110101000 : 11'b01110101011;
											assign node595 = (inp[8]) ? node599 : node596;
												assign node596 = (inp[6]) ? 11'b01011101001 : 11'b01010101001;
												assign node599 = (inp[6]) ? 11'b01010001010 : 11'b01010101011;
									assign node602 = (inp[6]) ? node616 : node603;
										assign node603 = (inp[8]) ? node611 : node604;
											assign node604 = (inp[11]) ? node608 : node605;
												assign node605 = (inp[9]) ? 11'b01010101000 : 11'b01000101000;
												assign node608 = (inp[9]) ? 11'b01000101010 : 11'b01110101010;
											assign node611 = (inp[11]) ? node613 : 11'b01011101000;
												assign node613 = (inp[9]) ? 11'b01001101010 : 11'b01101101000;
										assign node616 = (inp[11]) ? node622 : node617;
											assign node617 = (inp[8]) ? node619 : 11'b01000001011;
												assign node619 = (inp[9]) ? 11'b01011001011 : 11'b01011101011;
											assign node622 = (inp[9]) ? 11'b01001101010 : node623;
												assign node623 = (inp[8]) ? 11'b01100101011 : 11'b01111001001;
								assign node627 = (inp[9]) ? node651 : node628;
									assign node628 = (inp[11]) ? node638 : node629;
										assign node629 = (inp[8]) ? node633 : node630;
											assign node630 = (inp[6]) ? 11'b01100000010 : 11'b01100001001;
											assign node633 = (inp[5]) ? node635 : 11'b01111101010;
												assign node635 = (inp[6]) ? 11'b01100001001 : 11'b01101001010;
										assign node638 = (inp[8]) ? node646 : node639;
											assign node639 = (inp[5]) ? node643 : node640;
												assign node640 = (inp[6]) ? 11'b01011001011 : 11'b01010001001;
												assign node643 = (inp[6]) ? 11'b01010101000 : 11'b01010001010;
											assign node646 = (inp[6]) ? 11'b01000001010 : node647;
												assign node647 = (inp[5]) ? 11'b01001001010 : 11'b01001001001;
									assign node651 = (inp[11]) ? node665 : node652;
										assign node652 = (inp[6]) ? node658 : node653;
											assign node653 = (inp[5]) ? 11'b01000001010 : node654;
												assign node654 = (inp[8]) ? 11'b01000001011 : 11'b01000001001;
											assign node658 = (inp[5]) ? node662 : node659;
												assign node659 = (inp[8]) ? 11'b01001101010 : 11'b01001000000;
												assign node662 = (inp[8]) ? 11'b01000001001 : 11'b01001001011;
										assign node665 = (inp[5]) ? node671 : node666;
											assign node666 = (inp[8]) ? node668 : 11'b01000001001;
												assign node668 = (inp[6]) ? 11'b01001101001 : 11'b01001001001;
											assign node671 = (inp[8]) ? node673 : 11'b01000101000;
												assign node673 = (inp[6]) ? 11'b01000001001 : 11'b01000001000;
				assign node676 = (inp[0]) ? node1014 : node677;
					assign node677 = (inp[8]) ? node849 : node678;
						assign node678 = (inp[6]) ? node768 : node679;
							assign node679 = (inp[5]) ? node723 : node680;
								assign node680 = (inp[4]) ? node698 : node681;
									assign node681 = (inp[9]) ? node687 : node682;
										assign node682 = (inp[11]) ? 11'b01100010111 : node683;
											assign node683 = (inp[3]) ? 11'b11101001010 : 11'b01101001010;
										assign node687 = (inp[3]) ? node691 : node688;
											assign node688 = (inp[10]) ? 11'b11110110111 : 11'b01010010011;
											assign node691 = (inp[10]) ? node695 : node692;
												assign node692 = (inp[11]) ? 11'b11011100111 : 11'b11101100111;
												assign node695 = (inp[11]) ? 11'b01101110101 : 11'b01110110111;
									assign node698 = (inp[9]) ? node710 : node699;
										assign node699 = (inp[10]) ? node705 : node700;
											assign node700 = (inp[3]) ? 11'b11000100101 : node701;
												assign node701 = (inp[11]) ? 11'b01110100101 : 11'b01100100101;
											assign node705 = (inp[3]) ? node707 : 11'b11001110101;
												assign node707 = (inp[11]) ? 11'b01011110001 : 11'b01000100001;
										assign node710 = (inp[10]) ? node716 : node711;
											assign node711 = (inp[3]) ? node713 : 11'b01000100101;
												assign node713 = (inp[11]) ? 11'b11100110011 : 11'b11011010001;
											assign node716 = (inp[3]) ? node720 : node717;
												assign node717 = (inp[11]) ? 11'b11011010011 : 11'b11011000001;
												assign node720 = (inp[11]) ? 11'b01011010011 : 11'b01000010011;
								assign node723 = (inp[4]) ? node741 : node724;
									assign node724 = (inp[3]) ? node732 : node725;
										assign node725 = (inp[10]) ? 11'b11011010011 : node726;
											assign node726 = (inp[11]) ? 11'b01101010000 : node727;
												assign node727 = (inp[9]) ? 11'b01101010001 : 11'b01100010011;
										assign node732 = (inp[10]) ? node738 : node733;
											assign node733 = (inp[9]) ? node735 : 11'b11011000000;
												assign node735 = (inp[11]) ? 11'b11101010110 : 11'b11110010101;
											assign node738 = (inp[9]) ? 11'b01110000110 : 11'b01100000100;
									assign node741 = (inp[9]) ? node755 : node742;
										assign node742 = (inp[10]) ? node750 : node743;
											assign node743 = (inp[3]) ? node747 : node744;
												assign node744 = (inp[11]) ? 11'b01101110110 : 11'b01111110100;
												assign node747 = (inp[11]) ? 11'b11011110110 : 11'b11000110110;
											assign node750 = (inp[3]) ? 11'b01111110010 : node751;
												assign node751 = (inp[11]) ? 11'b11110100110 : 11'b11100100110;
										assign node755 = (inp[11]) ? node763 : node756;
											assign node756 = (inp[3]) ? node760 : node757;
												assign node757 = (inp[10]) ? 11'b11110110010 : 11'b01001110110;
												assign node760 = (inp[10]) ? 11'b01000100000 : 11'b11100100010;
											assign node763 = (inp[10]) ? node765 : 11'b01110100100;
												assign node765 = (inp[3]) ? 11'b01010100000 : 11'b11101100000;
							assign node768 = (inp[5]) ? node808 : node769;
								assign node769 = (inp[4]) ? node791 : node770;
									assign node770 = (inp[9]) ? node780 : node771;
										assign node771 = (inp[3]) ? node777 : node772;
											assign node772 = (inp[10]) ? node774 : 11'b01111001010;
												assign node774 = (inp[11]) ? 11'b11100001000 : 11'b11110001011;
											assign node777 = (inp[10]) ? 11'b01110011100 : 11'b11100011010;
										assign node780 = (inp[11]) ? node788 : node781;
											assign node781 = (inp[10]) ? node785 : node782;
												assign node782 = (inp[3]) ? 11'b11101101110 : 11'b01100001001;
												assign node785 = (inp[3]) ? 11'b01110111110 : 11'b11111111110;
											assign node788 = (inp[10]) ? 11'b11000011110 : 11'b11011001110;
									assign node791 = (inp[10]) ? node799 : node792;
										assign node792 = (inp[11]) ? node794 : 11'b01010101110;
											assign node794 = (inp[9]) ? node796 : 11'b01110001100;
												assign node796 = (inp[3]) ? 11'b11110111000 : 11'b01100111100;
										assign node799 = (inp[3]) ? node801 : 11'b11011111110;
											assign node801 = (inp[9]) ? node805 : node802;
												assign node802 = (inp[11]) ? 11'b01000111010 : 11'b01011101010;
												assign node805 = (inp[11]) ? 11'b01011111010 : 11'b01011011000;
								assign node808 = (inp[11]) ? node828 : node809;
									assign node809 = (inp[9]) ? node819 : node810;
										assign node810 = (inp[3]) ? node814 : node811;
											assign node811 = (inp[10]) ? 11'b11110001110 : 11'b01111011100;
											assign node814 = (inp[10]) ? node816 : 11'b11100111000;
												assign node816 = (inp[4]) ? 11'b01100011000 : 11'b01011011100;
										assign node819 = (inp[4]) ? node823 : node820;
											assign node820 = (inp[3]) ? 11'b01100001100 : 11'b11000001100;
											assign node823 = (inp[3]) ? 11'b11101100011 : node824;
												assign node824 = (inp[10]) ? 11'b11111110011 : 11'b01000011100;
									assign node828 = (inp[4]) ? node838 : node829;
										assign node829 = (inp[10]) ? node835 : node830;
											assign node830 = (inp[3]) ? 11'b11110110101 : node831;
												assign node831 = (inp[9]) ? 11'b01001100001 : 11'b01110110001;
											assign node835 = (inp[9]) ? 11'b01111000111 : 11'b01101100111;
										assign node838 = (inp[3]) ? node846 : node839;
											assign node839 = (inp[10]) ? node843 : node840;
												assign node840 = (inp[9]) ? 11'b01111000111 : 11'b01101010111;
												assign node843 = (inp[9]) ? 11'b11111000001 : 11'b11100000101;
											assign node846 = (inp[9]) ? 11'b01010000001 : 11'b01000000011;
						assign node849 = (inp[5]) ? node933 : node850;
							assign node850 = (inp[11]) ? node896 : node851;
								assign node851 = (inp[10]) ? node873 : node852;
									assign node852 = (inp[3]) ? node864 : node853;
										assign node853 = (inp[4]) ? node861 : node854;
											assign node854 = (inp[9]) ? node858 : node855;
												assign node855 = (inp[6]) ? 11'b01100000011 : 11'b01100100010;
												assign node858 = (inp[6]) ? 11'b01110100001 : 11'b01110000010;
											assign node861 = (inp[9]) ? 11'b01010100111 : 11'b01000000100;
										assign node864 = (inp[6]) ? node870 : node865;
											assign node865 = (inp[9]) ? 11'b11000000100 : node866;
												assign node866 = (inp[4]) ? 11'b11110000100 : 11'b11011000010;
											assign node870 = (inp[4]) ? 11'b11100100111 : 11'b11001100011;
									assign node873 = (inp[3]) ? node883 : node874;
										assign node874 = (inp[4]) ? node878 : node875;
											assign node875 = (inp[6]) ? 11'b11101100001 : 11'b11101010100;
											assign node878 = (inp[9]) ? node880 : 11'b11001110111;
												assign node880 = (inp[6]) ? 11'b11110000011 : 11'b11111100011;
										assign node883 = (inp[9]) ? node889 : node884;
											assign node884 = (inp[4]) ? 11'b01101100011 : node885;
												assign node885 = (inp[6]) ? 11'b01001100101 : 11'b01000000110;
											assign node889 = (inp[4]) ? node893 : node890;
												assign node890 = (inp[6]) ? 11'b01011110101 : 11'b01011010100;
												assign node893 = (inp[6]) ? 11'b01010010011 : 11'b01001110001;
								assign node896 = (inp[4]) ? node914 : node897;
									assign node897 = (inp[3]) ? node905 : node898;
										assign node898 = (inp[6]) ? node902 : node899;
											assign node899 = (inp[10]) ? 11'b11000100001 : 11'b01101100001;
											assign node902 = (inp[9]) ? 11'b01000010001 : 11'b01110000001;
										assign node905 = (inp[10]) ? node911 : node906;
											assign node906 = (inp[9]) ? 11'b11010000111 : node907;
												assign node907 = (inp[6]) ? 11'b11011010001 : 11'b11010110001;
											assign node911 = (inp[9]) ? 11'b01001010111 : 11'b01100010111;
									assign node914 = (inp[10]) ? node926 : node915;
										assign node915 = (inp[9]) ? node919 : node916;
											assign node916 = (inp[6]) ? 11'b11110100100 : 11'b11101000101;
											assign node919 = (inp[3]) ? node923 : node920;
												assign node920 = (inp[6]) ? 11'b01111110110 : 11'b01101110101;
												assign node923 = (inp[6]) ? 11'b11111110000 : 11'b11111110001;
										assign node926 = (inp[3]) ? node930 : node927;
											assign node927 = (inp[6]) ? 11'b11010110100 : 11'b11010010101;
											assign node930 = (inp[9]) ? 11'b01010110011 : 11'b01011110010;
							assign node933 = (inp[11]) ? node979 : node934;
								assign node934 = (inp[6]) ? node962 : node935;
									assign node935 = (inp[3]) ? node949 : node936;
										assign node936 = (inp[10]) ? node942 : node937;
											assign node937 = (inp[4]) ? node939 : 11'b01110110001;
												assign node939 = (inp[9]) ? 11'b01010010101 : 11'b01010010111;
											assign node942 = (inp[4]) ? node946 : node943;
												assign node943 = (inp[9]) ? 11'b11111000101 : 11'b11001110001;
												assign node946 = (inp[9]) ? 11'b11011110000 : 11'b11111000111;
										assign node949 = (inp[10]) ? node955 : node950;
											assign node950 = (inp[9]) ? node952 : 11'b11101010111;
												assign node952 = (inp[4]) ? 11'b11000000001 : 11'b11101010101;
											assign node955 = (inp[9]) ? node959 : node956;
												assign node956 = (inp[4]) ? 11'b01101010001 : 11'b01010110101;
												assign node959 = (inp[4]) ? 11'b01001100010 : 11'b01000000111;
									assign node962 = (inp[4]) ? node970 : node963;
										assign node963 = (inp[3]) ? node965 : 11'b11101000100;
											assign node965 = (inp[10]) ? 11'b01000010110 : node966;
												assign node966 = (inp[9]) ? 11'b11100010100 : 11'b11101010000;
										assign node970 = (inp[9]) ? node972 : 11'b01000010110;
											assign node972 = (inp[10]) ? node976 : node973;
												assign node973 = (inp[3]) ? 11'b11010100010 : 11'b01011110110;
												assign node976 = (inp[3]) ? 11'b01010100000 : 11'b11010110000;
								assign node979 = (inp[4]) ? node995 : node980;
									assign node980 = (inp[3]) ? node988 : node981;
										assign node981 = (inp[6]) ? node985 : node982;
											assign node982 = (inp[9]) ? 11'b01101100000 : 11'b11101110010;
											assign node985 = (inp[10]) ? 11'b11011000100 : 11'b01110100010;
										assign node988 = (inp[9]) ? node992 : node989;
											assign node989 = (inp[6]) ? 11'b01110100100 : 11'b01111100110;
											assign node992 = (inp[10]) ? 11'b01011000100 : 11'b11011010110;
									assign node995 = (inp[9]) ? node1003 : node996;
										assign node996 = (inp[10]) ? node1000 : node997;
											assign node997 = (inp[6]) ? 11'b01010010110 : 11'b11010010110;
											assign node1000 = (inp[3]) ? 11'b01011000010 : 11'b11000000110;
										assign node1003 = (inp[10]) ? node1009 : node1004;
											assign node1004 = (inp[3]) ? node1006 : 11'b01011000110;
												assign node1006 = (inp[6]) ? 11'b11010000010 : 11'b11011000000;
											assign node1009 = (inp[3]) ? 11'b01010000000 : node1010;
												assign node1010 = (inp[6]) ? 11'b11010000000 : 11'b11000000000;
					assign node1014 = (inp[3]) ? node1204 : node1015;
						assign node1015 = (inp[6]) ? node1111 : node1016;
							assign node1016 = (inp[5]) ? node1066 : node1017;
								assign node1017 = (inp[11]) ? node1041 : node1018;
									assign node1018 = (inp[9]) ? node1028 : node1019;
										assign node1019 = (inp[8]) ? node1023 : node1020;
											assign node1020 = (inp[10]) ? 11'b01010001100 : 11'b01001001000;
											assign node1023 = (inp[10]) ? 11'b01101000100 : node1024;
												assign node1024 = (inp[4]) ? 11'b01100000010 : 11'b01100100000;
										assign node1028 = (inp[10]) ? node1034 : node1029;
											assign node1029 = (inp[8]) ? 11'b01110000100 : node1030;
												assign node1030 = (inp[4]) ? 11'b01101010111 : 11'b01001100101;
											assign node1034 = (inp[8]) ? node1038 : node1035;
												assign node1035 = (inp[4]) ? 11'b01110010011 : 11'b01010110001;
												assign node1038 = (inp[4]) ? 11'b01011110001 : 11'b01111010010;
									assign node1041 = (inp[9]) ? node1055 : node1042;
										assign node1042 = (inp[10]) ? node1050 : node1043;
											assign node1043 = (inp[8]) ? node1047 : node1044;
												assign node1044 = (inp[4]) ? 11'b01010110011 : 11'b01010010001;
												assign node1047 = (inp[4]) ? 11'b01111010001 : 11'b01110110011;
											assign node1050 = (inp[4]) ? 11'b01010000111 : node1051;
												assign node1051 = (inp[8]) ? 11'b01101010111 : 11'b01001010101;
										assign node1055 = (inp[10]) ? node1059 : node1056;
											assign node1056 = (inp[8]) ? 11'b01001010101 : 11'b01000100101;
											assign node1059 = (inp[8]) ? node1063 : node1060;
												assign node1060 = (inp[4]) ? 11'b01111000001 : 11'b01001100011;
												assign node1063 = (inp[4]) ? 11'b01010100001 : 11'b01100000001;
								assign node1066 = (inp[11]) ? node1090 : node1067;
									assign node1067 = (inp[4]) ? node1079 : node1068;
										assign node1068 = (inp[8]) ? node1074 : node1069;
											assign node1069 = (inp[10]) ? 11'b01111000101 : node1070;
												assign node1070 = (inp[9]) ? 11'b01010000111 : 11'b01000000001;
											assign node1074 = (inp[10]) ? 11'b01001010001 : node1075;
												assign node1075 = (inp[9]) ? 11'b01101000111 : 11'b01101100001;
										assign node1079 = (inp[8]) ? node1083 : node1080;
											assign node1080 = (inp[10]) ? 11'b01010110100 : 11'b01101110100;
											assign node1083 = (inp[9]) ? node1087 : node1084;
												assign node1084 = (inp[10]) ? 11'b01111010101 : 11'b01000000001;
												assign node1087 = (inp[10]) ? 11'b01011110010 : 11'b01010010111;
									assign node1090 = (inp[10]) ? node1102 : node1091;
										assign node1091 = (inp[9]) ? node1097 : node1092;
											assign node1092 = (inp[8]) ? node1094 : 11'b01101110000;
												assign node1094 = (inp[4]) ? 11'b01011010000 : 11'b01110110000;
											assign node1097 = (inp[8]) ? 11'b01010110110 : node1098;
												assign node1098 = (inp[4]) ? 11'b01111100110 : 11'b01111010110;
										assign node1102 = (inp[9]) ? node1106 : node1103;
											assign node1103 = (inp[4]) ? 11'b01010000100 : 11'b01000010110;
											assign node1106 = (inp[8]) ? node1108 : 11'b01110000000;
												assign node1108 = (inp[4]) ? 11'b01010000010 : 11'b01011000010;
							assign node1111 = (inp[8]) ? node1155 : node1112;
								assign node1112 = (inp[5]) ? node1134 : node1113;
									assign node1113 = (inp[4]) ? node1121 : node1114;
										assign node1114 = (inp[9]) ? node1118 : node1115;
											assign node1115 = (inp[11]) ? 11'b01001011000 : 11'b01011001001;
											assign node1118 = (inp[10]) ? 11'b01001111000 : 11'b01011101110;
										assign node1121 = (inp[10]) ? node1129 : node1122;
											assign node1122 = (inp[9]) ? node1126 : node1123;
												assign node1123 = (inp[11]) ? 11'b01001111010 : 11'b01010101010;
												assign node1126 = (inp[11]) ? 11'b01010101110 : 11'b01110111100;
											assign node1129 = (inp[9]) ? 11'b01101011010 : node1130;
												assign node1130 = (inp[11]) ? 11'b01111101100 : 11'b01001111100;
									assign node1134 = (inp[11]) ? node1146 : node1135;
										assign node1135 = (inp[4]) ? node1141 : node1136;
											assign node1136 = (inp[10]) ? 11'b01110011010 : node1137;
												assign node1137 = (inp[9]) ? 11'b01001001100 : 11'b01010101000;
											assign node1141 = (inp[9]) ? node1143 : 11'b01000011110;
												assign node1143 = (inp[10]) ? 11'b01101110001 : 11'b01111110111;
										assign node1146 = (inp[4]) ? node1152 : node1147;
											assign node1147 = (inp[10]) ? 11'b01100100001 : node1148;
												assign node1148 = (inp[9]) ? 11'b01100110111 : 11'b01000110011;
											assign node1152 = (inp[9]) ? 11'b01100000011 : 11'b01111010001;
								assign node1155 = (inp[5]) ? node1179 : node1156;
									assign node1156 = (inp[4]) ? node1170 : node1157;
										assign node1157 = (inp[10]) ? node1163 : node1158;
											assign node1158 = (inp[11]) ? 11'b01101010011 : node1159;
												assign node1159 = (inp[9]) ? 11'b01100100101 : 11'b01110000001;
											assign node1163 = (inp[11]) ? node1167 : node1164;
												assign node1164 = (inp[9]) ? 11'b01101110011 : 11'b01111100111;
												assign node1167 = (inp[9]) ? 11'b01111100000 : 11'b01111010101;
										assign node1170 = (inp[9]) ? node1176 : node1171;
											assign node1171 = (inp[10]) ? 11'b01110110101 : node1172;
												assign node1172 = (inp[11]) ? 11'b01100110010 : 11'b01110100011;
											assign node1176 = (inp[10]) ? 11'b01000010001 : 11'b01011010111;
									assign node1179 = (inp[10]) ? node1195 : node1180;
										assign node1180 = (inp[9]) ? node1188 : node1181;
											assign node1181 = (inp[11]) ? node1185 : node1182;
												assign node1182 = (inp[4]) ? 11'b01010000000 : 11'b01111000000;
												assign node1185 = (inp[4]) ? 11'b01000010000 : 11'b01101110000;
											assign node1188 = (inp[4]) ? node1192 : node1189;
												assign node1189 = (inp[11]) ? 11'b01000110100 : 11'b01110000100;
												assign node1192 = (inp[11]) ? 11'b01001000100 : 11'b01001110100;
										assign node1195 = (inp[11]) ? node1201 : node1196;
											assign node1196 = (inp[9]) ? node1198 : 11'b01101110110;
												assign node1198 = (inp[4]) ? 11'b01000110010 : 11'b01011010010;
											assign node1201 = (inp[4]) ? 11'b01001000110 : 11'b01001000010;
						assign node1204 = (inp[10]) ? node1292 : node1205;
							assign node1205 = (inp[8]) ? node1241 : node1206;
								assign node1206 = (inp[11]) ? node1222 : node1207;
									assign node1207 = (inp[5]) ? node1219 : node1208;
										assign node1208 = (inp[4]) ? node1216 : node1209;
											assign node1209 = (inp[9]) ? node1213 : node1210;
												assign node1210 = (inp[6]) ? 11'b01011001001 : 11'b01011001000;
												assign node1213 = (inp[6]) ? 11'b01011111000 : 11'b01011110001;
											assign node1216 = (inp[6]) ? 11'b01011111010 : 11'b01011110011;
										assign node1219 = (inp[4]) ? 11'b01101011000 : 11'b01110101010;
									assign node1222 = (inp[5]) ? node1230 : node1223;
										assign node1223 = (inp[6]) ? node1225 : 11'b01100100001;
											assign node1225 = (inp[4]) ? node1227 : 11'b01111011000;
												assign node1227 = (inp[9]) ? 11'b01101101010 : 11'b01101111000;
										assign node1230 = (inp[9]) ? node1236 : node1231;
											assign node1231 = (inp[4]) ? 11'b01011110000 : node1232;
												assign node1232 = (inp[6]) ? 11'b01111100011 : 11'b01110000010;
											assign node1236 = (inp[4]) ? node1238 : 11'b01001010000;
												assign node1238 = (inp[6]) ? 11'b01001000011 : 11'b01001100010;
								assign node1241 = (inp[5]) ? node1265 : node1242;
									assign node1242 = (inp[9]) ? node1252 : node1243;
										assign node1243 = (inp[11]) ? node1249 : node1244;
											assign node1244 = (inp[4]) ? 11'b01011110011 : node1245;
												assign node1245 = (inp[6]) ? 11'b01011100001 : 11'b01011000000;
											assign node1249 = (inp[4]) ? 11'b01100110010 : 11'b01000100011;
										assign node1252 = (inp[4]) ? node1260 : node1253;
											assign node1253 = (inp[11]) ? node1257 : node1254;
												assign node1254 = (inp[6]) ? 11'b01000110001 : 11'b01001010010;
												assign node1257 = (inp[6]) ? 11'b01111110010 : 11'b01110010001;
											assign node1260 = (inp[6]) ? 11'b01101000001 : node1261;
												assign node1261 = (inp[11]) ? 11'b01101100001 : 11'b01100100001;
									assign node1265 = (inp[11]) ? node1281 : node1266;
										assign node1266 = (inp[4]) ? node1274 : node1267;
											assign node1267 = (inp[9]) ? node1271 : node1268;
												assign node1268 = (inp[6]) ? 11'b01111000010 : 11'b01111100001;
												assign node1271 = (inp[6]) ? 11'b01111010010 : 11'b01111010011;
											assign node1274 = (inp[9]) ? node1278 : node1275;
												assign node1275 = (inp[6]) ? 11'b01100010010 : 11'b01101010001;
												assign node1278 = (inp[6]) ? 11'b01000100010 : 11'b01001100010;
										assign node1281 = (inp[4]) ? node1287 : node1282;
											assign node1282 = (inp[9]) ? node1284 : 11'b01101100010;
												assign node1284 = (inp[6]) ? 11'b01001010010 : 11'b01000110010;
											assign node1287 = (inp[6]) ? node1289 : 11'b01000010000;
												assign node1289 = (inp[9]) ? 11'b01000000010 : 11'b01000010010;
							assign node1292 = (inp[9]) ? node1328 : node1293;
								assign node1293 = (inp[6]) ? node1313 : node1294;
									assign node1294 = (inp[4]) ? node1304 : node1295;
										assign node1295 = (inp[11]) ? node1299 : node1296;
											assign node1296 = (inp[5]) ? 11'b01001000011 : 11'b01010000000;
											assign node1299 = (inp[5]) ? node1301 : 11'b01111000011;
												assign node1301 = (inp[8]) ? 11'b01101100010 : 11'b01111000010;
										assign node1304 = (inp[11]) ? node1310 : node1305;
											assign node1305 = (inp[8]) ? 11'b01100000011 : node1306;
												assign node1306 = (inp[5]) ? 11'b01111100000 : 11'b01100100011;
											assign node1310 = (inp[5]) ? 11'b01010100010 : 11'b01010100011;
									assign node1313 = (inp[8]) ? node1323 : node1314;
										assign node1314 = (inp[4]) ? node1320 : node1315;
											assign node1315 = (inp[11]) ? 11'b01101001010 : node1316;
												assign node1316 = (inp[5]) ? 11'b01001001000 : 11'b01000001011;
											assign node1320 = (inp[5]) ? 11'b01110001010 : 11'b01010101000;
										assign node1323 = (inp[11]) ? 11'b01001100000 : node1324;
											assign node1324 = (inp[5]) ? 11'b01101100000 : 11'b01111000011;
								assign node1328 = (inp[5]) ? node1350 : node1329;
									assign node1329 = (inp[11]) ? node1343 : node1330;
										assign node1330 = (inp[8]) ? node1336 : node1331;
											assign node1331 = (inp[6]) ? 11'b01001001000 : node1332;
												assign node1332 = (inp[4]) ? 11'b01000000001 : 11'b01000100011;
											assign node1336 = (inp[6]) ? node1340 : node1337;
												assign node1337 = (inp[4]) ? 11'b01001100011 : 11'b01000000010;
												assign node1340 = (inp[4]) ? 11'b01000000011 : 11'b01001100011;
										assign node1343 = (inp[4]) ? node1347 : node1344;
											assign node1344 = (inp[8]) ? 11'b01011000001 : 11'b01010100011;
											assign node1347 = (inp[6]) ? 11'b01000100000 : 11'b01000100001;
									assign node1350 = (inp[11]) ? node1360 : node1351;
										assign node1351 = (inp[8]) ? node1357 : node1352;
											assign node1352 = (inp[6]) ? 11'b01011001010 : node1353;
												assign node1353 = (inp[4]) ? 11'b01001000010 : 11'b01011100010;
											assign node1357 = (inp[6]) ? 11'b01000100000 : 11'b01010000001;
										assign node1360 = (inp[4]) ? node1364 : node1361;
											assign node1361 = (inp[8]) ? 11'b01001000000 : 11'b01000000000;
											assign node1364 = (inp[6]) ? node1368 : node1365;
												assign node1365 = (inp[8]) ? 11'b01000000000 : 11'b01000100000;
												assign node1368 = (inp[8]) ? 11'b01000000000 : 11'b01000000001;
			assign node1371 = (inp[6]) ? node2025 : node1372;
				assign node1372 = (inp[2]) ? node1710 : node1373;
					assign node1373 = (inp[8]) ? node1553 : node1374;
						assign node1374 = (inp[5]) ? node1468 : node1375;
							assign node1375 = (inp[0]) ? node1421 : node1376;
								assign node1376 = (inp[10]) ? node1398 : node1377;
									assign node1377 = (inp[3]) ? node1389 : node1378;
										assign node1378 = (inp[4]) ? node1384 : node1379;
											assign node1379 = (inp[11]) ? 11'b01110010011 : node1380;
												assign node1380 = (inp[9]) ? 11'b01010100011 : 11'b01011100011;
											assign node1384 = (inp[9]) ? 11'b01111000111 : node1385;
												assign node1385 = (inp[11]) ? 11'b01000100111 : 11'b01010100111;
										assign node1389 = (inp[4]) ? node1393 : node1390;
											assign node1390 = (inp[11]) ? 11'b11111100111 : 11'b11011100011;
											assign node1393 = (inp[11]) ? 11'b11001110001 : node1394;
												assign node1394 = (inp[9]) ? 11'b11110010011 : 11'b11010100111;
									assign node1398 = (inp[4]) ? node1410 : node1399;
										assign node1399 = (inp[3]) ? node1407 : node1400;
											assign node1400 = (inp[9]) ? node1404 : node1401;
												assign node1401 = (inp[11]) ? 11'b11011000001 : 11'b11011100001;
												assign node1404 = (inp[11]) ? 11'b11111110101 : 11'b11011110101;
											assign node1407 = (inp[11]) ? 11'b01010010101 : 11'b01010100101;
										assign node1410 = (inp[11]) ? node1416 : node1411;
											assign node1411 = (inp[9]) ? node1413 : 11'b11010110101;
												assign node1413 = (inp[3]) ? 11'b01110010001 : 11'b11110000001;
											assign node1416 = (inp[3]) ? 11'b01100110011 : node1417;
												assign node1417 = (inp[9]) ? 11'b11100110001 : 11'b11100110101;
								assign node1421 = (inp[11]) ? node1443 : node1422;
									assign node1422 = (inp[4]) ? node1430 : node1423;
										assign node1423 = (inp[9]) ? node1425 : 11'b01000100111;
											assign node1425 = (inp[10]) ? node1427 : 11'b01001110011;
												assign node1427 = (inp[3]) ? 11'b01001100001 : 11'b01001110011;
										assign node1430 = (inp[10]) ? node1436 : node1431;
											assign node1431 = (inp[9]) ? 11'b01101010101 : node1432;
												assign node1432 = (inp[3]) ? 11'b01000110011 : 11'b01000100001;
											assign node1436 = (inp[3]) ? node1440 : node1437;
												assign node1437 = (inp[9]) ? 11'b01100010011 : 11'b01001010111;
												assign node1440 = (inp[9]) ? 11'b01000000001 : 11'b01101000001;
									assign node1443 = (inp[4]) ? node1455 : node1444;
										assign node1444 = (inp[3]) ? node1450 : node1445;
											assign node1445 = (inp[9]) ? 11'b01100010101 : node1446;
												assign node1446 = (inp[10]) ? 11'b01000010111 : 11'b01001010001;
											assign node1450 = (inp[10]) ? node1452 : 11'b01101110011;
												assign node1452 = (inp[9]) ? 11'b01011100001 : 11'b01100000001;
										assign node1455 = (inp[3]) ? node1463 : node1456;
											assign node1456 = (inp[10]) ? node1460 : node1457;
												assign node1457 = (inp[9]) ? 11'b01011100101 : 11'b01010110001;
												assign node1460 = (inp[9]) ? 11'b01110100011 : 11'b01111100111;
											assign node1463 = (inp[10]) ? 11'b01000100001 : node1464;
												assign node1464 = (inp[9]) ? 11'b01110100011 : 11'b01110110011;
							assign node1468 = (inp[11]) ? node1510 : node1469;
								assign node1469 = (inp[4]) ? node1491 : node1470;
									assign node1470 = (inp[0]) ? node1480 : node1471;
										assign node1471 = (inp[10]) ? node1477 : node1472;
											assign node1472 = (inp[3]) ? 11'b11011010001 : node1473;
												assign node1473 = (inp[9]) ? 11'b01010010011 : 11'b01011010011;
											assign node1477 = (inp[3]) ? 11'b01110010111 : 11'b11111000101;
										assign node1480 = (inp[10]) ? node1486 : node1481;
											assign node1481 = (inp[3]) ? 11'b01101010011 : node1482;
												assign node1482 = (inp[9]) ? 11'b01000000111 : 11'b01001000011;
											assign node1486 = (inp[3]) ? 11'b01000000001 : node1487;
												assign node1487 = (inp[9]) ? 11'b01101010001 : 11'b01101000101;
									assign node1491 = (inp[9]) ? node1501 : node1492;
										assign node1492 = (inp[0]) ? node1496 : node1493;
											assign node1493 = (inp[10]) ? 11'b11000000111 : 11'b11100010101;
											assign node1496 = (inp[3]) ? node1498 : 11'b01010010101;
												assign node1498 = (inp[10]) ? 11'b01111100000 : 11'b01110010011;
										assign node1501 = (inp[3]) ? node1507 : node1502;
											assign node1502 = (inp[10]) ? 11'b11010110010 : node1503;
												assign node1503 = (inp[0]) ? 11'b01111110110 : 11'b01101110100;
											assign node1507 = (inp[0]) ? 11'b01001100000 : 11'b11011100000;
								assign node1510 = (inp[4]) ? node1530 : node1511;
									assign node1511 = (inp[3]) ? node1519 : node1512;
										assign node1512 = (inp[0]) ? node1516 : node1513;
											assign node1513 = (inp[9]) ? 11'b01100100000 : 11'b01010110000;
											assign node1516 = (inp[9]) ? 11'b01110110110 : 11'b01001110010;
										assign node1519 = (inp[9]) ? node1527 : node1520;
											assign node1520 = (inp[10]) ? node1524 : node1521;
												assign node1521 = (inp[0]) ? 11'b01101100000 : 11'b11111100000;
												assign node1524 = (inp[0]) ? 11'b01110100010 : 11'b01001100100;
											assign node1527 = (inp[0]) ? 11'b01001000010 : 11'b01011000100;
									assign node1530 = (inp[10]) ? node1542 : node1531;
										assign node1531 = (inp[3]) ? node1539 : node1532;
											assign node1532 = (inp[9]) ? node1536 : node1533;
												assign node1533 = (inp[0]) ? 11'b01101010000 : 11'b01011010100;
												assign node1536 = (inp[0]) ? 11'b01111000100 : 11'b01001000110;
											assign node1539 = (inp[9]) ? 11'b11101000010 : 11'b11110010110;
										assign node1542 = (inp[3]) ? node1546 : node1543;
											assign node1543 = (inp[9]) ? 11'b01110000010 : 11'b11010000110;
											assign node1546 = (inp[9]) ? node1550 : node1547;
												assign node1547 = (inp[0]) ? 11'b01011000010 : 11'b01110000000;
												assign node1550 = (inp[0]) ? 11'b01000000000 : 11'b01100000000;
						assign node1553 = (inp[5]) ? node1629 : node1554;
							assign node1554 = (inp[11]) ? node1600 : node1555;
								assign node1555 = (inp[0]) ? node1579 : node1556;
									assign node1556 = (inp[9]) ? node1568 : node1557;
										assign node1557 = (inp[4]) ? node1565 : node1558;
											assign node1558 = (inp[3]) ? node1562 : node1559;
												assign node1559 = (inp[10]) ? 11'b11011100000 : 11'b01010000010;
												assign node1562 = (inp[10]) ? 11'b01111100100 : 11'b11111100010;
											assign node1565 = (inp[3]) ? 11'b11011100100 : 11'b11110110100;
										assign node1568 = (inp[4]) ? node1574 : node1569;
											assign node1569 = (inp[10]) ? node1571 : 11'b01000100010;
												assign node1571 = (inp[3]) ? 11'b01101110110 : 11'b11000110100;
											assign node1574 = (inp[10]) ? node1576 : 11'b11001010000;
												assign node1576 = (inp[3]) ? 11'b01110010010 : 11'b11011000010;
									assign node1579 = (inp[3]) ? node1591 : node1580;
										assign node1580 = (inp[10]) ? node1584 : node1581;
											assign node1581 = (inp[9]) ? 11'b01110100100 : 11'b01100000000;
											assign node1584 = (inp[4]) ? node1588 : node1585;
												assign node1585 = (inp[9]) ? 11'b01111110010 : 11'b01101100110;
												assign node1588 = (inp[9]) ? 11'b01001010000 : 11'b01100110100;
										assign node1591 = (inp[4]) ? node1597 : node1592;
											assign node1592 = (inp[10]) ? 11'b01001100000 : node1593;
												assign node1593 = (inp[9]) ? 11'b01010110010 : 11'b01001100010;
											assign node1597 = (inp[10]) ? 11'b01000000010 : 11'b01111000010;
								assign node1600 = (inp[4]) ? node1614 : node1601;
									assign node1601 = (inp[3]) ? node1609 : node1602;
										assign node1602 = (inp[10]) ? node1606 : node1603;
											assign node1603 = (inp[0]) ? 11'b01001010100 : 11'b01101010000;
											assign node1606 = (inp[9]) ? 11'b01100000010 : 11'b11101000010;
										assign node1609 = (inp[9]) ? node1611 : 11'b01010000000;
											assign node1611 = (inp[10]) ? 11'b01110010100 : 11'b01100010000;
									assign node1614 = (inp[0]) ? node1622 : node1615;
										assign node1615 = (inp[10]) ? node1619 : node1616;
											assign node1616 = (inp[3]) ? 11'b10001101111 : 11'b00101101111;
											assign node1619 = (inp[9]) ? 11'b00101111011 : 11'b10101111101;
										assign node1622 = (inp[10]) ? node1624 : 11'b00111111001;
											assign node1624 = (inp[9]) ? 11'b00011101011 : node1625;
												assign node1625 = (inp[3]) ? 11'b00000101001 : 11'b00000101111;
							assign node1629 = (inp[0]) ? node1673 : node1630;
								assign node1630 = (inp[9]) ? node1652 : node1631;
									assign node1631 = (inp[4]) ? node1643 : node1632;
										assign node1632 = (inp[11]) ? node1640 : node1633;
											assign node1633 = (inp[10]) ? node1637 : node1634;
												assign node1634 = (inp[3]) ? 11'b10010111001 : 11'b00010111011;
												assign node1637 = (inp[3]) ? 11'b00101011111 : 11'b10110111001;
											assign node1640 = (inp[3]) ? 11'b10001101001 : 11'b10000111001;
										assign node1643 = (inp[11]) ? 11'b10101001111 : node1644;
											assign node1644 = (inp[10]) ? node1648 : node1645;
												assign node1645 = (inp[3]) ? 11'b10001011111 : 11'b00100011101;
												assign node1648 = (inp[3]) ? 11'b00011011001 : 11'b10011001111;
									assign node1652 = (inp[4]) ? node1660 : node1653;
										assign node1653 = (inp[10]) ? node1657 : node1654;
											assign node1654 = (inp[11]) ? 11'b10111111101 : 11'b10011011101;
											assign node1657 = (inp[11]) ? 11'b00100101111 : 11'b00110001111;
										assign node1660 = (inp[3]) ? node1666 : node1661;
											assign node1661 = (inp[10]) ? 11'b10100011001 : node1662;
												assign node1662 = (inp[11]) ? 11'b00111001101 : 11'b00110011101;
											assign node1666 = (inp[10]) ? node1670 : node1667;
												assign node1667 = (inp[11]) ? 11'b10110001011 : 11'b10100001011;
												assign node1670 = (inp[11]) ? 11'b00100001001 : 11'b00111101001;
								assign node1673 = (inp[9]) ? node1691 : node1674;
									assign node1674 = (inp[11]) ? node1684 : node1675;
										assign node1675 = (inp[3]) ? node1679 : node1676;
											assign node1676 = (inp[10]) ? 11'b00010101101 : 11'b00011001011;
											assign node1679 = (inp[10]) ? node1681 : 11'b00100101011;
												assign node1681 = (inp[4]) ? 11'b00100001011 : 11'b00011001001;
										assign node1684 = (inp[4]) ? node1688 : node1685;
											assign node1685 = (inp[3]) ? 11'b00110101011 : 11'b00101111001;
											assign node1688 = (inp[3]) ? 11'b00010111001 : 11'b00000111011;
									assign node1691 = (inp[10]) ? node1701 : node1692;
										assign node1692 = (inp[4]) ? node1696 : node1693;
											assign node1693 = (inp[11]) ? 11'b00011111011 : 11'b00101011001;
											assign node1696 = (inp[3]) ? 11'b00010001001 : node1697;
												assign node1697 = (inp[11]) ? 11'b00001001101 : 11'b00010011101;
										assign node1701 = (inp[11]) ? node1707 : node1702;
											assign node1702 = (inp[4]) ? node1704 : 11'b00010001011;
												assign node1704 = (inp[3]) ? 11'b00001101001 : 11'b00001111011;
											assign node1707 = (inp[3]) ? 11'b00000001001 : 11'b00010001011;
					assign node1710 = (inp[0]) ? node1876 : node1711;
						assign node1711 = (inp[8]) ? node1797 : node1712;
							assign node1712 = (inp[9]) ? node1754 : node1713;
								assign node1713 = (inp[10]) ? node1731 : node1714;
									assign node1714 = (inp[5]) ? node1722 : node1715;
										assign node1715 = (inp[4]) ? node1719 : node1716;
											assign node1716 = (inp[3]) ? 11'b10111001011 : 11'b00111001011;
											assign node1719 = (inp[3]) ? 11'b10110101100 : 11'b00111101100;
										assign node1722 = (inp[4]) ? node1728 : node1723;
											assign node1723 = (inp[11]) ? 11'b00111011000 : node1724;
												assign node1724 = (inp[3]) ? 11'b10110111000 : 11'b00110111010;
											assign node1728 = (inp[11]) ? 11'b00110111111 : 11'b00100111110;
									assign node1731 = (inp[3]) ? node1739 : node1732;
										assign node1732 = (inp[11]) ? node1734 : 11'b10111001100;
											assign node1734 = (inp[4]) ? 11'b10010011110 : node1735;
												assign node1735 = (inp[5]) ? 11'b10010011010 : 11'b10101001000;
										assign node1739 = (inp[4]) ? node1747 : node1740;
											assign node1740 = (inp[5]) ? node1744 : node1741;
												assign node1741 = (inp[11]) ? 11'b00111011110 : 11'b00100001111;
												assign node1744 = (inp[11]) ? 11'b00110001100 : 11'b00011111110;
											assign node1747 = (inp[5]) ? node1751 : node1748;
												assign node1748 = (inp[11]) ? 11'b00000011000 : 11'b00010101000;
												assign node1751 = (inp[11]) ? 11'b00011101011 : 11'b00101011010;
								assign node1754 = (inp[5]) ? node1776 : node1755;
									assign node1755 = (inp[4]) ? node1767 : node1756;
										assign node1756 = (inp[10]) ? node1762 : node1757;
											assign node1757 = (inp[11]) ? node1759 : 11'b00110001011;
												assign node1759 = (inp[3]) ? 11'b10000001100 : 11'b00001011000;
											assign node1762 = (inp[11]) ? node1764 : 11'b10101111110;
												assign node1764 = (inp[3]) ? 11'b00111011110 : 11'b10010011110;
										assign node1767 = (inp[3]) ? node1771 : node1768;
											assign node1768 = (inp[10]) ? 11'b10001101000 : 11'b00011101100;
											assign node1771 = (inp[10]) ? 11'b00001111010 : node1772;
												assign node1772 = (inp[11]) ? 11'b10111111010 : 11'b10001111010;
									assign node1776 = (inp[11]) ? node1788 : node1777;
										assign node1777 = (inp[4]) ? node1783 : node1778;
											assign node1778 = (inp[10]) ? 11'b00110101100 : node1779;
												assign node1779 = (inp[3]) ? 11'b10101111110 : 11'b00111111000;
											assign node1783 = (inp[3]) ? node1785 : 11'b00010011110;
												assign node1785 = (inp[10]) ? 11'b00011001010 : 11'b10110001000;
										assign node1788 = (inp[4]) ? node1792 : node1789;
											assign node1789 = (inp[3]) ? 11'b00101101111 : 11'b10001101101;
											assign node1792 = (inp[10]) ? node1794 : 11'b00101101101;
												assign node1794 = (inp[3]) ? 11'b00000101001 : 11'b10110101011;
							assign node1797 = (inp[5]) ? node1837 : node1798;
								assign node1798 = (inp[9]) ? node1820 : node1799;
									assign node1799 = (inp[4]) ? node1811 : node1800;
										assign node1800 = (inp[3]) ? node1806 : node1801;
											assign node1801 = (inp[10]) ? 11'b10010101011 : node1802;
												assign node1802 = (inp[11]) ? 11'b00111101001 : 11'b00110101011;
											assign node1806 = (inp[10]) ? 11'b00100111101 : node1807;
												assign node1807 = (inp[11]) ? 11'b10000111011 : 11'b10000101001;
										assign node1811 = (inp[10]) ? node1817 : node1812;
											assign node1812 = (inp[11]) ? node1814 : 11'b00011001101;
												assign node1814 = (inp[3]) ? 11'b10110101101 : 11'b00000101101;
											assign node1817 = (inp[11]) ? 11'b00011011001 : 11'b00110001001;
									assign node1820 = (inp[4]) ? node1828 : node1821;
										assign node1821 = (inp[10]) ? node1823 : 11'b10010001101;
											assign node1823 = (inp[3]) ? node1825 : 11'b10110011111;
												assign node1825 = (inp[11]) ? 11'b00010111111 : 11'b00000011101;
										assign node1828 = (inp[3]) ? node1832 : node1829;
											assign node1829 = (inp[11]) ? 11'b00111011101 : 11'b00000001111;
											assign node1832 = (inp[11]) ? node1834 : 11'b10110011001;
												assign node1834 = (inp[10]) ? 11'b00000011011 : 11'b10100011011;
								assign node1837 = (inp[4]) ? node1855 : node1838;
									assign node1838 = (inp[11]) ? node1848 : node1839;
										assign node1839 = (inp[9]) ? node1843 : node1840;
											assign node1840 = (inp[3]) ? 11'b00001011101 : 11'b10011011011;
											assign node1843 = (inp[3]) ? 11'b10110011111 : node1844;
												assign node1844 = (inp[10]) ? 11'b10100001101 : 11'b00100011001;
										assign node1848 = (inp[9]) ? 11'b00111001000 : node1849;
											assign node1849 = (inp[3]) ? 11'b10100101000 : node1850;
												assign node1850 = (inp[10]) ? 11'b10110111000 : 11'b00110111010;
									assign node1855 = (inp[11]) ? node1865 : node1856;
										assign node1856 = (inp[9]) ? node1860 : node1857;
											assign node1857 = (inp[10]) ? 11'b00110111010 : 11'b00001111110;
											assign node1860 = (inp[3]) ? node1862 : 11'b10001111000;
												assign node1862 = (inp[10]) ? 11'b00011101000 : 11'b10011101010;
										assign node1865 = (inp[3]) ? node1873 : node1866;
											assign node1866 = (inp[10]) ? node1870 : node1867;
												assign node1867 = (inp[9]) ? 11'b00011001100 : 11'b00010011110;
												assign node1870 = (inp[9]) ? 11'b10010001010 : 11'b10011001100;
											assign node1873 = (inp[9]) ? 11'b10000001010 : 11'b10000011100;
						assign node1876 = (inp[3]) ? node1954 : node1877;
							assign node1877 = (inp[5]) ? node1911 : node1878;
								assign node1878 = (inp[8]) ? node1896 : node1879;
									assign node1879 = (inp[4]) ? node1889 : node1880;
										assign node1880 = (inp[11]) ? node1886 : node1881;
											assign node1881 = (inp[10]) ? 11'b00010001111 : node1882;
												assign node1882 = (inp[9]) ? 11'b00000001111 : 11'b00001001001;
											assign node1886 = (inp[9]) ? 11'b00110011110 : 11'b00001011100;
										assign node1889 = (inp[9]) ? node1891 : 11'b00011011010;
											assign node1891 = (inp[10]) ? node1893 : 11'b00101111100;
												assign node1893 = (inp[11]) ? 11'b00111101010 : 11'b00110111010;
									assign node1896 = (inp[10]) ? node1906 : node1897;
										assign node1897 = (inp[9]) ? node1903 : node1898;
											assign node1898 = (inp[11]) ? 11'b00110111011 : node1899;
												assign node1899 = (inp[4]) ? 11'b00101001001 : 11'b00100101001;
											assign node1903 = (inp[11]) ? 11'b00001111101 : 11'b00000011111;
										assign node1906 = (inp[11]) ? node1908 : 11'b00110011001;
											assign node1908 = (inp[9]) ? 11'b00010001011 : 11'b00011001101;
								assign node1911 = (inp[9]) ? node1933 : node1912;
									assign node1912 = (inp[10]) ? node1924 : node1913;
										assign node1913 = (inp[11]) ? node1919 : node1914;
											assign node1914 = (inp[8]) ? node1916 : 11'b00110101000;
												assign node1916 = (inp[4]) ? 11'b00001101010 : 11'b00101001011;
											assign node1919 = (inp[8]) ? node1921 : 11'b00011011010;
												assign node1921 = (inp[4]) ? 11'b00010011000 : 11'b00110111000;
										assign node1924 = (inp[11]) ? node1930 : node1925;
											assign node1925 = (inp[4]) ? node1927 : 11'b00110101100;
												assign node1927 = (inp[8]) ? 11'b00110111100 : 11'b00011011110;
											assign node1930 = (inp[4]) ? 11'b00100101101 : 11'b00000011110;
									assign node1933 = (inp[10]) ? node1947 : node1934;
										assign node1934 = (inp[4]) ? node1942 : node1935;
											assign node1935 = (inp[11]) ? node1939 : node1936;
												assign node1936 = (inp[8]) ? 11'b00100001101 : 11'b00011101110;
												assign node1939 = (inp[8]) ? 11'b00011011110 : 11'b00110011100;
											assign node1942 = (inp[11]) ? 11'b00111101111 : node1943;
												assign node1943 = (inp[8]) ? 11'b00011111110 : 11'b00100011110;
										assign node1947 = (inp[8]) ? node1951 : node1948;
											assign node1948 = (inp[4]) ? 11'b00110011000 : 11'b00111101011;
											assign node1951 = (inp[4]) ? 11'b00011111010 : 11'b00010001010;
							assign node1954 = (inp[10]) ? node1988 : node1955;
								assign node1955 = (inp[8]) ? node1971 : node1956;
									assign node1956 = (inp[5]) ? node1968 : node1957;
										assign node1957 = (inp[11]) ? node1961 : node1958;
											assign node1958 = (inp[9]) ? 11'b00111101000 : 11'b00010111000;
											assign node1961 = (inp[4]) ? node1965 : node1962;
												assign node1962 = (inp[9]) ? 11'b00110011010 : 11'b00011001010;
												assign node1965 = (inp[9]) ? 11'b00101101010 : 11'b00101011000;
										assign node1968 = (inp[9]) ? 11'b00001111011 : 11'b00010111011;
									assign node1971 = (inp[4]) ? node1979 : node1972;
										assign node1972 = (inp[9]) ? node1974 : 11'b00000101001;
											assign node1974 = (inp[11]) ? 11'b00001011000 : node1975;
												assign node1975 = (inp[5]) ? 11'b00110011001 : 11'b00000011001;
										assign node1979 = (inp[9]) ? node1983 : node1980;
											assign node1980 = (inp[11]) ? 11'b00100111001 : 11'b00100111010;
											assign node1983 = (inp[5]) ? 11'b00000001000 : node1984;
												assign node1984 = (inp[11]) ? 11'b00100001011 : 11'b00101101011;
								assign node1988 = (inp[8]) ? node2008 : node1989;
									assign node1989 = (inp[5]) ? node1999 : node1990;
										assign node1990 = (inp[9]) ? node1992 : 11'b00000001001;
											assign node1992 = (inp[4]) ? node1996 : node1993;
												assign node1993 = (inp[11]) ? 11'b00011001010 : 11'b00001101010;
												assign node1996 = (inp[11]) ? 11'b00001101000 : 11'b00000101000;
										assign node1999 = (inp[11]) ? 11'b00011101011 : node2000;
											assign node2000 = (inp[4]) ? node2004 : node2001;
												assign node2001 = (inp[9]) ? 11'b00010101010 : 11'b00001101010;
												assign node2004 = (inp[9]) ? 11'b00001001010 : 11'b00111001000;
									assign node2008 = (inp[5]) ? node2018 : node2009;
										assign node2009 = (inp[4]) ? node2015 : node2010;
											assign node2010 = (inp[11]) ? 11'b00010101001 : node2011;
												assign node2011 = (inp[9]) ? 11'b00001001011 : 11'b00011001001;
											assign node2015 = (inp[11]) ? 11'b00001001011 : 11'b00110001001;
										assign node2018 = (inp[9]) ? 11'b00000001000 : node2019;
											assign node2019 = (inp[11]) ? 11'b00101001010 : node2020;
												assign node2020 = (inp[4]) ? 11'b00100101010 : 11'b00010001011;
				assign node2025 = (inp[8]) ? node2361 : node2026;
					assign node2026 = (inp[5]) ? node2182 : node2027;
						assign node2027 = (inp[2]) ? node2103 : node2028;
							assign node2028 = (inp[11]) ? node2070 : node2029;
								assign node2029 = (inp[3]) ? node2051 : node2030;
									assign node2030 = (inp[9]) ? node2038 : node2031;
										assign node2031 = (inp[10]) ? node2035 : node2032;
											assign node2032 = (inp[0]) ? 11'b00011101000 : 11'b00011101110;
											assign node2035 = (inp[0]) ? 11'b00010111100 : 11'b10010111100;
										assign node2038 = (inp[4]) ? node2046 : node2039;
											assign node2039 = (inp[10]) ? node2043 : node2040;
												assign node2040 = (inp[0]) ? 11'b00010101110 : 11'b00010101000;
												assign node2043 = (inp[0]) ? 11'b00011111010 : 11'b10011111110;
											assign node2046 = (inp[0]) ? node2048 : 11'b10111001010;
												assign node2048 = (inp[10]) ? 11'b00111011010 : 11'b00111011110;
									assign node2051 = (inp[4]) ? node2061 : node2052;
										assign node2052 = (inp[0]) ? node2058 : node2053;
											assign node2053 = (inp[10]) ? node2055 : 11'b10000101110;
												assign node2055 = (inp[9]) ? 11'b00001111100 : 11'b00000101110;
											assign node2058 = (inp[10]) ? 11'b00000101010 : 11'b00000111000;
										assign node2061 = (inp[9]) ? node2065 : node2062;
											assign node2062 = (inp[0]) ? 11'b00000111010 : 11'b10001101100;
											assign node2065 = (inp[0]) ? node2067 : 11'b00101011000;
												assign node2067 = (inp[10]) ? 11'b00001001000 : 11'b00101001000;
								assign node2070 = (inp[4]) ? node2090 : node2071;
									assign node2071 = (inp[0]) ? node2077 : node2072;
										assign node2072 = (inp[10]) ? node2074 : 11'b10010011000;
											assign node2074 = (inp[9]) ? 11'b10101011100 : 11'b00011011110;
										assign node2077 = (inp[3]) ? node2085 : node2078;
											assign node2078 = (inp[9]) ? node2082 : node2079;
												assign node2079 = (inp[10]) ? 11'b00010011100 : 11'b00010011000;
												assign node2082 = (inp[10]) ? 11'b00000001010 : 11'b00111011110;
											assign node2085 = (inp[9]) ? 11'b00101011000 : node2086;
												assign node2086 = (inp[10]) ? 11'b00101001010 : 11'b00000001010;
									assign node2090 = (inp[9]) ? node2098 : node2091;
										assign node2091 = (inp[10]) ? node2095 : node2092;
											assign node2092 = (inp[0]) ? 11'b00111110011 : 11'b10110001100;
											assign node2095 = (inp[0]) ? 11'b00011100011 : 11'b00111110011;
										assign node2098 = (inp[3]) ? node2100 : 11'b10110110001;
											assign node2100 = (inp[10]) ? 11'b00100110011 : 11'b10000110011;
							assign node2103 = (inp[11]) ? node2143 : node2104;
								assign node2104 = (inp[4]) ? node2122 : node2105;
									assign node2105 = (inp[10]) ? node2115 : node2106;
										assign node2106 = (inp[9]) ? node2112 : node2107;
											assign node2107 = (inp[0]) ? node2109 : 11'b00111000010;
												assign node2109 = (inp[3]) ? 11'b00011000010 : 11'b00011000000;
											assign node2112 = (inp[0]) ? 11'b00010000100 : 11'b00110000000;
										assign node2115 = (inp[3]) ? 11'b00101110111 : node2116;
											assign node2116 = (inp[9]) ? 11'b10100010100 : node2117;
												assign node2117 = (inp[0]) ? 11'b00001000100 : 11'b10101000010;
									assign node2122 = (inp[3]) ? node2132 : node2123;
										assign node2123 = (inp[0]) ? node2129 : node2124;
											assign node2124 = (inp[9]) ? 11'b10011100011 : node2125;
												assign node2125 = (inp[10]) ? 11'b10101110101 : 11'b00111100101;
											assign node2129 = (inp[10]) ? 11'b00101110011 : 11'b00110110111;
										assign node2132 = (inp[10]) ? node2138 : node2133;
											assign node2133 = (inp[0]) ? node2135 : 11'b10010110001;
												assign node2135 = (inp[9]) ? 11'b00110100001 : 11'b00011110001;
											assign node2138 = (inp[9]) ? 11'b00001110001 : node2139;
												assign node2139 = (inp[0]) ? 11'b00100100001 : 11'b00000100011;
								assign node2143 = (inp[4]) ? node2161 : node2144;
									assign node2144 = (inp[9]) ? node2154 : node2145;
										assign node2145 = (inp[10]) ? node2147 : 11'b10111110001;
											assign node2147 = (inp[3]) ? node2151 : node2148;
												assign node2148 = (inp[0]) ? 11'b00010110101 : 11'b10110100011;
												assign node2151 = (inp[0]) ? 11'b00100100011 : 11'b00100110101;
										assign node2154 = (inp[10]) ? node2158 : node2155;
											assign node2155 = (inp[0]) ? 11'b00100110101 : 11'b00000110011;
											assign node2158 = (inp[0]) ? 11'b00011000001 : 11'b00111010111;
									assign node2161 = (inp[10]) ? node2171 : node2162;
										assign node2162 = (inp[3]) ? node2166 : node2163;
											assign node2163 = (inp[9]) ? 11'b00110010101 : 11'b00101000101;
											assign node2166 = (inp[0]) ? node2168 : 11'b10000000111;
												assign node2168 = (inp[9]) ? 11'b00101000001 : 11'b00100010011;
										assign node2171 = (inp[3]) ? node2175 : node2172;
											assign node2172 = (inp[9]) ? 11'b10001010001 : 11'b10000010101;
											assign node2175 = (inp[9]) ? node2179 : node2176;
												assign node2176 = (inp[0]) ? 11'b00010000001 : 11'b00010010011;
												assign node2179 = (inp[0]) ? 11'b00001000001 : 11'b00001010011;
						assign node2182 = (inp[0]) ? node2274 : node2183;
							assign node2183 = (inp[9]) ? node2237 : node2184;
								assign node2184 = (inp[10]) ? node2208 : node2185;
									assign node2185 = (inp[3]) ? node2201 : node2186;
										assign node2186 = (inp[2]) ? node2194 : node2187;
											assign node2187 = (inp[4]) ? node2191 : node2188;
												assign node2188 = (inp[11]) ? 11'b00001010001 : 11'b00011110011;
												assign node2191 = (inp[11]) ? 11'b00010110101 : 11'b00001010101;
											assign node2194 = (inp[4]) ? node2198 : node2195;
												assign node2195 = (inp[11]) ? 11'b00100110001 : 11'b00110010011;
												assign node2198 = (inp[11]) ? 11'b00110010111 : 11'b00100110111;
										assign node2201 = (inp[4]) ? node2203 : 11'b10000100011;
											assign node2203 = (inp[2]) ? node2205 : 11'b10100110111;
												assign node2205 = (inp[11]) ? 11'b10010010101 : 11'b10000110101;
									assign node2208 = (inp[3]) ? node2222 : node2209;
										assign node2209 = (inp[4]) ? node2215 : node2210;
											assign node2210 = (inp[2]) ? node2212 : 11'b10100010001;
												assign node2212 = (inp[11]) ? 11'b10010110001 : 11'b10010010011;
											assign node2215 = (inp[2]) ? node2219 : node2216;
												assign node2216 = (inp[11]) ? 11'b10000100101 : 11'b10010000111;
												assign node2219 = (inp[11]) ? 11'b10111000111 : 11'b10100100111;
										assign node2222 = (inp[11]) ? node2230 : node2223;
											assign node2223 = (inp[4]) ? node2227 : node2224;
												assign node2224 = (inp[2]) ? 11'b00000010101 : 11'b00101110101;
												assign node2227 = (inp[2]) ? 11'b00111110011 : 11'b00000010001;
											assign node2230 = (inp[4]) ? node2234 : node2231;
												assign node2231 = (inp[2]) ? 11'b00111000111 : 11'b00010000101;
												assign node2234 = (inp[2]) ? 11'b00011000001 : 11'b00111100011;
								assign node2237 = (inp[4]) ? node2255 : node2238;
									assign node2238 = (inp[10]) ? node2248 : node2239;
										assign node2239 = (inp[3]) ? node2245 : node2240;
											assign node2240 = (inp[11]) ? 11'b00101100011 : node2241;
												assign node2241 = (inp[2]) ? 11'b00101110011 : 11'b00000110011;
											assign node2245 = (inp[2]) ? 11'b10111110101 : 11'b10001110101;
										assign node2248 = (inp[3]) ? node2250 : 11'b10100100101;
											assign node2250 = (inp[2]) ? 11'b00100000111 : node2251;
												assign node2251 = (inp[11]) ? 11'b00001100101 : 11'b00011000111;
									assign node2255 = (inp[10]) ? node2265 : node2256;
										assign node2256 = (inp[3]) ? node2260 : node2257;
											assign node2257 = (inp[11]) ? 11'b00101000111 : 11'b00011110101;
											assign node2260 = (inp[11]) ? node2262 : 11'b10000000001;
												assign node2262 = (inp[2]) ? 11'b10001000001 : 11'b10111100001;
										assign node2265 = (inp[3]) ? node2269 : node2266;
											assign node2266 = (inp[11]) ? 11'b10010100011 : 11'b10101110001;
											assign node2269 = (inp[2]) ? 11'b00000100011 : node2270;
												assign node2270 = (inp[11]) ? 11'b00100100001 : 11'b00101000011;
							assign node2274 = (inp[3]) ? node2316 : node2275;
								assign node2275 = (inp[4]) ? node2293 : node2276;
									assign node2276 = (inp[10]) ? node2284 : node2277;
										assign node2277 = (inp[9]) ? 11'b00001100111 : node2278;
											assign node2278 = (inp[11]) ? node2280 : 11'b00010000011;
												assign node2280 = (inp[2]) ? 11'b00000110001 : 11'b00010010011;
										assign node2284 = (inp[11]) ? node2290 : node2285;
											assign node2285 = (inp[9]) ? node2287 : 11'b00111100101;
												assign node2287 = (inp[2]) ? 11'b00111110001 : 11'b00111010011;
											assign node2290 = (inp[9]) ? 11'b00100000011 : 11'b00011010111;
									assign node2293 = (inp[11]) ? node2307 : node2294;
										assign node2294 = (inp[2]) ? node2302 : node2295;
											assign node2295 = (inp[9]) ? node2299 : node2296;
												assign node2296 = (inp[10]) ? 11'b00000010111 : 11'b00101000011;
												assign node2299 = (inp[10]) ? 11'b00111010001 : 11'b00100010101;
											assign node2302 = (inp[9]) ? 11'b00101110001 : node2303;
												assign node2303 = (inp[10]) ? 11'b00000110101 : 11'b00100100001;
										assign node2307 = (inp[9]) ? node2311 : node2308;
											assign node2308 = (inp[10]) ? 11'b00111100111 : 11'b00110110001;
											assign node2311 = (inp[10]) ? 11'b00100100011 : node2312;
												assign node2312 = (inp[2]) ? 11'b00101000111 : 11'b00101100111;
								assign node2316 = (inp[10]) ? node2342 : node2317;
									assign node2317 = (inp[9]) ? node2329 : node2318;
										assign node2318 = (inp[4]) ? node2324 : node2319;
											assign node2319 = (inp[2]) ? node2321 : 11'b00101100001;
												assign node2321 = (inp[11]) ? 11'b00110100001 : 11'b00110000001;
											assign node2324 = (inp[11]) ? node2326 : 11'b00111010001;
												assign node2326 = (inp[2]) ? 11'b00010010001 : 11'b00000110011;
										assign node2329 = (inp[4]) ? node2337 : node2330;
											assign node2330 = (inp[11]) ? node2334 : node2331;
												assign node2331 = (inp[2]) ? 11'b00111110011 : 11'b00100110011;
												assign node2334 = (inp[2]) ? 11'b00001010001 : 11'b00011110011;
											assign node2337 = (inp[11]) ? 11'b00001000001 : node2338;
												assign node2338 = (inp[2]) ? 11'b00011100011 : 11'b00001000011;
									assign node2342 = (inp[4]) ? node2354 : node2343;
										assign node2343 = (inp[11]) ? node2351 : node2344;
											assign node2344 = (inp[9]) ? node2348 : node2345;
												assign node2345 = (inp[2]) ? 11'b00000000001 : 11'b00000100011;
												assign node2348 = (inp[2]) ? 11'b00010100011 : 11'b00011000001;
											assign node2351 = (inp[9]) ? 11'b00000000001 : 11'b00110000001;
										assign node2354 = (inp[9]) ? 11'b00000100011 : node2355;
											assign node2355 = (inp[11]) ? 11'b00011100001 : node2356;
												assign node2356 = (inp[2]) ? 11'b00111100011 : 11'b00110000011;
					assign node2361 = (inp[0]) ? node2513 : node2362;
						assign node2362 = (inp[9]) ? node2448 : node2363;
							assign node2363 = (inp[11]) ? node2411 : node2364;
								assign node2364 = (inp[5]) ? node2384 : node2365;
									assign node2365 = (inp[4]) ? node2375 : node2366;
										assign node2366 = (inp[10]) ? node2372 : node2367;
											assign node2367 = (inp[3]) ? 11'b10100100001 : node2368;
												assign node2368 = (inp[2]) ? 11'b00110000011 : 11'b00010100011;
											assign node2372 = (inp[3]) ? 11'b00111000111 : 11'b10001000011;
										assign node2375 = (inp[2]) ? node2381 : node2376;
											assign node2376 = (inp[3]) ? node2378 : 11'b10101010111;
												assign node2378 = (inp[10]) ? 11'b00011000001 : 11'b10011000101;
											assign node2381 = (inp[3]) ? 11'b00111100010 : 11'b10011110100;
									assign node2384 = (inp[2]) ? node2400 : node2385;
										assign node2385 = (inp[4]) ? node2393 : node2386;
											assign node2386 = (inp[3]) ? node2390 : node2387;
												assign node2387 = (inp[10]) ? 11'b10100010010 : 11'b00010010010;
												assign node2390 = (inp[10]) ? 11'b00110010100 : 11'b10010010000;
											assign node2393 = (inp[3]) ? node2397 : node2394;
												assign node2394 = (inp[10]) ? 11'b10010000100 : 11'b00100010100;
												assign node2397 = (inp[10]) ? 11'b00011110010 : 11'b10000010110;
										assign node2400 = (inp[4]) ? node2408 : node2401;
											assign node2401 = (inp[10]) ? node2405 : node2402;
												assign node2402 = (inp[3]) ? 11'b10111110000 : 11'b00111110010;
												assign node2405 = (inp[3]) ? 11'b00011110100 : 11'b10011110010;
											assign node2408 = (inp[10]) ? 11'b00101110000 : 11'b10101110100;
								assign node2411 = (inp[2]) ? node2431 : node2412;
									assign node2412 = (inp[4]) ? node2422 : node2413;
										assign node2413 = (inp[5]) ? node2419 : node2414;
											assign node2414 = (inp[3]) ? 11'b10111110010 : node2415;
												assign node2415 = (inp[10]) ? 11'b10101100000 : 11'b00001100000;
											assign node2419 = (inp[10]) ? 11'b00001100100 : 11'b10010100000;
										assign node2422 = (inp[5]) ? node2428 : node2423;
											assign node2423 = (inp[10]) ? node2425 : 11'b10001100100;
												assign node2425 = (inp[3]) ? 11'b00100110010 : 11'b10110110100;
											assign node2428 = (inp[10]) ? 11'b10101000100 : 11'b10111010110;
									assign node2431 = (inp[4]) ? node2437 : node2432;
										assign node2432 = (inp[3]) ? 11'b00101000100 : node2433;
											assign node2433 = (inp[5]) ? 11'b10101010010 : 11'b10001000000;
										assign node2437 = (inp[3]) ? node2443 : node2438;
											assign node2438 = (inp[5]) ? 11'b00001010110 : node2439;
												assign node2439 = (inp[10]) ? 11'b10001010100 : 11'b00010000100;
											assign node2443 = (inp[10]) ? 11'b00001010010 : node2444;
												assign node2444 = (inp[5]) ? 11'b10001010100 : 11'b10101000110;
							assign node2448 = (inp[2]) ? node2482 : node2449;
								assign node2449 = (inp[4]) ? node2463 : node2450;
									assign node2450 = (inp[11]) ? node2460 : node2451;
										assign node2451 = (inp[3]) ? node2455 : node2452;
											assign node2452 = (inp[10]) ? 11'b10001000110 : 11'b00001000001;
											assign node2455 = (inp[5]) ? 11'b00110000110 : node2456;
												assign node2456 = (inp[10]) ? 11'b00100010111 : 11'b10110000111;
										assign node2460 = (inp[3]) ? 11'b10100100100 : 11'b00110110010;
									assign node2463 = (inp[5]) ? node2473 : node2464;
										assign node2464 = (inp[11]) ? node2468 : node2465;
											assign node2465 = (inp[10]) ? 11'b10010000001 : 11'b10000010001;
											assign node2468 = (inp[10]) ? node2470 : 11'b00000110100;
												assign node2470 = (inp[3]) ? 11'b00101010010 : 11'b10101010000;
										assign node2473 = (inp[11]) ? node2479 : node2474;
											assign node2474 = (inp[3]) ? node2476 : 11'b00101110100;
												assign node2476 = (inp[10]) ? 11'b00100100000 : 11'b10111100000;
											assign node2479 = (inp[3]) ? 11'b10110000000 : 11'b10100000010;
								assign node2482 = (inp[11]) ? node2502 : node2483;
									assign node2483 = (inp[10]) ? node2495 : node2484;
										assign node2484 = (inp[5]) ? node2490 : node2485;
											assign node2485 = (inp[3]) ? node2487 : 11'b00011100100;
												assign node2487 = (inp[4]) ? 11'b10100110010 : 11'b10001100100;
											assign node2490 = (inp[4]) ? 11'b00000110110 : node2491;
												assign node2491 = (inp[3]) ? 11'b10110110100 : 11'b00110110010;
										assign node2495 = (inp[3]) ? node2499 : node2496;
											assign node2496 = (inp[5]) ? 11'b10000110010 : 11'b10100100000;
											assign node2499 = (inp[5]) ? 11'b00000100000 : 11'b00000110100;
									assign node2502 = (inp[5]) ? node2506 : node2503;
										assign node2503 = (inp[4]) ? 11'b00000010010 : 11'b10010000110;
										assign node2506 = (inp[3]) ? node2508 : 11'b00000000110;
											assign node2508 = (inp[4]) ? node2510 : 11'b00000000100;
												assign node2510 = (inp[10]) ? 11'b00000000000 : 11'b10000000000;
						assign node2513 = (inp[3]) ? node2591 : node2514;
							assign node2514 = (inp[9]) ? node2552 : node2515;
								assign node2515 = (inp[10]) ? node2533 : node2516;
									assign node2516 = (inp[11]) ? node2526 : node2517;
										assign node2517 = (inp[5]) ? node2521 : node2518;
											assign node2518 = (inp[4]) ? 11'b00111000011 : 11'b00110100001;
											assign node2521 = (inp[4]) ? 11'b00000000000 : node2522;
												assign node2522 = (inp[2]) ? 11'b00111100010 : 11'b00110000010;
										assign node2526 = (inp[2]) ? 11'b00101010010 : node2527;
											assign node2527 = (inp[4]) ? 11'b00101110000 : node2528;
												assign node2528 = (inp[5]) ? 11'b00110110000 : 11'b00111110010;
									assign node2533 = (inp[5]) ? node2541 : node2534;
										assign node2534 = (inp[11]) ? node2538 : node2535;
											assign node2535 = (inp[2]) ? 11'b00111100100 : 11'b00111000101;
											assign node2538 = (inp[4]) ? 11'b00001000110 : 11'b00111010110;
										assign node2541 = (inp[11]) ? node2547 : node2542;
											assign node2542 = (inp[4]) ? 11'b00101110110 : node2543;
												assign node2543 = (inp[2]) ? 11'b00011100110 : 11'b00000000110;
											assign node2547 = (inp[4]) ? 11'b00001000110 : node2548;
												assign node2548 = (inp[2]) ? 11'b00101010110 : 11'b00101110100;
								assign node2552 = (inp[10]) ? node2574 : node2553;
									assign node2553 = (inp[11]) ? node2565 : node2554;
										assign node2554 = (inp[4]) ? node2562 : node2555;
											assign node2555 = (inp[2]) ? node2559 : node2556;
												assign node2556 = (inp[5]) ? 11'b00101000100 : 11'b00101000101;
												assign node2559 = (inp[5]) ? 11'b00110100110 : 11'b00101100100;
											assign node2562 = (inp[5]) ? 11'b00001110110 : 11'b00000010101;
										assign node2565 = (inp[4]) ? node2571 : node2566;
											assign node2566 = (inp[5]) ? 11'b00011110100 : node2567;
												assign node2567 = (inp[2]) ? 11'b00010010110 : 11'b00010110110;
											assign node2571 = (inp[5]) ? 11'b00000000110 : 11'b00111000110;
									assign node2574 = (inp[11]) ? node2582 : node2575;
										assign node2575 = (inp[2]) ? 11'b00000110000 : node2576;
											assign node2576 = (inp[5]) ? 11'b00011010000 : node2577;
												assign node2577 = (inp[4]) ? 11'b00010010001 : 11'b00100010011;
										assign node2582 = (inp[2]) ? node2586 : node2583;
											assign node2583 = (inp[4]) ? 11'b00000000010 : 11'b00000100000;
											assign node2586 = (inp[5]) ? 11'b00000000010 : node2587;
												assign node2587 = (inp[4]) ? 11'b00000000010 : 11'b00110000010;
							assign node2591 = (inp[9]) ? node2631 : node2592;
								assign node2592 = (inp[11]) ? node2614 : node2593;
									assign node2593 = (inp[2]) ? node2605 : node2594;
										assign node2594 = (inp[10]) ? node2600 : node2595;
											assign node2595 = (inp[5]) ? node2597 : 11'b00001010001;
												assign node2597 = (inp[4]) ? 11'b00110010000 : 11'b00100000000;
											assign node2600 = (inp[5]) ? node2602 : 11'b00110000011;
												assign node2602 = (inp[4]) ? 11'b00101100000 : 11'b00011000010;
										assign node2605 = (inp[5]) ? node2611 : node2606;
											assign node2606 = (inp[10]) ? 11'b00111100010 : node2607;
												assign node2607 = (inp[4]) ? 11'b00011110010 : 11'b00011100010;
											assign node2611 = (inp[4]) ? 11'b00101100000 : 11'b00111100000;
									assign node2614 = (inp[2]) ? node2620 : node2615;
										assign node2615 = (inp[5]) ? 11'b00001000000 : node2616;
											assign node2616 = (inp[4]) ? 11'b00000100010 : 11'b00110100000;
										assign node2620 = (inp[4]) ? node2626 : node2621;
											assign node2621 = (inp[10]) ? node2623 : 11'b00001000010;
												assign node2623 = (inp[5]) ? 11'b00101000000 : 11'b00111000000;
											assign node2626 = (inp[10]) ? 11'b00001000000 : node2627;
												assign node2627 = (inp[5]) ? 11'b00001010000 : 11'b00101010000;
								assign node2631 = (inp[10]) ? node2653 : node2632;
									assign node2632 = (inp[4]) ? node2642 : node2633;
										assign node2633 = (inp[11]) ? node2635 : 11'b00010010001;
											assign node2635 = (inp[2]) ? node2639 : node2636;
												assign node2636 = (inp[5]) ? 11'b00010110010 : 11'b00100110000;
												assign node2639 = (inp[5]) ? 11'b00000010000 : 11'b00110010000;
										assign node2642 = (inp[5]) ? node2648 : node2643;
											assign node2643 = (inp[11]) ? node2645 : 11'b00110000011;
												assign node2645 = (inp[2]) ? 11'b00100000000 : 11'b00111000000;
											assign node2648 = (inp[11]) ? node2650 : 11'b00011100000;
												assign node2650 = (inp[2]) ? 11'b00000000000 : 11'b00010000000;
									assign node2653 = (inp[4]) ? node2669 : node2654;
										assign node2654 = (inp[2]) ? node2662 : node2655;
											assign node2655 = (inp[11]) ? node2659 : node2656;
												assign node2656 = (inp[5]) ? 11'b00010000010 : 11'b00000000001;
												assign node2659 = (inp[5]) ? 11'b00000100010 : 11'b00011100010;
											assign node2662 = (inp[11]) ? node2666 : node2663;
												assign node2663 = (inp[5]) ? 11'b00010100000 : 11'b00000100010;
												assign node2666 = (inp[5]) ? 11'b00000000000 : 11'b00010000000;
										assign node2669 = (inp[11]) ? 11'b00000000000 : node2670;
											assign node2670 = (inp[5]) ? 11'b00000100000 : node2671;
												assign node2671 = (inp[2]) ? 11'b00000100010 : 11'b00001100010;
		assign node2676 = (inp[7]) ? node4012 : node2677;
			assign node2677 = (inp[6]) ? node3347 : node2678;
				assign node2678 = (inp[8]) ? node2992 : node2679;
					assign node2679 = (inp[0]) ? node2845 : node2680;
						assign node2680 = (inp[9]) ? node2766 : node2681;
							assign node2681 = (inp[4]) ? node2721 : node2682;
								assign node2682 = (inp[10]) ? node2706 : node2683;
									assign node2683 = (inp[3]) ? node2697 : node2684;
										assign node2684 = (inp[5]) ? node2690 : node2685;
											assign node2685 = (inp[2]) ? 11'b00100101011 : node2686;
												assign node2686 = (inp[11]) ? 11'b00001001011 : 11'b00001101011;
											assign node2690 = (inp[2]) ? node2694 : node2691;
												assign node2691 = (inp[11]) ? 11'b00000111001 : 11'b00000011001;
												assign node2694 = (inp[11]) ? 11'b00101111001 : 11'b00101011001;
										assign node2697 = (inp[5]) ? node2701 : node2698;
											assign node2698 = (inp[11]) ? 11'b10110111001 : 11'b10101001000;
											assign node2701 = (inp[11]) ? node2703 : 11'b10100011011;
												assign node2703 = (inp[2]) ? 11'b10011101011 : 11'b10101001011;
									assign node2706 = (inp[3]) ? node2714 : node2707;
										assign node2707 = (inp[5]) ? node2711 : node2708;
											assign node2708 = (inp[11]) ? 11'b10001001011 : 11'b10001101011;
											assign node2711 = (inp[2]) ? 11'b10001111011 : 11'b10101011001;
										assign node2714 = (inp[2]) ? 11'b00101111111 : node2715;
											assign node2715 = (inp[11]) ? 11'b00011001111 : node2716;
												assign node2716 = (inp[5]) ? 11'b00101111111 : 11'b00001101101;
								assign node2721 = (inp[3]) ? node2745 : node2722;
									assign node2722 = (inp[10]) ? node2732 : node2723;
										assign node2723 = (inp[2]) ? node2727 : node2724;
											assign node2724 = (inp[5]) ? 11'b00000011111 : 11'b00001101111;
											assign node2727 = (inp[5]) ? 11'b00111011111 : node2728;
												assign node2728 = (inp[11]) ? 11'b00110101101 : 11'b00100001100;
										assign node2732 = (inp[5]) ? node2740 : node2733;
											assign node2733 = (inp[11]) ? node2737 : node2734;
												assign node2734 = (inp[2]) ? 11'b10111111101 : 11'b10001111111;
												assign node2737 = (inp[2]) ? 11'b10000111111 : 11'b10111011111;
											assign node2740 = (inp[2]) ? 11'b10100001111 : node2741;
												assign node2741 = (inp[11]) ? 11'b10001001111 : 11'b10011101101;
									assign node2745 = (inp[10]) ? node2757 : node2746;
										assign node2746 = (inp[5]) ? node2752 : node2747;
											assign node2747 = (inp[11]) ? 11'b10111001101 : node2748;
												assign node2748 = (inp[2]) ? 11'b10101101111 : 11'b10001101101;
											assign node2752 = (inp[2]) ? node2754 : 11'b10111111111;
												assign node2754 = (inp[11]) ? 11'b10011111111 : 11'b10001011101;
										assign node2757 = (inp[2]) ? node2761 : node2758;
											assign node2758 = (inp[5]) ? 11'b00101001001 : 11'b00101101001;
											assign node2761 = (inp[5]) ? 11'b00001101011 : node2762;
												assign node2762 = (inp[11]) ? 11'b00010111001 : 11'b00001101001;
							assign node2766 = (inp[11]) ? node2808 : node2767;
								assign node2767 = (inp[2]) ? node2785 : node2768;
									assign node2768 = (inp[4]) ? node2776 : node2769;
										assign node2769 = (inp[3]) ? node2773 : node2770;
											assign node2770 = (inp[5]) ? 11'b00001111001 : 11'b00000101011;
											assign node2773 = (inp[10]) ? 11'b00010101111 : 11'b10000111111;
										assign node2776 = (inp[10]) ? node2782 : node2777;
											assign node2777 = (inp[3]) ? node2779 : 11'b00111111101;
												assign node2779 = (inp[5]) ? 11'b10000101011 : 11'b10100111001;
											assign node2782 = (inp[5]) ? 11'b00100101011 : 11'b10100101011;
									assign node2785 = (inp[4]) ? node2797 : node2786;
										assign node2786 = (inp[5]) ? node2790 : node2787;
											assign node2787 = (inp[10]) ? 11'b10110011100 : 11'b10100001110;
											assign node2790 = (inp[10]) ? node2794 : node2791;
												assign node2791 = (inp[3]) ? 11'b10111011111 : 11'b00100011001;
												assign node2794 = (inp[3]) ? 11'b00101001101 : 11'b10001001111;
										assign node2797 = (inp[3]) ? node2803 : node2798;
											assign node2798 = (inp[5]) ? node2800 : 11'b10010101011;
												assign node2800 = (inp[10]) ? 11'b10110011001 : 11'b00000011101;
											assign node2803 = (inp[10]) ? node2805 : 11'b10100001011;
												assign node2805 = (inp[5]) ? 11'b00001101011 : 11'b00000111001;
								assign node2808 = (inp[2]) ? node2828 : node2809;
									assign node2809 = (inp[5]) ? node2817 : node2810;
										assign node2810 = (inp[4]) ? node2814 : node2811;
											assign node2811 = (inp[10]) ? 11'b10100011111 : 11'b10100001101;
											assign node2814 = (inp[10]) ? 11'b00110011001 : 11'b10010011001;
										assign node2817 = (inp[10]) ? node2823 : node2818;
											assign node2818 = (inp[3]) ? 11'b10111001001 : node2819;
												assign node2819 = (inp[4]) ? 11'b00011001111 : 11'b00111001001;
											assign node2823 = (inp[4]) ? 11'b10010001011 : node2824;
												assign node2824 = (inp[3]) ? 11'b00000001101 : 11'b10110001101;
									assign node2828 = (inp[5]) ? node2836 : node2829;
										assign node2829 = (inp[4]) ? node2831 : 11'b10011101111;
											assign node2831 = (inp[10]) ? node2833 : 11'b00111011111;
												assign node2833 = (inp[3]) ? 11'b00011011001 : 11'b10011011011;
										assign node2836 = (inp[4]) ? node2840 : node2837;
											assign node2837 = (inp[10]) ? 11'b10010101111 : 11'b00010101011;
											assign node2840 = (inp[3]) ? node2842 : 11'b00111101101;
												assign node2842 = (inp[10]) ? 11'b00010101001 : 11'b10001101001;
						assign node2845 = (inp[9]) ? node2917 : node2846;
							assign node2846 = (inp[3]) ? node2880 : node2847;
								assign node2847 = (inp[10]) ? node2865 : node2848;
									assign node2848 = (inp[11]) ? node2858 : node2849;
										assign node2849 = (inp[2]) ? node2851 : 11'b00001101011;
											assign node2851 = (inp[5]) ? node2855 : node2852;
												assign node2852 = (inp[4]) ? 11'b00000001000 : 11'b00001001010;
												assign node2855 = (inp[4]) ? 11'b00111001001 : 11'b00000001011;
										assign node2858 = (inp[4]) ? 11'b00101111011 : node2859;
											assign node2859 = (inp[5]) ? 11'b00000111001 : node2860;
												assign node2860 = (inp[2]) ? 11'b00010111011 : 11'b00001011011;
									assign node2865 = (inp[11]) ? node2875 : node2866;
										assign node2866 = (inp[2]) ? node2872 : node2867;
											assign node2867 = (inp[4]) ? node2869 : 11'b00101101111;
												assign node2869 = (inp[5]) ? 11'b00011111111 : 11'b00001111111;
											assign node2872 = (inp[5]) ? 11'b00110001111 : 11'b00011001110;
										assign node2875 = (inp[5]) ? node2877 : 11'b00001011111;
											assign node2877 = (inp[2]) ? 11'b00001111101 : 11'b00011011101;
								assign node2880 = (inp[4]) ? node2902 : node2881;
									assign node2881 = (inp[2]) ? node2891 : node2882;
										assign node2882 = (inp[11]) ? node2886 : node2883;
											assign node2883 = (inp[10]) ? 11'b00001101001 : 11'b00101101001;
											assign node2886 = (inp[5]) ? node2888 : 11'b00101001001;
												assign node2888 = (inp[10]) ? 11'b00111001011 : 11'b00101001011;
										assign node2891 = (inp[5]) ? node2899 : node2892;
											assign node2892 = (inp[11]) ? node2896 : node2893;
												assign node2893 = (inp[10]) ? 11'b00001001000 : 11'b00011001000;
												assign node2896 = (inp[10]) ? 11'b00101101001 : 11'b00010101001;
											assign node2899 = (inp[10]) ? 11'b00000001011 : 11'b00110001001;
									assign node2902 = (inp[10]) ? node2912 : node2903;
										assign node2903 = (inp[2]) ? node2909 : node2904;
											assign node2904 = (inp[11]) ? node2906 : 11'b00111111001;
												assign node2906 = (inp[5]) ? 11'b00001011011 : 11'b00111011001;
											assign node2909 = (inp[11]) ? 11'b00011111001 : 11'b00011111011;
										assign node2912 = (inp[11]) ? node2914 : 11'b00101101001;
											assign node2914 = (inp[2]) ? 11'b00011001011 : 11'b00011001001;
							assign node2917 = (inp[3]) ? node2959 : node2918;
								assign node2918 = (inp[10]) ? node2936 : node2919;
									assign node2919 = (inp[11]) ? node2929 : node2920;
										assign node2920 = (inp[4]) ? node2922 : 11'b00000101111;
											assign node2922 = (inp[5]) ? node2926 : node2923;
												assign node2923 = (inp[2]) ? 11'b00101111101 : 11'b00100111111;
												assign node2926 = (inp[2]) ? 11'b00100011111 : 11'b00110111111;
										assign node2929 = (inp[5]) ? node2933 : node2930;
											assign node2930 = (inp[4]) ? 11'b00010001111 : 11'b00100011111;
											assign node2933 = (inp[2]) ? 11'b00110111101 : 11'b00111001101;
									assign node2936 = (inp[11]) ? node2948 : node2937;
										assign node2937 = (inp[2]) ? node2943 : node2938;
											assign node2938 = (inp[4]) ? 11'b00100111001 : node2939;
												assign node2939 = (inp[5]) ? 11'b00100111011 : 11'b00000111011;
											assign node2943 = (inp[4]) ? node2945 : 11'b00101011001;
												assign node2945 = (inp[5]) ? 11'b00111111011 : 11'b00110111001;
										assign node2948 = (inp[5]) ? node2954 : node2949;
											assign node2949 = (inp[2]) ? node2951 : 11'b00010001011;
												assign node2951 = (inp[4]) ? 11'b00111001011 : 11'b00001101001;
											assign node2954 = (inp[2]) ? node2956 : 11'b00110001001;
												assign node2956 = (inp[4]) ? 11'b00110101001 : 11'b00110101011;
								assign node2959 = (inp[4]) ? node2975 : node2960;
									assign node2960 = (inp[10]) ? node2970 : node2961;
										assign node2961 = (inp[5]) ? node2965 : node2962;
											assign node2962 = (inp[2]) ? 11'b00010011000 : 11'b00000111001;
											assign node2965 = (inp[11]) ? node2967 : 11'b00111011011;
												assign node2967 = (inp[2]) ? 11'b00000111001 : 11'b00010011011;
										assign node2970 = (inp[11]) ? 11'b00000001011 : node2971;
											assign node2971 = (inp[5]) ? 11'b00010101001 : 11'b00000101001;
									assign node2975 = (inp[5]) ? node2983 : node2976;
										assign node2976 = (inp[11]) ? node2980 : node2977;
											assign node2977 = (inp[2]) ? 11'b00110101011 : 11'b00100101001;
											assign node2980 = (inp[10]) ? 11'b00000001001 : 11'b00101001001;
										assign node2983 = (inp[10]) ? node2989 : node2984;
											assign node2984 = (inp[2]) ? node2986 : 11'b00000101011;
												assign node2986 = (inp[11]) ? 11'b00000101011 : 11'b00010001001;
											assign node2989 = (inp[11]) ? 11'b00000101001 : 11'b00001101011;
					assign node2992 = (inp[0]) ? node3174 : node2993;
						assign node2993 = (inp[11]) ? node3083 : node2994;
							assign node2994 = (inp[2]) ? node3036 : node2995;
								assign node2995 = (inp[10]) ? node3013 : node2996;
									assign node2996 = (inp[3]) ? node3002 : node2997;
										assign node2997 = (inp[4]) ? 11'b00111111100 : node2998;
											assign node2998 = (inp[9]) ? 11'b00011101010 : 11'b00000001011;
										assign node3002 = (inp[4]) ? node3006 : node3003;
											assign node3003 = (inp[9]) ? 11'b10001111110 : 11'b10000011010;
											assign node3006 = (inp[9]) ? node3010 : node3007;
												assign node3007 = (inp[5]) ? 11'b10010111110 : 11'b10000101110;
												assign node3010 = (inp[5]) ? 11'b10110101000 : 11'b10011111010;
									assign node3013 = (inp[3]) ? node3025 : node3014;
										assign node3014 = (inp[5]) ? node3022 : node3015;
											assign node3015 = (inp[4]) ? node3019 : node3016;
												assign node3016 = (inp[9]) ? 11'b10010111110 : 11'b10001101010;
												assign node3019 = (inp[9]) ? 11'b10001101000 : 11'b10100111100;
											assign node3022 = (inp[9]) ? 11'b10001101100 : 11'b10000101110;
										assign node3025 = (inp[4]) ? node3033 : node3026;
											assign node3026 = (inp[5]) ? node3030 : node3027;
												assign node3027 = (inp[9]) ? 11'b00110111100 : 11'b00101101100;
												assign node3030 = (inp[9]) ? 11'b00101101110 : 11'b00110011110;
											assign node3033 = (inp[9]) ? 11'b00101101000 : 11'b00011101010;
								assign node3036 = (inp[5]) ? node3060 : node3037;
									assign node3037 = (inp[9]) ? node3049 : node3038;
										assign node3038 = (inp[3]) ? node3042 : node3039;
											assign node3039 = (inp[4]) ? 11'b00000001111 : 11'b00100101011;
											assign node3042 = (inp[10]) ? node3046 : node3043;
												assign node3043 = (inp[4]) ? 11'b10110001101 : 11'b10010101001;
												assign node3046 = (inp[4]) ? 11'b00100001001 : 11'b00001001111;
										assign node3049 = (inp[3]) ? node3057 : node3050;
											assign node3050 = (inp[10]) ? node3054 : node3051;
												assign node3051 = (inp[4]) ? 11'b00011001111 : 11'b00111001001;
												assign node3054 = (inp[4]) ? 11'b10111001001 : 11'b10101011101;
											assign node3057 = (inp[10]) ? 11'b00010011111 : 11'b10101011011;
									assign node3060 = (inp[3]) ? node3072 : node3061;
										assign node3061 = (inp[10]) ? node3065 : node3062;
											assign node3062 = (inp[4]) ? 11'b00010111110 : 11'b00111111000;
											assign node3065 = (inp[9]) ? node3069 : node3066;
												assign node3066 = (inp[4]) ? 11'b10110101100 : 11'b10001111000;
												assign node3069 = (inp[4]) ? 11'b10011011010 : 11'b10110101110;
										assign node3072 = (inp[9]) ? node3078 : node3073;
											assign node3073 = (inp[10]) ? node3075 : 11'b10100111110;
												assign node3075 = (inp[4]) ? 11'b00101011010 : 11'b00011111110;
											assign node3078 = (inp[4]) ? node3080 : 11'b00000101100;
												assign node3080 = (inp[10]) ? 11'b00001001000 : 11'b10001001000;
							assign node3083 = (inp[5]) ? node3129 : node3084;
								assign node3084 = (inp[2]) ? node3108 : node3085;
									assign node3085 = (inp[9]) ? node3099 : node3086;
										assign node3086 = (inp[4]) ? node3092 : node3087;
											assign node3087 = (inp[3]) ? 11'b10100111010 : node3088;
												assign node3088 = (inp[10]) ? 11'b10110101000 : 11'b00000101000;
											assign node3092 = (inp[10]) ? node3096 : node3093;
												assign node3093 = (inp[3]) ? 11'b10010001100 : 11'b00110001110;
												assign node3096 = (inp[3]) ? 11'b00100011000 : 11'b10110011110;
										assign node3099 = (inp[3]) ? node3103 : node3100;
											assign node3100 = (inp[4]) ? 11'b00001011110 : 11'b00111011000;
											assign node3103 = (inp[4]) ? node3105 : 11'b10101001100;
												assign node3105 = (inp[10]) ? 11'b00111011000 : 11'b10011011000;
									assign node3108 = (inp[4]) ? node3118 : node3109;
										assign node3109 = (inp[9]) ? node3115 : node3110;
											assign node3110 = (inp[3]) ? 11'b10010011011 : node3111;
												assign node3111 = (inp[10]) ? 11'b10000001011 : 11'b00101001001;
											assign node3115 = (inp[10]) ? 11'b00001111110 : 11'b00000011011;
										assign node3118 = (inp[9]) ? node3122 : node3119;
											assign node3119 = (inp[10]) ? 11'b10011111100 : 11'b00011101100;
											assign node3122 = (inp[3]) ? node3126 : node3123;
												assign node3123 = (inp[10]) ? 11'b10000111010 : 11'b00100111110;
												assign node3126 = (inp[10]) ? 11'b00010111000 : 11'b10110111000;
								assign node3129 = (inp[3]) ? node3155 : node3130;
									assign node3130 = (inp[10]) ? node3142 : node3131;
										assign node3131 = (inp[9]) ? node3137 : node3132;
											assign node3132 = (inp[4]) ? 11'b00101011100 : node3133;
												assign node3133 = (inp[2]) ? 11'b00100011010 : 11'b00001111010;
											assign node3137 = (inp[4]) ? node3139 : 11'b00100001000;
												assign node3139 = (inp[2]) ? 11'b00000001100 : 11'b00100001110;
										assign node3142 = (inp[2]) ? node3148 : node3143;
											assign node3143 = (inp[9]) ? node3145 : 11'b10010111010;
												assign node3145 = (inp[4]) ? 11'b10110001010 : 11'b10110101100;
											assign node3148 = (inp[9]) ? node3152 : node3149;
												assign node3149 = (inp[4]) ? 11'b10001001100 : 11'b10100011000;
												assign node3152 = (inp[4]) ? 11'b10000001010 : 11'b10001001110;
									assign node3155 = (inp[4]) ? node3161 : node3156;
										assign node3156 = (inp[9]) ? node3158 : 11'b00110001110;
											assign node3158 = (inp[2]) ? 11'b00011001100 : 11'b00111001110;
										assign node3161 = (inp[10]) ? node3167 : node3162;
											assign node3162 = (inp[9]) ? node3164 : 11'b10011011100;
												assign node3164 = (inp[2]) ? 11'b10010001010 : 11'b10100001000;
											assign node3167 = (inp[9]) ? node3171 : node3168;
												assign node3168 = (inp[2]) ? 11'b00010001010 : 11'b00110001010;
												assign node3171 = (inp[2]) ? 11'b00010001000 : 11'b00110001000;
						assign node3174 = (inp[3]) ? node3260 : node3175;
							assign node3175 = (inp[9]) ? node3221 : node3176;
								assign node3176 = (inp[10]) ? node3202 : node3177;
									assign node3177 = (inp[11]) ? node3191 : node3178;
										assign node3178 = (inp[5]) ? node3186 : node3179;
											assign node3179 = (inp[4]) ? node3183 : node3180;
												assign node3180 = (inp[2]) ? 11'b00100101011 : 11'b00100001011;
												assign node3183 = (inp[2]) ? 11'b00100001001 : 11'b00100101010;
											assign node3186 = (inp[2]) ? node3188 : 11'b00011101000;
												assign node3188 = (inp[4]) ? 11'b00000101010 : 11'b00101101010;
										assign node3191 = (inp[2]) ? node3197 : node3192;
											assign node3192 = (inp[5]) ? 11'b00101111010 : node3193;
												assign node3193 = (inp[4]) ? 11'b00110011000 : 11'b00100111000;
											assign node3197 = (inp[4]) ? 11'b00111111010 : node3198;
												assign node3198 = (inp[5]) ? 11'b00110011010 : 11'b00111011001;
									assign node3202 = (inp[2]) ? node3210 : node3203;
										assign node3203 = (inp[4]) ? node3207 : node3204;
											assign node3204 = (inp[5]) ? 11'b00110111110 : 11'b00110111100;
											assign node3207 = (inp[5]) ? 11'b00100111100 : 11'b00101111110;
										assign node3210 = (inp[11]) ? node3216 : node3211;
											assign node3211 = (inp[5]) ? 11'b00111011110 : node3212;
												assign node3212 = (inp[4]) ? 11'b00100011111 : 11'b00101001111;
											assign node3216 = (inp[4]) ? node3218 : 11'b00100011101;
												assign node3218 = (inp[5]) ? 11'b00010001110 : 11'b00011101100;
								assign node3221 = (inp[10]) ? node3239 : node3222;
									assign node3222 = (inp[2]) ? node3230 : node3223;
										assign node3223 = (inp[5]) ? 11'b00000111110 : node3224;
											assign node3224 = (inp[11]) ? node3226 : 11'b00011111110;
												assign node3226 = (inp[4]) ? 11'b00101001110 : 11'b00001011100;
										assign node3230 = (inp[11]) ? node3232 : 11'b00101101100;
											assign node3232 = (inp[4]) ? node3236 : node3233;
												assign node3233 = (inp[5]) ? 11'b00010011100 : 11'b00000011111;
												assign node3236 = (inp[5]) ? 11'b00010001100 : 11'b00110101100;
									assign node3239 = (inp[11]) ? node3249 : node3240;
										assign node3240 = (inp[4]) ? node3246 : node3241;
											assign node3241 = (inp[5]) ? 11'b00000111010 : node3242;
												assign node3242 = (inp[2]) ? 11'b00111011001 : 11'b00110111010;
											assign node3246 = (inp[5]) ? 11'b00011011000 : 11'b00001111000;
										assign node3249 = (inp[4]) ? node3255 : node3250;
											assign node3250 = (inp[5]) ? 11'b00011001010 : node3251;
												assign node3251 = (inp[2]) ? 11'b00101101010 : 11'b00101001000;
											assign node3255 = (inp[5]) ? 11'b00010001000 : node3256;
												assign node3256 = (inp[2]) ? 11'b00010101010 : 11'b00011001010;
							assign node3260 = (inp[11]) ? node3304 : node3261;
								assign node3261 = (inp[5]) ? node3285 : node3262;
									assign node3262 = (inp[2]) ? node3274 : node3263;
										assign node3263 = (inp[10]) ? node3269 : node3264;
											assign node3264 = (inp[9]) ? 11'b00011111000 : node3265;
												assign node3265 = (inp[4]) ? 11'b00000111000 : 11'b00000001001;
											assign node3269 = (inp[9]) ? 11'b00000101000 : node3270;
												assign node3270 = (inp[4]) ? 11'b00111101000 : 11'b00011101000;
										assign node3274 = (inp[9]) ? node3282 : node3275;
											assign node3275 = (inp[4]) ? node3279 : node3276;
												assign node3276 = (inp[10]) ? 11'b00011001001 : 11'b00010101001;
												assign node3279 = (inp[10]) ? 11'b00110001001 : 11'b00010011011;
											assign node3282 = (inp[4]) ? 11'b00001001011 : 11'b00000001011;
									assign node3285 = (inp[10]) ? node3293 : node3286;
										assign node3286 = (inp[9]) ? 11'b00101111010 : node3287;
											assign node3287 = (inp[2]) ? node3289 : 11'b00100001000;
												assign node3289 = (inp[4]) ? 11'b00100111000 : 11'b00111101000;
										assign node3293 = (inp[4]) ? node3299 : node3294;
											assign node3294 = (inp[2]) ? node3296 : 11'b00011101010;
												assign node3296 = (inp[9]) ? 11'b00010101000 : 11'b00011101010;
											assign node3299 = (inp[9]) ? 11'b00001101000 : node3300;
												assign node3300 = (inp[2]) ? 11'b00101001010 : 11'b00100101010;
								assign node3304 = (inp[5]) ? node3328 : node3305;
									assign node3305 = (inp[4]) ? node3319 : node3306;
										assign node3306 = (inp[2]) ? node3314 : node3307;
											assign node3307 = (inp[9]) ? node3311 : node3308;
												assign node3308 = (inp[10]) ? 11'b00111001010 : 11'b00010101010;
												assign node3311 = (inp[10]) ? 11'b00010001010 : 11'b00101011010;
											assign node3314 = (inp[9]) ? node3316 : 11'b00110001011;
												assign node3316 = (inp[10]) ? 11'b00011101000 : 11'b00110011001;
										assign node3319 = (inp[10]) ? node3323 : node3320;
											assign node3320 = (inp[2]) ? 11'b00100101000 : 11'b00111001000;
											assign node3323 = (inp[2]) ? node3325 : 11'b00000001000;
												assign node3325 = (inp[9]) ? 11'b00000101000 : 11'b00000101010;
									assign node3328 = (inp[4]) ? node3338 : node3329;
										assign node3329 = (inp[9]) ? node3335 : node3330;
											assign node3330 = (inp[2]) ? node3332 : 11'b00100101000;
												assign node3332 = (inp[10]) ? 11'b00100001010 : 11'b00100001000;
											assign node3335 = (inp[2]) ? 11'b00001001000 : 11'b00001001010;
										assign node3338 = (inp[10]) ? node3344 : node3339;
											assign node3339 = (inp[9]) ? node3341 : 11'b00001011000;
												assign node3341 = (inp[2]) ? 11'b00000001010 : 11'b00010001010;
											assign node3344 = (inp[9]) ? 11'b00000001000 : 11'b00000001010;
				assign node3347 = (inp[2]) ? node3699 : node3348;
					assign node3348 = (inp[8]) ? node3516 : node3349;
						assign node3349 = (inp[5]) ? node3433 : node3350;
							assign node3350 = (inp[11]) ? node3392 : node3351;
								assign node3351 = (inp[0]) ? node3373 : node3352;
									assign node3352 = (inp[3]) ? node3364 : node3353;
										assign node3353 = (inp[10]) ? node3359 : node3354;
											assign node3354 = (inp[9]) ? 11'b00101101100 : node3355;
												assign node3355 = (inp[4]) ? 11'b00000101110 : 11'b00001101010;
											assign node3359 = (inp[9]) ? 11'b10000111110 : node3360;
												assign node3360 = (inp[4]) ? 11'b10000111100 : 11'b10001101000;
										assign node3364 = (inp[10]) ? 11'b00111101010 : node3365;
											assign node3365 = (inp[9]) ? node3369 : node3366;
												assign node3366 = (inp[4]) ? 11'b10010101100 : 11'b10011101000;
												assign node3369 = (inp[4]) ? 11'b10111111010 : 11'b10010101110;
									assign node3373 = (inp[3]) ? node3381 : node3374;
										assign node3374 = (inp[10]) ? node3378 : node3375;
											assign node3375 = (inp[9]) ? 11'b00011101100 : 11'b00011101010;
											assign node3378 = (inp[4]) ? 11'b00111111000 : 11'b00010111000;
										assign node3381 = (inp[4]) ? node3385 : node3382;
											assign node3382 = (inp[10]) ? 11'b00000101000 : 11'b00000111010;
											assign node3385 = (inp[9]) ? node3389 : node3386;
												assign node3386 = (inp[10]) ? 11'b00101101010 : 11'b00000111000;
												assign node3389 = (inp[10]) ? 11'b00001101000 : 11'b00101101010;
								assign node3392 = (inp[4]) ? node3406 : node3393;
									assign node3393 = (inp[9]) ? node3401 : node3394;
										assign node3394 = (inp[10]) ? 11'b10010101000 : node3395;
											assign node3395 = (inp[0]) ? node3397 : 11'b10000111010;
												assign node3397 = (inp[3]) ? 11'b00000101000 : 11'b00010111010;
										assign node3401 = (inp[10]) ? 11'b00001011100 : node3402;
											assign node3402 = (inp[0]) ? 11'b00110111100 : 11'b00110111000;
									assign node3406 = (inp[9]) ? node3420 : node3407;
										assign node3407 = (inp[3]) ? node3413 : node3408;
											assign node3408 = (inp[10]) ? 11'b00101001100 : node3409;
												assign node3409 = (inp[0]) ? 11'b00001011010 : 11'b00011001110;
											assign node3413 = (inp[10]) ? node3417 : node3414;
												assign node3414 = (inp[0]) ? 11'b00111011000 : 11'b10101001110;
												assign node3417 = (inp[0]) ? 11'b00010001010 : 11'b00100011010;
										assign node3420 = (inp[0]) ? node3428 : node3421;
											assign node3421 = (inp[3]) ? node3425 : node3422;
												assign node3422 = (inp[10]) ? 11'b10100011010 : 11'b00000011110;
												assign node3425 = (inp[10]) ? 11'b00110011000 : 11'b10010011000;
											assign node3428 = (inp[10]) ? node3430 : 11'b00110001010;
												assign node3430 = (inp[3]) ? 11'b00000001000 : 11'b00100001010;
							assign node3433 = (inp[11]) ? node3469 : node3434;
								assign node3434 = (inp[9]) ? node3450 : node3435;
									assign node3435 = (inp[4]) ? node3441 : node3436;
										assign node3436 = (inp[0]) ? node3438 : 11'b00000011000;
											assign node3438 = (inp[3]) ? 11'b00101001010 : 11'b00011001010;
										assign node3441 = (inp[3]) ? node3445 : node3442;
											assign node3442 = (inp[0]) ? 11'b00000011100 : 11'b10000001110;
											assign node3445 = (inp[10]) ? 11'b00010011000 : node3446;
												assign node3446 = (inp[0]) ? 11'b00110011010 : 11'b10100011110;
									assign node3450 = (inp[4]) ? node3460 : node3451;
										assign node3451 = (inp[10]) ? 11'b10110001110 : node3452;
											assign node3452 = (inp[3]) ? node3456 : node3453;
												assign node3453 = (inp[0]) ? 11'b00011001100 : 11'b00011011010;
												assign node3456 = (inp[0]) ? 11'b00101011000 : 11'b10001011100;
										assign node3460 = (inp[3]) ? node3464 : node3461;
											assign node3461 = (inp[10]) ? 11'b10001110001 : 11'b00101110111;
											assign node3464 = (inp[0]) ? node3466 : 11'b10011100001;
												assign node3466 = (inp[10]) ? 11'b00001100011 : 11'b00001100001;
								assign node3469 = (inp[0]) ? node3493 : node3470;
									assign node3470 = (inp[9]) ? node3480 : node3471;
										assign node3471 = (inp[4]) ? node3473 : 11'b00000100101;
											assign node3473 = (inp[10]) ? node3477 : node3474;
												assign node3474 = (inp[3]) ? 11'b10111110101 : 11'b00001110111;
												assign node3477 = (inp[3]) ? 11'b00101100011 : 11'b10011100111;
										assign node3480 = (inp[4]) ? node3486 : node3481;
											assign node3481 = (inp[3]) ? 11'b00011100111 : node3482;
												assign node3482 = (inp[10]) ? 11'b10100100101 : 11'b00110100011;
											assign node3486 = (inp[3]) ? node3490 : node3487;
												assign node3487 = (inp[10]) ? 11'b10000100011 : 11'b00011100101;
												assign node3490 = (inp[10]) ? 11'b00110100001 : 11'b10100100011;
									assign node3493 = (inp[3]) ? node3503 : node3494;
										assign node3494 = (inp[9]) ? node3500 : node3495;
											assign node3495 = (inp[10]) ? 11'b00111100111 : node3496;
												assign node3496 = (inp[4]) ? 11'b00111110001 : 11'b00011110001;
											assign node3500 = (inp[4]) ? 11'b00101100101 : 11'b00100110111;
										assign node3503 = (inp[10]) ? node3509 : node3504;
											assign node3504 = (inp[9]) ? node3506 : 11'b00001110001;
												assign node3506 = (inp[4]) ? 11'b00010100011 : 11'b00010110001;
											assign node3509 = (inp[9]) ? node3513 : node3510;
												assign node3510 = (inp[4]) ? 11'b00011100001 : 11'b00110100001;
												assign node3513 = (inp[4]) ? 11'b00000100001 : 11'b00001100011;
						assign node3516 = (inp[0]) ? node3600 : node3517;
							assign node3517 = (inp[5]) ? node3561 : node3518;
								assign node3518 = (inp[11]) ? node3540 : node3519;
									assign node3519 = (inp[9]) ? node3529 : node3520;
										assign node3520 = (inp[4]) ? node3526 : node3521;
											assign node3521 = (inp[3]) ? node3523 : 11'b10010100001;
												assign node3523 = (inp[10]) ? 11'b00101000111 : 11'b10110100001;
											assign node3526 = (inp[3]) ? 11'b00000000001 : 11'b00101000101;
										assign node3529 = (inp[4]) ? node3535 : node3530;
											assign node3530 = (inp[10]) ? node3532 : 11'b00011000001;
												assign node3532 = (inp[3]) ? 11'b00111010101 : 11'b10001010111;
											assign node3535 = (inp[3]) ? 11'b10010010001 : node3536;
												assign node3536 = (inp[10]) ? 11'b10000000001 : 11'b00110000111;
									assign node3540 = (inp[4]) ? node3554 : node3541;
										assign node3541 = (inp[9]) ? node3547 : node3542;
											assign node3542 = (inp[3]) ? node3544 : 11'b10111000011;
												assign node3544 = (inp[10]) ? 11'b00011010101 : 11'b10101010001;
											assign node3547 = (inp[10]) ? node3551 : node3548;
												assign node3548 = (inp[3]) ? 11'b10110000111 : 11'b00101010001;
												assign node3551 = (inp[3]) ? 11'b00100010101 : 11'b10010010101;
										assign node3554 = (inp[9]) ? node3558 : node3555;
											assign node3555 = (inp[3]) ? 11'b10010000101 : 11'b00110000111;
											assign node3558 = (inp[10]) ? 11'b10111110011 : 11'b00011110101;
								assign node3561 = (inp[11]) ? node3581 : node3562;
									assign node3562 = (inp[10]) ? node3572 : node3563;
										assign node3563 = (inp[4]) ? 11'b00111110101 : node3564;
											assign node3564 = (inp[3]) ? node3568 : node3565;
												assign node3565 = (inp[9]) ? 11'b00000110011 : 11'b00001110001;
												assign node3568 = (inp[9]) ? 11'b10010110101 : 11'b10000110011;
										assign node3572 = (inp[3]) ? node3578 : node3573;
											assign node3573 = (inp[4]) ? node3575 : 11'b10110110001;
												assign node3575 = (inp[9]) ? 11'b10100110011 : 11'b10001100111;
											assign node3578 = (inp[4]) ? 11'b00110100001 : 11'b00101100111;
									assign node3581 = (inp[4]) ? node3593 : node3582;
										assign node3582 = (inp[9]) ? node3590 : node3583;
											assign node3583 = (inp[3]) ? node3587 : node3584;
												assign node3584 = (inp[10]) ? 11'b10000110001 : 11'b00010110011;
												assign node3587 = (inp[10]) ? 11'b00011000111 : 11'b10000100011;
											assign node3590 = (inp[10]) ? 11'b00111000111 : 11'b00011000011;
										assign node3593 = (inp[10]) ? node3597 : node3594;
											assign node3594 = (inp[9]) ? 11'b00100000101 : 11'b00101010101;
											assign node3597 = (inp[3]) ? 11'b00110000001 : 11'b10110000001;
							assign node3600 = (inp[3]) ? node3648 : node3601;
								assign node3601 = (inp[5]) ? node3621 : node3602;
									assign node3602 = (inp[9]) ? node3614 : node3603;
										assign node3603 = (inp[11]) ? node3609 : node3604;
											assign node3604 = (inp[10]) ? 11'b00110010101 : node3605;
												assign node3605 = (inp[4]) ? 11'b00110000011 : 11'b00110100011;
											assign node3609 = (inp[10]) ? 11'b00101010111 : node3610;
												assign node3610 = (inp[4]) ? 11'b00100010011 : 11'b00111010001;
										assign node3614 = (inp[10]) ? node3618 : node3615;
											assign node3615 = (inp[4]) ? 11'b00000010111 : 11'b00010010111;
											assign node3618 = (inp[4]) ? 11'b00011010011 : 11'b00110000001;
									assign node3621 = (inp[11]) ? node3635 : node3622;
										assign node3622 = (inp[4]) ? node3630 : node3623;
											assign node3623 = (inp[10]) ? node3627 : node3624;
												assign node3624 = (inp[9]) ? 11'b00100100111 : 11'b00110100011;
												assign node3627 = (inp[9]) ? 11'b00011110011 : 11'b00000100101;
											assign node3630 = (inp[10]) ? 11'b00111110111 : node3631;
												assign node3631 = (inp[9]) ? 11'b00001110101 : 11'b00001100001;
										assign node3635 = (inp[4]) ? node3641 : node3636;
											assign node3636 = (inp[9]) ? 11'b00011010101 : node3637;
												assign node3637 = (inp[10]) ? 11'b00100110101 : 11'b00110110011;
											assign node3641 = (inp[10]) ? node3645 : node3642;
												assign node3642 = (inp[9]) ? 11'b00010000111 : 11'b00011010001;
												assign node3645 = (inp[9]) ? 11'b00000000001 : 11'b00000000111;
								assign node3648 = (inp[10]) ? node3676 : node3649;
									assign node3649 = (inp[4]) ? node3661 : node3650;
										assign node3650 = (inp[9]) ? node3654 : node3651;
											assign node3651 = (inp[11]) ? 11'b00011000011 : 11'b00000100001;
											assign node3654 = (inp[5]) ? node3658 : node3655;
												assign node3655 = (inp[11]) ? 11'b00100010011 : 11'b00011010011;
												assign node3658 = (inp[11]) ? 11'b00011010001 : 11'b00100110001;
										assign node3661 = (inp[9]) ? node3669 : node3662;
											assign node3662 = (inp[11]) ? node3666 : node3663;
												assign node3663 = (inp[5]) ? 11'b00111110011 : 11'b00000010011;
												assign node3666 = (inp[5]) ? 11'b00010010011 : 11'b00110010001;
											assign node3669 = (inp[5]) ? node3673 : node3670;
												assign node3670 = (inp[11]) ? 11'b00111100011 : 11'b00110000001;
												assign node3673 = (inp[11]) ? 11'b00010000011 : 11'b00010100011;
									assign node3676 = (inp[4]) ? node3690 : node3677;
										assign node3677 = (inp[5]) ? node3685 : node3678;
											assign node3678 = (inp[9]) ? node3682 : node3679;
												assign node3679 = (inp[11]) ? 11'b00111000001 : 11'b00011000011;
												assign node3682 = (inp[11]) ? 11'b00010000011 : 11'b00001000001;
											assign node3685 = (inp[11]) ? 11'b00001000011 : node3686;
												assign node3686 = (inp[9]) ? 11'b00011100011 : 11'b00010100011;
										assign node3690 = (inp[5]) ? node3696 : node3691;
											assign node3691 = (inp[11]) ? node3693 : 11'b00001000011;
												assign node3693 = (inp[9]) ? 11'b00001100001 : 11'b00001100011;
											assign node3696 = (inp[11]) ? 11'b00000000001 : 11'b00101100001;
					assign node3699 = (inp[5]) ? node3857 : node3700;
						assign node3700 = (inp[11]) ? node3766 : node3701;
							assign node3701 = (inp[8]) ? node3737 : node3702;
								assign node3702 = (inp[9]) ? node3724 : node3703;
									assign node3703 = (inp[4]) ? node3713 : node3704;
										assign node3704 = (inp[0]) ? node3710 : node3705;
											assign node3705 = (inp[10]) ? node3707 : 11'b00101000011;
												assign node3707 = (inp[3]) ? 11'b00111000111 : 11'b10111000001;
											assign node3710 = (inp[3]) ? 11'b00001000011 : 11'b00001000101;
										assign node3713 = (inp[0]) ? node3717 : node3714;
											assign node3714 = (inp[3]) ? 11'b00010000001 : 11'b00100000101;
											assign node3717 = (inp[10]) ? node3721 : node3718;
												assign node3718 = (inp[3]) ? 11'b00010010011 : 11'b00010000001;
												assign node3721 = (inp[3]) ? 11'b00100000001 : 11'b00000010111;
									assign node3724 = (inp[4]) ? node3730 : node3725;
										assign node3725 = (inp[0]) ? node3727 : 11'b10110010111;
											assign node3727 = (inp[3]) ? 11'b00000000011 : 11'b00000010011;
										assign node3730 = (inp[0]) ? node3734 : node3731;
											assign node3731 = (inp[10]) ? 11'b10001100010 : 11'b10001110010;
											assign node3734 = (inp[3]) ? 11'b00111100010 : 11'b00101110000;
								assign node3737 = (inp[4]) ? node3753 : node3738;
									assign node3738 = (inp[9]) ? node3748 : node3739;
										assign node3739 = (inp[0]) ? node3745 : node3740;
											assign node3740 = (inp[3]) ? 11'b10000000010 : node3741;
												assign node3741 = (inp[10]) ? 11'b10100000000 : 11'b00100000010;
											assign node3745 = (inp[3]) ? 11'b00011100010 : 11'b00110000010;
										assign node3748 = (inp[3]) ? 11'b00001100010 : node3749;
											assign node3749 = (inp[0]) ? 11'b00101100110 : 11'b00111100010;
									assign node3753 = (inp[9]) ? node3763 : node3754;
										assign node3754 = (inp[0]) ? node3760 : node3755;
											assign node3755 = (inp[3]) ? node3757 : 11'b10001110100;
												assign node3757 = (inp[10]) ? 11'b00100100010 : 11'b10101100100;
											assign node3760 = (inp[10]) ? 11'b00110110110 : 11'b00011110000;
										assign node3763 = (inp[10]) ? 11'b10110100010 : 11'b10110110000;
							assign node3766 = (inp[0]) ? node3816 : node3767;
								assign node3767 = (inp[10]) ? node3789 : node3768;
									assign node3768 = (inp[3]) ? node3778 : node3769;
										assign node3769 = (inp[9]) ? node3775 : node3770;
											assign node3770 = (inp[4]) ? 11'b00001100100 : node3771;
												assign node3771 = (inp[8]) ? 11'b00110100000 : 11'b00111100010;
											assign node3775 = (inp[8]) ? 11'b00001110000 : 11'b00101110100;
										assign node3778 = (inp[8]) ? node3786 : node3779;
											assign node3779 = (inp[9]) ? node3783 : node3780;
												assign node3780 = (inp[4]) ? 11'b10010100100 : 11'b10101110010;
												assign node3783 = (inp[4]) ? 11'b10111110010 : 11'b10010100100;
											assign node3786 = (inp[4]) ? 11'b10110110010 : 11'b10010110000;
									assign node3789 = (inp[3]) ? node3805 : node3790;
										assign node3790 = (inp[4]) ? node3798 : node3791;
											assign node3791 = (inp[9]) ? node3795 : node3792;
												assign node3792 = (inp[8]) ? 11'b10011100010 : 11'b10101100000;
												assign node3795 = (inp[8]) ? 11'b10101110110 : 11'b10000110100;
											assign node3798 = (inp[8]) ? node3802 : node3799;
												assign node3799 = (inp[9]) ? 11'b10011110010 : 11'b10011110110;
												assign node3802 = (inp[9]) ? 11'b10010110010 : 11'b10010110110;
										assign node3805 = (inp[4]) ? node3811 : node3806;
											assign node3806 = (inp[8]) ? node3808 : 11'b00110110110;
												assign node3808 = (inp[9]) ? 11'b00001110110 : 11'b00101110110;
											assign node3811 = (inp[9]) ? node3813 : 11'b00001110010;
												assign node3813 = (inp[8]) ? 11'b00010110000 : 11'b00011110000;
								assign node3816 = (inp[10]) ? node3838 : node3817;
									assign node3817 = (inp[9]) ? node3829 : node3818;
										assign node3818 = (inp[4]) ? node3824 : node3819;
											assign node3819 = (inp[3]) ? node3821 : 11'b00001110010;
												assign node3821 = (inp[8]) ? 11'b00000100000 : 11'b00011100000;
											assign node3824 = (inp[8]) ? 11'b00101110000 : node3825;
												assign node3825 = (inp[3]) ? 11'b00100110000 : 11'b00000110000;
										assign node3829 = (inp[3]) ? node3835 : node3830;
											assign node3830 = (inp[4]) ? node3832 : 11'b00011110100;
												assign node3832 = (inp[8]) ? 11'b00100100100 : 11'b00011100100;
											assign node3835 = (inp[8]) ? 11'b00111110010 : 11'b00110110000;
									assign node3838 = (inp[4]) ? node3848 : node3839;
										assign node3839 = (inp[8]) ? node3843 : node3840;
											assign node3840 = (inp[3]) ? 11'b00100100010 : 11'b00011110100;
											assign node3843 = (inp[3]) ? node3845 : 11'b00111100010;
												assign node3845 = (inp[9]) ? 11'b00011100000 : 11'b00111100000;
										assign node3848 = (inp[8]) ? node3852 : node3849;
											assign node3849 = (inp[9]) ? 11'b00101100010 : 11'b00111100110;
											assign node3852 = (inp[3]) ? 11'b00000100000 : node3853;
												assign node3853 = (inp[9]) ? 11'b00000100010 : 11'b00000100110;
						assign node3857 = (inp[10]) ? node3927 : node3858;
							assign node3858 = (inp[9]) ? node3884 : node3859;
								assign node3859 = (inp[0]) ? node3871 : node3860;
									assign node3860 = (inp[8]) ? node3866 : node3861;
										assign node3861 = (inp[3]) ? node3863 : 11'b00110010000;
											assign node3863 = (inp[11]) ? 11'b10010000000 : 11'b10011010100;
										assign node3866 = (inp[11]) ? node3868 : 11'b10101010010;
											assign node3868 = (inp[3]) ? 11'b10111000010 : 11'b00111010010;
									assign node3871 = (inp[4]) ? node3877 : node3872;
										assign node3872 = (inp[8]) ? node3874 : 11'b00110000010;
											assign node3874 = (inp[11]) ? 11'b00101000010 : 11'b00111000010;
										assign node3877 = (inp[11]) ? node3879 : 11'b00101000010;
											assign node3879 = (inp[8]) ? 11'b00000010010 : node3880;
												assign node3880 = (inp[3]) ? 11'b00011010010 : 11'b00111010010;
								assign node3884 = (inp[4]) ? node3908 : node3885;
									assign node3885 = (inp[8]) ? node3897 : node3886;
										assign node3886 = (inp[11]) ? node3894 : node3887;
											assign node3887 = (inp[3]) ? node3891 : node3888;
												assign node3888 = (inp[0]) ? 11'b00000100110 : 11'b00110110010;
												assign node3891 = (inp[0]) ? 11'b00110110000 : 11'b10100110110;
											assign node3894 = (inp[0]) ? 11'b00100010100 : 11'b00000000000;
										assign node3897 = (inp[3]) ? node3903 : node3898;
											assign node3898 = (inp[0]) ? 11'b00111000110 : node3899;
												assign node3899 = (inp[11]) ? 11'b00111000010 : 11'b00101010000;
											assign node3903 = (inp[0]) ? 11'b00111010010 : node3904;
												assign node3904 = (inp[11]) ? 11'b10011010110 : 11'b10101010110;
									assign node3908 = (inp[3]) ? node3922 : node3909;
										assign node3909 = (inp[11]) ? node3917 : node3910;
											assign node3910 = (inp[8]) ? node3914 : node3911;
												assign node3911 = (inp[0]) ? 11'b00111010100 : 11'b00001010110;
												assign node3914 = (inp[0]) ? 11'b00000010110 : 11'b00010010110;
											assign node3917 = (inp[8]) ? 11'b00000000110 : node3918;
												assign node3918 = (inp[0]) ? 11'b00100000110 : 11'b00110000110;
										assign node3922 = (inp[0]) ? node3924 : 11'b10010000010;
											assign node3924 = (inp[8]) ? 11'b00000000010 : 11'b00011000000;
							assign node3927 = (inp[3]) ? node3969 : node3928;
								assign node3928 = (inp[0]) ? node3950 : node3929;
									assign node3929 = (inp[4]) ? node3941 : node3930;
										assign node3930 = (inp[9]) ? node3936 : node3931;
											assign node3931 = (inp[8]) ? 11'b10111010000 : node3932;
												assign node3932 = (inp[11]) ? 11'b10000010010 : 11'b10000110010;
											assign node3936 = (inp[11]) ? 11'b10011000110 : node3937;
												assign node3937 = (inp[8]) ? 11'b10101000110 : 11'b10000100100;
										assign node3941 = (inp[9]) ? node3945 : node3942;
											assign node3942 = (inp[8]) ? 11'b10110000100 : 11'b10111000100;
											assign node3945 = (inp[8]) ? node3947 : 11'b10110010010;
												assign node3947 = (inp[11]) ? 11'b10010000000 : 11'b10010010000;
									assign node3950 = (inp[9]) ? node3958 : node3951;
										assign node3951 = (inp[11]) ? node3953 : 11'b00100100100;
											assign node3953 = (inp[4]) ? node3955 : 11'b00010010110;
												assign node3955 = (inp[8]) ? 11'b00000000100 : 11'b00111000100;
										assign node3958 = (inp[8]) ? node3964 : node3959;
											assign node3959 = (inp[4]) ? node3961 : 11'b00101000010;
												assign node3961 = (inp[11]) ? 11'b00100000000 : 11'b00100010010;
											assign node3964 = (inp[4]) ? 11'b00000010000 : node3965;
												assign node3965 = (inp[11]) ? 11'b00001000000 : 11'b00011010000;
								assign node3969 = (inp[4]) ? node3991 : node3970;
									assign node3970 = (inp[0]) ? node3982 : node3971;
										assign node3971 = (inp[8]) ? node3977 : node3972;
											assign node3972 = (inp[9]) ? node3974 : 11'b00100000110;
												assign node3974 = (inp[11]) ? 11'b00111000100 : 11'b00100100100;
											assign node3977 = (inp[11]) ? node3979 : 11'b00001010100;
												assign node3979 = (inp[9]) ? 11'b00011000100 : 11'b00111000100;
										assign node3982 = (inp[11]) ? node3986 : node3983;
											assign node3983 = (inp[8]) ? 11'b00011000000 : 11'b00000100000;
											assign node3986 = (inp[9]) ? 11'b00001000000 : node3987;
												assign node3987 = (inp[8]) ? 11'b00101000000 : 11'b00110000000;
									assign node3991 = (inp[9]) ? node4003 : node3992;
										assign node3992 = (inp[11]) ? node3998 : node3993;
											assign node3993 = (inp[8]) ? node3995 : 11'b00101010010;
												assign node3995 = (inp[0]) ? 11'b00100000000 : 11'b00110010000;
											assign node3998 = (inp[8]) ? 11'b00010000000 : node3999;
												assign node3999 = (inp[0]) ? 11'b00011000000 : 11'b00001000000;
										assign node4003 = (inp[0]) ? node4009 : node4004;
											assign node4004 = (inp[8]) ? 11'b00010000000 : node4005;
												assign node4005 = (inp[11]) ? 11'b00010000000 : 11'b00010000010;
											assign node4009 = (inp[11]) ? 11'b00000000000 : 11'b00000000010;
			assign node4012 = (inp[6]) ? node4670 : node4013;
				assign node4013 = (inp[2]) ? node4329 : node4014;
					assign node4014 = (inp[5]) ? node4158 : node4015;
						assign node4015 = (inp[0]) ? node4083 : node4016;
							assign node4016 = (inp[10]) ? node4056 : node4017;
								assign node4017 = (inp[3]) ? node4039 : node4018;
									assign node4018 = (inp[4]) ? node4026 : node4019;
										assign node4019 = (inp[8]) ? node4023 : node4020;
											assign node4020 = (inp[11]) ? 11'b00111110011 : 11'b00011100011;
											assign node4023 = (inp[11]) ? 11'b00100110011 : 11'b00000000001;
										assign node4026 = (inp[8]) ? node4032 : node4027;
											assign node4027 = (inp[11]) ? 11'b00001100101 : node4028;
												assign node4028 = (inp[9]) ? 11'b00110100111 : 11'b00010100111;
											assign node4032 = (inp[11]) ? node4036 : node4033;
												assign node4033 = (inp[9]) ? 11'b00101100101 : 11'b00111100101;
												assign node4036 = (inp[9]) ? 11'b00011110111 : 11'b00101100111;
									assign node4039 = (inp[4]) ? node4049 : node4040;
										assign node4040 = (inp[9]) ? node4044 : node4041;
											assign node4041 = (inp[11]) ? 11'b10011110011 : 11'b10011100011;
											assign node4044 = (inp[11]) ? node4046 : 11'b10101100111;
												assign node4046 = (inp[8]) ? 11'b10110100101 : 11'b10111100111;
										assign node4049 = (inp[9]) ? node4051 : 11'b10010100111;
											assign node4051 = (inp[11]) ? node4053 : 11'b10001110001;
												assign node4053 = (inp[8]) ? 11'b10001110011 : 11'b10000110011;
								assign node4056 = (inp[3]) ? node4068 : node4057;
									assign node4057 = (inp[4]) ? node4063 : node4058;
										assign node4058 = (inp[9]) ? 11'b10001110111 : node4059;
											assign node4059 = (inp[8]) ? 11'b10100100001 : 11'b10011100001;
										assign node4063 = (inp[8]) ? node4065 : 11'b10100110111;
											assign node4065 = (inp[9]) ? 11'b10101110011 : 11'b10101110101;
									assign node4068 = (inp[4]) ? node4076 : node4069;
										assign node4069 = (inp[9]) ? node4073 : node4070;
											assign node4070 = (inp[8]) ? 11'b00110000101 : 11'b00011100101;
											assign node4073 = (inp[11]) ? 11'b00001110101 : 11'b00101110101;
										assign node4076 = (inp[8]) ? node4080 : node4077;
											assign node4077 = (inp[11]) ? 11'b00100110001 : 11'b00110110001;
											assign node4080 = (inp[9]) ? 11'b00110110011 : 11'b00111110001;
							assign node4083 = (inp[10]) ? node4123 : node4084;
								assign node4084 = (inp[9]) ? node4104 : node4085;
									assign node4085 = (inp[11]) ? node4097 : node4086;
										assign node4086 = (inp[4]) ? node4090 : node4087;
											assign node4087 = (inp[3]) ? 11'b00000000011 : 11'b00100000011;
											assign node4090 = (inp[8]) ? node4094 : node4091;
												assign node4091 = (inp[3]) ? 11'b00000110011 : 11'b00000100011;
												assign node4094 = (inp[3]) ? 11'b00001110011 : 11'b00101100001;
										assign node4097 = (inp[8]) ? node4101 : node4098;
											assign node4098 = (inp[4]) ? 11'b00010110011 : 11'b00001110011;
											assign node4101 = (inp[3]) ? 11'b00111110001 : 11'b00100110001;
									assign node4104 = (inp[3]) ? node4116 : node4105;
										assign node4105 = (inp[4]) ? node4111 : node4106;
											assign node4106 = (inp[11]) ? 11'b00000110111 : node4107;
												assign node4107 = (inp[8]) ? 11'b00111100111 : 11'b00001100111;
											assign node4111 = (inp[8]) ? 11'b00101100111 : node4112;
												assign node4112 = (inp[11]) ? 11'b00010100111 : 11'b00100110111;
										assign node4116 = (inp[11]) ? 11'b00100110001 : node4117;
											assign node4117 = (inp[4]) ? 11'b00100100011 : node4118;
												assign node4118 = (inp[8]) ? 11'b00011110011 : 11'b00001110011;
								assign node4123 = (inp[3]) ? node4143 : node4124;
									assign node4124 = (inp[9]) ? node4136 : node4125;
										assign node4125 = (inp[8]) ? node4129 : node4126;
											assign node4126 = (inp[4]) ? 11'b00000110101 : 11'b00001100101;
											assign node4129 = (inp[4]) ? node4133 : node4130;
												assign node4130 = (inp[11]) ? 11'b00110110111 : 11'b00100000101;
												assign node4133 = (inp[11]) ? 11'b00001100101 : 11'b00101110111;
										assign node4136 = (inp[4]) ? node4140 : node4137;
											assign node4137 = (inp[11]) ? 11'b00011100001 : 11'b00111110001;
											assign node4140 = (inp[8]) ? 11'b00000110011 : 11'b00110100001;
									assign node4143 = (inp[8]) ? node4151 : node4144;
										assign node4144 = (inp[4]) ? node4148 : node4145;
											assign node4145 = (inp[11]) ? 11'b00101100001 : 11'b00001100001;
											assign node4148 = (inp[9]) ? 11'b00000100001 : 11'b00100100001;
										assign node4151 = (inp[9]) ? node4155 : node4152;
											assign node4152 = (inp[4]) ? 11'b00111100001 : 11'b00110100011;
											assign node4155 = (inp[4]) ? 11'b00001100001 : 11'b00011100011;
						assign node4158 = (inp[0]) ? node4244 : node4159;
							assign node4159 = (inp[11]) ? node4205 : node4160;
								assign node4160 = (inp[10]) ? node4182 : node4161;
									assign node4161 = (inp[3]) ? node4171 : node4162;
										assign node4162 = (inp[4]) ? 11'b00100110111 : node4163;
											assign node4163 = (inp[9]) ? node4167 : node4164;
												assign node4164 = (inp[8]) ? 11'b00011110001 : 11'b00010110001;
												assign node4167 = (inp[8]) ? 11'b00000110001 : 11'b00011010001;
										assign node4171 = (inp[8]) ? node4177 : node4172;
											assign node4172 = (inp[9]) ? node4174 : 11'b10101010101;
												assign node4174 = (inp[4]) ? 11'b10010000001 : 11'b10011010111;
											assign node4177 = (inp[4]) ? 11'b10000110101 : node4178;
												assign node4178 = (inp[9]) ? 11'b10010110101 : 11'b10010110011;
									assign node4182 = (inp[3]) ? node4192 : node4183;
										assign node4183 = (inp[4]) ? node4189 : node4184;
											assign node4184 = (inp[9]) ? 11'b10010100111 : node4185;
												assign node4185 = (inp[8]) ? 11'b10110110011 : 11'b10111010011;
											assign node4189 = (inp[9]) ? 11'b10101010001 : 11'b10000000111;
										assign node4192 = (inp[9]) ? node4198 : node4193;
											assign node4193 = (inp[4]) ? node4195 : 11'b00111010101;
												assign node4195 = (inp[8]) ? 11'b00011010011 : 11'b00000010011;
											assign node4198 = (inp[4]) ? node4202 : node4199;
												assign node4199 = (inp[8]) ? 11'b00110100111 : 11'b00001000111;
												assign node4202 = (inp[8]) ? 11'b00111000001 : 11'b00110000011;
								assign node4205 = (inp[9]) ? node4229 : node4206;
									assign node4206 = (inp[3]) ? node4214 : node4207;
										assign node4207 = (inp[10]) ? node4211 : node4208;
											assign node4208 = (inp[8]) ? 11'b00011010011 : 11'b00011010111;
											assign node4211 = (inp[8]) ? 11'b10001010011 : 11'b10111010011;
										assign node4214 = (inp[10]) ? node4222 : node4215;
											assign node4215 = (inp[4]) ? node4219 : node4216;
												assign node4216 = (inp[8]) ? 11'b10001000011 : 11'b10110000001;
												assign node4219 = (inp[8]) ? 11'b10110010101 : 11'b10111010101;
											assign node4222 = (inp[4]) ? node4226 : node4223;
												assign node4223 = (inp[8]) ? 11'b00011000101 : 11'b00001000111;
												assign node4226 = (inp[8]) ? 11'b00100000011 : 11'b00110000011;
									assign node4229 = (inp[4]) ? node4237 : node4230;
										assign node4230 = (inp[3]) ? 11'b00011000111 : node4231;
											assign node4231 = (inp[10]) ? node4233 : 11'b00101000011;
												assign node4233 = (inp[8]) ? 11'b10100000111 : 11'b10101000101;
										assign node4237 = (inp[10]) ? node4241 : node4238;
											assign node4238 = (inp[3]) ? 11'b10100000011 : 11'b00000000111;
											assign node4241 = (inp[3]) ? 11'b00100000001 : 11'b10100000001;
							assign node4244 = (inp[3]) ? node4292 : node4245;
								assign node4245 = (inp[11]) ? node4271 : node4246;
									assign node4246 = (inp[4]) ? node4260 : node4247;
										assign node4247 = (inp[10]) ? node4255 : node4248;
											assign node4248 = (inp[8]) ? node4252 : node4249;
												assign node4249 = (inp[9]) ? 11'b00001000101 : 11'b00000100001;
												assign node4252 = (inp[9]) ? 11'b00110100101 : 11'b00101100001;
											assign node4255 = (inp[8]) ? node4257 : 11'b00101000111;
												assign node4257 = (inp[9]) ? 11'b00000110011 : 11'b00010100111;
										assign node4260 = (inp[9]) ? node4266 : node4261;
											assign node4261 = (inp[10]) ? node4263 : 11'b00010100001;
												assign node4263 = (inp[8]) ? 11'b00100110101 : 11'b00010010111;
											assign node4266 = (inp[8]) ? 11'b00011010111 : node4267;
												assign node4267 = (inp[10]) ? 11'b00100010011 : 11'b00110010101;
									assign node4271 = (inp[4]) ? node4283 : node4272;
										assign node4272 = (inp[10]) ? node4276 : node4273;
											assign node4273 = (inp[9]) ? 11'b00001010101 : 11'b00000010001;
											assign node4276 = (inp[9]) ? node4280 : node4277;
												assign node4277 = (inp[8]) ? 11'b00111010101 : 11'b00011010111;
												assign node4280 = (inp[8]) ? 11'b00010000011 : 11'b00111000011;
										assign node4283 = (inp[8]) ? node4289 : node4284;
											assign node4284 = (inp[9]) ? 11'b00110000111 : node4285;
												assign node4285 = (inp[10]) ? 11'b00101000101 : 11'b00101010011;
											assign node4289 = (inp[10]) ? 11'b00010000111 : 11'b00000000111;
								assign node4292 = (inp[10]) ? node4310 : node4293;
									assign node4293 = (inp[4]) ? node4303 : node4294;
										assign node4294 = (inp[8]) ? node4300 : node4295;
											assign node4295 = (inp[11]) ? 11'b00100000001 : node4296;
												assign node4296 = (inp[9]) ? 11'b00101010011 : 11'b00101000011;
											assign node4300 = (inp[9]) ? 11'b00100110001 : 11'b00100100011;
										assign node4303 = (inp[9]) ? node4307 : node4304;
											assign node4304 = (inp[8]) ? 11'b00110110001 : 11'b00001010001;
											assign node4307 = (inp[8]) ? 11'b00011000001 : 11'b00000000001;
									assign node4310 = (inp[9]) ? node4318 : node4311;
										assign node4311 = (inp[4]) ? node4313 : 11'b00010100001;
											assign node4313 = (inp[8]) ? 11'b00101000011 : node4314;
												assign node4314 = (inp[11]) ? 11'b00010000011 : 11'b00110000001;
										assign node4318 = (inp[4]) ? node4324 : node4319;
											assign node4319 = (inp[11]) ? node4321 : 11'b00011000001;
												assign node4321 = (inp[8]) ? 11'b00000000011 : 11'b00001000011;
											assign node4324 = (inp[8]) ? 11'b00001000001 : node4325;
												assign node4325 = (inp[11]) ? 11'b00000000001 : 11'b00000000011;
					assign node4329 = (inp[8]) ? node4497 : node4330;
						assign node4330 = (inp[5]) ? node4420 : node4331;
							assign node4331 = (inp[11]) ? node4371 : node4332;
								assign node4332 = (inp[4]) ? node4352 : node4333;
									assign node4333 = (inp[0]) ? node4345 : node4334;
										assign node4334 = (inp[10]) ? node4340 : node4335;
											assign node4335 = (inp[3]) ? 11'b10111000111 : node4336;
												assign node4336 = (inp[9]) ? 11'b00111000001 : 11'b00111000011;
											assign node4340 = (inp[3]) ? node4342 : 11'b10101000011;
												assign node4342 = (inp[9]) ? 11'b00101010111 : 11'b00101000101;
										assign node4345 = (inp[10]) ? 11'b00011010011 : node4346;
											assign node4346 = (inp[9]) ? 11'b00001000101 : node4347;
												assign node4347 = (inp[3]) ? 11'b00011000011 : 11'b00001000011;
									assign node4352 = (inp[9]) ? node4360 : node4353;
										assign node4353 = (inp[0]) ? node4357 : node4354;
											assign node4354 = (inp[10]) ? 11'b10101010101 : 11'b00111000101;
											assign node4357 = (inp[10]) ? 11'b00100000011 : 11'b00001000001;
										assign node4360 = (inp[0]) ? node4368 : node4361;
											assign node4361 = (inp[10]) ? node4365 : node4362;
												assign node4362 = (inp[3]) ? 11'b10000010011 : 11'b00010000111;
												assign node4365 = (inp[3]) ? 11'b00010010001 : 11'b10000000001;
											assign node4368 = (inp[3]) ? 11'b00110000001 : 11'b00110010001;
								assign node4371 = (inp[4]) ? node4399 : node4372;
									assign node4372 = (inp[9]) ? node4384 : node4373;
										assign node4373 = (inp[0]) ? node4381 : node4374;
											assign node4374 = (inp[3]) ? node4378 : node4375;
												assign node4375 = (inp[10]) ? 11'b10100000011 : 11'b00110000011;
												assign node4378 = (inp[10]) ? 11'b00110010101 : 11'b10100010011;
											assign node4381 = (inp[3]) ? 11'b00100000001 : 11'b00000010111;
										assign node4384 = (inp[10]) ? node4392 : node4385;
											assign node4385 = (inp[0]) ? node4389 : node4386;
												assign node4386 = (inp[3]) ? 11'b10000000101 : 11'b00000010001;
												assign node4389 = (inp[3]) ? 11'b00111110010 : 11'b00110010101;
											assign node4392 = (inp[0]) ? node4396 : node4393;
												assign node4393 = (inp[3]) ? 11'b00111110110 : 11'b10011110110;
												assign node4396 = (inp[3]) ? 11'b00011100010 : 11'b00001100010;
									assign node4399 = (inp[9]) ? node4409 : node4400;
										assign node4400 = (inp[0]) ? node4404 : node4401;
											assign node4401 = (inp[10]) ? 11'b00001110000 : 11'b10011100100;
											assign node4404 = (inp[10]) ? 11'b00011100010 : node4405;
												assign node4405 = (inp[3]) ? 11'b00101110000 : 11'b00011110000;
										assign node4409 = (inp[0]) ? node4417 : node4410;
											assign node4410 = (inp[10]) ? node4414 : node4411;
												assign node4411 = (inp[3]) ? 11'b10111110010 : 11'b00101110110;
												assign node4414 = (inp[3]) ? 11'b00001110000 : 11'b10001110010;
											assign node4417 = (inp[3]) ? 11'b00101100010 : 11'b00001100110;
							assign node4420 = (inp[0]) ? node4462 : node4421;
								assign node4421 = (inp[11]) ? node4437 : node4422;
									assign node4422 = (inp[4]) ? node4430 : node4423;
										assign node4423 = (inp[10]) ? node4425 : 11'b10100110100;
											assign node4425 = (inp[3]) ? node4427 : 11'b10010100100;
												assign node4427 = (inp[9]) ? 11'b00110100110 : 11'b00010110110;
										assign node4430 = (inp[9]) ? node4434 : node4431;
											assign node4431 = (inp[3]) ? 11'b00100110000 : 11'b00100110110;
											assign node4434 = (inp[10]) ? 11'b10101110010 : 11'b10111100010;
									assign node4437 = (inp[4]) ? node4449 : node4438;
										assign node4438 = (inp[9]) ? node4442 : node4439;
											assign node4439 = (inp[3]) ? 11'b10001100000 : 11'b00111110000;
											assign node4442 = (inp[3]) ? node4446 : node4443;
												assign node4443 = (inp[10]) ? 11'b10001100110 : 11'b00001100010;
												assign node4446 = (inp[10]) ? 11'b00101100100 : 11'b10111110110;
										assign node4449 = (inp[3]) ? node4455 : node4450;
											assign node4450 = (inp[10]) ? 11'b10100100110 : node4451;
												assign node4451 = (inp[9]) ? 11'b00100100110 : 11'b00111110100;
											assign node4455 = (inp[10]) ? node4459 : node4456;
												assign node4456 = (inp[9]) ? 11'b10010100000 : 11'b10001110100;
												assign node4459 = (inp[9]) ? 11'b00000100000 : 11'b00010100010;
								assign node4462 = (inp[3]) ? node4480 : node4463;
									assign node4463 = (inp[9]) ? node4469 : node4464;
										assign node4464 = (inp[10]) ? 11'b00010110100 : node4465;
											assign node4465 = (inp[4]) ? 11'b00101110000 : 11'b00011110000;
										assign node4469 = (inp[10]) ? node4475 : node4470;
											assign node4470 = (inp[4]) ? node4472 : 11'b00010100100;
												assign node4472 = (inp[11]) ? 11'b00110100100 : 11'b00100110100;
											assign node4475 = (inp[4]) ? 11'b00111110010 : node4476;
												assign node4476 = (inp[11]) ? 11'b00111100000 : 11'b00100110000;
									assign node4480 = (inp[9]) ? node4490 : node4481;
										assign node4481 = (inp[10]) ? node4485 : node4482;
											assign node4482 = (inp[11]) ? 11'b00111100000 : 11'b00110100010;
											assign node4485 = (inp[4]) ? node4487 : 11'b00000100010;
												assign node4487 = (inp[11]) ? 11'b00010100010 : 11'b00110100000;
										assign node4490 = (inp[4]) ? node4494 : node4491;
											assign node4491 = (inp[10]) ? 11'b00001100000 : 11'b00001110010;
											assign node4494 = (inp[11]) ? 11'b00000100000 : 11'b00001100010;
						assign node4497 = (inp[11]) ? node4589 : node4498;
							assign node4498 = (inp[4]) ? node4544 : node4499;
								assign node4499 = (inp[5]) ? node4523 : node4500;
									assign node4500 = (inp[3]) ? node4514 : node4501;
										assign node4501 = (inp[9]) ? node4509 : node4502;
											assign node4502 = (inp[10]) ? node4506 : node4503;
												assign node4503 = (inp[0]) ? 11'b00100100010 : 11'b00110100010;
												assign node4506 = (inp[0]) ? 11'b00100100110 : 11'b10100100010;
											assign node4509 = (inp[10]) ? 11'b00111010010 : node4510;
												assign node4510 = (inp[0]) ? 11'b00110100100 : 11'b00100100000;
										assign node4514 = (inp[0]) ? node4520 : node4515;
											assign node4515 = (inp[10]) ? 11'b00001010110 : node4516;
												assign node4516 = (inp[9]) ? 11'b10010100100 : 11'b10000100010;
											assign node4520 = (inp[10]) ? 11'b00010100000 : 11'b00000110000;
									assign node4523 = (inp[10]) ? node4537 : node4524;
										assign node4524 = (inp[9]) ? node4530 : node4525;
											assign node4525 = (inp[0]) ? 11'b00100000000 : node4526;
												assign node4526 = (inp[3]) ? 11'b10100010000 : 11'b00110010000;
											assign node4530 = (inp[3]) ? node4534 : node4531;
												assign node4531 = (inp[0]) ? 11'b00101000110 : 11'b00101010010;
												assign node4534 = (inp[0]) ? 11'b00111010000 : 11'b10111010100;
										assign node4537 = (inp[9]) ? 11'b00011000100 : node4538;
											assign node4538 = (inp[0]) ? 11'b00001000110 : node4539;
												assign node4539 = (inp[3]) ? 11'b00001010110 : 11'b10011010010;
								assign node4544 = (inp[3]) ? node4570 : node4545;
									assign node4545 = (inp[10]) ? node4561 : node4546;
										assign node4546 = (inp[9]) ? node4554 : node4547;
											assign node4547 = (inp[0]) ? node4551 : node4548;
												assign node4548 = (inp[5]) ? 11'b00001010100 : 11'b00011000110;
												assign node4551 = (inp[5]) ? 11'b00001000000 : 11'b00101000010;
											assign node4554 = (inp[5]) ? node4558 : node4555;
												assign node4555 = (inp[0]) ? 11'b00001010100 : 11'b00001000100;
												assign node4558 = (inp[0]) ? 11'b00011010100 : 11'b00001010110;
										assign node4561 = (inp[0]) ? node4565 : node4562;
											assign node4562 = (inp[5]) ? 11'b10001010000 : 11'b10011010100;
											assign node4565 = (inp[9]) ? node4567 : 11'b00111010110;
												assign node4567 = (inp[5]) ? 11'b00011010000 : 11'b00011010010;
									assign node4570 = (inp[0]) ? node4580 : node4571;
										assign node4571 = (inp[10]) ? node4577 : node4572;
											assign node4572 = (inp[9]) ? 11'b10111010010 : node4573;
												assign node4573 = (inp[5]) ? 11'b10111010110 : 11'b10101000110;
											assign node4577 = (inp[5]) ? 11'b00111010010 : 11'b00111000000;
										assign node4580 = (inp[9]) ? node4586 : node4581;
											assign node4581 = (inp[5]) ? 11'b00101010010 : node4582;
												assign node4582 = (inp[10]) ? 11'b00111000000 : 11'b00011010000;
											assign node4586 = (inp[5]) ? 11'b00001000000 : 11'b00001000010;
							assign node4589 = (inp[3]) ? node4631 : node4590;
								assign node4590 = (inp[4]) ? node4610 : node4591;
									assign node4591 = (inp[9]) ? node4599 : node4592;
										assign node4592 = (inp[5]) ? node4594 : 11'b00111010000;
											assign node4594 = (inp[10]) ? node4596 : 11'b00110010010;
												assign node4596 = (inp[0]) ? 11'b00110010110 : 11'b10110010010;
										assign node4599 = (inp[5]) ? node4607 : node4600;
											assign node4600 = (inp[10]) ? node4604 : node4601;
												assign node4601 = (inp[0]) ? 11'b00000010110 : 11'b00010010010;
												assign node4604 = (inp[0]) ? 11'b00100000010 : 11'b10100010110;
											assign node4607 = (inp[10]) ? 11'b10010000100 : 11'b00010010100;
									assign node4610 = (inp[10]) ? node4624 : node4611;
										assign node4611 = (inp[0]) ? node4619 : node4612;
											assign node4612 = (inp[9]) ? node4616 : node4613;
												assign node4613 = (inp[5]) ? 11'b00010010110 : 11'b00000000100;
												assign node4616 = (inp[5]) ? 11'b00010000100 : 11'b00110010110;
											assign node4619 = (inp[9]) ? 11'b00110000110 : node4620;
												assign node4620 = (inp[5]) ? 11'b00010010010 : 11'b00110010000;
										assign node4624 = (inp[9]) ? node4628 : node4625;
											assign node4625 = (inp[5]) ? 11'b00010000110 : 11'b10000010100;
											assign node4628 = (inp[0]) ? 11'b00010000000 : 11'b10010000000;
								assign node4631 = (inp[0]) ? node4649 : node4632;
									assign node4632 = (inp[10]) ? node4640 : node4633;
										assign node4633 = (inp[4]) ? node4635 : 11'b10100000010;
											assign node4635 = (inp[9]) ? node4637 : 11'b10000010110;
												assign node4637 = (inp[5]) ? 11'b10000000000 : 11'b10100010010;
										assign node4640 = (inp[5]) ? node4644 : node4641;
											assign node4641 = (inp[9]) ? 11'b00010010100 : 11'b00010010010;
											assign node4644 = (inp[4]) ? 11'b00000000010 : node4645;
												assign node4645 = (inp[9]) ? 11'b00000000100 : 11'b00100000110;
									assign node4649 = (inp[10]) ? node4665 : node4650;
										assign node4650 = (inp[5]) ? node4658 : node4651;
											assign node4651 = (inp[9]) ? node4655 : node4652;
												assign node4652 = (inp[4]) ? 11'b00100010000 : 11'b00001000000;
												assign node4655 = (inp[4]) ? 11'b00100000010 : 11'b00110010010;
											assign node4658 = (inp[9]) ? node4662 : node4659;
												assign node4659 = (inp[4]) ? 11'b00000010010 : 11'b00100000010;
												assign node4662 = (inp[4]) ? 11'b00000000000 : 11'b00000010000;
										assign node4665 = (inp[9]) ? 11'b00000000000 : node4666;
											assign node4666 = (inp[4]) ? 11'b00000000010 : 11'b00110000010;
				assign node4670 = (inp[2]) ? node4982 : node4671;
					assign node4671 = (inp[8]) ? node4833 : node4672;
						assign node4672 = (inp[11]) ? node4746 : node4673;
							assign node4673 = (inp[0]) ? node4713 : node4674;
								assign node4674 = (inp[10]) ? node4694 : node4675;
									assign node4675 = (inp[5]) ? node4685 : node4676;
										assign node4676 = (inp[9]) ? node4682 : node4677;
											assign node4677 = (inp[3]) ? node4679 : 11'b00011100110;
												assign node4679 = (inp[4]) ? 11'b10001100110 : 11'b10001100010;
											assign node4682 = (inp[4]) ? 11'b10101110000 : 11'b10001100100;
										assign node4685 = (inp[9]) ? 11'b10011110110 : node4686;
											assign node4686 = (inp[4]) ? node4690 : node4687;
												assign node4687 = (inp[3]) ? 11'b10000110000 : 11'b00010110000;
												assign node4690 = (inp[3]) ? 11'b10111110100 : 11'b00001110100;
									assign node4694 = (inp[3]) ? node4704 : node4695;
										assign node4695 = (inp[9]) ? node4701 : node4696;
											assign node4696 = (inp[4]) ? 11'b10011110110 : node4697;
												assign node4697 = (inp[5]) ? 11'b10111110010 : 11'b10011100010;
											assign node4701 = (inp[4]) ? 11'b10111100000 : 11'b10101100110;
										assign node4704 = (inp[4]) ? node4708 : node4705;
											assign node4705 = (inp[9]) ? 11'b00001110100 : 11'b00001100110;
											assign node4708 = (inp[5]) ? 11'b00101100010 : node4709;
												assign node4709 = (inp[9]) ? 11'b00101110000 : 11'b00101100010;
								assign node4713 = (inp[3]) ? node4731 : node4714;
									assign node4714 = (inp[9]) ? node4720 : node4715;
										assign node4715 = (inp[5]) ? 11'b00001110100 : node4716;
											assign node4716 = (inp[10]) ? 11'b00011100110 : 11'b00011100010;
										assign node4720 = (inp[10]) ? node4724 : node4721;
											assign node4721 = (inp[4]) ? 11'b00111110100 : 11'b00011100110;
											assign node4724 = (inp[4]) ? node4728 : node4725;
												assign node4725 = (inp[5]) ? 11'b00111110000 : 11'b00011110000;
												assign node4728 = (inp[5]) ? 11'b00111110010 : 11'b00111110000;
									assign node4731 = (inp[4]) ? node4737 : node4732;
										assign node4732 = (inp[9]) ? node4734 : 11'b00001100010;
											assign node4734 = (inp[5]) ? 11'b00101110010 : 11'b00001100000;
										assign node4737 = (inp[10]) ? node4741 : node4738;
											assign node4738 = (inp[9]) ? 11'b00101100000 : 11'b00111110000;
											assign node4741 = (inp[9]) ? 11'b00001100010 : node4742;
												assign node4742 = (inp[5]) ? 11'b00111100010 : 11'b00101100010;
							assign node4746 = (inp[0]) ? node4792 : node4747;
								assign node4747 = (inp[4]) ? node4771 : node4748;
									assign node4748 = (inp[3]) ? node4762 : node4749;
										assign node4749 = (inp[10]) ? node4757 : node4750;
											assign node4750 = (inp[9]) ? node4754 : node4751;
												assign node4751 = (inp[5]) ? 11'b00001110010 : 11'b00001100000;
												assign node4754 = (inp[5]) ? 11'b00101100000 : 11'b00100110010;
											assign node4757 = (inp[5]) ? 11'b10101110000 : node4758;
												assign node4758 = (inp[9]) ? 11'b10100110100 : 11'b10000100010;
										assign node4762 = (inp[10]) ? node4768 : node4763;
											assign node4763 = (inp[5]) ? node4765 : 11'b10110100100;
												assign node4765 = (inp[9]) ? 11'b10001110100 : 11'b10111100000;
											assign node4768 = (inp[5]) ? 11'b00000100110 : 11'b00010110100;
									assign node4771 = (inp[9]) ? node4781 : node4772;
										assign node4772 = (inp[3]) ? node4776 : node4773;
											assign node4773 = (inp[5]) ? 11'b10000100110 : 11'b10100110110;
											assign node4776 = (inp[10]) ? 11'b00110100000 : node4777;
												assign node4777 = (inp[5]) ? 11'b10100110110 : 11'b10110100110;
										assign node4781 = (inp[5]) ? node4787 : node4782;
											assign node4782 = (inp[3]) ? node4784 : 11'b00010110110;
												assign node4784 = (inp[10]) ? 11'b00100110000 : 11'b10000110010;
											assign node4787 = (inp[3]) ? node4789 : 11'b10010100000;
												assign node4789 = (inp[10]) ? 11'b00100100000 : 11'b10110100000;
								assign node4792 = (inp[9]) ? node4808 : node4793;
									assign node4793 = (inp[4]) ? node4801 : node4794;
										assign node4794 = (inp[5]) ? node4796 : 11'b00010110110;
											assign node4796 = (inp[3]) ? 11'b00101100000 : node4797;
												assign node4797 = (inp[10]) ? 11'b00001110100 : 11'b00011110000;
										assign node4801 = (inp[10]) ? 11'b00010100000 : node4802;
											assign node4802 = (inp[3]) ? node4804 : 11'b00110110010;
												assign node4804 = (inp[5]) ? 11'b00000110010 : 11'b00110110010;
									assign node4808 = (inp[10]) ? node4822 : node4809;
										assign node4809 = (inp[3]) ? node4817 : node4810;
											assign node4810 = (inp[4]) ? node4814 : node4811;
												assign node4811 = (inp[5]) ? 11'b00101110100 : 11'b00110110100;
												assign node4814 = (inp[5]) ? 11'b00100100100 : 11'b00000100110;
											assign node4817 = (inp[5]) ? node4819 : 11'b00100110000;
												assign node4819 = (inp[4]) ? 11'b00010100000 : 11'b00010110010;
										assign node4822 = (inp[3]) ? node4828 : node4823;
											assign node4823 = (inp[4]) ? 11'b00100100000 : node4824;
												assign node4824 = (inp[5]) ? 11'b00100100010 : 11'b00000100000;
											assign node4828 = (inp[4]) ? 11'b00000100000 : node4829;
												assign node4829 = (inp[5]) ? 11'b00000100010 : 11'b00010100000;
						assign node4833 = (inp[5]) ? node4917 : node4834;
							assign node4834 = (inp[11]) ? node4880 : node4835;
								assign node4835 = (inp[4]) ? node4859 : node4836;
									assign node4836 = (inp[9]) ? node4848 : node4837;
										assign node4837 = (inp[10]) ? node4845 : node4838;
											assign node4838 = (inp[3]) ? node4842 : node4839;
												assign node4839 = (inp[0]) ? 11'b00110100010 : 11'b00010100010;
												assign node4842 = (inp[0]) ? 11'b00000100010 : 11'b10100100010;
											assign node4845 = (inp[0]) ? 11'b00010100010 : 11'b00110100110;
										assign node4848 = (inp[0]) ? node4854 : node4849;
											assign node4849 = (inp[3]) ? 11'b10110100100 : node4850;
												assign node4850 = (inp[10]) ? 11'b10010110100 : 11'b00000100010;
											assign node4854 = (inp[3]) ? 11'b00010110000 : node4855;
												assign node4855 = (inp[10]) ? 11'b00100110000 : 11'b00100100110;
									assign node4859 = (inp[9]) ? node4869 : node4860;
										assign node4860 = (inp[0]) ? node4864 : node4861;
											assign node4861 = (inp[10]) ? 11'b10100110100 : 11'b00110100100;
											assign node4864 = (inp[10]) ? node4866 : 11'b00000110000;
												assign node4866 = (inp[3]) ? 11'b00111000010 : 11'b00111010110;
										assign node4869 = (inp[10]) ? node4877 : node4870;
											assign node4870 = (inp[3]) ? node4874 : node4871;
												assign node4871 = (inp[0]) ? 11'b00001010110 : 11'b00101000110;
												assign node4874 = (inp[0]) ? 11'b00111000010 : 11'b10001010010;
											assign node4877 = (inp[0]) ? 11'b00011010010 : 11'b10011000010;
								assign node4880 = (inp[0]) ? node4900 : node4881;
									assign node4881 = (inp[9]) ? node4889 : node4882;
										assign node4882 = (inp[4]) ? node4886 : node4883;
											assign node4883 = (inp[3]) ? 11'b00001010100 : 11'b00001000010;
											assign node4886 = (inp[10]) ? 11'b10111010110 : 11'b10001000110;
										assign node4889 = (inp[4]) ? node4895 : node4890;
											assign node4890 = (inp[3]) ? node4892 : 11'b00111010000;
												assign node4892 = (inp[10]) ? 11'b00111010110 : 11'b10101000100;
											assign node4895 = (inp[10]) ? 11'b10101010000 : node4896;
												assign node4896 = (inp[3]) ? 11'b10011010000 : 11'b00001010110;
									assign node4900 = (inp[10]) ? node4910 : node4901;
										assign node4901 = (inp[3]) ? node4907 : node4902;
											assign node4902 = (inp[9]) ? node4904 : 11'b00111010000;
												assign node4904 = (inp[4]) ? 11'b00111000100 : 11'b00011010100;
											assign node4907 = (inp[9]) ? 11'b00111000000 : 11'b00011000000;
										assign node4910 = (inp[9]) ? node4914 : node4911;
											assign node4911 = (inp[4]) ? 11'b00011000110 : 11'b00101010100;
											assign node4914 = (inp[4]) ? 11'b00001000000 : 11'b00111000010;
							assign node4917 = (inp[4]) ? node4949 : node4918;
								assign node4918 = (inp[9]) ? node4932 : node4919;
									assign node4919 = (inp[10]) ? node4929 : node4920;
										assign node4920 = (inp[11]) ? node4924 : node4921;
											assign node4921 = (inp[0]) ? 11'b00101000000 : 11'b10011010000;
											assign node4924 = (inp[3]) ? 11'b10010000010 : node4925;
												assign node4925 = (inp[0]) ? 11'b00110010010 : 11'b00000010000;
										assign node4929 = (inp[3]) ? 11'b00110010110 : 11'b00100010110;
									assign node4932 = (inp[0]) ? node4940 : node4933;
										assign node4933 = (inp[10]) ? node4935 : 11'b00000000010;
											assign node4935 = (inp[11]) ? node4937 : 11'b00110000110;
												assign node4937 = (inp[3]) ? 11'b00100000110 : 11'b10100000110;
										assign node4940 = (inp[10]) ? node4944 : node4941;
											assign node4941 = (inp[3]) ? 11'b00100010010 : 11'b00100000110;
											assign node4944 = (inp[3]) ? node4946 : 11'b00010010010;
												assign node4946 = (inp[11]) ? 11'b00000000010 : 11'b00010000010;
								assign node4949 = (inp[0]) ? node4967 : node4950;
									assign node4950 = (inp[9]) ? node4960 : node4951;
										assign node4951 = (inp[11]) ? node4955 : node4952;
											assign node4952 = (inp[3]) ? 11'b10000010110 : 11'b10010000100;
											assign node4955 = (inp[10]) ? 11'b00100000000 : node4956;
												assign node4956 = (inp[3]) ? 11'b10110010100 : 11'b00110010100;
										assign node4960 = (inp[10]) ? node4964 : node4961;
											assign node4961 = (inp[3]) ? 11'b10110000000 : 11'b00110000100;
											assign node4964 = (inp[3]) ? 11'b00100000000 : 11'b10100000000;
									assign node4967 = (inp[10]) ? node4977 : node4968;
										assign node4968 = (inp[9]) ? 11'b00010000000 : node4969;
											assign node4969 = (inp[3]) ? node4973 : node4970;
												assign node4970 = (inp[11]) ? 11'b00010010000 : 11'b00000000010;
												assign node4973 = (inp[11]) ? 11'b00010010000 : 11'b00110010000;
										assign node4977 = (inp[11]) ? 11'b00000000100 : node4978;
											assign node4978 = (inp[3]) ? 11'b00100000000 : 11'b00110010100;
					assign node4982 = (inp[8]) ? node5142 : node4983;
						assign node4983 = (inp[5]) ? node5059 : node4984;
							assign node4984 = (inp[4]) ? node5024 : node4985;
								assign node4985 = (inp[0]) ? node5007 : node4986;
									assign node4986 = (inp[11]) ? node4994 : node4987;
										assign node4987 = (inp[10]) ? 11'b00101000110 : node4988;
											assign node4988 = (inp[3]) ? node4990 : 11'b00111000010;
												assign node4990 = (inp[9]) ? 11'b10111000110 : 11'b10111000010;
										assign node4994 = (inp[10]) ? node5002 : node4995;
											assign node4995 = (inp[9]) ? node4999 : node4996;
												assign node4996 = (inp[3]) ? 11'b10111010010 : 11'b00101000000;
												assign node4999 = (inp[3]) ? 11'b10001000110 : 11'b00001010010;
											assign node5002 = (inp[3]) ? node5004 : 11'b10011010110;
												assign node5004 = (inp[9]) ? 11'b00111010110 : 11'b00101010110;
									assign node5007 = (inp[3]) ? node5015 : node5008;
										assign node5008 = (inp[10]) ? node5010 : 11'b00101010110;
											assign node5010 = (inp[9]) ? 11'b00011000010 : node5011;
												assign node5011 = (inp[11]) ? 11'b00011010110 : 11'b00001000110;
										assign node5015 = (inp[10]) ? node5019 : node5016;
											assign node5016 = (inp[9]) ? 11'b00111010010 : 11'b00011000010;
											assign node5019 = (inp[9]) ? node5021 : 11'b00101000010;
												assign node5021 = (inp[11]) ? 11'b00011000010 : 11'b00001000010;
								assign node5024 = (inp[9]) ? node5040 : node5025;
									assign node5025 = (inp[10]) ? node5033 : node5026;
										assign node5026 = (inp[0]) ? node5030 : node5027;
											assign node5027 = (inp[3]) ? 11'b10001000110 : 11'b00101000110;
											assign node5030 = (inp[3]) ? 11'b00101010010 : 11'b00001010010;
										assign node5033 = (inp[3]) ? node5037 : node5034;
											assign node5034 = (inp[0]) ? 11'b00001010100 : 11'b10001010110;
											assign node5037 = (inp[0]) ? 11'b00011000000 : 11'b00001000000;
									assign node5040 = (inp[10]) ? node5048 : node5041;
										assign node5041 = (inp[3]) ? node5043 : 11'b00111010100;
											assign node5043 = (inp[0]) ? 11'b00111000000 : node5044;
												assign node5044 = (inp[11]) ? 11'b10101010000 : 11'b10011010000;
										assign node5048 = (inp[0]) ? node5054 : node5049;
											assign node5049 = (inp[3]) ? 11'b00001010000 : node5050;
												assign node5050 = (inp[11]) ? 11'b10001010000 : 11'b10011000000;
											assign node5054 = (inp[3]) ? 11'b00001000000 : node5055;
												assign node5055 = (inp[11]) ? 11'b00101000000 : 11'b00101010000;
							assign node5059 = (inp[11]) ? node5101 : node5060;
								assign node5060 = (inp[9]) ? node5080 : node5061;
									assign node5061 = (inp[4]) ? node5073 : node5062;
										assign node5062 = (inp[10]) ? node5068 : node5063;
											assign node5063 = (inp[0]) ? 11'b00011000000 : node5064;
												assign node5064 = (inp[3]) ? 11'b10111010000 : 11'b00111010000;
											assign node5068 = (inp[0]) ? node5070 : 11'b00001010100;
												assign node5070 = (inp[3]) ? 11'b00001000000 : 11'b00101000100;
										assign node5073 = (inp[10]) ? node5077 : node5074;
											assign node5074 = (inp[3]) ? 11'b10000010110 : 11'b00100010110;
											assign node5077 = (inp[0]) ? 11'b00000010110 : 11'b00110010010;
									assign node5080 = (inp[0]) ? node5094 : node5081;
										assign node5081 = (inp[4]) ? node5087 : node5082;
											assign node5082 = (inp[3]) ? node5084 : 11'b10010000110;
												assign node5084 = (inp[10]) ? 11'b00110000110 : 11'b10110010110;
											assign node5087 = (inp[10]) ? node5091 : node5088;
												assign node5088 = (inp[3]) ? 11'b10110000010 : 11'b00010010110;
												assign node5091 = (inp[3]) ? 11'b00000000010 : 11'b10100010010;
										assign node5094 = (inp[4]) ? 11'b00100010010 : node5095;
											assign node5095 = (inp[3]) ? node5097 : 11'b00110010010;
												assign node5097 = (inp[10]) ? 11'b00010000010 : 11'b00110010010;
								assign node5101 = (inp[9]) ? node5121 : node5102;
									assign node5102 = (inp[0]) ? node5112 : node5103;
										assign node5103 = (inp[10]) ? node5105 : 11'b10000000010;
											assign node5105 = (inp[3]) ? node5109 : node5106;
												assign node5106 = (inp[4]) ? 11'b10110000100 : 11'b10010010000;
												assign node5109 = (inp[4]) ? 11'b00010000000 : 11'b00110000100;
										assign node5112 = (inp[3]) ? node5118 : node5113;
											assign node5113 = (inp[10]) ? node5115 : 11'b00110010000;
												assign node5115 = (inp[4]) ? 11'b00110000100 : 11'b00010010100;
											assign node5118 = (inp[10]) ? 11'b00010000000 : 11'b00010010000;
									assign node5121 = (inp[0]) ? node5135 : node5122;
										assign node5122 = (inp[4]) ? node5130 : node5123;
											assign node5123 = (inp[3]) ? node5127 : node5124;
												assign node5124 = (inp[10]) ? 11'b10000000100 : 11'b00010000000;
												assign node5127 = (inp[10]) ? 11'b00100000100 : 11'b10100010100;
											assign node5130 = (inp[3]) ? node5132 : 11'b00100000100;
												assign node5132 = (inp[10]) ? 11'b00000000000 : 11'b10000000000;
										assign node5135 = (inp[10]) ? node5139 : node5136;
											assign node5136 = (inp[4]) ? 11'b00100000100 : 11'b00100010100;
											assign node5139 = (inp[4]) ? 11'b00100000000 : 11'b00000000000;
						assign node5142 = (inp[5]) ? node5210 : node5143;
							assign node5143 = (inp[11]) ? node5177 : node5144;
								assign node5144 = (inp[9]) ? node5162 : node5145;
									assign node5145 = (inp[0]) ? node5155 : node5146;
										assign node5146 = (inp[3]) ? node5150 : node5147;
											assign node5147 = (inp[4]) ? 11'b00000000110 : 11'b00110000010;
											assign node5150 = (inp[4]) ? node5152 : 11'b00010000110;
												assign node5152 = (inp[10]) ? 11'b00110000010 : 11'b10110000110;
										assign node5155 = (inp[4]) ? node5157 : 11'b00010000010;
											assign node5157 = (inp[3]) ? node5159 : 11'b00110000010;
												assign node5159 = (inp[10]) ? 11'b00110000010 : 11'b00010010010;
									assign node5162 = (inp[10]) ? node5172 : node5163;
										assign node5163 = (inp[3]) ? node5167 : node5164;
											assign node5164 = (inp[0]) ? 11'b00010010110 : 11'b00100000010;
											assign node5167 = (inp[4]) ? node5169 : 11'b10000000110;
												assign node5169 = (inp[0]) ? 11'b00100000010 : 11'b10100010010;
										assign node5172 = (inp[3]) ? node5174 : 11'b00100010010;
											assign node5174 = (inp[0]) ? 11'b00000000010 : 11'b00000010010;
								assign node5177 = (inp[4]) ? node5195 : node5178;
									assign node5178 = (inp[9]) ? node5190 : node5179;
										assign node5179 = (inp[10]) ? node5185 : node5180;
											assign node5180 = (inp[3]) ? 11'b00000000010 : node5181;
												assign node5181 = (inp[0]) ? 11'b00100010010 : 11'b00100000010;
											assign node5185 = (inp[0]) ? node5187 : 11'b10000000010;
												assign node5187 = (inp[3]) ? 11'b00110000000 : 11'b00110010100;
										assign node5190 = (inp[0]) ? 11'b00110010000 : node5191;
											assign node5191 = (inp[3]) ? 11'b00010010100 : 11'b00010010000;
									assign node5195 = (inp[10]) ? node5203 : node5196;
										assign node5196 = (inp[3]) ? node5198 : 11'b00010000100;
											assign node5198 = (inp[0]) ? 11'b00100010000 : node5199;
												assign node5199 = (inp[9]) ? 11'b10100010000 : 11'b10100000100;
										assign node5203 = (inp[3]) ? node5207 : node5204;
											assign node5204 = (inp[9]) ? 11'b10000010000 : 11'b10000010100;
											assign node5207 = (inp[0]) ? 11'b00000000000 : 11'b00000010000;
							assign node5210 = (inp[4]) ? node5254 : node5211;
								assign node5211 = (inp[11]) ? node5235 : node5212;
									assign node5212 = (inp[10]) ? node5226 : node5213;
										assign node5213 = (inp[0]) ? node5219 : node5214;
											assign node5214 = (inp[9]) ? 11'b10110010100 : node5215;
												assign node5215 = (inp[3]) ? 11'b10110010000 : 11'b00110010000;
											assign node5219 = (inp[3]) ? node5223 : node5220;
												assign node5220 = (inp[9]) ? 11'b00110000100 : 11'b00110000000;
												assign node5223 = (inp[9]) ? 11'b00110010000 : 11'b00110000000;
										assign node5226 = (inp[0]) ? node5230 : node5227;
											assign node5227 = (inp[9]) ? 11'b00010000100 : 11'b00010010100;
											assign node5230 = (inp[9]) ? 11'b00010010000 : node5231;
												assign node5231 = (inp[3]) ? 11'b00010000000 : 11'b00010000100;
									assign node5235 = (inp[9]) ? node5247 : node5236;
										assign node5236 = (inp[3]) ? node5244 : node5237;
											assign node5237 = (inp[0]) ? node5241 : node5238;
												assign node5238 = (inp[10]) ? 11'b10100010000 : 11'b00100010000;
												assign node5241 = (inp[10]) ? 11'b00100010100 : 11'b00100010000;
											assign node5244 = (inp[0]) ? 11'b00100000000 : 11'b00100000100;
										assign node5247 = (inp[0]) ? node5249 : 11'b00100000000;
											assign node5249 = (inp[10]) ? 11'b00000000000 : node5250;
												assign node5250 = (inp[3]) ? 11'b00000010000 : 11'b00000010100;
								assign node5254 = (inp[0]) ? node5268 : node5255;
									assign node5255 = (inp[9]) ? node5263 : node5256;
										assign node5256 = (inp[10]) ? node5260 : node5257;
											assign node5257 = (inp[3]) ? 11'b10100010100 : 11'b00010010100;
											assign node5260 = (inp[11]) ? 11'b10000000100 : 11'b10100000100;
										assign node5263 = (inp[3]) ? node5265 : 11'b10000010000;
											assign node5265 = (inp[10]) ? 11'b00000000000 : 11'b10000000000;
									assign node5268 = (inp[10]) ? node5280 : node5269;
										assign node5269 = (inp[9]) ? node5277 : node5270;
											assign node5270 = (inp[3]) ? node5274 : node5271;
												assign node5271 = (inp[11]) ? 11'b00000010000 : 11'b00010000000;
												assign node5274 = (inp[11]) ? 11'b00000010000 : 11'b00100010000;
											assign node5277 = (inp[3]) ? 11'b00000000000 : 11'b00000010100;
										assign node5280 = (inp[11]) ? node5282 : 11'b00000010000;
											assign node5282 = (inp[9]) ? 11'b00000000000 : 11'b00000000100;

endmodule