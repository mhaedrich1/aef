module dtc_split25_bm82 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node114;

	assign outp = (inp[0]) ? node56 : node1;
		assign node1 = (inp[3]) ? node31 : node2;
			assign node2 = (inp[6]) ? node16 : node3;
				assign node3 = (inp[7]) ? node9 : node4;
					assign node4 = (inp[4]) ? node6 : 3'b001;
						assign node6 = (inp[1]) ? 3'b101 : 3'b111;
					assign node9 = (inp[1]) ? node13 : node10;
						assign node10 = (inp[4]) ? 3'b111 : 3'b111;
						assign node13 = (inp[8]) ? 3'b101 : 3'b001;
				assign node16 = (inp[1]) ? node24 : node17;
					assign node17 = (inp[11]) ? node21 : node18;
						assign node18 = (inp[7]) ? 3'b110 : 3'b001;
						assign node21 = (inp[10]) ? 3'b011 : 3'b101;
					assign node24 = (inp[9]) ? node28 : node25;
						assign node25 = (inp[4]) ? 3'b100 : 3'b000;
						assign node28 = (inp[4]) ? 3'b001 : 3'b010;
			assign node31 = (inp[6]) ? node41 : node32;
				assign node32 = (inp[9]) ? 3'b111 : node33;
					assign node33 = (inp[1]) ? node37 : node34;
						assign node34 = (inp[8]) ? 3'b111 : 3'b111;
						assign node37 = (inp[7]) ? 3'b111 : 3'b111;
				assign node41 = (inp[9]) ? node49 : node42;
					assign node42 = (inp[1]) ? node46 : node43;
						assign node43 = (inp[7]) ? 3'b101 : 3'b111;
						assign node46 = (inp[7]) ? 3'b110 : 3'b101;
					assign node49 = (inp[1]) ? node53 : node50;
						assign node50 = (inp[11]) ? 3'b111 : 3'b111;
						assign node53 = (inp[7]) ? 3'b101 : 3'b111;
		assign node56 = (inp[6]) ? node88 : node57;
			assign node57 = (inp[3]) ? node73 : node58;
				assign node58 = (inp[1]) ? node66 : node59;
					assign node59 = (inp[4]) ? node63 : node60;
						assign node60 = (inp[9]) ? 3'b000 : 3'b100;
						assign node63 = (inp[7]) ? 3'b100 : 3'b011;
					assign node66 = (inp[7]) ? node70 : node67;
						assign node67 = (inp[4]) ? 3'b110 : 3'b010;
						assign node70 = (inp[9]) ? 3'b100 : 3'b000;
				assign node73 = (inp[7]) ? node81 : node74;
					assign node74 = (inp[9]) ? node78 : node75;
						assign node75 = (inp[1]) ? 3'b101 : 3'b011;
						assign node78 = (inp[1]) ? 3'b111 : 3'b111;
					assign node81 = (inp[1]) ? node85 : node82;
						assign node82 = (inp[9]) ? 3'b011 : 3'b001;
						assign node85 = (inp[10]) ? 3'b011 : 3'b110;
			assign node88 = (inp[3]) ? node102 : node89;
				assign node89 = (inp[9]) ? node95 : node90;
					assign node90 = (inp[4]) ? node92 : 3'b000;
						assign node92 = (inp[5]) ? 3'b000 : 3'b000;
					assign node95 = (inp[1]) ? node99 : node96;
						assign node96 = (inp[7]) ? 3'b000 : 3'b010;
						assign node99 = (inp[7]) ? 3'b000 : 3'b000;
				assign node102 = (inp[9]) ? node110 : node103;
					assign node103 = (inp[7]) ? node107 : node104;
						assign node104 = (inp[1]) ? 3'b000 : 3'b110;
						assign node107 = (inp[1]) ? 3'b000 : 3'b000;
					assign node110 = (inp[1]) ? node114 : node111;
						assign node111 = (inp[7]) ? 3'b110 : 3'b101;
						assign node114 = (inp[7]) ? 3'b000 : 3'b010;

endmodule