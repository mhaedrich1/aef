module dtc_split75_bm96 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node212;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node224;
	wire [3-1:0] node227;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node245;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node252;
	wire [3-1:0] node254;
	wire [3-1:0] node255;

	assign outp = (inp[7]) ? node18 : node1;
		assign node1 = (inp[6]) ? node3 : 3'b000;
			assign node3 = (inp[3]) ? node5 : 3'b000;
				assign node5 = (inp[1]) ? node7 : 3'b000;
					assign node7 = (inp[2]) ? node9 : 3'b000;
						assign node9 = (inp[8]) ? node11 : 3'b000;
							assign node11 = (inp[9]) ? 3'b000 : node12;
								assign node12 = (inp[10]) ? 3'b000 : node13;
									assign node13 = (inp[4]) ? 3'b100 : 3'b000;
		assign node18 = (inp[6]) ? node20 : 3'b000;
			assign node20 = (inp[3]) ? node122 : node21;
				assign node21 = (inp[4]) ? node33 : node22;
					assign node22 = (inp[9]) ? node24 : 3'b011;
						assign node24 = (inp[1]) ? 3'b011 : node25;
							assign node25 = (inp[5]) ? node29 : node26;
								assign node26 = (inp[10]) ? 3'b011 : 3'b111;
								assign node29 = (inp[10]) ? 3'b101 : 3'b011;
					assign node33 = (inp[1]) ? node93 : node34;
						assign node34 = (inp[0]) ? node66 : node35;
							assign node35 = (inp[9]) ? node45 : node36;
								assign node36 = (inp[11]) ? 3'b010 : node37;
									assign node37 = (inp[10]) ? node41 : node38;
										assign node38 = (inp[8]) ? 3'b010 : 3'b001;
										assign node41 = (inp[8]) ? 3'b001 : 3'b010;
								assign node45 = (inp[5]) ? node51 : node46;
									assign node46 = (inp[11]) ? 3'b001 : node47;
										assign node47 = (inp[10]) ? 3'b001 : 3'b010;
									assign node51 = (inp[2]) ? node59 : node52;
										assign node52 = (inp[10]) ? node56 : node53;
											assign node53 = (inp[11]) ? 3'b001 : 3'b010;
											assign node56 = (inp[11]) ? 3'b010 : 3'b001;
										assign node59 = (inp[8]) ? node63 : node60;
											assign node60 = (inp[11]) ? 3'b000 : 3'b001;
											assign node63 = (inp[10]) ? 3'b000 : 3'b000;
							assign node66 = (inp[9]) ? node76 : node67;
								assign node67 = (inp[10]) ? node69 : 3'b001;
									assign node69 = (inp[5]) ? node71 : 3'b001;
										assign node71 = (inp[11]) ? node73 : 3'b001;
											assign node73 = (inp[8]) ? 3'b010 : 3'b001;
								assign node76 = (inp[11]) ? node82 : node77;
									assign node77 = (inp[10]) ? node79 : 3'b110;
										assign node79 = (inp[5]) ? 3'b001 : 3'b101;
									assign node82 = (inp[10]) ? node88 : node83;
										assign node83 = (inp[5]) ? 3'b001 : node84;
											assign node84 = (inp[8]) ? 3'b101 : 3'b001;
										assign node88 = (inp[5]) ? node90 : 3'b001;
											assign node90 = (inp[8]) ? 3'b110 : 3'b010;
						assign node93 = (inp[9]) ? node111 : node94;
							assign node94 = (inp[0]) ? node96 : 3'b010;
								assign node96 = (inp[11]) ? node104 : node97;
									assign node97 = (inp[8]) ? node101 : node98;
										assign node98 = (inp[10]) ? 3'b001 : 3'b010;
										assign node101 = (inp[10]) ? 3'b010 : 3'b001;
									assign node104 = (inp[2]) ? node106 : 3'b001;
										assign node106 = (inp[8]) ? node108 : 3'b001;
											assign node108 = (inp[10]) ? 3'b001 : 3'b010;
							assign node111 = (inp[0]) ? 3'b010 : node112;
								assign node112 = (inp[10]) ? node114 : 3'b010;
									assign node114 = (inp[2]) ? 3'b010 : node115;
										assign node115 = (inp[8]) ? node117 : 3'b010;
											assign node117 = (inp[5]) ? 3'b000 : 3'b010;
				assign node122 = (inp[1]) ? node190 : node123;
					assign node123 = (inp[4]) ? node145 : node124;
						assign node124 = (inp[9]) ? node130 : node125;
							assign node125 = (inp[0]) ? 3'b111 : node126;
								assign node126 = (inp[10]) ? 3'b110 : 3'b111;
							assign node130 = (inp[10]) ? node138 : node131;
								assign node131 = (inp[11]) ? node135 : node132;
									assign node132 = (inp[0]) ? 3'b111 : 3'b110;
									assign node135 = (inp[0]) ? 3'b110 : 3'b111;
								assign node138 = (inp[5]) ? node142 : node139;
									assign node139 = (inp[0]) ? 3'b110 : 3'b111;
									assign node142 = (inp[0]) ? 3'b010 : 3'b011;
						assign node145 = (inp[0]) ? node171 : node146;
							assign node146 = (inp[9]) ? node162 : node147;
								assign node147 = (inp[10]) ? node157 : node148;
									assign node148 = (inp[5]) ? 3'b011 : node149;
										assign node149 = (inp[11]) ? node153 : node150;
											assign node150 = (inp[8]) ? 3'b011 : 3'b111;
											assign node153 = (inp[2]) ? 3'b011 : 3'b011;
									assign node157 = (inp[11]) ? 3'b001 : node158;
										assign node158 = (inp[8]) ? 3'b101 : 3'b001;
								assign node162 = (inp[11]) ? node166 : node163;
									assign node163 = (inp[10]) ? 3'b110 : 3'b001;
									assign node166 = (inp[10]) ? node168 : 3'b110;
										assign node168 = (inp[5]) ? 3'b010 : 3'b110;
							assign node171 = (inp[9]) ? node181 : node172;
								assign node172 = (inp[5]) ? node174 : 3'b110;
									assign node174 = (inp[10]) ? node176 : 3'b110;
										assign node176 = (inp[2]) ? node178 : 3'b110;
											assign node178 = (inp[11]) ? 3'b010 : 3'b110;
								assign node181 = (inp[11]) ? node185 : node182;
									assign node182 = (inp[10]) ? 3'b100 : 3'b010;
									assign node185 = (inp[10]) ? node187 : 3'b100;
										assign node187 = (inp[5]) ? 3'b000 : 3'b100;
					assign node190 = (inp[4]) ? node216 : node191;
						assign node191 = (inp[9]) ? node207 : node192;
							assign node192 = (inp[0]) ? node194 : 3'b100;
								assign node194 = (inp[11]) ? node200 : node195;
									assign node195 = (inp[8]) ? 3'b101 : node196;
										assign node196 = (inp[10]) ? 3'b100 : 3'b101;
									assign node200 = (inp[10]) ? 3'b100 : node201;
										assign node201 = (inp[8]) ? node203 : 3'b100;
											assign node203 = (inp[5]) ? 3'b100 : 3'b101;
							assign node207 = (inp[0]) ? 3'b100 : node208;
								assign node208 = (inp[8]) ? node210 : 3'b101;
									assign node210 = (inp[10]) ? node212 : 3'b101;
										assign node212 = (inp[11]) ? 3'b100 : 3'b101;
						assign node216 = (inp[0]) ? node234 : node217;
							assign node217 = (inp[9]) ? node227 : node218;
								assign node218 = (inp[11]) ? node220 : 3'b001;
									assign node220 = (inp[5]) ? node222 : 3'b001;
										assign node222 = (inp[10]) ? node224 : 3'b001;
											assign node224 = (inp[8]) ? 3'b000 : 3'b001;
								assign node227 = (inp[8]) ? node229 : 3'b010;
									assign node229 = (inp[5]) ? node231 : 3'b010;
										assign node231 = (inp[11]) ? 3'b100 : 3'b010;
							assign node234 = (inp[9]) ? node250 : node235;
								assign node235 = (inp[8]) ? node241 : node236;
									assign node236 = (inp[10]) ? 3'b100 : node237;
										assign node237 = (inp[11]) ? 3'b100 : 3'b010;
									assign node241 = (inp[11]) ? node245 : node242;
										assign node242 = (inp[10]) ? 3'b010 : 3'b110;
										assign node245 = (inp[2]) ? node247 : 3'b100;
											assign node247 = (inp[10]) ? 3'b100 : 3'b010;
								assign node250 = (inp[8]) ? node252 : 3'b000;
									assign node252 = (inp[2]) ? node254 : 3'b000;
										assign node254 = (inp[10]) ? 3'b000 : node255;
											assign node255 = (inp[11]) ? 3'b000 : 3'b100;

endmodule