module dtc_split66_bm24 (
	input  wire [13-1:0] inp,
	output wire [13-1:0] outp
);

	wire [13-1:0] node1;
	wire [13-1:0] node2;
	wire [13-1:0] node3;
	wire [13-1:0] node4;
	wire [13-1:0] node5;
	wire [13-1:0] node6;
	wire [13-1:0] node7;
	wire [13-1:0] node8;
	wire [13-1:0] node11;
	wire [13-1:0] node14;
	wire [13-1:0] node15;
	wire [13-1:0] node18;
	wire [13-1:0] node21;
	wire [13-1:0] node22;
	wire [13-1:0] node23;
	wire [13-1:0] node26;
	wire [13-1:0] node29;
	wire [13-1:0] node30;
	wire [13-1:0] node33;
	wire [13-1:0] node36;
	wire [13-1:0] node37;
	wire [13-1:0] node38;
	wire [13-1:0] node39;
	wire [13-1:0] node42;
	wire [13-1:0] node45;
	wire [13-1:0] node46;
	wire [13-1:0] node49;
	wire [13-1:0] node52;
	wire [13-1:0] node53;
	wire [13-1:0] node54;
	wire [13-1:0] node57;
	wire [13-1:0] node60;
	wire [13-1:0] node61;
	wire [13-1:0] node64;
	wire [13-1:0] node67;
	wire [13-1:0] node68;
	wire [13-1:0] node69;
	wire [13-1:0] node70;
	wire [13-1:0] node71;
	wire [13-1:0] node74;
	wire [13-1:0] node77;
	wire [13-1:0] node78;
	wire [13-1:0] node81;
	wire [13-1:0] node84;
	wire [13-1:0] node85;
	wire [13-1:0] node86;
	wire [13-1:0] node89;
	wire [13-1:0] node92;
	wire [13-1:0] node93;
	wire [13-1:0] node96;
	wire [13-1:0] node99;
	wire [13-1:0] node100;
	wire [13-1:0] node101;
	wire [13-1:0] node102;
	wire [13-1:0] node105;
	wire [13-1:0] node108;
	wire [13-1:0] node109;
	wire [13-1:0] node112;
	wire [13-1:0] node115;
	wire [13-1:0] node116;
	wire [13-1:0] node117;
	wire [13-1:0] node120;
	wire [13-1:0] node123;
	wire [13-1:0] node124;
	wire [13-1:0] node127;
	wire [13-1:0] node130;
	wire [13-1:0] node131;
	wire [13-1:0] node132;
	wire [13-1:0] node133;
	wire [13-1:0] node134;
	wire [13-1:0] node135;
	wire [13-1:0] node138;
	wire [13-1:0] node141;
	wire [13-1:0] node142;
	wire [13-1:0] node145;
	wire [13-1:0] node148;
	wire [13-1:0] node149;
	wire [13-1:0] node150;
	wire [13-1:0] node153;
	wire [13-1:0] node156;
	wire [13-1:0] node157;
	wire [13-1:0] node160;
	wire [13-1:0] node163;
	wire [13-1:0] node164;
	wire [13-1:0] node165;
	wire [13-1:0] node166;
	wire [13-1:0] node169;
	wire [13-1:0] node172;
	wire [13-1:0] node173;
	wire [13-1:0] node176;
	wire [13-1:0] node179;
	wire [13-1:0] node180;
	wire [13-1:0] node181;
	wire [13-1:0] node184;
	wire [13-1:0] node187;
	wire [13-1:0] node188;
	wire [13-1:0] node191;
	wire [13-1:0] node194;
	wire [13-1:0] node195;
	wire [13-1:0] node196;
	wire [13-1:0] node197;
	wire [13-1:0] node198;
	wire [13-1:0] node201;
	wire [13-1:0] node204;
	wire [13-1:0] node205;
	wire [13-1:0] node208;
	wire [13-1:0] node211;
	wire [13-1:0] node212;
	wire [13-1:0] node213;
	wire [13-1:0] node216;
	wire [13-1:0] node219;
	wire [13-1:0] node220;
	wire [13-1:0] node223;
	wire [13-1:0] node226;
	wire [13-1:0] node227;
	wire [13-1:0] node228;
	wire [13-1:0] node229;
	wire [13-1:0] node232;
	wire [13-1:0] node235;
	wire [13-1:0] node236;
	wire [13-1:0] node239;
	wire [13-1:0] node242;
	wire [13-1:0] node243;
	wire [13-1:0] node244;
	wire [13-1:0] node247;
	wire [13-1:0] node250;
	wire [13-1:0] node251;
	wire [13-1:0] node254;
	wire [13-1:0] node257;
	wire [13-1:0] node258;
	wire [13-1:0] node259;
	wire [13-1:0] node260;
	wire [13-1:0] node261;
	wire [13-1:0] node262;
	wire [13-1:0] node263;
	wire [13-1:0] node266;
	wire [13-1:0] node269;
	wire [13-1:0] node270;
	wire [13-1:0] node273;
	wire [13-1:0] node276;
	wire [13-1:0] node277;
	wire [13-1:0] node278;
	wire [13-1:0] node281;
	wire [13-1:0] node284;
	wire [13-1:0] node285;
	wire [13-1:0] node288;
	wire [13-1:0] node291;
	wire [13-1:0] node292;
	wire [13-1:0] node293;
	wire [13-1:0] node294;
	wire [13-1:0] node297;
	wire [13-1:0] node300;
	wire [13-1:0] node301;
	wire [13-1:0] node304;
	wire [13-1:0] node307;
	wire [13-1:0] node308;
	wire [13-1:0] node309;
	wire [13-1:0] node312;
	wire [13-1:0] node315;
	wire [13-1:0] node316;
	wire [13-1:0] node319;
	wire [13-1:0] node322;
	wire [13-1:0] node323;
	wire [13-1:0] node324;
	wire [13-1:0] node325;
	wire [13-1:0] node326;
	wire [13-1:0] node329;
	wire [13-1:0] node332;
	wire [13-1:0] node333;
	wire [13-1:0] node336;
	wire [13-1:0] node339;
	wire [13-1:0] node340;
	wire [13-1:0] node341;
	wire [13-1:0] node344;
	wire [13-1:0] node347;
	wire [13-1:0] node348;
	wire [13-1:0] node351;
	wire [13-1:0] node354;
	wire [13-1:0] node355;
	wire [13-1:0] node356;
	wire [13-1:0] node357;
	wire [13-1:0] node360;
	wire [13-1:0] node363;
	wire [13-1:0] node364;
	wire [13-1:0] node367;
	wire [13-1:0] node370;
	wire [13-1:0] node371;
	wire [13-1:0] node372;
	wire [13-1:0] node375;
	wire [13-1:0] node378;
	wire [13-1:0] node379;
	wire [13-1:0] node382;
	wire [13-1:0] node385;
	wire [13-1:0] node386;
	wire [13-1:0] node387;
	wire [13-1:0] node388;
	wire [13-1:0] node389;
	wire [13-1:0] node390;
	wire [13-1:0] node393;
	wire [13-1:0] node396;
	wire [13-1:0] node397;
	wire [13-1:0] node400;
	wire [13-1:0] node403;
	wire [13-1:0] node404;
	wire [13-1:0] node405;
	wire [13-1:0] node408;
	wire [13-1:0] node411;
	wire [13-1:0] node412;
	wire [13-1:0] node415;
	wire [13-1:0] node418;
	wire [13-1:0] node419;
	wire [13-1:0] node420;
	wire [13-1:0] node421;
	wire [13-1:0] node424;
	wire [13-1:0] node427;
	wire [13-1:0] node428;
	wire [13-1:0] node431;
	wire [13-1:0] node434;
	wire [13-1:0] node435;
	wire [13-1:0] node436;
	wire [13-1:0] node439;
	wire [13-1:0] node442;
	wire [13-1:0] node443;
	wire [13-1:0] node446;
	wire [13-1:0] node449;
	wire [13-1:0] node450;
	wire [13-1:0] node451;
	wire [13-1:0] node452;
	wire [13-1:0] node453;
	wire [13-1:0] node456;
	wire [13-1:0] node459;
	wire [13-1:0] node460;
	wire [13-1:0] node463;
	wire [13-1:0] node466;
	wire [13-1:0] node467;
	wire [13-1:0] node468;
	wire [13-1:0] node471;
	wire [13-1:0] node474;
	wire [13-1:0] node475;
	wire [13-1:0] node478;
	wire [13-1:0] node481;
	wire [13-1:0] node482;
	wire [13-1:0] node483;
	wire [13-1:0] node484;
	wire [13-1:0] node487;
	wire [13-1:0] node490;
	wire [13-1:0] node491;
	wire [13-1:0] node494;
	wire [13-1:0] node497;
	wire [13-1:0] node498;
	wire [13-1:0] node499;
	wire [13-1:0] node502;
	wire [13-1:0] node505;
	wire [13-1:0] node506;
	wire [13-1:0] node509;
	wire [13-1:0] node512;
	wire [13-1:0] node513;
	wire [13-1:0] node514;
	wire [13-1:0] node515;
	wire [13-1:0] node516;
	wire [13-1:0] node517;
	wire [13-1:0] node518;
	wire [13-1:0] node519;
	wire [13-1:0] node522;
	wire [13-1:0] node525;
	wire [13-1:0] node526;
	wire [13-1:0] node529;
	wire [13-1:0] node532;
	wire [13-1:0] node533;
	wire [13-1:0] node534;
	wire [13-1:0] node537;
	wire [13-1:0] node540;
	wire [13-1:0] node541;
	wire [13-1:0] node544;
	wire [13-1:0] node547;
	wire [13-1:0] node548;
	wire [13-1:0] node549;
	wire [13-1:0] node550;
	wire [13-1:0] node553;
	wire [13-1:0] node556;
	wire [13-1:0] node557;
	wire [13-1:0] node560;
	wire [13-1:0] node563;
	wire [13-1:0] node564;
	wire [13-1:0] node565;
	wire [13-1:0] node568;
	wire [13-1:0] node571;
	wire [13-1:0] node572;
	wire [13-1:0] node575;
	wire [13-1:0] node578;
	wire [13-1:0] node579;
	wire [13-1:0] node580;
	wire [13-1:0] node581;
	wire [13-1:0] node582;
	wire [13-1:0] node585;
	wire [13-1:0] node588;
	wire [13-1:0] node589;
	wire [13-1:0] node592;
	wire [13-1:0] node595;
	wire [13-1:0] node596;
	wire [13-1:0] node597;
	wire [13-1:0] node600;
	wire [13-1:0] node603;
	wire [13-1:0] node604;
	wire [13-1:0] node607;
	wire [13-1:0] node610;
	wire [13-1:0] node611;
	wire [13-1:0] node612;
	wire [13-1:0] node613;
	wire [13-1:0] node616;
	wire [13-1:0] node619;
	wire [13-1:0] node620;
	wire [13-1:0] node623;
	wire [13-1:0] node626;
	wire [13-1:0] node627;
	wire [13-1:0] node628;
	wire [13-1:0] node631;
	wire [13-1:0] node634;
	wire [13-1:0] node635;
	wire [13-1:0] node638;
	wire [13-1:0] node641;
	wire [13-1:0] node642;
	wire [13-1:0] node643;
	wire [13-1:0] node644;
	wire [13-1:0] node645;
	wire [13-1:0] node646;
	wire [13-1:0] node649;
	wire [13-1:0] node652;
	wire [13-1:0] node653;
	wire [13-1:0] node656;
	wire [13-1:0] node659;
	wire [13-1:0] node660;
	wire [13-1:0] node661;
	wire [13-1:0] node664;
	wire [13-1:0] node667;
	wire [13-1:0] node668;
	wire [13-1:0] node671;
	wire [13-1:0] node674;
	wire [13-1:0] node675;
	wire [13-1:0] node676;
	wire [13-1:0] node677;
	wire [13-1:0] node680;
	wire [13-1:0] node683;
	wire [13-1:0] node684;
	wire [13-1:0] node687;
	wire [13-1:0] node690;
	wire [13-1:0] node691;
	wire [13-1:0] node692;
	wire [13-1:0] node695;
	wire [13-1:0] node698;
	wire [13-1:0] node699;
	wire [13-1:0] node702;
	wire [13-1:0] node705;
	wire [13-1:0] node706;
	wire [13-1:0] node707;
	wire [13-1:0] node708;
	wire [13-1:0] node709;
	wire [13-1:0] node712;
	wire [13-1:0] node715;
	wire [13-1:0] node716;
	wire [13-1:0] node719;
	wire [13-1:0] node722;
	wire [13-1:0] node723;
	wire [13-1:0] node724;
	wire [13-1:0] node727;
	wire [13-1:0] node730;
	wire [13-1:0] node731;
	wire [13-1:0] node734;
	wire [13-1:0] node737;
	wire [13-1:0] node738;
	wire [13-1:0] node739;
	wire [13-1:0] node740;
	wire [13-1:0] node743;
	wire [13-1:0] node746;
	wire [13-1:0] node747;
	wire [13-1:0] node750;
	wire [13-1:0] node753;
	wire [13-1:0] node754;
	wire [13-1:0] node755;
	wire [13-1:0] node758;
	wire [13-1:0] node761;
	wire [13-1:0] node762;
	wire [13-1:0] node765;
	wire [13-1:0] node768;
	wire [13-1:0] node769;
	wire [13-1:0] node770;
	wire [13-1:0] node771;
	wire [13-1:0] node772;
	wire [13-1:0] node773;
	wire [13-1:0] node774;
	wire [13-1:0] node777;
	wire [13-1:0] node780;
	wire [13-1:0] node781;
	wire [13-1:0] node784;
	wire [13-1:0] node787;
	wire [13-1:0] node788;
	wire [13-1:0] node789;
	wire [13-1:0] node792;
	wire [13-1:0] node795;
	wire [13-1:0] node796;
	wire [13-1:0] node799;
	wire [13-1:0] node802;
	wire [13-1:0] node803;
	wire [13-1:0] node804;
	wire [13-1:0] node805;
	wire [13-1:0] node808;
	wire [13-1:0] node811;
	wire [13-1:0] node812;
	wire [13-1:0] node815;
	wire [13-1:0] node818;
	wire [13-1:0] node819;
	wire [13-1:0] node820;
	wire [13-1:0] node823;
	wire [13-1:0] node826;
	wire [13-1:0] node827;
	wire [13-1:0] node830;
	wire [13-1:0] node833;
	wire [13-1:0] node834;
	wire [13-1:0] node835;
	wire [13-1:0] node836;
	wire [13-1:0] node837;
	wire [13-1:0] node840;
	wire [13-1:0] node843;
	wire [13-1:0] node844;
	wire [13-1:0] node847;
	wire [13-1:0] node850;
	wire [13-1:0] node851;
	wire [13-1:0] node852;
	wire [13-1:0] node855;
	wire [13-1:0] node858;
	wire [13-1:0] node859;
	wire [13-1:0] node862;
	wire [13-1:0] node865;
	wire [13-1:0] node866;
	wire [13-1:0] node867;
	wire [13-1:0] node868;
	wire [13-1:0] node871;
	wire [13-1:0] node874;
	wire [13-1:0] node875;
	wire [13-1:0] node878;
	wire [13-1:0] node881;
	wire [13-1:0] node882;
	wire [13-1:0] node883;
	wire [13-1:0] node886;
	wire [13-1:0] node889;
	wire [13-1:0] node890;
	wire [13-1:0] node893;
	wire [13-1:0] node896;
	wire [13-1:0] node897;
	wire [13-1:0] node898;
	wire [13-1:0] node899;
	wire [13-1:0] node900;
	wire [13-1:0] node901;
	wire [13-1:0] node904;
	wire [13-1:0] node907;
	wire [13-1:0] node908;
	wire [13-1:0] node911;
	wire [13-1:0] node914;
	wire [13-1:0] node915;
	wire [13-1:0] node916;
	wire [13-1:0] node919;
	wire [13-1:0] node922;
	wire [13-1:0] node923;
	wire [13-1:0] node926;
	wire [13-1:0] node929;
	wire [13-1:0] node930;
	wire [13-1:0] node931;
	wire [13-1:0] node932;
	wire [13-1:0] node935;
	wire [13-1:0] node938;
	wire [13-1:0] node939;
	wire [13-1:0] node942;
	wire [13-1:0] node945;
	wire [13-1:0] node946;
	wire [13-1:0] node947;
	wire [13-1:0] node950;
	wire [13-1:0] node953;
	wire [13-1:0] node954;
	wire [13-1:0] node957;
	wire [13-1:0] node960;
	wire [13-1:0] node961;
	wire [13-1:0] node962;
	wire [13-1:0] node963;
	wire [13-1:0] node964;
	wire [13-1:0] node967;
	wire [13-1:0] node970;
	wire [13-1:0] node971;
	wire [13-1:0] node974;
	wire [13-1:0] node977;
	wire [13-1:0] node978;
	wire [13-1:0] node979;
	wire [13-1:0] node982;
	wire [13-1:0] node985;
	wire [13-1:0] node986;
	wire [13-1:0] node989;
	wire [13-1:0] node992;
	wire [13-1:0] node993;
	wire [13-1:0] node994;
	wire [13-1:0] node995;
	wire [13-1:0] node998;
	wire [13-1:0] node1001;
	wire [13-1:0] node1002;
	wire [13-1:0] node1005;
	wire [13-1:0] node1008;
	wire [13-1:0] node1009;
	wire [13-1:0] node1010;
	wire [13-1:0] node1013;
	wire [13-1:0] node1016;
	wire [13-1:0] node1017;
	wire [13-1:0] node1020;

	assign outp = (inp[1]) ? node512 : node1;
		assign node1 = (inp[9]) ? node257 : node2;
			assign node2 = (inp[10]) ? node130 : node3;
				assign node3 = (inp[11]) ? node67 : node4;
					assign node4 = (inp[6]) ? node36 : node5;
						assign node5 = (inp[2]) ? node21 : node6;
							assign node6 = (inp[7]) ? node14 : node7;
								assign node7 = (inp[3]) ? node11 : node8;
									assign node8 = (inp[5]) ? 13'b0001111111111 : 13'b0011111111111;
									assign node11 = (inp[0]) ? 13'b0000111111111 : 13'b0001111111111;
								assign node14 = (inp[5]) ? node18 : node15;
									assign node15 = (inp[4]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node18 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
							assign node21 = (inp[4]) ? node29 : node22;
								assign node22 = (inp[12]) ? node26 : node23;
									assign node23 = (inp[8]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node26 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node29 = (inp[3]) ? node33 : node30;
									assign node30 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node33 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
						assign node36 = (inp[12]) ? node52 : node37;
							assign node37 = (inp[0]) ? node45 : node38;
								assign node38 = (inp[3]) ? node42 : node39;
									assign node39 = (inp[5]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node42 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node45 = (inp[3]) ? node49 : node46;
									assign node46 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node49 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node52 = (inp[5]) ? node60 : node53;
								assign node53 = (inp[2]) ? node57 : node54;
									assign node54 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node57 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node60 = (inp[3]) ? node64 : node61;
									assign node61 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node64 = (inp[0]) ? 13'b0000000011111 : 13'b0000001111111;
					assign node67 = (inp[4]) ? node99 : node68;
						assign node68 = (inp[2]) ? node84 : node69;
							assign node69 = (inp[7]) ? node77 : node70;
								assign node70 = (inp[0]) ? node74 : node71;
									assign node71 = (inp[3]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node74 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node77 = (inp[5]) ? node81 : node78;
									assign node78 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node81 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node84 = (inp[0]) ? node92 : node85;
								assign node85 = (inp[6]) ? node89 : node86;
									assign node86 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node89 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node92 = (inp[7]) ? node96 : node93;
									assign node93 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node96 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node99 = (inp[3]) ? node115 : node100;
							assign node100 = (inp[6]) ? node108 : node101;
								assign node101 = (inp[12]) ? node105 : node102;
									assign node102 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node105 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node108 = (inp[5]) ? node112 : node109;
									assign node109 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node112 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node115 = (inp[12]) ? node123 : node116;
								assign node116 = (inp[2]) ? node120 : node117;
									assign node117 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node120 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node123 = (inp[6]) ? node127 : node124;
									assign node124 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node127 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
				assign node130 = (inp[5]) ? node194 : node131;
					assign node131 = (inp[3]) ? node163 : node132;
						assign node132 = (inp[11]) ? node148 : node133;
							assign node133 = (inp[2]) ? node141 : node134;
								assign node134 = (inp[12]) ? node138 : node135;
									assign node135 = (inp[4]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node138 = (inp[7]) ? 13'b0000011111111 : 13'b0001111111111;
								assign node141 = (inp[4]) ? node145 : node142;
									assign node142 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node145 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node148 = (inp[6]) ? node156 : node149;
								assign node149 = (inp[0]) ? node153 : node150;
									assign node150 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node153 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node156 = (inp[4]) ? node160 : node157;
									assign node157 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node160 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node163 = (inp[2]) ? node179 : node164;
							assign node164 = (inp[6]) ? node172 : node165;
								assign node165 = (inp[12]) ? node169 : node166;
									assign node166 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node169 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node172 = (inp[8]) ? node176 : node173;
									assign node173 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node176 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node179 = (inp[12]) ? node187 : node180;
								assign node180 = (inp[6]) ? node184 : node181;
									assign node181 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node184 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node187 = (inp[11]) ? node191 : node188;
									assign node188 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node191 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
					assign node194 = (inp[7]) ? node226 : node195;
						assign node195 = (inp[4]) ? node211 : node196;
							assign node196 = (inp[12]) ? node204 : node197;
								assign node197 = (inp[3]) ? node201 : node198;
									assign node198 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node201 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node204 = (inp[11]) ? node208 : node205;
									assign node205 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node208 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node211 = (inp[6]) ? node219 : node212;
								assign node212 = (inp[2]) ? node216 : node213;
									assign node213 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node216 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node219 = (inp[2]) ? node223 : node220;
									assign node220 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node223 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node226 = (inp[6]) ? node242 : node227;
							assign node227 = (inp[11]) ? node235 : node228;
								assign node228 = (inp[3]) ? node232 : node229;
									assign node229 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node232 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node235 = (inp[0]) ? node239 : node236;
									assign node236 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node239 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node242 = (inp[4]) ? node250 : node243;
								assign node243 = (inp[2]) ? node247 : node244;
									assign node244 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node247 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node250 = (inp[3]) ? node254 : node251;
									assign node251 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node254 = (inp[12]) ? 13'b0000000001111 : 13'b0000000011111;
			assign node257 = (inp[3]) ? node385 : node258;
				assign node258 = (inp[11]) ? node322 : node259;
					assign node259 = (inp[12]) ? node291 : node260;
						assign node260 = (inp[0]) ? node276 : node261;
							assign node261 = (inp[5]) ? node269 : node262;
								assign node262 = (inp[8]) ? node266 : node263;
									assign node263 = (inp[7]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node266 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node269 = (inp[6]) ? node273 : node270;
									assign node270 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node273 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node276 = (inp[8]) ? node284 : node277;
								assign node277 = (inp[7]) ? node281 : node278;
									assign node278 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node281 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node284 = (inp[4]) ? node288 : node285;
									assign node285 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node288 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node291 = (inp[8]) ? node307 : node292;
							assign node292 = (inp[7]) ? node300 : node293;
								assign node293 = (inp[5]) ? node297 : node294;
									assign node294 = (inp[4]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node297 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node300 = (inp[5]) ? node304 : node301;
									assign node301 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node304 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node307 = (inp[0]) ? node315 : node308;
								assign node308 = (inp[4]) ? node312 : node309;
									assign node309 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node312 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node315 = (inp[10]) ? node319 : node316;
									assign node316 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node319 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
					assign node322 = (inp[7]) ? node354 : node323;
						assign node323 = (inp[10]) ? node339 : node324;
							assign node324 = (inp[2]) ? node332 : node325;
								assign node325 = (inp[6]) ? node329 : node326;
									assign node326 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node329 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node332 = (inp[6]) ? node336 : node333;
									assign node333 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node336 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node339 = (inp[0]) ? node347 : node340;
								assign node340 = (inp[5]) ? node344 : node341;
									assign node341 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node344 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node347 = (inp[12]) ? node351 : node348;
									assign node348 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node351 = (inp[4]) ? 13'b0000000001111 : 13'b0000000111111;
						assign node354 = (inp[4]) ? node370 : node355;
							assign node355 = (inp[5]) ? node363 : node356;
								assign node356 = (inp[12]) ? node360 : node357;
									assign node357 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node360 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node363 = (inp[12]) ? node367 : node364;
									assign node364 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node367 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node370 = (inp[0]) ? node378 : node371;
								assign node371 = (inp[10]) ? node375 : node372;
									assign node372 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node375 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node378 = (inp[5]) ? node382 : node379;
									assign node379 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node382 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
				assign node385 = (inp[12]) ? node449 : node386;
					assign node386 = (inp[8]) ? node418 : node387;
						assign node387 = (inp[4]) ? node403 : node388;
							assign node388 = (inp[7]) ? node396 : node389;
								assign node389 = (inp[10]) ? node393 : node390;
									assign node390 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node393 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node396 = (inp[5]) ? node400 : node397;
									assign node397 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node400 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node403 = (inp[5]) ? node411 : node404;
								assign node404 = (inp[11]) ? node408 : node405;
									assign node405 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node408 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node411 = (inp[11]) ? node415 : node412;
									assign node412 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node415 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node418 = (inp[7]) ? node434 : node419;
							assign node419 = (inp[10]) ? node427 : node420;
								assign node420 = (inp[4]) ? node424 : node421;
									assign node421 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node424 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node427 = (inp[2]) ? node431 : node428;
									assign node428 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node431 = (inp[5]) ? 13'b0000000001111 : 13'b0000000111111;
							assign node434 = (inp[6]) ? node442 : node435;
								assign node435 = (inp[10]) ? node439 : node436;
									assign node436 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node439 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node442 = (inp[5]) ? node446 : node443;
									assign node443 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node446 = (inp[10]) ? 13'b0000000000111 : 13'b0000000011111;
					assign node449 = (inp[5]) ? node481 : node450;
						assign node450 = (inp[11]) ? node466 : node451;
							assign node451 = (inp[2]) ? node459 : node452;
								assign node452 = (inp[6]) ? node456 : node453;
									assign node453 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node456 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node459 = (inp[10]) ? node463 : node460;
									assign node460 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node463 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node466 = (inp[7]) ? node474 : node467;
								assign node467 = (inp[4]) ? node471 : node468;
									assign node468 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node471 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node474 = (inp[6]) ? node478 : node475;
									assign node475 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node478 = (inp[4]) ? 13'b0000000000111 : 13'b0000000011111;
						assign node481 = (inp[7]) ? node497 : node482;
							assign node482 = (inp[8]) ? node490 : node483;
								assign node483 = (inp[11]) ? node487 : node484;
									assign node484 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node487 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node490 = (inp[0]) ? node494 : node491;
									assign node491 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node494 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node497 = (inp[6]) ? node505 : node498;
								assign node498 = (inp[11]) ? node502 : node499;
									assign node499 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node502 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node505 = (inp[0]) ? node509 : node506;
									assign node506 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node509 = (inp[2]) ? 13'b0000000000111 : 13'b0000000001111;
		assign node512 = (inp[2]) ? node768 : node513;
			assign node513 = (inp[12]) ? node641 : node514;
				assign node514 = (inp[8]) ? node578 : node515;
					assign node515 = (inp[7]) ? node547 : node516;
						assign node516 = (inp[6]) ? node532 : node517;
							assign node517 = (inp[4]) ? node525 : node518;
								assign node518 = (inp[0]) ? node522 : node519;
									assign node519 = (inp[10]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node522 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node525 = (inp[5]) ? node529 : node526;
									assign node526 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node529 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node532 = (inp[0]) ? node540 : node533;
								assign node533 = (inp[5]) ? node537 : node534;
									assign node534 = (inp[4]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node537 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node540 = (inp[3]) ? node544 : node541;
									assign node541 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node544 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node547 = (inp[9]) ? node563 : node548;
							assign node548 = (inp[10]) ? node556 : node549;
								assign node549 = (inp[4]) ? node553 : node550;
									assign node550 = (inp[5]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node553 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node556 = (inp[11]) ? node560 : node557;
									assign node557 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node560 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node563 = (inp[3]) ? node571 : node564;
								assign node564 = (inp[11]) ? node568 : node565;
									assign node565 = (inp[4]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node568 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node571 = (inp[10]) ? node575 : node572;
									assign node572 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node575 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
					assign node578 = (inp[3]) ? node610 : node579;
						assign node579 = (inp[10]) ? node595 : node580;
							assign node580 = (inp[6]) ? node588 : node581;
								assign node581 = (inp[4]) ? node585 : node582;
									assign node582 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node585 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node588 = (inp[11]) ? node592 : node589;
									assign node589 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node592 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node595 = (inp[9]) ? node603 : node596;
								assign node596 = (inp[5]) ? node600 : node597;
									assign node597 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node600 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node603 = (inp[6]) ? node607 : node604;
									assign node604 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node607 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node610 = (inp[0]) ? node626 : node611;
							assign node611 = (inp[10]) ? node619 : node612;
								assign node612 = (inp[5]) ? node616 : node613;
									assign node613 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node616 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node619 = (inp[9]) ? node623 : node620;
									assign node620 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node623 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node626 = (inp[4]) ? node634 : node627;
								assign node627 = (inp[6]) ? node631 : node628;
									assign node628 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node631 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node634 = (inp[7]) ? node638 : node635;
									assign node635 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node638 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
				assign node641 = (inp[3]) ? node705 : node642;
					assign node642 = (inp[9]) ? node674 : node643;
						assign node643 = (inp[10]) ? node659 : node644;
							assign node644 = (inp[4]) ? node652 : node645;
								assign node645 = (inp[5]) ? node649 : node646;
									assign node646 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node649 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node652 = (inp[11]) ? node656 : node653;
									assign node653 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node656 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node659 = (inp[7]) ? node667 : node660;
								assign node660 = (inp[11]) ? node664 : node661;
									assign node661 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node664 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node667 = (inp[8]) ? node671 : node668;
									assign node668 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node671 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node674 = (inp[11]) ? node690 : node675;
							assign node675 = (inp[5]) ? node683 : node676;
								assign node676 = (inp[10]) ? node680 : node677;
									assign node677 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node680 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node683 = (inp[8]) ? node687 : node684;
									assign node684 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node687 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node690 = (inp[4]) ? node698 : node691;
								assign node691 = (inp[10]) ? node695 : node692;
									assign node692 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node695 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node698 = (inp[8]) ? node702 : node699;
									assign node699 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node702 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
					assign node705 = (inp[11]) ? node737 : node706;
						assign node706 = (inp[8]) ? node722 : node707;
							assign node707 = (inp[10]) ? node715 : node708;
								assign node708 = (inp[5]) ? node712 : node709;
									assign node709 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node712 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node715 = (inp[5]) ? node719 : node716;
									assign node716 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node719 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node722 = (inp[0]) ? node730 : node723;
								assign node723 = (inp[9]) ? node727 : node724;
									assign node724 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node727 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node730 = (inp[4]) ? node734 : node731;
									assign node731 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node734 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node737 = (inp[5]) ? node753 : node738;
							assign node738 = (inp[0]) ? node746 : node739;
								assign node739 = (inp[7]) ? node743 : node740;
									assign node740 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node743 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node746 = (inp[9]) ? node750 : node747;
									assign node747 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node750 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node753 = (inp[4]) ? node761 : node754;
								assign node754 = (inp[10]) ? node758 : node755;
									assign node755 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node758 = (inp[8]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node761 = (inp[8]) ? node765 : node762;
									assign node762 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node765 = (inp[7]) ? 13'b0000000000111 : 13'b0000000001111;
			assign node768 = (inp[7]) ? node896 : node769;
				assign node769 = (inp[11]) ? node833 : node770;
					assign node770 = (inp[9]) ? node802 : node771;
						assign node771 = (inp[4]) ? node787 : node772;
							assign node772 = (inp[12]) ? node780 : node773;
								assign node773 = (inp[5]) ? node777 : node774;
									assign node774 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node777 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node780 = (inp[3]) ? node784 : node781;
									assign node781 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node784 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node787 = (inp[10]) ? node795 : node788;
								assign node788 = (inp[6]) ? node792 : node789;
									assign node789 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node792 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node795 = (inp[12]) ? node799 : node796;
									assign node796 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node799 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node802 = (inp[10]) ? node818 : node803;
							assign node803 = (inp[0]) ? node811 : node804;
								assign node804 = (inp[3]) ? node808 : node805;
									assign node805 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node808 = (inp[4]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node811 = (inp[4]) ? node815 : node812;
									assign node812 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node815 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node818 = (inp[8]) ? node826 : node819;
								assign node819 = (inp[5]) ? node823 : node820;
									assign node820 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node823 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node826 = (inp[0]) ? node830 : node827;
									assign node827 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node830 = (inp[4]) ? 13'b0000000001111 : 13'b0000000011111;
					assign node833 = (inp[4]) ? node865 : node834;
						assign node834 = (inp[9]) ? node850 : node835;
							assign node835 = (inp[3]) ? node843 : node836;
								assign node836 = (inp[10]) ? node840 : node837;
									assign node837 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node840 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node843 = (inp[6]) ? node847 : node844;
									assign node844 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node847 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node850 = (inp[0]) ? node858 : node851;
								assign node851 = (inp[5]) ? node855 : node852;
									assign node852 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node855 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node858 = (inp[10]) ? node862 : node859;
									assign node859 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node862 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node865 = (inp[5]) ? node881 : node866;
							assign node866 = (inp[3]) ? node874 : node867;
								assign node867 = (inp[8]) ? node871 : node868;
									assign node868 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node871 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node874 = (inp[9]) ? node878 : node875;
									assign node875 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node878 = (inp[8]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node881 = (inp[12]) ? node889 : node882;
								assign node882 = (inp[10]) ? node886 : node883;
									assign node883 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node886 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node889 = (inp[3]) ? node893 : node890;
									assign node890 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node893 = (inp[10]) ? 13'b0000000000111 : 13'b0000000001111;
				assign node896 = (inp[4]) ? node960 : node897;
					assign node897 = (inp[11]) ? node929 : node898;
						assign node898 = (inp[3]) ? node914 : node899;
							assign node899 = (inp[0]) ? node907 : node900;
								assign node900 = (inp[9]) ? node904 : node901;
									assign node901 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node904 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node907 = (inp[5]) ? node911 : node908;
									assign node908 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node911 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node914 = (inp[0]) ? node922 : node915;
								assign node915 = (inp[6]) ? node919 : node916;
									assign node916 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node919 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node922 = (inp[6]) ? node926 : node923;
									assign node923 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node926 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node929 = (inp[5]) ? node945 : node930;
							assign node930 = (inp[0]) ? node938 : node931;
								assign node931 = (inp[12]) ? node935 : node932;
									assign node932 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node935 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node938 = (inp[3]) ? node942 : node939;
									assign node939 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node942 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node945 = (inp[9]) ? node953 : node946;
								assign node946 = (inp[6]) ? node950 : node947;
									assign node947 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node950 = (inp[12]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node953 = (inp[3]) ? node957 : node954;
									assign node954 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node957 = (inp[10]) ? 13'b0000000000111 : 13'b0000000001111;
					assign node960 = (inp[8]) ? node992 : node961;
						assign node961 = (inp[11]) ? node977 : node962;
							assign node962 = (inp[0]) ? node970 : node963;
								assign node963 = (inp[10]) ? node967 : node964;
									assign node964 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node967 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node970 = (inp[3]) ? node974 : node971;
									assign node971 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node974 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node977 = (inp[9]) ? node985 : node978;
								assign node978 = (inp[5]) ? node982 : node979;
									assign node979 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node982 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node985 = (inp[12]) ? node989 : node986;
									assign node986 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node989 = (inp[10]) ? 13'b0000000000111 : 13'b0000000001111;
						assign node992 = (inp[10]) ? node1008 : node993;
							assign node993 = (inp[9]) ? node1001 : node994;
								assign node994 = (inp[0]) ? node998 : node995;
									assign node995 = (inp[11]) ? 13'b0000000011111 : 13'b0000000011111;
									assign node998 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1001 = (inp[12]) ? node1005 : node1002;
									assign node1002 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1005 = (inp[0]) ? 13'b0000000000111 : 13'b0000000001111;
							assign node1008 = (inp[9]) ? node1016 : node1009;
								assign node1009 = (inp[3]) ? node1013 : node1010;
									assign node1010 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1013 = (inp[12]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node1016 = (inp[5]) ? node1020 : node1017;
									assign node1017 = (inp[11]) ? 13'b0000000000111 : 13'b0000000001111;
									assign node1020 = (inp[11]) ? 13'b0000000000011 : 13'b0000000000111;

endmodule