module dtc_split75_bm15 (
	input  wire [15-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node6;
	wire [1-1:0] node8;
	wire [1-1:0] node10;
	wire [1-1:0] node13;
	wire [1-1:0] node14;
	wire [1-1:0] node16;
	wire [1-1:0] node19;
	wire [1-1:0] node20;
	wire [1-1:0] node23;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node28;
	wire [1-1:0] node30;
	wire [1-1:0] node33;
	wire [1-1:0] node34;
	wire [1-1:0] node37;
	wire [1-1:0] node40;
	wire [1-1:0] node41;
	wire [1-1:0] node42;
	wire [1-1:0] node45;
	wire [1-1:0] node48;
	wire [1-1:0] node49;
	wire [1-1:0] node52;
	wire [1-1:0] node55;
	wire [1-1:0] node56;
	wire [1-1:0] node57;
	wire [1-1:0] node58;
	wire [1-1:0] node60;
	wire [1-1:0] node63;
	wire [1-1:0] node64;
	wire [1-1:0] node67;
	wire [1-1:0] node70;
	wire [1-1:0] node71;
	wire [1-1:0] node72;
	wire [1-1:0] node75;
	wire [1-1:0] node78;
	wire [1-1:0] node79;
	wire [1-1:0] node82;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node87;
	wire [1-1:0] node88;
	wire [1-1:0] node91;
	wire [1-1:0] node94;
	wire [1-1:0] node95;
	wire [1-1:0] node98;
	wire [1-1:0] node101;
	wire [1-1:0] node102;
	wire [1-1:0] node103;
	wire [1-1:0] node106;
	wire [1-1:0] node109;
	wire [1-1:0] node110;
	wire [1-1:0] node113;
	wire [1-1:0] node116;
	wire [1-1:0] node117;
	wire [1-1:0] node118;
	wire [1-1:0] node119;
	wire [1-1:0] node120;
	wire [1-1:0] node122;
	wire [1-1:0] node125;
	wire [1-1:0] node126;
	wire [1-1:0] node129;
	wire [1-1:0] node132;
	wire [1-1:0] node133;
	wire [1-1:0] node134;
	wire [1-1:0] node137;
	wire [1-1:0] node140;
	wire [1-1:0] node141;
	wire [1-1:0] node144;
	wire [1-1:0] node147;
	wire [1-1:0] node148;
	wire [1-1:0] node149;
	wire [1-1:0] node150;
	wire [1-1:0] node153;
	wire [1-1:0] node156;
	wire [1-1:0] node157;
	wire [1-1:0] node160;
	wire [1-1:0] node163;
	wire [1-1:0] node164;
	wire [1-1:0] node165;
	wire [1-1:0] node168;
	wire [1-1:0] node171;
	wire [1-1:0] node172;
	wire [1-1:0] node175;
	wire [1-1:0] node178;
	wire [1-1:0] node179;
	wire [1-1:0] node180;
	wire [1-1:0] node181;
	wire [1-1:0] node182;
	wire [1-1:0] node185;
	wire [1-1:0] node188;
	wire [1-1:0] node189;
	wire [1-1:0] node192;
	wire [1-1:0] node195;
	wire [1-1:0] node196;
	wire [1-1:0] node197;
	wire [1-1:0] node200;
	wire [1-1:0] node203;
	wire [1-1:0] node204;
	wire [1-1:0] node207;
	wire [1-1:0] node210;
	wire [1-1:0] node211;
	wire [1-1:0] node212;
	wire [1-1:0] node213;
	wire [1-1:0] node216;
	wire [1-1:0] node219;
	wire [1-1:0] node220;
	wire [1-1:0] node223;
	wire [1-1:0] node226;
	wire [1-1:0] node227;
	wire [1-1:0] node228;
	wire [1-1:0] node231;
	wire [1-1:0] node234;
	wire [1-1:0] node235;
	wire [1-1:0] node238;
	wire [1-1:0] node241;
	wire [1-1:0] node242;
	wire [1-1:0] node243;
	wire [1-1:0] node244;
	wire [1-1:0] node245;
	wire [1-1:0] node246;
	wire [1-1:0] node248;
	wire [1-1:0] node251;
	wire [1-1:0] node252;
	wire [1-1:0] node255;
	wire [1-1:0] node258;
	wire [1-1:0] node259;
	wire [1-1:0] node260;
	wire [1-1:0] node263;
	wire [1-1:0] node266;
	wire [1-1:0] node267;
	wire [1-1:0] node270;
	wire [1-1:0] node273;
	wire [1-1:0] node274;
	wire [1-1:0] node275;
	wire [1-1:0] node276;
	wire [1-1:0] node279;
	wire [1-1:0] node282;
	wire [1-1:0] node283;
	wire [1-1:0] node286;
	wire [1-1:0] node289;
	wire [1-1:0] node290;
	wire [1-1:0] node291;
	wire [1-1:0] node294;
	wire [1-1:0] node297;
	wire [1-1:0] node298;
	wire [1-1:0] node301;
	wire [1-1:0] node304;
	wire [1-1:0] node305;
	wire [1-1:0] node306;
	wire [1-1:0] node307;
	wire [1-1:0] node308;
	wire [1-1:0] node311;
	wire [1-1:0] node314;
	wire [1-1:0] node315;
	wire [1-1:0] node318;
	wire [1-1:0] node321;
	wire [1-1:0] node322;
	wire [1-1:0] node323;
	wire [1-1:0] node326;
	wire [1-1:0] node329;
	wire [1-1:0] node330;
	wire [1-1:0] node333;
	wire [1-1:0] node336;
	wire [1-1:0] node337;
	wire [1-1:0] node338;
	wire [1-1:0] node339;
	wire [1-1:0] node342;
	wire [1-1:0] node345;
	wire [1-1:0] node346;
	wire [1-1:0] node349;
	wire [1-1:0] node352;
	wire [1-1:0] node353;
	wire [1-1:0] node354;
	wire [1-1:0] node357;
	wire [1-1:0] node360;
	wire [1-1:0] node361;
	wire [1-1:0] node364;
	wire [1-1:0] node367;
	wire [1-1:0] node368;
	wire [1-1:0] node369;
	wire [1-1:0] node370;
	wire [1-1:0] node371;
	wire [1-1:0] node372;
	wire [1-1:0] node375;
	wire [1-1:0] node378;
	wire [1-1:0] node379;
	wire [1-1:0] node382;
	wire [1-1:0] node385;
	wire [1-1:0] node386;
	wire [1-1:0] node387;
	wire [1-1:0] node390;
	wire [1-1:0] node393;
	wire [1-1:0] node394;
	wire [1-1:0] node397;
	wire [1-1:0] node400;
	wire [1-1:0] node401;
	wire [1-1:0] node402;
	wire [1-1:0] node403;
	wire [1-1:0] node406;
	wire [1-1:0] node409;
	wire [1-1:0] node410;
	wire [1-1:0] node413;
	wire [1-1:0] node416;
	wire [1-1:0] node417;
	wire [1-1:0] node418;
	wire [1-1:0] node421;
	wire [1-1:0] node424;
	wire [1-1:0] node425;
	wire [1-1:0] node428;
	wire [1-1:0] node431;
	wire [1-1:0] node432;
	wire [1-1:0] node433;
	wire [1-1:0] node434;
	wire [1-1:0] node435;
	wire [1-1:0] node438;
	wire [1-1:0] node441;
	wire [1-1:0] node442;
	wire [1-1:0] node445;
	wire [1-1:0] node448;
	wire [1-1:0] node449;
	wire [1-1:0] node450;
	wire [1-1:0] node453;
	wire [1-1:0] node456;
	wire [1-1:0] node457;
	wire [1-1:0] node460;
	wire [1-1:0] node463;
	wire [1-1:0] node464;
	wire [1-1:0] node465;
	wire [1-1:0] node466;
	wire [1-1:0] node469;
	wire [1-1:0] node472;
	wire [1-1:0] node473;
	wire [1-1:0] node476;
	wire [1-1:0] node479;
	wire [1-1:0] node480;
	wire [1-1:0] node481;
	wire [1-1:0] node484;
	wire [1-1:0] node487;
	wire [1-1:0] node488;
	wire [1-1:0] node492;
	wire [1-1:0] node493;
	wire [1-1:0] node494;
	wire [1-1:0] node495;
	wire [1-1:0] node496;
	wire [1-1:0] node497;
	wire [1-1:0] node498;
	wire [1-1:0] node500;
	wire [1-1:0] node503;
	wire [1-1:0] node504;
	wire [1-1:0] node507;
	wire [1-1:0] node510;
	wire [1-1:0] node511;
	wire [1-1:0] node512;
	wire [1-1:0] node515;
	wire [1-1:0] node518;
	wire [1-1:0] node519;
	wire [1-1:0] node522;
	wire [1-1:0] node525;
	wire [1-1:0] node526;
	wire [1-1:0] node527;
	wire [1-1:0] node528;
	wire [1-1:0] node531;
	wire [1-1:0] node534;
	wire [1-1:0] node535;
	wire [1-1:0] node538;
	wire [1-1:0] node541;
	wire [1-1:0] node542;
	wire [1-1:0] node543;
	wire [1-1:0] node546;
	wire [1-1:0] node549;
	wire [1-1:0] node550;
	wire [1-1:0] node553;
	wire [1-1:0] node556;
	wire [1-1:0] node557;
	wire [1-1:0] node558;
	wire [1-1:0] node559;
	wire [1-1:0] node560;
	wire [1-1:0] node563;
	wire [1-1:0] node566;
	wire [1-1:0] node567;
	wire [1-1:0] node570;
	wire [1-1:0] node573;
	wire [1-1:0] node574;
	wire [1-1:0] node575;
	wire [1-1:0] node578;
	wire [1-1:0] node581;
	wire [1-1:0] node582;
	wire [1-1:0] node585;
	wire [1-1:0] node588;
	wire [1-1:0] node589;
	wire [1-1:0] node590;
	wire [1-1:0] node591;
	wire [1-1:0] node594;
	wire [1-1:0] node597;
	wire [1-1:0] node598;
	wire [1-1:0] node601;
	wire [1-1:0] node604;
	wire [1-1:0] node605;
	wire [1-1:0] node606;
	wire [1-1:0] node609;
	wire [1-1:0] node612;
	wire [1-1:0] node613;
	wire [1-1:0] node616;
	wire [1-1:0] node619;
	wire [1-1:0] node620;
	wire [1-1:0] node621;
	wire [1-1:0] node622;
	wire [1-1:0] node623;
	wire [1-1:0] node624;
	wire [1-1:0] node627;
	wire [1-1:0] node630;
	wire [1-1:0] node631;
	wire [1-1:0] node634;
	wire [1-1:0] node637;
	wire [1-1:0] node638;
	wire [1-1:0] node639;
	wire [1-1:0] node642;
	wire [1-1:0] node645;
	wire [1-1:0] node646;
	wire [1-1:0] node649;
	wire [1-1:0] node652;
	wire [1-1:0] node653;
	wire [1-1:0] node654;
	wire [1-1:0] node655;
	wire [1-1:0] node658;
	wire [1-1:0] node661;
	wire [1-1:0] node662;
	wire [1-1:0] node665;
	wire [1-1:0] node668;
	wire [1-1:0] node669;
	wire [1-1:0] node670;
	wire [1-1:0] node673;
	wire [1-1:0] node676;
	wire [1-1:0] node677;
	wire [1-1:0] node680;
	wire [1-1:0] node683;
	wire [1-1:0] node684;
	wire [1-1:0] node685;
	wire [1-1:0] node686;
	wire [1-1:0] node687;
	wire [1-1:0] node690;
	wire [1-1:0] node693;
	wire [1-1:0] node694;
	wire [1-1:0] node697;
	wire [1-1:0] node700;
	wire [1-1:0] node701;
	wire [1-1:0] node702;
	wire [1-1:0] node705;
	wire [1-1:0] node708;
	wire [1-1:0] node709;
	wire [1-1:0] node712;
	wire [1-1:0] node715;
	wire [1-1:0] node716;
	wire [1-1:0] node717;
	wire [1-1:0] node718;
	wire [1-1:0] node721;
	wire [1-1:0] node724;
	wire [1-1:0] node725;
	wire [1-1:0] node728;
	wire [1-1:0] node731;
	wire [1-1:0] node732;
	wire [1-1:0] node733;
	wire [1-1:0] node736;
	wire [1-1:0] node739;
	wire [1-1:0] node740;
	wire [1-1:0] node744;
	wire [1-1:0] node745;
	wire [1-1:0] node746;
	wire [1-1:0] node747;
	wire [1-1:0] node748;
	wire [1-1:0] node749;
	wire [1-1:0] node750;
	wire [1-1:0] node753;
	wire [1-1:0] node756;
	wire [1-1:0] node757;
	wire [1-1:0] node760;
	wire [1-1:0] node763;
	wire [1-1:0] node764;
	wire [1-1:0] node765;
	wire [1-1:0] node768;
	wire [1-1:0] node771;
	wire [1-1:0] node772;
	wire [1-1:0] node775;
	wire [1-1:0] node778;
	wire [1-1:0] node779;
	wire [1-1:0] node780;
	wire [1-1:0] node781;
	wire [1-1:0] node784;
	wire [1-1:0] node787;
	wire [1-1:0] node788;
	wire [1-1:0] node791;
	wire [1-1:0] node794;
	wire [1-1:0] node795;
	wire [1-1:0] node796;
	wire [1-1:0] node799;
	wire [1-1:0] node802;
	wire [1-1:0] node803;
	wire [1-1:0] node806;
	wire [1-1:0] node809;
	wire [1-1:0] node810;
	wire [1-1:0] node811;
	wire [1-1:0] node812;
	wire [1-1:0] node813;
	wire [1-1:0] node816;
	wire [1-1:0] node819;
	wire [1-1:0] node820;
	wire [1-1:0] node823;
	wire [1-1:0] node826;
	wire [1-1:0] node827;
	wire [1-1:0] node828;
	wire [1-1:0] node831;
	wire [1-1:0] node834;
	wire [1-1:0] node835;
	wire [1-1:0] node838;
	wire [1-1:0] node841;
	wire [1-1:0] node842;
	wire [1-1:0] node843;
	wire [1-1:0] node844;
	wire [1-1:0] node847;
	wire [1-1:0] node850;
	wire [1-1:0] node851;
	wire [1-1:0] node854;
	wire [1-1:0] node857;
	wire [1-1:0] node858;
	wire [1-1:0] node859;
	wire [1-1:0] node862;
	wire [1-1:0] node865;
	wire [1-1:0] node866;
	wire [1-1:0] node870;
	wire [1-1:0] node871;
	wire [1-1:0] node872;
	wire [1-1:0] node873;
	wire [1-1:0] node874;
	wire [1-1:0] node875;
	wire [1-1:0] node878;
	wire [1-1:0] node881;
	wire [1-1:0] node882;
	wire [1-1:0] node885;
	wire [1-1:0] node888;
	wire [1-1:0] node889;
	wire [1-1:0] node890;
	wire [1-1:0] node893;
	wire [1-1:0] node896;
	wire [1-1:0] node897;
	wire [1-1:0] node900;
	wire [1-1:0] node903;
	wire [1-1:0] node904;
	wire [1-1:0] node905;
	wire [1-1:0] node906;
	wire [1-1:0] node909;
	wire [1-1:0] node912;
	wire [1-1:0] node913;
	wire [1-1:0] node916;
	wire [1-1:0] node919;
	wire [1-1:0] node920;
	wire [1-1:0] node921;
	wire [1-1:0] node924;
	wire [1-1:0] node927;
	wire [1-1:0] node928;
	wire [1-1:0] node932;
	wire [1-1:0] node933;
	wire [1-1:0] node934;
	wire [1-1:0] node935;
	wire [1-1:0] node936;
	wire [1-1:0] node939;
	wire [1-1:0] node942;
	wire [1-1:0] node943;
	wire [1-1:0] node946;
	wire [1-1:0] node949;
	wire [1-1:0] node950;
	wire [1-1:0] node951;
	wire [1-1:0] node954;
	wire [1-1:0] node957;
	wire [1-1:0] node958;
	wire [1-1:0] node962;
	wire [1-1:0] node963;
	wire [1-1:0] node964;
	wire [1-1:0] node965;
	wire [1-1:0] node968;
	wire [1-1:0] node971;
	wire [1-1:0] node972;
	wire [1-1:0] node976;
	wire [1-1:0] node977;
	wire [1-1:0] node978;

	assign outp = (inp[12]) ? node492 : node1;
		assign node1 = (inp[1]) ? node241 : node2;
			assign node2 = (inp[13]) ? node116 : node3;
				assign node3 = (inp[11]) ? node55 : node4;
					assign node4 = (inp[5]) ? node26 : node5;
						assign node5 = (inp[10]) ? node13 : node6;
							assign node6 = (inp[3]) ? node8 : 1'b1;
								assign node8 = (inp[7]) ? node10 : 1'b1;
									assign node10 = (inp[2]) ? 1'b1 : 1'b1;
							assign node13 = (inp[8]) ? node19 : node14;
								assign node14 = (inp[14]) ? node16 : 1'b1;
									assign node16 = (inp[0]) ? 1'b1 : 1'b1;
								assign node19 = (inp[7]) ? node23 : node20;
									assign node20 = (inp[3]) ? 1'b1 : 1'b1;
									assign node23 = (inp[2]) ? 1'b1 : 1'b1;
						assign node26 = (inp[3]) ? node40 : node27;
							assign node27 = (inp[10]) ? node33 : node28;
								assign node28 = (inp[7]) ? node30 : 1'b1;
									assign node30 = (inp[9]) ? 1'b1 : 1'b1;
								assign node33 = (inp[0]) ? node37 : node34;
									assign node34 = (inp[2]) ? 1'b1 : 1'b1;
									assign node37 = (inp[14]) ? 1'b1 : 1'b1;
							assign node40 = (inp[8]) ? node48 : node41;
								assign node41 = (inp[14]) ? node45 : node42;
									assign node42 = (inp[2]) ? 1'b1 : 1'b1;
									assign node45 = (inp[10]) ? 1'b1 : 1'b1;
								assign node48 = (inp[7]) ? node52 : node49;
									assign node49 = (inp[9]) ? 1'b1 : 1'b1;
									assign node52 = (inp[4]) ? 1'b0 : 1'b1;
					assign node55 = (inp[4]) ? node85 : node56;
						assign node56 = (inp[2]) ? node70 : node57;
							assign node57 = (inp[9]) ? node63 : node58;
								assign node58 = (inp[6]) ? node60 : 1'b1;
									assign node60 = (inp[7]) ? 1'b1 : 1'b1;
								assign node63 = (inp[6]) ? node67 : node64;
									assign node64 = (inp[14]) ? 1'b1 : 1'b1;
									assign node67 = (inp[0]) ? 1'b1 : 1'b1;
							assign node70 = (inp[8]) ? node78 : node71;
								assign node71 = (inp[9]) ? node75 : node72;
									assign node72 = (inp[7]) ? 1'b1 : 1'b1;
									assign node75 = (inp[14]) ? 1'b1 : 1'b1;
								assign node78 = (inp[3]) ? node82 : node79;
									assign node79 = (inp[14]) ? 1'b1 : 1'b1;
									assign node82 = (inp[9]) ? 1'b0 : 1'b1;
						assign node85 = (inp[2]) ? node101 : node86;
							assign node86 = (inp[3]) ? node94 : node87;
								assign node87 = (inp[9]) ? node91 : node88;
									assign node88 = (inp[10]) ? 1'b1 : 1'b1;
									assign node91 = (inp[7]) ? 1'b1 : 1'b1;
								assign node94 = (inp[9]) ? node98 : node95;
									assign node95 = (inp[6]) ? 1'b1 : 1'b1;
									assign node98 = (inp[5]) ? 1'b0 : 1'b1;
							assign node101 = (inp[5]) ? node109 : node102;
								assign node102 = (inp[9]) ? node106 : node103;
									assign node103 = (inp[14]) ? 1'b1 : 1'b1;
									assign node106 = (inp[10]) ? 1'b0 : 1'b1;
								assign node109 = (inp[8]) ? node113 : node110;
									assign node110 = (inp[9]) ? 1'b0 : 1'b1;
									assign node113 = (inp[14]) ? 1'b0 : 1'b0;
				assign node116 = (inp[0]) ? node178 : node117;
					assign node117 = (inp[10]) ? node147 : node118;
						assign node118 = (inp[9]) ? node132 : node119;
							assign node119 = (inp[6]) ? node125 : node120;
								assign node120 = (inp[3]) ? node122 : 1'b1;
									assign node122 = (inp[7]) ? 1'b1 : 1'b1;
								assign node125 = (inp[2]) ? node129 : node126;
									assign node126 = (inp[8]) ? 1'b1 : 1'b1;
									assign node129 = (inp[3]) ? 1'b1 : 1'b1;
							assign node132 = (inp[3]) ? node140 : node133;
								assign node133 = (inp[8]) ? node137 : node134;
									assign node134 = (inp[5]) ? 1'b1 : 1'b1;
									assign node137 = (inp[2]) ? 1'b1 : 1'b1;
								assign node140 = (inp[7]) ? node144 : node141;
									assign node141 = (inp[14]) ? 1'b1 : 1'b1;
									assign node144 = (inp[5]) ? 1'b0 : 1'b1;
						assign node147 = (inp[5]) ? node163 : node148;
							assign node148 = (inp[8]) ? node156 : node149;
								assign node149 = (inp[6]) ? node153 : node150;
									assign node150 = (inp[11]) ? 1'b1 : 1'b1;
									assign node153 = (inp[4]) ? 1'b1 : 1'b1;
								assign node156 = (inp[9]) ? node160 : node157;
									assign node157 = (inp[6]) ? 1'b1 : 1'b1;
									assign node160 = (inp[14]) ? 1'b0 : 1'b1;
							assign node163 = (inp[6]) ? node171 : node164;
								assign node164 = (inp[8]) ? node168 : node165;
									assign node165 = (inp[2]) ? 1'b1 : 1'b1;
									assign node168 = (inp[7]) ? 1'b0 : 1'b1;
								assign node171 = (inp[3]) ? node175 : node172;
									assign node172 = (inp[2]) ? 1'b0 : 1'b1;
									assign node175 = (inp[14]) ? 1'b0 : 1'b0;
					assign node178 = (inp[9]) ? node210 : node179;
						assign node179 = (inp[4]) ? node195 : node180;
							assign node180 = (inp[7]) ? node188 : node181;
								assign node181 = (inp[10]) ? node185 : node182;
									assign node182 = (inp[14]) ? 1'b1 : 1'b1;
									assign node185 = (inp[8]) ? 1'b1 : 1'b1;
								assign node188 = (inp[11]) ? node192 : node189;
									assign node189 = (inp[6]) ? 1'b1 : 1'b1;
									assign node192 = (inp[10]) ? 1'b0 : 1'b1;
							assign node195 = (inp[6]) ? node203 : node196;
								assign node196 = (inp[3]) ? node200 : node197;
									assign node197 = (inp[2]) ? 1'b1 : 1'b1;
									assign node200 = (inp[5]) ? 1'b0 : 1'b1;
								assign node203 = (inp[7]) ? node207 : node204;
									assign node204 = (inp[2]) ? 1'b0 : 1'b1;
									assign node207 = (inp[8]) ? 1'b0 : 1'b0;
						assign node210 = (inp[2]) ? node226 : node211;
							assign node211 = (inp[4]) ? node219 : node212;
								assign node212 = (inp[10]) ? node216 : node213;
									assign node213 = (inp[5]) ? 1'b1 : 1'b1;
									assign node216 = (inp[3]) ? 1'b0 : 1'b1;
								assign node219 = (inp[7]) ? node223 : node220;
									assign node220 = (inp[5]) ? 1'b0 : 1'b1;
									assign node223 = (inp[11]) ? 1'b0 : 1'b0;
							assign node226 = (inp[5]) ? node234 : node227;
								assign node227 = (inp[7]) ? node231 : node228;
									assign node228 = (inp[3]) ? 1'b0 : 1'b1;
									assign node231 = (inp[10]) ? 1'b0 : 1'b0;
								assign node234 = (inp[8]) ? node238 : node235;
									assign node235 = (inp[6]) ? 1'b0 : 1'b0;
									assign node238 = (inp[11]) ? 1'b0 : 1'b0;
			assign node241 = (inp[3]) ? node367 : node242;
				assign node242 = (inp[5]) ? node304 : node243;
					assign node243 = (inp[6]) ? node273 : node244;
						assign node244 = (inp[8]) ? node258 : node245;
							assign node245 = (inp[7]) ? node251 : node246;
								assign node246 = (inp[4]) ? node248 : 1'b1;
									assign node248 = (inp[13]) ? 1'b1 : 1'b1;
								assign node251 = (inp[0]) ? node255 : node252;
									assign node252 = (inp[4]) ? 1'b1 : 1'b1;
									assign node255 = (inp[14]) ? 1'b1 : 1'b1;
							assign node258 = (inp[10]) ? node266 : node259;
								assign node259 = (inp[9]) ? node263 : node260;
									assign node260 = (inp[13]) ? 1'b1 : 1'b1;
									assign node263 = (inp[14]) ? 1'b1 : 1'b1;
								assign node266 = (inp[4]) ? node270 : node267;
									assign node267 = (inp[0]) ? 1'b1 : 1'b1;
									assign node270 = (inp[13]) ? 1'b0 : 1'b1;
						assign node273 = (inp[10]) ? node289 : node274;
							assign node274 = (inp[8]) ? node282 : node275;
								assign node275 = (inp[7]) ? node279 : node276;
									assign node276 = (inp[13]) ? 1'b1 : 1'b1;
									assign node279 = (inp[11]) ? 1'b1 : 1'b1;
								assign node282 = (inp[11]) ? node286 : node283;
									assign node283 = (inp[2]) ? 1'b1 : 1'b1;
									assign node286 = (inp[2]) ? 1'b0 : 1'b1;
							assign node289 = (inp[14]) ? node297 : node290;
								assign node290 = (inp[11]) ? node294 : node291;
									assign node291 = (inp[0]) ? 1'b1 : 1'b1;
									assign node294 = (inp[8]) ? 1'b0 : 1'b1;
								assign node297 = (inp[11]) ? node301 : node298;
									assign node298 = (inp[8]) ? 1'b0 : 1'b1;
									assign node301 = (inp[13]) ? 1'b0 : 1'b0;
					assign node304 = (inp[7]) ? node336 : node305;
						assign node305 = (inp[0]) ? node321 : node306;
							assign node306 = (inp[13]) ? node314 : node307;
								assign node307 = (inp[8]) ? node311 : node308;
									assign node308 = (inp[11]) ? 1'b1 : 1'b1;
									assign node311 = (inp[2]) ? 1'b1 : 1'b1;
								assign node314 = (inp[14]) ? node318 : node315;
									assign node315 = (inp[10]) ? 1'b1 : 1'b1;
									assign node318 = (inp[6]) ? 1'b0 : 1'b1;
							assign node321 = (inp[10]) ? node329 : node322;
								assign node322 = (inp[14]) ? node326 : node323;
									assign node323 = (inp[4]) ? 1'b1 : 1'b1;
									assign node326 = (inp[11]) ? 1'b0 : 1'b1;
								assign node329 = (inp[9]) ? node333 : node330;
									assign node330 = (inp[2]) ? 1'b0 : 1'b1;
									assign node333 = (inp[11]) ? 1'b0 : 1'b0;
						assign node336 = (inp[10]) ? node352 : node337;
							assign node337 = (inp[9]) ? node345 : node338;
								assign node338 = (inp[6]) ? node342 : node339;
									assign node339 = (inp[0]) ? 1'b1 : 1'b1;
									assign node342 = (inp[2]) ? 1'b0 : 1'b1;
								assign node345 = (inp[13]) ? node349 : node346;
									assign node346 = (inp[14]) ? 1'b0 : 1'b1;
									assign node349 = (inp[2]) ? 1'b0 : 1'b0;
							assign node352 = (inp[0]) ? node360 : node353;
								assign node353 = (inp[14]) ? node357 : node354;
									assign node354 = (inp[8]) ? 1'b0 : 1'b1;
									assign node357 = (inp[9]) ? 1'b0 : 1'b0;
								assign node360 = (inp[8]) ? node364 : node361;
									assign node361 = (inp[4]) ? 1'b0 : 1'b0;
									assign node364 = (inp[11]) ? 1'b0 : 1'b0;
				assign node367 = (inp[13]) ? node431 : node368;
					assign node368 = (inp[5]) ? node400 : node369;
						assign node369 = (inp[7]) ? node385 : node370;
							assign node370 = (inp[10]) ? node378 : node371;
								assign node371 = (inp[11]) ? node375 : node372;
									assign node372 = (inp[4]) ? 1'b1 : 1'b1;
									assign node375 = (inp[14]) ? 1'b1 : 1'b1;
								assign node378 = (inp[9]) ? node382 : node379;
									assign node379 = (inp[6]) ? 1'b1 : 1'b1;
									assign node382 = (inp[2]) ? 1'b0 : 1'b1;
							assign node385 = (inp[0]) ? node393 : node386;
								assign node386 = (inp[8]) ? node390 : node387;
									assign node387 = (inp[10]) ? 1'b1 : 1'b1;
									assign node390 = (inp[14]) ? 1'b0 : 1'b1;
								assign node393 = (inp[14]) ? node397 : node394;
									assign node394 = (inp[2]) ? 1'b0 : 1'b1;
									assign node397 = (inp[9]) ? 1'b0 : 1'b0;
						assign node400 = (inp[8]) ? node416 : node401;
							assign node401 = (inp[4]) ? node409 : node402;
								assign node402 = (inp[10]) ? node406 : node403;
									assign node403 = (inp[0]) ? 1'b1 : 1'b1;
									assign node406 = (inp[2]) ? 1'b0 : 1'b1;
								assign node409 = (inp[6]) ? node413 : node410;
									assign node410 = (inp[2]) ? 1'b0 : 1'b1;
									assign node413 = (inp[14]) ? 1'b0 : 1'b0;
							assign node416 = (inp[9]) ? node424 : node417;
								assign node417 = (inp[14]) ? node421 : node418;
									assign node418 = (inp[11]) ? 1'b0 : 1'b1;
									assign node421 = (inp[10]) ? 1'b0 : 1'b0;
								assign node424 = (inp[0]) ? node428 : node425;
									assign node425 = (inp[4]) ? 1'b0 : 1'b0;
									assign node428 = (inp[14]) ? 1'b0 : 1'b0;
					assign node431 = (inp[2]) ? node463 : node432;
						assign node432 = (inp[11]) ? node448 : node433;
							assign node433 = (inp[7]) ? node441 : node434;
								assign node434 = (inp[6]) ? node438 : node435;
									assign node435 = (inp[9]) ? 1'b1 : 1'b1;
									assign node438 = (inp[10]) ? 1'b0 : 1'b1;
								assign node441 = (inp[8]) ? node445 : node442;
									assign node442 = (inp[5]) ? 1'b0 : 1'b1;
									assign node445 = (inp[9]) ? 1'b0 : 1'b0;
							assign node448 = (inp[4]) ? node456 : node449;
								assign node449 = (inp[0]) ? node453 : node450;
									assign node450 = (inp[7]) ? 1'b0 : 1'b1;
									assign node453 = (inp[14]) ? 1'b0 : 1'b0;
								assign node456 = (inp[14]) ? node460 : node457;
									assign node457 = (inp[8]) ? 1'b0 : 1'b0;
									assign node460 = (inp[10]) ? 1'b0 : 1'b0;
						assign node463 = (inp[8]) ? node479 : node464;
							assign node464 = (inp[9]) ? node472 : node465;
								assign node465 = (inp[0]) ? node469 : node466;
									assign node466 = (inp[5]) ? 1'b0 : 1'b1;
									assign node469 = (inp[14]) ? 1'b0 : 1'b0;
								assign node472 = (inp[14]) ? node476 : node473;
									assign node473 = (inp[0]) ? 1'b0 : 1'b0;
									assign node476 = (inp[4]) ? 1'b0 : 1'b0;
							assign node479 = (inp[14]) ? node487 : node480;
								assign node480 = (inp[4]) ? node484 : node481;
									assign node481 = (inp[7]) ? 1'b0 : 1'b0;
									assign node484 = (inp[6]) ? 1'b0 : 1'b0;
								assign node487 = (inp[9]) ? 1'b0 : node488;
									assign node488 = (inp[11]) ? 1'b0 : 1'b0;
		assign node492 = (inp[6]) ? node744 : node493;
			assign node493 = (inp[7]) ? node619 : node494;
				assign node494 = (inp[3]) ? node556 : node495;
					assign node495 = (inp[1]) ? node525 : node496;
						assign node496 = (inp[2]) ? node510 : node497;
							assign node497 = (inp[10]) ? node503 : node498;
								assign node498 = (inp[9]) ? node500 : 1'b1;
									assign node500 = (inp[11]) ? 1'b1 : 1'b1;
								assign node503 = (inp[8]) ? node507 : node504;
									assign node504 = (inp[4]) ? 1'b1 : 1'b1;
									assign node507 = (inp[13]) ? 1'b1 : 1'b1;
							assign node510 = (inp[4]) ? node518 : node511;
								assign node511 = (inp[13]) ? node515 : node512;
									assign node512 = (inp[0]) ? 1'b1 : 1'b1;
									assign node515 = (inp[10]) ? 1'b1 : 1'b1;
								assign node518 = (inp[11]) ? node522 : node519;
									assign node519 = (inp[0]) ? 1'b1 : 1'b1;
									assign node522 = (inp[9]) ? 1'b0 : 1'b1;
						assign node525 = (inp[11]) ? node541 : node526;
							assign node526 = (inp[5]) ? node534 : node527;
								assign node527 = (inp[2]) ? node531 : node528;
									assign node528 = (inp[8]) ? 1'b1 : 1'b1;
									assign node531 = (inp[9]) ? 1'b1 : 1'b1;
								assign node534 = (inp[4]) ? node538 : node535;
									assign node535 = (inp[9]) ? 1'b1 : 1'b1;
									assign node538 = (inp[0]) ? 1'b0 : 1'b1;
							assign node541 = (inp[13]) ? node549 : node542;
								assign node542 = (inp[4]) ? node546 : node543;
									assign node543 = (inp[9]) ? 1'b1 : 1'b1;
									assign node546 = (inp[14]) ? 1'b0 : 1'b1;
								assign node549 = (inp[4]) ? node553 : node550;
									assign node550 = (inp[2]) ? 1'b0 : 1'b1;
									assign node553 = (inp[9]) ? 1'b0 : 1'b0;
					assign node556 = (inp[5]) ? node588 : node557;
						assign node557 = (inp[0]) ? node573 : node558;
							assign node558 = (inp[1]) ? node566 : node559;
								assign node559 = (inp[8]) ? node563 : node560;
									assign node560 = (inp[2]) ? 1'b1 : 1'b1;
									assign node563 = (inp[14]) ? 1'b1 : 1'b1;
								assign node566 = (inp[4]) ? node570 : node567;
									assign node567 = (inp[14]) ? 1'b1 : 1'b1;
									assign node570 = (inp[2]) ? 1'b0 : 1'b1;
							assign node573 = (inp[4]) ? node581 : node574;
								assign node574 = (inp[13]) ? node578 : node575;
									assign node575 = (inp[10]) ? 1'b1 : 1'b1;
									assign node578 = (inp[2]) ? 1'b0 : 1'b1;
								assign node581 = (inp[9]) ? node585 : node582;
									assign node582 = (inp[13]) ? 1'b0 : 1'b1;
									assign node585 = (inp[11]) ? 1'b0 : 1'b0;
						assign node588 = (inp[9]) ? node604 : node589;
							assign node589 = (inp[1]) ? node597 : node590;
								assign node590 = (inp[11]) ? node594 : node591;
									assign node591 = (inp[0]) ? 1'b1 : 1'b1;
									assign node594 = (inp[2]) ? 1'b0 : 1'b1;
								assign node597 = (inp[13]) ? node601 : node598;
									assign node598 = (inp[10]) ? 1'b0 : 1'b1;
									assign node601 = (inp[4]) ? 1'b0 : 1'b0;
							assign node604 = (inp[2]) ? node612 : node605;
								assign node605 = (inp[1]) ? node609 : node606;
									assign node606 = (inp[4]) ? 1'b0 : 1'b1;
									assign node609 = (inp[14]) ? 1'b0 : 1'b0;
								assign node612 = (inp[13]) ? node616 : node613;
									assign node613 = (inp[8]) ? 1'b0 : 1'b0;
									assign node616 = (inp[10]) ? 1'b0 : 1'b0;
				assign node619 = (inp[5]) ? node683 : node620;
					assign node620 = (inp[0]) ? node652 : node621;
						assign node621 = (inp[9]) ? node637 : node622;
							assign node622 = (inp[10]) ? node630 : node623;
								assign node623 = (inp[13]) ? node627 : node624;
									assign node624 = (inp[3]) ? 1'b1 : 1'b1;
									assign node627 = (inp[8]) ? 1'b1 : 1'b1;
								assign node630 = (inp[14]) ? node634 : node631;
									assign node631 = (inp[3]) ? 1'b1 : 1'b1;
									assign node634 = (inp[13]) ? 1'b0 : 1'b1;
							assign node637 = (inp[4]) ? node645 : node638;
								assign node638 = (inp[8]) ? node642 : node639;
									assign node639 = (inp[2]) ? 1'b1 : 1'b1;
									assign node642 = (inp[1]) ? 1'b0 : 1'b1;
								assign node645 = (inp[11]) ? node649 : node646;
									assign node646 = (inp[2]) ? 1'b0 : 1'b1;
									assign node649 = (inp[3]) ? 1'b0 : 1'b0;
						assign node652 = (inp[2]) ? node668 : node653;
							assign node653 = (inp[1]) ? node661 : node654;
								assign node654 = (inp[3]) ? node658 : node655;
									assign node655 = (inp[13]) ? 1'b1 : 1'b1;
									assign node658 = (inp[11]) ? 1'b0 : 1'b1;
								assign node661 = (inp[4]) ? node665 : node662;
									assign node662 = (inp[3]) ? 1'b0 : 1'b1;
									assign node665 = (inp[10]) ? 1'b0 : 1'b0;
							assign node668 = (inp[4]) ? node676 : node669;
								assign node669 = (inp[3]) ? node673 : node670;
									assign node670 = (inp[14]) ? 1'b0 : 1'b1;
									assign node673 = (inp[9]) ? 1'b0 : 1'b0;
								assign node676 = (inp[14]) ? node680 : node677;
									assign node677 = (inp[11]) ? 1'b0 : 1'b0;
									assign node680 = (inp[3]) ? 1'b0 : 1'b0;
					assign node683 = (inp[14]) ? node715 : node684;
						assign node684 = (inp[9]) ? node700 : node685;
							assign node685 = (inp[2]) ? node693 : node686;
								assign node686 = (inp[4]) ? node690 : node687;
									assign node687 = (inp[10]) ? 1'b1 : 1'b1;
									assign node690 = (inp[1]) ? 1'b0 : 1'b1;
								assign node693 = (inp[10]) ? node697 : node694;
									assign node694 = (inp[3]) ? 1'b0 : 1'b1;
									assign node697 = (inp[0]) ? 1'b0 : 1'b0;
							assign node700 = (inp[0]) ? node708 : node701;
								assign node701 = (inp[1]) ? node705 : node702;
									assign node702 = (inp[8]) ? 1'b0 : 1'b1;
									assign node705 = (inp[13]) ? 1'b0 : 1'b0;
								assign node708 = (inp[4]) ? node712 : node709;
									assign node709 = (inp[8]) ? 1'b0 : 1'b0;
									assign node712 = (inp[1]) ? 1'b0 : 1'b0;
						assign node715 = (inp[10]) ? node731 : node716;
							assign node716 = (inp[8]) ? node724 : node717;
								assign node717 = (inp[4]) ? node721 : node718;
									assign node718 = (inp[1]) ? 1'b0 : 1'b1;
									assign node721 = (inp[3]) ? 1'b0 : 1'b0;
								assign node724 = (inp[11]) ? node728 : node725;
									assign node725 = (inp[9]) ? 1'b0 : 1'b0;
									assign node728 = (inp[1]) ? 1'b0 : 1'b0;
							assign node731 = (inp[4]) ? node739 : node732;
								assign node732 = (inp[11]) ? node736 : node733;
									assign node733 = (inp[3]) ? 1'b0 : 1'b0;
									assign node736 = (inp[13]) ? 1'b0 : 1'b0;
								assign node739 = (inp[13]) ? 1'b0 : node740;
									assign node740 = (inp[3]) ? 1'b0 : 1'b0;
			assign node744 = (inp[13]) ? node870 : node745;
				assign node745 = (inp[8]) ? node809 : node746;
					assign node746 = (inp[5]) ? node778 : node747;
						assign node747 = (inp[10]) ? node763 : node748;
							assign node748 = (inp[2]) ? node756 : node749;
								assign node749 = (inp[9]) ? node753 : node750;
									assign node750 = (inp[3]) ? 1'b1 : 1'b1;
									assign node753 = (inp[1]) ? 1'b1 : 1'b1;
								assign node756 = (inp[3]) ? node760 : node757;
									assign node757 = (inp[9]) ? 1'b1 : 1'b1;
									assign node760 = (inp[14]) ? 1'b0 : 1'b1;
							assign node763 = (inp[14]) ? node771 : node764;
								assign node764 = (inp[0]) ? node768 : node765;
									assign node765 = (inp[4]) ? 1'b1 : 1'b1;
									assign node768 = (inp[7]) ? 1'b0 : 1'b1;
								assign node771 = (inp[11]) ? node775 : node772;
									assign node772 = (inp[3]) ? 1'b0 : 1'b1;
									assign node775 = (inp[9]) ? 1'b0 : 1'b0;
						assign node778 = (inp[4]) ? node794 : node779;
							assign node779 = (inp[11]) ? node787 : node780;
								assign node780 = (inp[10]) ? node784 : node781;
									assign node781 = (inp[0]) ? 1'b1 : 1'b1;
									assign node784 = (inp[3]) ? 1'b0 : 1'b1;
								assign node787 = (inp[3]) ? node791 : node788;
									assign node788 = (inp[9]) ? 1'b0 : 1'b1;
									assign node791 = (inp[1]) ? 1'b0 : 1'b0;
							assign node794 = (inp[0]) ? node802 : node795;
								assign node795 = (inp[7]) ? node799 : node796;
									assign node796 = (inp[9]) ? 1'b0 : 1'b1;
									assign node799 = (inp[10]) ? 1'b0 : 1'b0;
								assign node802 = (inp[14]) ? node806 : node803;
									assign node803 = (inp[7]) ? 1'b0 : 1'b0;
									assign node806 = (inp[3]) ? 1'b0 : 1'b0;
					assign node809 = (inp[0]) ? node841 : node810;
						assign node810 = (inp[9]) ? node826 : node811;
							assign node811 = (inp[14]) ? node819 : node812;
								assign node812 = (inp[11]) ? node816 : node813;
									assign node813 = (inp[3]) ? 1'b1 : 1'b1;
									assign node816 = (inp[2]) ? 1'b0 : 1'b1;
								assign node819 = (inp[2]) ? node823 : node820;
									assign node820 = (inp[4]) ? 1'b0 : 1'b1;
									assign node823 = (inp[5]) ? 1'b0 : 1'b0;
							assign node826 = (inp[10]) ? node834 : node827;
								assign node827 = (inp[1]) ? node831 : node828;
									assign node828 = (inp[2]) ? 1'b0 : 1'b1;
									assign node831 = (inp[4]) ? 1'b0 : 1'b0;
								assign node834 = (inp[1]) ? node838 : node835;
									assign node835 = (inp[3]) ? 1'b0 : 1'b0;
									assign node838 = (inp[7]) ? 1'b0 : 1'b0;
						assign node841 = (inp[4]) ? node857 : node842;
							assign node842 = (inp[5]) ? node850 : node843;
								assign node843 = (inp[11]) ? node847 : node844;
									assign node844 = (inp[7]) ? 1'b0 : 1'b1;
									assign node847 = (inp[3]) ? 1'b0 : 1'b0;
								assign node850 = (inp[10]) ? node854 : node851;
									assign node851 = (inp[14]) ? 1'b0 : 1'b0;
									assign node854 = (inp[11]) ? 1'b0 : 1'b0;
							assign node857 = (inp[7]) ? node865 : node858;
								assign node858 = (inp[9]) ? node862 : node859;
									assign node859 = (inp[3]) ? 1'b0 : 1'b0;
									assign node862 = (inp[2]) ? 1'b0 : 1'b0;
								assign node865 = (inp[1]) ? 1'b0 : node866;
									assign node866 = (inp[11]) ? 1'b0 : 1'b0;
				assign node870 = (inp[8]) ? node932 : node871;
					assign node871 = (inp[11]) ? node903 : node872;
						assign node872 = (inp[0]) ? node888 : node873;
							assign node873 = (inp[3]) ? node881 : node874;
								assign node874 = (inp[5]) ? node878 : node875;
									assign node875 = (inp[9]) ? 1'b1 : 1'b1;
									assign node878 = (inp[14]) ? 1'b0 : 1'b1;
								assign node881 = (inp[4]) ? node885 : node882;
									assign node882 = (inp[14]) ? 1'b0 : 1'b1;
									assign node885 = (inp[9]) ? 1'b0 : 1'b0;
							assign node888 = (inp[1]) ? node896 : node889;
								assign node889 = (inp[10]) ? node893 : node890;
									assign node890 = (inp[14]) ? 1'b0 : 1'b1;
									assign node893 = (inp[2]) ? 1'b0 : 1'b0;
								assign node896 = (inp[2]) ? node900 : node897;
									assign node897 = (inp[14]) ? 1'b0 : 1'b0;
									assign node900 = (inp[3]) ? 1'b0 : 1'b0;
						assign node903 = (inp[9]) ? node919 : node904;
							assign node904 = (inp[10]) ? node912 : node905;
								assign node905 = (inp[3]) ? node909 : node906;
									assign node906 = (inp[14]) ? 1'b0 : 1'b1;
									assign node909 = (inp[5]) ? 1'b0 : 1'b0;
								assign node912 = (inp[14]) ? node916 : node913;
									assign node913 = (inp[4]) ? 1'b0 : 1'b0;
									assign node916 = (inp[5]) ? 1'b0 : 1'b0;
							assign node919 = (inp[0]) ? node927 : node920;
								assign node920 = (inp[14]) ? node924 : node921;
									assign node921 = (inp[5]) ? 1'b0 : 1'b0;
									assign node924 = (inp[4]) ? 1'b0 : 1'b0;
								assign node927 = (inp[1]) ? 1'b0 : node928;
									assign node928 = (inp[10]) ? 1'b0 : 1'b0;
					assign node932 = (inp[9]) ? node962 : node933;
						assign node933 = (inp[2]) ? node949 : node934;
							assign node934 = (inp[7]) ? node942 : node935;
								assign node935 = (inp[4]) ? node939 : node936;
									assign node936 = (inp[1]) ? 1'b0 : 1'b1;
									assign node939 = (inp[0]) ? 1'b0 : 1'b0;
								assign node942 = (inp[4]) ? node946 : node943;
									assign node943 = (inp[3]) ? 1'b0 : 1'b0;
									assign node946 = (inp[0]) ? 1'b0 : 1'b0;
							assign node949 = (inp[14]) ? node957 : node950;
								assign node950 = (inp[1]) ? node954 : node951;
									assign node951 = (inp[11]) ? 1'b0 : 1'b0;
									assign node954 = (inp[10]) ? 1'b0 : 1'b0;
								assign node957 = (inp[10]) ? 1'b0 : node958;
									assign node958 = (inp[0]) ? 1'b0 : 1'b0;
						assign node962 = (inp[0]) ? node976 : node963;
							assign node963 = (inp[4]) ? node971 : node964;
								assign node964 = (inp[10]) ? node968 : node965;
									assign node965 = (inp[7]) ? 1'b0 : 1'b0;
									assign node968 = (inp[11]) ? 1'b0 : 1'b0;
								assign node971 = (inp[1]) ? 1'b0 : node972;
									assign node972 = (inp[14]) ? 1'b0 : 1'b0;
							assign node976 = (inp[10]) ? 1'b0 : node977;
								assign node977 = (inp[7]) ? 1'b0 : node978;
									assign node978 = (inp[3]) ? 1'b0 : 1'b0;

endmodule