module dtc_split66_bm84 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node171;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node247;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node260;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node273;
	wire [3-1:0] node275;
	wire [3-1:0] node278;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;

	assign outp = (inp[9]) ? node214 : node1;
		assign node1 = (inp[6]) ? node127 : node2;
			assign node2 = (inp[10]) ? node50 : node3;
				assign node3 = (inp[7]) ? node11 : node4;
					assign node4 = (inp[3]) ? node6 : 3'b111;
						assign node6 = (inp[11]) ? node8 : 3'b111;
							assign node8 = (inp[8]) ? 3'b011 : 3'b111;
					assign node11 = (inp[11]) ? node27 : node12;
						assign node12 = (inp[3]) ? node20 : node13;
							assign node13 = (inp[8]) ? node15 : 3'b111;
								assign node15 = (inp[1]) ? node17 : 3'b111;
									assign node17 = (inp[2]) ? 3'b111 : 3'b011;
							assign node20 = (inp[8]) ? 3'b011 : node21;
								assign node21 = (inp[4]) ? node23 : 3'b111;
									assign node23 = (inp[5]) ? 3'b011 : 3'b111;
						assign node27 = (inp[3]) ? node37 : node28;
							assign node28 = (inp[2]) ? 3'b011 : node29;
								assign node29 = (inp[8]) ? node33 : node30;
									assign node30 = (inp[4]) ? 3'b011 : 3'b111;
									assign node33 = (inp[1]) ? 3'b001 : 3'b011;
							assign node37 = (inp[8]) ? node43 : node38;
								assign node38 = (inp[4]) ? node40 : 3'b011;
									assign node40 = (inp[5]) ? 3'b101 : 3'b111;
								assign node43 = (inp[0]) ? node45 : 3'b101;
									assign node45 = (inp[1]) ? node47 : 3'b101;
										assign node47 = (inp[2]) ? 3'b001 : 3'b101;
				assign node50 = (inp[11]) ? node98 : node51;
					assign node51 = (inp[8]) ? node73 : node52;
						assign node52 = (inp[3]) ? node60 : node53;
							assign node53 = (inp[7]) ? node55 : 3'b111;
								assign node55 = (inp[4]) ? 3'b101 : node56;
									assign node56 = (inp[2]) ? 3'b111 : 3'b011;
							assign node60 = (inp[4]) ? node70 : node61;
								assign node61 = (inp[7]) ? 3'b111 : node62;
									assign node62 = (inp[5]) ? 3'b011 : node63;
										assign node63 = (inp[1]) ? 3'b011 : node64;
											assign node64 = (inp[2]) ? 3'b011 : 3'b111;
								assign node70 = (inp[7]) ? 3'b001 : 3'b011;
						assign node73 = (inp[7]) ? node79 : node74;
							assign node74 = (inp[3]) ? node76 : 3'b011;
								assign node76 = (inp[4]) ? 3'b101 : 3'b001;
							assign node79 = (inp[2]) ? node91 : node80;
								assign node80 = (inp[3]) ? node86 : node81;
									assign node81 = (inp[5]) ? node83 : 3'b101;
										assign node83 = (inp[4]) ? 3'b001 : 3'b101;
									assign node86 = (inp[0]) ? node88 : 3'b001;
										assign node88 = (inp[1]) ? 3'b110 : 3'b001;
								assign node91 = (inp[1]) ? node93 : 3'b001;
									assign node93 = (inp[5]) ? node95 : 3'b001;
										assign node95 = (inp[0]) ? 3'b110 : 3'b001;
					assign node98 = (inp[7]) ? node108 : node99;
						assign node99 = (inp[3]) ? node103 : node100;
							assign node100 = (inp[8]) ? 3'b101 : 3'b011;
							assign node103 = (inp[8]) ? node105 : 3'b101;
								assign node105 = (inp[4]) ? 3'b001 : 3'b101;
						assign node108 = (inp[8]) ? node116 : node109;
							assign node109 = (inp[4]) ? node111 : 3'b101;
								assign node111 = (inp[3]) ? node113 : 3'b101;
									assign node113 = (inp[5]) ? 3'b110 : 3'b101;
							assign node116 = (inp[3]) ? node122 : node117;
								assign node117 = (inp[2]) ? 3'b101 : node118;
									assign node118 = (inp[1]) ? 3'b110 : 3'b101;
								assign node122 = (inp[4]) ? node124 : 3'b110;
									assign node124 = (inp[0]) ? 3'b010 : 3'b110;
			assign node127 = (inp[10]) ? node193 : node128;
				assign node128 = (inp[11]) ? node174 : node129;
					assign node129 = (inp[7]) ? node153 : node130;
						assign node130 = (inp[4]) ? node142 : node131;
							assign node131 = (inp[8]) ? node133 : 3'b011;
								assign node133 = (inp[5]) ? node135 : 3'b011;
									assign node135 = (inp[3]) ? 3'b001 : node136;
										assign node136 = (inp[2]) ? 3'b001 : node137;
											assign node137 = (inp[1]) ? 3'b001 : 3'b101;
							assign node142 = (inp[8]) ? node146 : node143;
								assign node143 = (inp[3]) ? 3'b101 : 3'b011;
								assign node146 = (inp[2]) ? 3'b001 : node147;
									assign node147 = (inp[3]) ? 3'b001 : node148;
										assign node148 = (inp[1]) ? 3'b001 : 3'b101;
						assign node153 = (inp[4]) ? node163 : node154;
							assign node154 = (inp[3]) ? node160 : node155;
								assign node155 = (inp[2]) ? 3'b001 : node156;
									assign node156 = (inp[8]) ? 3'b001 : 3'b101;
								assign node160 = (inp[8]) ? 3'b110 : 3'b001;
							assign node163 = (inp[3]) ? node167 : node164;
								assign node164 = (inp[8]) ? 3'b110 : 3'b001;
								assign node167 = (inp[8]) ? node169 : 3'b110;
									assign node169 = (inp[0]) ? node171 : 3'b110;
										assign node171 = (inp[5]) ? 3'b010 : 3'b110;
					assign node174 = (inp[7]) ? node178 : node175;
						assign node175 = (inp[8]) ? 3'b110 : 3'b001;
						assign node178 = (inp[8]) ? node184 : node179;
							assign node179 = (inp[3]) ? node181 : 3'b110;
								assign node181 = (inp[4]) ? 3'b010 : 3'b110;
							assign node184 = (inp[0]) ? node186 : 3'b010;
								assign node186 = (inp[3]) ? node188 : 3'b010;
									assign node188 = (inp[4]) ? node190 : 3'b010;
										assign node190 = (inp[5]) ? 3'b100 : 3'b010;
				assign node193 = (inp[7]) ? node201 : node194;
					assign node194 = (inp[11]) ? node198 : node195;
						assign node195 = (inp[8]) ? 3'b010 : 3'b110;
						assign node198 = (inp[8]) ? 3'b100 : 3'b010;
					assign node201 = (inp[11]) ? 3'b000 : node202;
						assign node202 = (inp[0]) ? node204 : 3'b100;
							assign node204 = (inp[8]) ? node206 : 3'b100;
								assign node206 = (inp[5]) ? node208 : 3'b100;
									assign node208 = (inp[3]) ? node210 : 3'b100;
										assign node210 = (inp[4]) ? 3'b000 : 3'b100;
		assign node214 = (inp[6]) ? node282 : node215;
			assign node215 = (inp[10]) ? node267 : node216;
				assign node216 = (inp[8]) ? node242 : node217;
					assign node217 = (inp[7]) ? node239 : node218;
						assign node218 = (inp[4]) ? node226 : node219;
							assign node219 = (inp[11]) ? 3'b001 : node220;
								assign node220 = (inp[3]) ? node222 : 3'b101;
									assign node222 = (inp[2]) ? 3'b001 : 3'b101;
							assign node226 = (inp[11]) ? node236 : node227;
								assign node227 = (inp[3]) ? node229 : 3'b101;
									assign node229 = (inp[2]) ? 3'b001 : node230;
										assign node230 = (inp[0]) ? node232 : 3'b101;
											assign node232 = (inp[5]) ? 3'b001 : 3'b101;
								assign node236 = (inp[3]) ? 3'b110 : 3'b101;
						assign node239 = (inp[11]) ? 3'b100 : 3'b010;
					assign node242 = (inp[7]) ? node254 : node243;
						assign node243 = (inp[11]) ? node245 : 3'b000;
							assign node245 = (inp[4]) ? node247 : 3'b010;
								assign node247 = (inp[0]) ? node249 : 3'b010;
									assign node249 = (inp[5]) ? node251 : 3'b010;
										assign node251 = (inp[3]) ? 3'b101 : 3'b110;
						assign node254 = (inp[11]) ? node264 : node255;
							assign node255 = (inp[3]) ? node257 : 3'b010;
								assign node257 = (inp[2]) ? 3'b100 : node258;
									assign node258 = (inp[5]) ? node260 : 3'b010;
										assign node260 = (inp[0]) ? 3'b100 : 3'b010;
							assign node264 = (inp[4]) ? 3'b000 : 3'b100;
				assign node267 = (inp[7]) ? 3'b000 : node268;
					assign node268 = (inp[8]) ? node278 : node269;
						assign node269 = (inp[11]) ? node271 : 3'b010;
							assign node271 = (inp[5]) ? node273 : 3'b100;
								assign node273 = (inp[0]) ? node275 : 3'b100;
									assign node275 = (inp[4]) ? 3'b000 : 3'b100;
						assign node278 = (inp[11]) ? 3'b000 : 3'b100;
			assign node282 = (inp[10]) ? 3'b000 : node283;
				assign node283 = (inp[11]) ? 3'b000 : node284;
					assign node284 = (inp[8]) ? 3'b000 : node285;
						assign node285 = (inp[7]) ? 3'b000 : 3'b100;

endmodule