module dtc_split66_bm55 (
	input  wire [8-1:0] inp,
	output wire [7-1:0] outp
);

	wire [7-1:0] node1;
	wire [7-1:0] node2;
	wire [7-1:0] node3;
	wire [7-1:0] node4;
	wire [7-1:0] node5;
	wire [7-1:0] node6;
	wire [7-1:0] node9;
	wire [7-1:0] node12;
	wire [7-1:0] node13;
	wire [7-1:0] node16;
	wire [7-1:0] node19;
	wire [7-1:0] node20;
	wire [7-1:0] node22;
	wire [7-1:0] node25;
	wire [7-1:0] node26;
	wire [7-1:0] node30;
	wire [7-1:0] node31;
	wire [7-1:0] node32;
	wire [7-1:0] node33;
	wire [7-1:0] node36;
	wire [7-1:0] node39;
	wire [7-1:0] node40;
	wire [7-1:0] node44;
	wire [7-1:0] node45;
	wire [7-1:0] node46;
	wire [7-1:0] node49;
	wire [7-1:0] node52;
	wire [7-1:0] node53;
	wire [7-1:0] node56;
	wire [7-1:0] node59;
	wire [7-1:0] node60;
	wire [7-1:0] node61;
	wire [7-1:0] node62;
	wire [7-1:0] node63;
	wire [7-1:0] node66;
	wire [7-1:0] node69;
	wire [7-1:0] node71;
	wire [7-1:0] node74;
	wire [7-1:0] node75;
	wire [7-1:0] node76;
	wire [7-1:0] node79;
	wire [7-1:0] node82;
	wire [7-1:0] node85;
	wire [7-1:0] node86;
	wire [7-1:0] node87;
	wire [7-1:0] node88;
	wire [7-1:0] node91;
	wire [7-1:0] node94;
	wire [7-1:0] node96;
	wire [7-1:0] node99;
	wire [7-1:0] node100;
	wire [7-1:0] node101;
	wire [7-1:0] node104;
	wire [7-1:0] node107;
	wire [7-1:0] node108;
	wire [7-1:0] node111;
	wire [7-1:0] node114;
	wire [7-1:0] node115;
	wire [7-1:0] node116;
	wire [7-1:0] node117;
	wire [7-1:0] node118;
	wire [7-1:0] node119;
	wire [7-1:0] node122;
	wire [7-1:0] node125;
	wire [7-1:0] node126;
	wire [7-1:0] node130;
	wire [7-1:0] node131;
	wire [7-1:0] node132;
	wire [7-1:0] node135;
	wire [7-1:0] node138;
	wire [7-1:0] node140;
	wire [7-1:0] node143;
	wire [7-1:0] node144;
	wire [7-1:0] node145;
	wire [7-1:0] node146;
	wire [7-1:0] node149;
	wire [7-1:0] node152;
	wire [7-1:0] node153;
	wire [7-1:0] node156;
	wire [7-1:0] node159;
	wire [7-1:0] node160;
	wire [7-1:0] node161;
	wire [7-1:0] node164;
	wire [7-1:0] node167;
	wire [7-1:0] node168;
	wire [7-1:0] node171;
	wire [7-1:0] node174;
	wire [7-1:0] node175;
	wire [7-1:0] node176;
	wire [7-1:0] node177;
	wire [7-1:0] node178;
	wire [7-1:0] node181;
	wire [7-1:0] node184;
	wire [7-1:0] node186;
	wire [7-1:0] node189;
	wire [7-1:0] node190;
	wire [7-1:0] node191;
	wire [7-1:0] node194;
	wire [7-1:0] node197;
	wire [7-1:0] node198;
	wire [7-1:0] node201;
	wire [7-1:0] node204;
	wire [7-1:0] node205;
	wire [7-1:0] node206;
	wire [7-1:0] node207;
	wire [7-1:0] node210;
	wire [7-1:0] node213;
	wire [7-1:0] node214;
	wire [7-1:0] node218;
	wire [7-1:0] node219;
	wire [7-1:0] node220;
	wire [7-1:0] node223;
	wire [7-1:0] node226;
	wire [7-1:0] node227;

	assign outp = (inp[2]) ? node114 : node1;
		assign node1 = (inp[6]) ? node59 : node2;
			assign node2 = (inp[4]) ? node30 : node3;
				assign node3 = (inp[5]) ? node19 : node4;
					assign node4 = (inp[0]) ? node12 : node5;
						assign node5 = (inp[3]) ? node9 : node6;
							assign node6 = (inp[7]) ? 7'b0110111 : 7'b0110101;
							assign node9 = (inp[7]) ? 7'b0111100 : 7'b0110110;
						assign node12 = (inp[1]) ? node16 : node13;
							assign node13 = (inp[7]) ? 7'b1110100 : 7'b0010100;
							assign node16 = (inp[3]) ? 7'b1101101 : 7'b1100100;
					assign node19 = (inp[1]) ? node25 : node20;
						assign node20 = (inp[3]) ? node22 : 7'b0100101;
							assign node22 = (inp[7]) ? 7'b0100100 : 7'b0101100;
						assign node25 = (inp[0]) ? 7'b1111100 : node26;
							assign node26 = (inp[7]) ? 7'b0100100 : 7'b1100100;
				assign node30 = (inp[3]) ? node44 : node31;
					assign node31 = (inp[0]) ? node39 : node32;
						assign node32 = (inp[5]) ? node36 : node33;
							assign node33 = (inp[1]) ? 7'b0001100 : 7'b0011101;
							assign node36 = (inp[1]) ? 7'b0010101 : 7'b0000101;
						assign node39 = (inp[5]) ? 7'b1100100 : node40;
							assign node40 = (inp[1]) ? 7'b1011101 : 7'b0111100;
					assign node44 = (inp[5]) ? node52 : node45;
						assign node45 = (inp[7]) ? node49 : node46;
							assign node46 = (inp[1]) ? 7'b0000110 : 7'b1011110;
							assign node49 = (inp[1]) ? 7'b1000100 : 7'b1000101;
						assign node52 = (inp[7]) ? node56 : node53;
							assign node53 = (inp[0]) ? 7'b0010100 : 7'b1001100;
							assign node56 = (inp[1]) ? 7'b0000100 : 7'b0000100;
			assign node59 = (inp[0]) ? node85 : node60;
				assign node60 = (inp[4]) ? node74 : node61;
					assign node61 = (inp[1]) ? node69 : node62;
						assign node62 = (inp[5]) ? node66 : node63;
							assign node63 = (inp[3]) ? 7'b1000100 : 7'b1010101;
							assign node66 = (inp[3]) ? 7'b0000100 : 7'b0000101;
						assign node69 = (inp[3]) ? node71 : 7'b1111011;
							assign node71 = (inp[5]) ? 7'b0100001 : 7'b0111001;
					assign node74 = (inp[1]) ? node82 : node75;
						assign node75 = (inp[3]) ? node79 : node76;
							assign node76 = (inp[5]) ? 7'b0110000 : 7'b1101010;
							assign node79 = (inp[5]) ? 7'b0110001 : 7'b1110001;
						assign node82 = (inp[7]) ? 7'b0100000 : 7'b1110000;
				assign node85 = (inp[1]) ? node99 : node86;
					assign node86 = (inp[3]) ? node94 : node87;
						assign node87 = (inp[4]) ? node91 : node88;
							assign node88 = (inp[7]) ? 7'b0100010 : 7'b1110000;
							assign node91 = (inp[5]) ? 7'b1000001 : 7'b1001011;
						assign node94 = (inp[7]) ? node96 : 7'b1001001;
							assign node96 = (inp[4]) ? 7'b0000001 : 7'b0010001;
					assign node99 = (inp[3]) ? node107 : node100;
						assign node100 = (inp[4]) ? node104 : node101;
							assign node101 = (inp[5]) ? 7'b1000000 : 7'b0000000;
							assign node104 = (inp[7]) ? 7'b0000000 : 7'b0011000;
						assign node107 = (inp[5]) ? node111 : node108;
							assign node108 = (inp[4]) ? 7'b0010010 : 7'b0011000;
							assign node111 = (inp[7]) ? 7'b0000000 : 7'b0010000;
		assign node114 = (inp[5]) ? node174 : node115;
			assign node115 = (inp[6]) ? node143 : node116;
				assign node116 = (inp[0]) ? node130 : node117;
					assign node117 = (inp[1]) ? node125 : node118;
						assign node118 = (inp[4]) ? node122 : node119;
							assign node119 = (inp[7]) ? 7'b0100001 : 7'b0110001;
							assign node122 = (inp[7]) ? 7'b0111011 : 7'b0101000;
						assign node125 = (inp[7]) ? 7'b1110010 : node126;
							assign node126 = (inp[3]) ? 7'b1111010 : 7'b0101001;
					assign node130 = (inp[1]) ? node138 : node131;
						assign node131 = (inp[7]) ? node135 : node132;
							assign node132 = (inp[4]) ? 7'b0001001 : 7'b0100010;
							assign node135 = (inp[4]) ? 7'b0011010 : 7'b1011001;
						assign node138 = (inp[4]) ? node140 : 7'b1011011;
							assign node140 = (inp[3]) ? 7'b1000000 : 7'b1011000;
				assign node143 = (inp[0]) ? node159 : node144;
					assign node144 = (inp[4]) ? node152 : node145;
						assign node145 = (inp[3]) ? node149 : node146;
							assign node146 = (inp[7]) ? 7'b1010011 : 7'b1010001;
							assign node149 = (inp[1]) ? 7'b0001001 : 7'b1000011;
						assign node152 = (inp[1]) ? node156 : node153;
							assign node153 = (inp[7]) ? 7'b1010000 : 7'b0001000;
							assign node156 = (inp[7]) ? 7'b0000000 : 7'b1000000;
					assign node159 = (inp[1]) ? node167 : node160;
						assign node160 = (inp[4]) ? node164 : node161;
							assign node161 = (inp[3]) ? 7'b1010010 : 7'b0010010;
							assign node164 = (inp[7]) ? 7'b1001010 : 7'b0001010;
						assign node167 = (inp[4]) ? node171 : node168;
							assign node168 = (inp[7]) ? 7'b0001000 : 7'b0001010;
							assign node171 = (inp[3]) ? 7'b0000000 : 7'b0000000;
			assign node174 = (inp[6]) ? node204 : node175;
				assign node175 = (inp[0]) ? node189 : node176;
					assign node176 = (inp[7]) ? node184 : node177;
						assign node177 = (inp[1]) ? node181 : node178;
							assign node178 = (inp[3]) ? 7'b0111001 : 7'b0110001;
							assign node181 = (inp[3]) ? 7'b1110000 : 7'b0111000;
						assign node184 = (inp[1]) ? node186 : 7'b0100001;
							assign node186 = (inp[3]) ? 7'b0100000 : 7'b0100000;
					assign node189 = (inp[4]) ? node197 : node190;
						assign node190 = (inp[3]) ? node194 : node191;
							assign node191 = (inp[1]) ? 7'b1000001 : 7'b0100000;
							assign node194 = (inp[1]) ? 7'b0000001 : 7'b0010001;
						assign node197 = (inp[3]) ? node201 : node198;
							assign node198 = (inp[1]) ? 7'b0010000 : 7'b1010000;
							assign node201 = (inp[7]) ? 7'b0000000 : 7'b0001000;
				assign node204 = (inp[4]) ? node218 : node205;
					assign node205 = (inp[0]) ? node213 : node206;
						assign node206 = (inp[3]) ? node210 : node207;
							assign node207 = (inp[1]) ? 7'b0010001 : 7'b0010001;
							assign node210 = (inp[7]) ? 7'b0000001 : 7'b0000001;
						assign node213 = (inp[1]) ? 7'b0000000 : node214;
							assign node214 = (inp[7]) ? 7'b0010000 : 7'b1011000;
					assign node218 = (inp[1]) ? node226 : node219;
						assign node219 = (inp[7]) ? node223 : node220;
							assign node220 = (inp[0]) ? 7'b1000000 : 7'b0000001;
							assign node223 = (inp[3]) ? 7'b0010000 : 7'b1010000;
						assign node226 = (inp[7]) ? 7'b0000000 : node227;
							assign node227 = (inp[3]) ? 7'b0000000 : 7'b0001000;

endmodule