module dtc_split875_bm73 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node104;

	assign outp = (inp[9]) ? node46 : node1;
		assign node1 = (inp[3]) ? node31 : node2;
			assign node2 = (inp[6]) ? node18 : node3;
				assign node3 = (inp[4]) ? node11 : node4;
					assign node4 = (inp[7]) ? node8 : node5;
						assign node5 = (inp[10]) ? 3'b111 : 3'b101;
						assign node8 = (inp[10]) ? 3'b101 : 3'b110;
					assign node11 = (inp[7]) ? node15 : node12;
						assign node12 = (inp[10]) ? 3'b101 : 3'b110;
						assign node15 = (inp[10]) ? 3'b010 : 3'b000;
				assign node18 = (inp[10]) ? node24 : node19;
					assign node19 = (inp[4]) ? 3'b000 : node20;
						assign node20 = (inp[7]) ? 3'b000 : 3'b000;
					assign node24 = (inp[7]) ? node28 : node25;
						assign node25 = (inp[4]) ? 3'b000 : 3'b010;
						assign node28 = (inp[4]) ? 3'b000 : 3'b000;
			assign node31 = (inp[6]) ? 3'b000 : node32;
				assign node32 = (inp[10]) ? node38 : node33;
					assign node33 = (inp[4]) ? 3'b000 : node34;
						assign node34 = (inp[7]) ? 3'b000 : 3'b000;
					assign node38 = (inp[4]) ? node42 : node39;
						assign node39 = (inp[7]) ? 3'b000 : 3'b010;
						assign node42 = (inp[7]) ? 3'b000 : 3'b000;
		assign node46 = (inp[3]) ? node76 : node47;
			assign node47 = (inp[6]) ? node61 : node48;
				assign node48 = (inp[10]) ? node56 : node49;
					assign node49 = (inp[4]) ? node53 : node50;
						assign node50 = (inp[7]) ? 3'b111 : 3'b111;
						assign node53 = (inp[7]) ? 3'b101 : 3'b111;
					assign node56 = (inp[4]) ? node58 : 3'b111;
						assign node58 = (inp[7]) ? 3'b111 : 3'b111;
				assign node61 = (inp[10]) ? node69 : node62;
					assign node62 = (inp[4]) ? node66 : node63;
						assign node63 = (inp[7]) ? 3'b010 : 3'b101;
						assign node66 = (inp[7]) ? 3'b000 : 3'b010;
					assign node69 = (inp[4]) ? node73 : node70;
						assign node70 = (inp[7]) ? 3'b001 : 3'b111;
						assign node73 = (inp[7]) ? 3'b110 : 3'b101;
			assign node76 = (inp[6]) ? node92 : node77;
				assign node77 = (inp[10]) ? node85 : node78;
					assign node78 = (inp[7]) ? node82 : node79;
						assign node79 = (inp[4]) ? 3'b110 : 3'b101;
						assign node82 = (inp[4]) ? 3'b000 : 3'b010;
					assign node85 = (inp[4]) ? node89 : node86;
						assign node86 = (inp[7]) ? 3'b001 : 3'b111;
						assign node89 = (inp[7]) ? 3'b110 : 3'b101;
				assign node92 = (inp[10]) ? node100 : node93;
					assign node93 = (inp[4]) ? node97 : node94;
						assign node94 = (inp[7]) ? 3'b000 : 3'b000;
						assign node97 = (inp[7]) ? 3'b000 : 3'b000;
					assign node100 = (inp[4]) ? node104 : node101;
						assign node101 = (inp[7]) ? 3'b100 : 3'b010;
						assign node104 = (inp[7]) ? 3'b000 : 3'b000;

endmodule