module dtc_split25_bm21 (
	input  wire [10-1:0] inp,
	output wire [10-1:0] outp
);

	wire [10-1:0] node1;
	wire [10-1:0] node2;
	wire [10-1:0] node3;
	wire [10-1:0] node4;
	wire [10-1:0] node5;
	wire [10-1:0] node6;
	wire [10-1:0] node7;
	wire [10-1:0] node10;
	wire [10-1:0] node13;
	wire [10-1:0] node15;
	wire [10-1:0] node18;
	wire [10-1:0] node19;
	wire [10-1:0] node20;
	wire [10-1:0] node24;
	wire [10-1:0] node27;
	wire [10-1:0] node28;
	wire [10-1:0] node29;
	wire [10-1:0] node30;
	wire [10-1:0] node34;
	wire [10-1:0] node37;
	wire [10-1:0] node38;
	wire [10-1:0] node42;
	wire [10-1:0] node43;
	wire [10-1:0] node44;
	wire [10-1:0] node45;
	wire [10-1:0] node47;
	wire [10-1:0] node50;
	wire [10-1:0] node51;
	wire [10-1:0] node55;
	wire [10-1:0] node56;
	wire [10-1:0] node57;
	wire [10-1:0] node60;
	wire [10-1:0] node63;
	wire [10-1:0] node64;
	wire [10-1:0] node68;
	wire [10-1:0] node69;
	wire [10-1:0] node70;
	wire [10-1:0] node71;
	wire [10-1:0] node74;
	wire [10-1:0] node77;
	wire [10-1:0] node78;
	wire [10-1:0] node82;
	wire [10-1:0] node83;
	wire [10-1:0] node84;
	wire [10-1:0] node88;
	wire [10-1:0] node89;
	wire [10-1:0] node93;
	wire [10-1:0] node94;
	wire [10-1:0] node95;
	wire [10-1:0] node96;
	wire [10-1:0] node97;
	wire [10-1:0] node99;
	wire [10-1:0] node103;
	wire [10-1:0] node104;
	wire [10-1:0] node105;
	wire [10-1:0] node109;
	wire [10-1:0] node112;
	wire [10-1:0] node113;
	wire [10-1:0] node114;
	wire [10-1:0] node117;
	wire [10-1:0] node119;
	wire [10-1:0] node122;
	wire [10-1:0] node123;
	wire [10-1:0] node124;
	wire [10-1:0] node127;
	wire [10-1:0] node130;
	wire [10-1:0] node131;
	wire [10-1:0] node134;
	wire [10-1:0] node137;
	wire [10-1:0] node138;
	wire [10-1:0] node139;
	wire [10-1:0] node141;
	wire [10-1:0] node142;
	wire [10-1:0] node145;
	wire [10-1:0] node148;
	wire [10-1:0] node150;
	wire [10-1:0] node151;
	wire [10-1:0] node155;
	wire [10-1:0] node156;
	wire [10-1:0] node157;
	wire [10-1:0] node158;
	wire [10-1:0] node162;
	wire [10-1:0] node163;
	wire [10-1:0] node166;
	wire [10-1:0] node169;
	wire [10-1:0] node170;
	wire [10-1:0] node174;
	wire [10-1:0] node175;
	wire [10-1:0] node176;
	wire [10-1:0] node177;
	wire [10-1:0] node178;
	wire [10-1:0] node179;
	wire [10-1:0] node180;
	wire [10-1:0] node183;
	wire [10-1:0] node186;
	wire [10-1:0] node187;
	wire [10-1:0] node191;
	wire [10-1:0] node192;
	wire [10-1:0] node195;
	wire [10-1:0] node196;
	wire [10-1:0] node200;
	wire [10-1:0] node201;
	wire [10-1:0] node202;
	wire [10-1:0] node205;
	wire [10-1:0] node206;
	wire [10-1:0] node209;
	wire [10-1:0] node212;
	wire [10-1:0] node214;
	wire [10-1:0] node216;
	wire [10-1:0] node219;
	wire [10-1:0] node220;
	wire [10-1:0] node221;
	wire [10-1:0] node224;
	wire [10-1:0] node225;
	wire [10-1:0] node226;
	wire [10-1:0] node229;
	wire [10-1:0] node232;
	wire [10-1:0] node233;
	wire [10-1:0] node236;
	wire [10-1:0] node239;
	wire [10-1:0] node240;
	wire [10-1:0] node241;
	wire [10-1:0] node243;
	wire [10-1:0] node247;
	wire [10-1:0] node248;
	wire [10-1:0] node250;
	wire [10-1:0] node253;
	wire [10-1:0] node254;
	wire [10-1:0] node258;
	wire [10-1:0] node259;
	wire [10-1:0] node260;
	wire [10-1:0] node261;
	wire [10-1:0] node262;
	wire [10-1:0] node264;
	wire [10-1:0] node267;
	wire [10-1:0] node269;
	wire [10-1:0] node272;
	wire [10-1:0] node273;
	wire [10-1:0] node276;
	wire [10-1:0] node279;
	wire [10-1:0] node280;
	wire [10-1:0] node281;
	wire [10-1:0] node282;
	wire [10-1:0] node285;
	wire [10-1:0] node288;
	wire [10-1:0] node289;
	wire [10-1:0] node292;
	wire [10-1:0] node295;
	wire [10-1:0] node296;
	wire [10-1:0] node298;
	wire [10-1:0] node301;
	wire [10-1:0] node302;
	wire [10-1:0] node305;
	wire [10-1:0] node308;
	wire [10-1:0] node309;
	wire [10-1:0] node310;
	wire [10-1:0] node311;
	wire [10-1:0] node314;
	wire [10-1:0] node315;
	wire [10-1:0] node319;
	wire [10-1:0] node320;
	wire [10-1:0] node321;
	wire [10-1:0] node325;
	wire [10-1:0] node328;
	wire [10-1:0] node329;
	wire [10-1:0] node332;
	wire [10-1:0] node333;

	assign outp = (inp[1]) ? node174 : node1;
		assign node1 = (inp[6]) ? node93 : node2;
			assign node2 = (inp[4]) ? node42 : node3;
				assign node3 = (inp[3]) ? node27 : node4;
					assign node4 = (inp[8]) ? node18 : node5;
						assign node5 = (inp[7]) ? node13 : node6;
							assign node6 = (inp[9]) ? node10 : node7;
								assign node7 = (inp[5]) ? 10'b0011111111 : 10'b0111111111;
								assign node10 = (inp[0]) ? 10'b0001111111 : 10'b0011111111;
							assign node13 = (inp[2]) ? node15 : 10'b0011111111;
								assign node15 = (inp[9]) ? 10'b0000111111 : 10'b0001111111;
						assign node18 = (inp[9]) ? node24 : node19;
							assign node19 = (inp[5]) ? 10'b0001111111 : node20;
								assign node20 = (inp[7]) ? 10'b0001111111 : 10'b0011111111;
							assign node24 = (inp[7]) ? 10'b0000011111 : 10'b0001111111;
					assign node27 = (inp[2]) ? node37 : node28;
						assign node28 = (inp[9]) ? node34 : node29;
							assign node29 = (inp[8]) ? 10'b0001111111 : node30;
								assign node30 = (inp[0]) ? 10'b0001111111 : 10'b0011111111;
							assign node34 = (inp[7]) ? 10'b0000111111 : 10'b0000011111;
						assign node37 = (inp[0]) ? 10'b0000011111 : node38;
							assign node38 = (inp[7]) ? 10'b0000011111 : 10'b0000111111;
				assign node42 = (inp[8]) ? node68 : node43;
					assign node43 = (inp[9]) ? node55 : node44;
						assign node44 = (inp[3]) ? node50 : node45;
							assign node45 = (inp[2]) ? node47 : 10'b0001111111;
								assign node47 = (inp[5]) ? 10'b0001111111 : 10'b0011111111;
							assign node50 = (inp[5]) ? 10'b0000011111 : node51;
								assign node51 = (inp[2]) ? 10'b0000111111 : 10'b0001111111;
						assign node55 = (inp[2]) ? node63 : node56;
							assign node56 = (inp[5]) ? node60 : node57;
								assign node57 = (inp[7]) ? 10'b0000111111 : 10'b0001111111;
								assign node60 = (inp[0]) ? 10'b0000011111 : 10'b0000111111;
							assign node63 = (inp[5]) ? 10'b0000011111 : node64;
								assign node64 = (inp[0]) ? 10'b0000011111 : 10'b0000111111;
					assign node68 = (inp[5]) ? node82 : node69;
						assign node69 = (inp[7]) ? node77 : node70;
							assign node70 = (inp[2]) ? node74 : node71;
								assign node71 = (inp[0]) ? 10'b0000111111 : 10'b0000111111;
								assign node74 = (inp[3]) ? 10'b0000011111 : 10'b0000111111;
							assign node77 = (inp[3]) ? 10'b0000011111 : node78;
								assign node78 = (inp[2]) ? 10'b0000011111 : 10'b0000111111;
						assign node82 = (inp[0]) ? node88 : node83;
							assign node83 = (inp[7]) ? 10'b0000001111 : node84;
								assign node84 = (inp[9]) ? 10'b0000011111 : 10'b0000011111;
							assign node88 = (inp[2]) ? 10'b0000000111 : node89;
								assign node89 = (inp[3]) ? 10'b0000000111 : 10'b0000001111;
			assign node93 = (inp[8]) ? node137 : node94;
				assign node94 = (inp[7]) ? node112 : node95;
					assign node95 = (inp[2]) ? node103 : node96;
						assign node96 = (inp[0]) ? 10'b0000111111 : node97;
							assign node97 = (inp[3]) ? node99 : 10'b0011111111;
								assign node99 = (inp[5]) ? 10'b0001111111 : 10'b0001111111;
						assign node103 = (inp[5]) ? node109 : node104;
							assign node104 = (inp[9]) ? 10'b0000111111 : node105;
								assign node105 = (inp[4]) ? 10'b0000111111 : 10'b0001111111;
							assign node109 = (inp[4]) ? 10'b0000011111 : 10'b0000111111;
					assign node112 = (inp[9]) ? node122 : node113;
						assign node113 = (inp[5]) ? node117 : node114;
							assign node114 = (inp[2]) ? 10'b0000111111 : 10'b0001111111;
							assign node117 = (inp[0]) ? node119 : 10'b0000111111;
								assign node119 = (inp[2]) ? 10'b0000001111 : 10'b0000011111;
						assign node122 = (inp[4]) ? node130 : node123;
							assign node123 = (inp[3]) ? node127 : node124;
								assign node124 = (inp[2]) ? 10'b0000011111 : 10'b0000111111;
								assign node127 = (inp[0]) ? 10'b0000001111 : 10'b0000011111;
							assign node130 = (inp[5]) ? node134 : node131;
								assign node131 = (inp[2]) ? 10'b0000001111 : 10'b0000011111;
								assign node134 = (inp[3]) ? 10'b0000000111 : 10'b0000001111;
				assign node137 = (inp[3]) ? node155 : node138;
					assign node138 = (inp[9]) ? node148 : node139;
						assign node139 = (inp[4]) ? node141 : 10'b0000111111;
							assign node141 = (inp[5]) ? node145 : node142;
								assign node142 = (inp[7]) ? 10'b0000011111 : 10'b0000111111;
								assign node145 = (inp[2]) ? 10'b0000000111 : 10'b0000001111;
						assign node148 = (inp[7]) ? node150 : 10'b0000011111;
							assign node150 = (inp[2]) ? 10'b0000001111 : node151;
								assign node151 = (inp[4]) ? 10'b0000001111 : 10'b0000011111;
					assign node155 = (inp[9]) ? node169 : node156;
						assign node156 = (inp[0]) ? node162 : node157;
							assign node157 = (inp[2]) ? 10'b0000001111 : node158;
								assign node158 = (inp[5]) ? 10'b0000011111 : 10'b0000111111;
							assign node162 = (inp[5]) ? node166 : node163;
								assign node163 = (inp[7]) ? 10'b0000001111 : 10'b0000011111;
								assign node166 = (inp[4]) ? 10'b0000000111 : 10'b0000001111;
						assign node169 = (inp[5]) ? 10'b0000000111 : node170;
							assign node170 = (inp[2]) ? 10'b0000000111 : 10'b0000001111;
		assign node174 = (inp[4]) ? node258 : node175;
			assign node175 = (inp[7]) ? node219 : node176;
				assign node176 = (inp[5]) ? node200 : node177;
					assign node177 = (inp[6]) ? node191 : node178;
						assign node178 = (inp[0]) ? node186 : node179;
							assign node179 = (inp[8]) ? node183 : node180;
								assign node180 = (inp[2]) ? 10'b0001111111 : 10'b0011111111;
								assign node183 = (inp[3]) ? 10'b0000111111 : 10'b0001111111;
							assign node186 = (inp[8]) ? 10'b0000111111 : node187;
								assign node187 = (inp[9]) ? 10'b0000111111 : 10'b0001111111;
						assign node191 = (inp[8]) ? node195 : node192;
							assign node192 = (inp[2]) ? 10'b0000111111 : 10'b0001111111;
							assign node195 = (inp[9]) ? 10'b0000001111 : node196;
								assign node196 = (inp[3]) ? 10'b0000111111 : 10'b0000011111;
					assign node200 = (inp[2]) ? node212 : node201;
						assign node201 = (inp[8]) ? node205 : node202;
							assign node202 = (inp[6]) ? 10'b0000111111 : 10'b0001111111;
							assign node205 = (inp[6]) ? node209 : node206;
								assign node206 = (inp[3]) ? 10'b0000011111 : 10'b0000111111;
								assign node209 = (inp[9]) ? 10'b0000001111 : 10'b0000011111;
						assign node212 = (inp[9]) ? node214 : 10'b0000011111;
							assign node214 = (inp[8]) ? node216 : 10'b0000011111;
								assign node216 = (inp[6]) ? 10'b0000001111 : 10'b0000000111;
				assign node219 = (inp[0]) ? node239 : node220;
					assign node220 = (inp[2]) ? node224 : node221;
						assign node221 = (inp[5]) ? 10'b0000111111 : 10'b0001111111;
						assign node224 = (inp[3]) ? node232 : node225;
							assign node225 = (inp[9]) ? node229 : node226;
								assign node226 = (inp[6]) ? 10'b0000011111 : 10'b0000111111;
								assign node229 = (inp[6]) ? 10'b0000001111 : 10'b0000011111;
							assign node232 = (inp[6]) ? node236 : node233;
								assign node233 = (inp[5]) ? 10'b0000001111 : 10'b0000001111;
								assign node236 = (inp[8]) ? 10'b0000000111 : 10'b0000001111;
					assign node239 = (inp[8]) ? node247 : node240;
						assign node240 = (inp[5]) ? 10'b0000001111 : node241;
							assign node241 = (inp[6]) ? node243 : 10'b0000111111;
								assign node243 = (inp[9]) ? 10'b0000001111 : 10'b0000011111;
						assign node247 = (inp[5]) ? node253 : node248;
							assign node248 = (inp[3]) ? node250 : 10'b0000001111;
								assign node250 = (inp[2]) ? 10'b0000000011 : 10'b0000001111;
							assign node253 = (inp[9]) ? 10'b0000000111 : node254;
								assign node254 = (inp[3]) ? 10'b0000000111 : 10'b0000011111;
			assign node258 = (inp[2]) ? node308 : node259;
				assign node259 = (inp[9]) ? node279 : node260;
					assign node260 = (inp[3]) ? node272 : node261;
						assign node261 = (inp[6]) ? node267 : node262;
							assign node262 = (inp[8]) ? node264 : 10'b0000111111;
								assign node264 = (inp[5]) ? 10'b0000011111 : 10'b0000111111;
							assign node267 = (inp[0]) ? node269 : 10'b0000111111;
								assign node269 = (inp[5]) ? 10'b0000001111 : 10'b0000011111;
						assign node272 = (inp[0]) ? node276 : node273;
							assign node273 = (inp[8]) ? 10'b0000011111 : 10'b0000001111;
							assign node276 = (inp[6]) ? 10'b0000000111 : 10'b0000001111;
					assign node279 = (inp[8]) ? node295 : node280;
						assign node280 = (inp[5]) ? node288 : node281;
							assign node281 = (inp[7]) ? node285 : node282;
								assign node282 = (inp[3]) ? 10'b0000011111 : 10'b0000111111;
								assign node285 = (inp[3]) ? 10'b0000001111 : 10'b0000011111;
							assign node288 = (inp[6]) ? node292 : node289;
								assign node289 = (inp[3]) ? 10'b0000001111 : 10'b0000011111;
								assign node292 = (inp[0]) ? 10'b0000000111 : 10'b0000001111;
						assign node295 = (inp[5]) ? node301 : node296;
							assign node296 = (inp[7]) ? node298 : 10'b0000001111;
								assign node298 = (inp[0]) ? 10'b0000000111 : 10'b0000001111;
							assign node301 = (inp[7]) ? node305 : node302;
								assign node302 = (inp[0]) ? 10'b0000000111 : 10'b0000001111;
								assign node305 = (inp[0]) ? 10'b0000000011 : 10'b0000000111;
				assign node308 = (inp[9]) ? node328 : node309;
					assign node309 = (inp[0]) ? node319 : node310;
						assign node310 = (inp[3]) ? node314 : node311;
							assign node311 = (inp[6]) ? 10'b0000001111 : 10'b0000011111;
							assign node314 = (inp[7]) ? 10'b0000001111 : node315;
								assign node315 = (inp[8]) ? 10'b0000000111 : 10'b0000011111;
						assign node319 = (inp[5]) ? node325 : node320;
							assign node320 = (inp[6]) ? 10'b0000011111 : node321;
								assign node321 = (inp[8]) ? 10'b0000000111 : 10'b0000001111;
							assign node325 = (inp[3]) ? 10'b0000000011 : 10'b0000000111;
					assign node328 = (inp[7]) ? node332 : node329;
						assign node329 = (inp[0]) ? 10'b0000000011 : 10'b0000000111;
						assign node332 = (inp[8]) ? 10'b0000000011 : node333;
							assign node333 = (inp[5]) ? 10'b0000000011 : 10'b0000001111;

endmodule