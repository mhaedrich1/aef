module dtc_split875_bm80 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node171;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node195;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node212;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node257;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node274;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node296;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node333;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node343;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node356;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node377;
	wire [3-1:0] node380;
	wire [3-1:0] node382;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node388;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node401;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node431;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node464;
	wire [3-1:0] node468;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node488;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node495;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node517;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node524;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node541;
	wire [3-1:0] node544;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node552;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node574;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node580;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node608;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node622;
	wire [3-1:0] node625;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node651;
	wire [3-1:0] node653;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node659;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node669;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node690;
	wire [3-1:0] node693;
	wire [3-1:0] node695;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node705;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node734;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node739;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node748;
	wire [3-1:0] node750;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node756;
	wire [3-1:0] node759;
	wire [3-1:0] node761;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node771;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node778;
	wire [3-1:0] node781;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node787;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node803;
	wire [3-1:0] node806;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node814;
	wire [3-1:0] node818;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node825;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node834;
	wire [3-1:0] node837;
	wire [3-1:0] node839;
	wire [3-1:0] node842;
	wire [3-1:0] node843;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node854;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node865;
	wire [3-1:0] node868;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node880;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node889;
	wire [3-1:0] node892;
	wire [3-1:0] node894;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node901;
	wire [3-1:0] node903;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node909;
	wire [3-1:0] node911;
	wire [3-1:0] node914;
	wire [3-1:0] node916;
	wire [3-1:0] node918;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node928;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node941;
	wire [3-1:0] node942;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node950;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node958;
	wire [3-1:0] node960;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node966;
	wire [3-1:0] node969;
	wire [3-1:0] node970;
	wire [3-1:0] node971;
	wire [3-1:0] node974;
	wire [3-1:0] node977;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node987;
	wire [3-1:0] node990;
	wire [3-1:0] node992;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node1001;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1008;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1016;
	wire [3-1:0] node1019;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1030;
	wire [3-1:0] node1032;
	wire [3-1:0] node1033;
	wire [3-1:0] node1036;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1043;
	wire [3-1:0] node1048;
	wire [3-1:0] node1049;
	wire [3-1:0] node1051;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1054;
	wire [3-1:0] node1057;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1067;
	wire [3-1:0] node1069;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1082;
	wire [3-1:0] node1083;
	wire [3-1:0] node1084;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1087;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1092;
	wire [3-1:0] node1095;
	wire [3-1:0] node1096;
	wire [3-1:0] node1100;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1105;
	wire [3-1:0] node1108;
	wire [3-1:0] node1109;
	wire [3-1:0] node1112;
	wire [3-1:0] node1115;
	wire [3-1:0] node1116;
	wire [3-1:0] node1117;
	wire [3-1:0] node1119;
	wire [3-1:0] node1122;
	wire [3-1:0] node1123;
	wire [3-1:0] node1126;
	wire [3-1:0] node1129;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1134;
	wire [3-1:0] node1137;
	wire [3-1:0] node1138;
	wire [3-1:0] node1142;
	wire [3-1:0] node1143;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1147;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1154;
	wire [3-1:0] node1157;
	wire [3-1:0] node1158;
	wire [3-1:0] node1159;
	wire [3-1:0] node1162;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1169;
	wire [3-1:0] node1172;
	wire [3-1:0] node1173;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1180;
	wire [3-1:0] node1181;
	wire [3-1:0] node1182;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1192;
	wire [3-1:0] node1194;
	wire [3-1:0] node1197;
	wire [3-1:0] node1198;
	wire [3-1:0] node1202;
	wire [3-1:0] node1203;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1210;
	wire [3-1:0] node1211;
	wire [3-1:0] node1215;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1219;
	wire [3-1:0] node1223;
	wire [3-1:0] node1225;
	wire [3-1:0] node1228;
	wire [3-1:0] node1229;
	wire [3-1:0] node1230;
	wire [3-1:0] node1234;
	wire [3-1:0] node1236;
	wire [3-1:0] node1239;
	wire [3-1:0] node1240;
	wire [3-1:0] node1241;
	wire [3-1:0] node1242;
	wire [3-1:0] node1246;
	wire [3-1:0] node1250;
	wire [3-1:0] node1251;
	wire [3-1:0] node1252;
	wire [3-1:0] node1253;
	wire [3-1:0] node1254;
	wire [3-1:0] node1256;
	wire [3-1:0] node1259;
	wire [3-1:0] node1260;
	wire [3-1:0] node1262;
	wire [3-1:0] node1267;
	wire [3-1:0] node1268;
	wire [3-1:0] node1269;
	wire [3-1:0] node1270;
	wire [3-1:0] node1273;
	wire [3-1:0] node1274;
	wire [3-1:0] node1278;
	wire [3-1:0] node1280;
	wire [3-1:0] node1281;
	wire [3-1:0] node1284;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1289;
	wire [3-1:0] node1293;
	wire [3-1:0] node1294;
	wire [3-1:0] node1295;
	wire [3-1:0] node1299;
	wire [3-1:0] node1302;
	wire [3-1:0] node1303;
	wire [3-1:0] node1304;
	wire [3-1:0] node1306;
	wire [3-1:0] node1307;
	wire [3-1:0] node1309;
	wire [3-1:0] node1315;
	wire [3-1:0] node1317;
	wire [3-1:0] node1318;
	wire [3-1:0] node1319;
	wire [3-1:0] node1320;
	wire [3-1:0] node1322;
	wire [3-1:0] node1325;
	wire [3-1:0] node1326;
	wire [3-1:0] node1327;
	wire [3-1:0] node1329;
	wire [3-1:0] node1330;
	wire [3-1:0] node1334;
	wire [3-1:0] node1336;
	wire [3-1:0] node1339;
	wire [3-1:0] node1341;
	wire [3-1:0] node1342;
	wire [3-1:0] node1346;
	wire [3-1:0] node1347;
	wire [3-1:0] node1348;
	wire [3-1:0] node1350;
	wire [3-1:0] node1352;
	wire [3-1:0] node1353;
	wire [3-1:0] node1360;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1363;
	wire [3-1:0] node1364;
	wire [3-1:0] node1365;
	wire [3-1:0] node1367;
	wire [3-1:0] node1368;
	wire [3-1:0] node1370;
	wire [3-1:0] node1372;
	wire [3-1:0] node1375;
	wire [3-1:0] node1376;
	wire [3-1:0] node1377;
	wire [3-1:0] node1381;
	wire [3-1:0] node1382;
	wire [3-1:0] node1384;
	wire [3-1:0] node1387;
	wire [3-1:0] node1389;
	wire [3-1:0] node1393;
	wire [3-1:0] node1394;
	wire [3-1:0] node1395;
	wire [3-1:0] node1396;
	wire [3-1:0] node1397;
	wire [3-1:0] node1399;
	wire [3-1:0] node1401;
	wire [3-1:0] node1404;
	wire [3-1:0] node1405;
	wire [3-1:0] node1407;
	wire [3-1:0] node1410;
	wire [3-1:0] node1411;
	wire [3-1:0] node1414;
	wire [3-1:0] node1417;
	wire [3-1:0] node1418;
	wire [3-1:0] node1419;
	wire [3-1:0] node1422;
	wire [3-1:0] node1424;
	wire [3-1:0] node1427;
	wire [3-1:0] node1428;
	wire [3-1:0] node1430;
	wire [3-1:0] node1433;
	wire [3-1:0] node1435;
	wire [3-1:0] node1438;
	wire [3-1:0] node1439;
	wire [3-1:0] node1440;
	wire [3-1:0] node1441;
	wire [3-1:0] node1442;
	wire [3-1:0] node1447;
	wire [3-1:0] node1448;
	wire [3-1:0] node1450;
	wire [3-1:0] node1454;
	wire [3-1:0] node1455;
	wire [3-1:0] node1456;
	wire [3-1:0] node1460;
	wire [3-1:0] node1461;
	wire [3-1:0] node1464;
	wire [3-1:0] node1466;
	wire [3-1:0] node1469;
	wire [3-1:0] node1471;
	wire [3-1:0] node1472;
	wire [3-1:0] node1473;
	wire [3-1:0] node1474;
	wire [3-1:0] node1478;
	wire [3-1:0] node1480;
	wire [3-1:0] node1483;
	wire [3-1:0] node1484;
	wire [3-1:0] node1486;
	wire [3-1:0] node1488;
	wire [3-1:0] node1491;
	wire [3-1:0] node1492;
	wire [3-1:0] node1496;
	wire [3-1:0] node1497;
	wire [3-1:0] node1498;
	wire [3-1:0] node1499;
	wire [3-1:0] node1500;
	wire [3-1:0] node1501;
	wire [3-1:0] node1503;
	wire [3-1:0] node1505;
	wire [3-1:0] node1508;
	wire [3-1:0] node1509;
	wire [3-1:0] node1510;
	wire [3-1:0] node1514;
	wire [3-1:0] node1517;
	wire [3-1:0] node1518;
	wire [3-1:0] node1519;
	wire [3-1:0] node1521;
	wire [3-1:0] node1524;
	wire [3-1:0] node1527;
	wire [3-1:0] node1528;
	wire [3-1:0] node1531;
	wire [3-1:0] node1533;
	wire [3-1:0] node1536;
	wire [3-1:0] node1537;
	wire [3-1:0] node1538;
	wire [3-1:0] node1539;
	wire [3-1:0] node1541;
	wire [3-1:0] node1544;
	wire [3-1:0] node1545;
	wire [3-1:0] node1549;
	wire [3-1:0] node1550;
	wire [3-1:0] node1552;
	wire [3-1:0] node1555;
	wire [3-1:0] node1557;
	wire [3-1:0] node1560;
	wire [3-1:0] node1561;
	wire [3-1:0] node1562;
	wire [3-1:0] node1564;
	wire [3-1:0] node1567;
	wire [3-1:0] node1570;
	wire [3-1:0] node1571;
	wire [3-1:0] node1573;
	wire [3-1:0] node1576;
	wire [3-1:0] node1579;
	wire [3-1:0] node1580;
	wire [3-1:0] node1582;
	wire [3-1:0] node1584;
	wire [3-1:0] node1586;
	wire [3-1:0] node1588;
	wire [3-1:0] node1591;
	wire [3-1:0] node1592;
	wire [3-1:0] node1593;
	wire [3-1:0] node1594;
	wire [3-1:0] node1595;
	wire [3-1:0] node1598;
	wire [3-1:0] node1601;
	wire [3-1:0] node1602;
	wire [3-1:0] node1606;
	wire [3-1:0] node1607;
	wire [3-1:0] node1608;
	wire [3-1:0] node1612;
	wire [3-1:0] node1613;
	wire [3-1:0] node1616;
	wire [3-1:0] node1619;
	wire [3-1:0] node1620;
	wire [3-1:0] node1622;
	wire [3-1:0] node1624;
	wire [3-1:0] node1627;
	wire [3-1:0] node1629;
	wire [3-1:0] node1631;
	wire [3-1:0] node1634;
	wire [3-1:0] node1635;
	wire [3-1:0] node1636;
	wire [3-1:0] node1637;
	wire [3-1:0] node1638;
	wire [3-1:0] node1639;
	wire [3-1:0] node1641;
	wire [3-1:0] node1645;
	wire [3-1:0] node1646;
	wire [3-1:0] node1648;
	wire [3-1:0] node1651;
	wire [3-1:0] node1653;
	wire [3-1:0] node1656;
	wire [3-1:0] node1657;
	wire [3-1:0] node1658;
	wire [3-1:0] node1662;
	wire [3-1:0] node1663;
	wire [3-1:0] node1665;
	wire [3-1:0] node1669;
	wire [3-1:0] node1670;
	wire [3-1:0] node1671;
	wire [3-1:0] node1672;
	wire [3-1:0] node1675;
	wire [3-1:0] node1676;
	wire [3-1:0] node1680;
	wire [3-1:0] node1681;
	wire [3-1:0] node1683;
	wire [3-1:0] node1686;
	wire [3-1:0] node1688;
	wire [3-1:0] node1691;
	wire [3-1:0] node1692;
	wire [3-1:0] node1693;
	wire [3-1:0] node1697;
	wire [3-1:0] node1698;
	wire [3-1:0] node1699;
	wire [3-1:0] node1703;
	wire [3-1:0] node1706;
	wire [3-1:0] node1707;
	wire [3-1:0] node1708;
	wire [3-1:0] node1709;
	wire [3-1:0] node1711;
	wire [3-1:0] node1713;
	wire [3-1:0] node1716;
	wire [3-1:0] node1717;
	wire [3-1:0] node1718;
	wire [3-1:0] node1722;
	wire [3-1:0] node1725;
	wire [3-1:0] node1726;
	wire [3-1:0] node1727;
	wire [3-1:0] node1730;
	wire [3-1:0] node1731;
	wire [3-1:0] node1735;
	wire [3-1:0] node1736;
	wire [3-1:0] node1737;
	wire [3-1:0] node1741;
	wire [3-1:0] node1743;
	wire [3-1:0] node1746;
	wire [3-1:0] node1747;
	wire [3-1:0] node1748;
	wire [3-1:0] node1749;
	wire [3-1:0] node1753;
	wire [3-1:0] node1756;
	wire [3-1:0] node1757;
	wire [3-1:0] node1758;
	wire [3-1:0] node1760;
	wire [3-1:0] node1763;
	wire [3-1:0] node1765;
	wire [3-1:0] node1768;
	wire [3-1:0] node1769;
	wire [3-1:0] node1770;
	wire [3-1:0] node1774;
	wire [3-1:0] node1777;
	wire [3-1:0] node1778;
	wire [3-1:0] node1779;
	wire [3-1:0] node1780;
	wire [3-1:0] node1781;
	wire [3-1:0] node1782;
	wire [3-1:0] node1783;
	wire [3-1:0] node1784;
	wire [3-1:0] node1786;
	wire [3-1:0] node1789;
	wire [3-1:0] node1790;
	wire [3-1:0] node1794;
	wire [3-1:0] node1795;
	wire [3-1:0] node1798;
	wire [3-1:0] node1800;
	wire [3-1:0] node1803;
	wire [3-1:0] node1804;
	wire [3-1:0] node1805;
	wire [3-1:0] node1807;
	wire [3-1:0] node1810;
	wire [3-1:0] node1811;
	wire [3-1:0] node1815;
	wire [3-1:0] node1817;
	wire [3-1:0] node1818;
	wire [3-1:0] node1822;
	wire [3-1:0] node1823;
	wire [3-1:0] node1824;
	wire [3-1:0] node1826;
	wire [3-1:0] node1827;
	wire [3-1:0] node1831;
	wire [3-1:0] node1832;
	wire [3-1:0] node1834;
	wire [3-1:0] node1837;
	wire [3-1:0] node1838;
	wire [3-1:0] node1842;
	wire [3-1:0] node1843;
	wire [3-1:0] node1844;
	wire [3-1:0] node1845;
	wire [3-1:0] node1849;
	wire [3-1:0] node1851;
	wire [3-1:0] node1854;
	wire [3-1:0] node1855;
	wire [3-1:0] node1856;
	wire [3-1:0] node1859;
	wire [3-1:0] node1863;
	wire [3-1:0] node1864;
	wire [3-1:0] node1865;
	wire [3-1:0] node1866;
	wire [3-1:0] node1868;
	wire [3-1:0] node1871;
	wire [3-1:0] node1872;
	wire [3-1:0] node1874;
	wire [3-1:0] node1877;
	wire [3-1:0] node1879;
	wire [3-1:0] node1882;
	wire [3-1:0] node1884;
	wire [3-1:0] node1886;
	wire [3-1:0] node1888;
	wire [3-1:0] node1891;
	wire [3-1:0] node1892;
	wire [3-1:0] node1893;
	wire [3-1:0] node1894;
	wire [3-1:0] node1895;
	wire [3-1:0] node1900;
	wire [3-1:0] node1902;
	wire [3-1:0] node1903;
	wire [3-1:0] node1907;
	wire [3-1:0] node1908;
	wire [3-1:0] node1909;
	wire [3-1:0] node1911;
	wire [3-1:0] node1915;
	wire [3-1:0] node1916;
	wire [3-1:0] node1919;
	wire [3-1:0] node1922;
	wire [3-1:0] node1923;
	wire [3-1:0] node1924;
	wire [3-1:0] node1925;
	wire [3-1:0] node1926;
	wire [3-1:0] node1928;
	wire [3-1:0] node1929;
	wire [3-1:0] node1934;
	wire [3-1:0] node1935;
	wire [3-1:0] node1936;
	wire [3-1:0] node1937;
	wire [3-1:0] node1942;
	wire [3-1:0] node1943;
	wire [3-1:0] node1946;
	wire [3-1:0] node1949;
	wire [3-1:0] node1950;
	wire [3-1:0] node1951;
	wire [3-1:0] node1953;
	wire [3-1:0] node1955;
	wire [3-1:0] node1958;
	wire [3-1:0] node1959;
	wire [3-1:0] node1960;
	wire [3-1:0] node1964;
	wire [3-1:0] node1965;
	wire [3-1:0] node1969;
	wire [3-1:0] node1970;
	wire [3-1:0] node1972;
	wire [3-1:0] node1974;
	wire [3-1:0] node1977;
	wire [3-1:0] node1978;
	wire [3-1:0] node1979;
	wire [3-1:0] node1983;
	wire [3-1:0] node1984;
	wire [3-1:0] node1988;
	wire [3-1:0] node1989;
	wire [3-1:0] node1990;
	wire [3-1:0] node1991;
	wire [3-1:0] node1992;
	wire [3-1:0] node1993;
	wire [3-1:0] node1996;
	wire [3-1:0] node1999;
	wire [3-1:0] node2000;
	wire [3-1:0] node2003;
	wire [3-1:0] node2006;
	wire [3-1:0] node2007;
	wire [3-1:0] node2010;
	wire [3-1:0] node2013;
	wire [3-1:0] node2014;
	wire [3-1:0] node2016;
	wire [3-1:0] node2019;
	wire [3-1:0] node2021;
	wire [3-1:0] node2022;
	wire [3-1:0] node2026;
	wire [3-1:0] node2027;
	wire [3-1:0] node2028;
	wire [3-1:0] node2030;
	wire [3-1:0] node2031;
	wire [3-1:0] node2035;
	wire [3-1:0] node2036;
	wire [3-1:0] node2038;
	wire [3-1:0] node2042;
	wire [3-1:0] node2043;
	wire [3-1:0] node2045;
	wire [3-1:0] node2048;
	wire [3-1:0] node2049;
	wire [3-1:0] node2051;
	wire [3-1:0] node2054;
	wire [3-1:0] node2057;
	wire [3-1:0] node2058;
	wire [3-1:0] node2059;
	wire [3-1:0] node2060;
	wire [3-1:0] node2061;
	wire [3-1:0] node2062;
	wire [3-1:0] node2064;
	wire [3-1:0] node2065;
	wire [3-1:0] node2069;
	wire [3-1:0] node2071;
	wire [3-1:0] node2074;
	wire [3-1:0] node2075;
	wire [3-1:0] node2076;
	wire [3-1:0] node2079;
	wire [3-1:0] node2080;
	wire [3-1:0] node2084;
	wire [3-1:0] node2085;
	wire [3-1:0] node2086;
	wire [3-1:0] node2090;
	wire [3-1:0] node2091;
	wire [3-1:0] node2094;
	wire [3-1:0] node2097;
	wire [3-1:0] node2098;
	wire [3-1:0] node2099;
	wire [3-1:0] node2100;
	wire [3-1:0] node2101;
	wire [3-1:0] node2105;
	wire [3-1:0] node2106;
	wire [3-1:0] node2109;
	wire [3-1:0] node2112;
	wire [3-1:0] node2114;
	wire [3-1:0] node2116;
	wire [3-1:0] node2119;
	wire [3-1:0] node2120;
	wire [3-1:0] node2122;
	wire [3-1:0] node2124;
	wire [3-1:0] node2127;
	wire [3-1:0] node2130;
	wire [3-1:0] node2131;
	wire [3-1:0] node2132;
	wire [3-1:0] node2133;
	wire [3-1:0] node2135;
	wire [3-1:0] node2137;
	wire [3-1:0] node2140;
	wire [3-1:0] node2141;
	wire [3-1:0] node2144;
	wire [3-1:0] node2145;
	wire [3-1:0] node2149;
	wire [3-1:0] node2150;
	wire [3-1:0] node2151;
	wire [3-1:0] node2152;
	wire [3-1:0] node2156;
	wire [3-1:0] node2157;
	wire [3-1:0] node2160;
	wire [3-1:0] node2163;
	wire [3-1:0] node2164;
	wire [3-1:0] node2166;
	wire [3-1:0] node2169;
	wire [3-1:0] node2172;
	wire [3-1:0] node2173;
	wire [3-1:0] node2174;
	wire [3-1:0] node2175;
	wire [3-1:0] node2177;
	wire [3-1:0] node2180;
	wire [3-1:0] node2182;
	wire [3-1:0] node2185;
	wire [3-1:0] node2186;
	wire [3-1:0] node2187;
	wire [3-1:0] node2192;
	wire [3-1:0] node2193;
	wire [3-1:0] node2195;
	wire [3-1:0] node2196;
	wire [3-1:0] node2200;
	wire [3-1:0] node2201;
	wire [3-1:0] node2205;
	wire [3-1:0] node2206;
	wire [3-1:0] node2207;
	wire [3-1:0] node2208;
	wire [3-1:0] node2209;
	wire [3-1:0] node2210;
	wire [3-1:0] node2211;
	wire [3-1:0] node2214;
	wire [3-1:0] node2218;
	wire [3-1:0] node2219;
	wire [3-1:0] node2221;
	wire [3-1:0] node2224;
	wire [3-1:0] node2226;
	wire [3-1:0] node2229;
	wire [3-1:0] node2230;
	wire [3-1:0] node2231;
	wire [3-1:0] node2233;
	wire [3-1:0] node2236;
	wire [3-1:0] node2237;
	wire [3-1:0] node2240;
	wire [3-1:0] node2243;
	wire [3-1:0] node2245;
	wire [3-1:0] node2248;
	wire [3-1:0] node2249;
	wire [3-1:0] node2250;
	wire [3-1:0] node2251;
	wire [3-1:0] node2252;
	wire [3-1:0] node2256;
	wire [3-1:0] node2257;
	wire [3-1:0] node2261;
	wire [3-1:0] node2262;
	wire [3-1:0] node2264;
	wire [3-1:0] node2267;
	wire [3-1:0] node2269;
	wire [3-1:0] node2272;
	wire [3-1:0] node2273;
	wire [3-1:0] node2274;
	wire [3-1:0] node2276;
	wire [3-1:0] node2279;
	wire [3-1:0] node2282;
	wire [3-1:0] node2283;
	wire [3-1:0] node2284;
	wire [3-1:0] node2288;
	wire [3-1:0] node2289;
	wire [3-1:0] node2293;
	wire [3-1:0] node2294;
	wire [3-1:0] node2295;
	wire [3-1:0] node2296;
	wire [3-1:0] node2297;
	wire [3-1:0] node2299;
	wire [3-1:0] node2302;
	wire [3-1:0] node2304;
	wire [3-1:0] node2307;
	wire [3-1:0] node2308;
	wire [3-1:0] node2309;
	wire [3-1:0] node2314;
	wire [3-1:0] node2315;
	wire [3-1:0] node2316;
	wire [3-1:0] node2319;
	wire [3-1:0] node2321;
	wire [3-1:0] node2324;
	wire [3-1:0] node2325;
	wire [3-1:0] node2328;
	wire [3-1:0] node2330;
	wire [3-1:0] node2333;
	wire [3-1:0] node2334;
	wire [3-1:0] node2335;
	wire [3-1:0] node2337;
	wire [3-1:0] node2340;
	wire [3-1:0] node2341;
	wire [3-1:0] node2342;
	wire [3-1:0] node2345;
	wire [3-1:0] node2348;
	wire [3-1:0] node2349;
	wire [3-1:0] node2353;
	wire [3-1:0] node2354;
	wire [3-1:0] node2355;
	wire [3-1:0] node2357;
	wire [3-1:0] node2360;
	wire [3-1:0] node2363;
	wire [3-1:0] node2364;
	wire [3-1:0] node2366;
	wire [3-1:0] node2369;
	wire [3-1:0] node2372;
	wire [3-1:0] node2373;
	wire [3-1:0] node2374;
	wire [3-1:0] node2375;
	wire [3-1:0] node2376;
	wire [3-1:0] node2377;
	wire [3-1:0] node2378;
	wire [3-1:0] node2379;
	wire [3-1:0] node2380;
	wire [3-1:0] node2383;
	wire [3-1:0] node2384;
	wire [3-1:0] node2388;
	wire [3-1:0] node2390;
	wire [3-1:0] node2393;
	wire [3-1:0] node2394;
	wire [3-1:0] node2395;
	wire [3-1:0] node2397;
	wire [3-1:0] node2400;
	wire [3-1:0] node2403;
	wire [3-1:0] node2404;
	wire [3-1:0] node2405;
	wire [3-1:0] node2408;
	wire [3-1:0] node2412;
	wire [3-1:0] node2413;
	wire [3-1:0] node2414;
	wire [3-1:0] node2417;
	wire [3-1:0] node2420;
	wire [3-1:0] node2421;
	wire [3-1:0] node2422;
	wire [3-1:0] node2424;
	wire [3-1:0] node2427;
	wire [3-1:0] node2430;
	wire [3-1:0] node2431;
	wire [3-1:0] node2433;
	wire [3-1:0] node2436;
	wire [3-1:0] node2439;
	wire [3-1:0] node2440;
	wire [3-1:0] node2441;
	wire [3-1:0] node2442;
	wire [3-1:0] node2443;
	wire [3-1:0] node2446;
	wire [3-1:0] node2449;
	wire [3-1:0] node2450;
	wire [3-1:0] node2454;
	wire [3-1:0] node2455;
	wire [3-1:0] node2457;
	wire [3-1:0] node2459;
	wire [3-1:0] node2462;
	wire [3-1:0] node2463;
	wire [3-1:0] node2464;
	wire [3-1:0] node2468;
	wire [3-1:0] node2471;
	wire [3-1:0] node2472;
	wire [3-1:0] node2473;
	wire [3-1:0] node2474;
	wire [3-1:0] node2477;
	wire [3-1:0] node2479;
	wire [3-1:0] node2482;
	wire [3-1:0] node2483;
	wire [3-1:0] node2486;
	wire [3-1:0] node2489;
	wire [3-1:0] node2490;
	wire [3-1:0] node2492;
	wire [3-1:0] node2493;
	wire [3-1:0] node2496;
	wire [3-1:0] node2499;
	wire [3-1:0] node2500;
	wire [3-1:0] node2503;
	wire [3-1:0] node2506;
	wire [3-1:0] node2507;
	wire [3-1:0] node2508;
	wire [3-1:0] node2509;
	wire [3-1:0] node2510;
	wire [3-1:0] node2511;
	wire [3-1:0] node2513;
	wire [3-1:0] node2516;
	wire [3-1:0] node2517;
	wire [3-1:0] node2521;
	wire [3-1:0] node2523;
	wire [3-1:0] node2525;
	wire [3-1:0] node2528;
	wire [3-1:0] node2529;
	wire [3-1:0] node2530;
	wire [3-1:0] node2531;
	wire [3-1:0] node2534;
	wire [3-1:0] node2537;
	wire [3-1:0] node2539;
	wire [3-1:0] node2542;
	wire [3-1:0] node2543;
	wire [3-1:0] node2545;
	wire [3-1:0] node2548;
	wire [3-1:0] node2551;
	wire [3-1:0] node2552;
	wire [3-1:0] node2553;
	wire [3-1:0] node2555;
	wire [3-1:0] node2557;
	wire [3-1:0] node2560;
	wire [3-1:0] node2563;
	wire [3-1:0] node2564;
	wire [3-1:0] node2565;
	wire [3-1:0] node2566;
	wire [3-1:0] node2570;
	wire [3-1:0] node2573;
	wire [3-1:0] node2574;
	wire [3-1:0] node2576;
	wire [3-1:0] node2579;
	wire [3-1:0] node2581;
	wire [3-1:0] node2584;
	wire [3-1:0] node2585;
	wire [3-1:0] node2586;
	wire [3-1:0] node2587;
	wire [3-1:0] node2588;
	wire [3-1:0] node2589;
	wire [3-1:0] node2594;
	wire [3-1:0] node2597;
	wire [3-1:0] node2598;
	wire [3-1:0] node2599;
	wire [3-1:0] node2600;
	wire [3-1:0] node2603;
	wire [3-1:0] node2606;
	wire [3-1:0] node2608;
	wire [3-1:0] node2611;
	wire [3-1:0] node2612;
	wire [3-1:0] node2616;
	wire [3-1:0] node2617;
	wire [3-1:0] node2618;
	wire [3-1:0] node2619;
	wire [3-1:0] node2622;
	wire [3-1:0] node2623;
	wire [3-1:0] node2627;
	wire [3-1:0] node2628;
	wire [3-1:0] node2630;
	wire [3-1:0] node2633;
	wire [3-1:0] node2636;
	wire [3-1:0] node2637;
	wire [3-1:0] node2639;
	wire [3-1:0] node2643;
	wire [3-1:0] node2644;
	wire [3-1:0] node2645;
	wire [3-1:0] node2646;
	wire [3-1:0] node2647;
	wire [3-1:0] node2649;
	wire [3-1:0] node2651;
	wire [3-1:0] node2654;
	wire [3-1:0] node2655;
	wire [3-1:0] node2656;
	wire [3-1:0] node2660;
	wire [3-1:0] node2661;
	wire [3-1:0] node2664;
	wire [3-1:0] node2667;
	wire [3-1:0] node2668;
	wire [3-1:0] node2669;
	wire [3-1:0] node2670;
	wire [3-1:0] node2671;
	wire [3-1:0] node2676;
	wire [3-1:0] node2677;
	wire [3-1:0] node2679;
	wire [3-1:0] node2683;
	wire [3-1:0] node2684;
	wire [3-1:0] node2685;
	wire [3-1:0] node2689;
	wire [3-1:0] node2690;
	wire [3-1:0] node2694;
	wire [3-1:0] node2695;
	wire [3-1:0] node2696;
	wire [3-1:0] node2697;
	wire [3-1:0] node2698;
	wire [3-1:0] node2702;
	wire [3-1:0] node2703;
	wire [3-1:0] node2706;
	wire [3-1:0] node2707;
	wire [3-1:0] node2711;
	wire [3-1:0] node2712;
	wire [3-1:0] node2713;
	wire [3-1:0] node2716;
	wire [3-1:0] node2720;
	wire [3-1:0] node2721;
	wire [3-1:0] node2722;
	wire [3-1:0] node2724;
	wire [3-1:0] node2725;
	wire [3-1:0] node2729;
	wire [3-1:0] node2730;
	wire [3-1:0] node2731;
	wire [3-1:0] node2735;
	wire [3-1:0] node2736;
	wire [3-1:0] node2740;
	wire [3-1:0] node2741;
	wire [3-1:0] node2742;
	wire [3-1:0] node2744;
	wire [3-1:0] node2747;
	wire [3-1:0] node2748;
	wire [3-1:0] node2752;
	wire [3-1:0] node2753;
	wire [3-1:0] node2756;
	wire [3-1:0] node2757;
	wire [3-1:0] node2761;
	wire [3-1:0] node2762;
	wire [3-1:0] node2763;
	wire [3-1:0] node2764;
	wire [3-1:0] node2765;
	wire [3-1:0] node2766;
	wire [3-1:0] node2769;
	wire [3-1:0] node2772;
	wire [3-1:0] node2773;
	wire [3-1:0] node2776;
	wire [3-1:0] node2779;
	wire [3-1:0] node2781;
	wire [3-1:0] node2782;
	wire [3-1:0] node2783;
	wire [3-1:0] node2787;
	wire [3-1:0] node2788;
	wire [3-1:0] node2792;
	wire [3-1:0] node2793;
	wire [3-1:0] node2794;
	wire [3-1:0] node2795;
	wire [3-1:0] node2797;
	wire [3-1:0] node2800;
	wire [3-1:0] node2801;
	wire [3-1:0] node2805;
	wire [3-1:0] node2806;
	wire [3-1:0] node2808;
	wire [3-1:0] node2811;
	wire [3-1:0] node2813;
	wire [3-1:0] node2816;
	wire [3-1:0] node2817;
	wire [3-1:0] node2819;
	wire [3-1:0] node2822;
	wire [3-1:0] node2823;
	wire [3-1:0] node2824;
	wire [3-1:0] node2829;
	wire [3-1:0] node2830;
	wire [3-1:0] node2831;
	wire [3-1:0] node2832;
	wire [3-1:0] node2833;
	wire [3-1:0] node2834;
	wire [3-1:0] node2838;
	wire [3-1:0] node2840;
	wire [3-1:0] node2843;
	wire [3-1:0] node2844;
	wire [3-1:0] node2847;
	wire [3-1:0] node2848;
	wire [3-1:0] node2852;
	wire [3-1:0] node2853;
	wire [3-1:0] node2854;
	wire [3-1:0] node2858;
	wire [3-1:0] node2859;
	wire [3-1:0] node2860;
	wire [3-1:0] node2864;
	wire [3-1:0] node2866;
	wire [3-1:0] node2869;
	wire [3-1:0] node2870;
	wire [3-1:0] node2871;
	wire [3-1:0] node2873;
	wire [3-1:0] node2875;
	wire [3-1:0] node2878;
	wire [3-1:0] node2879;
	wire [3-1:0] node2882;
	wire [3-1:0] node2883;
	wire [3-1:0] node2887;
	wire [3-1:0] node2888;
	wire [3-1:0] node2889;
	wire [3-1:0] node2890;
	wire [3-1:0] node2893;
	wire [3-1:0] node2896;
	wire [3-1:0] node2897;
	wire [3-1:0] node2900;
	wire [3-1:0] node2903;
	wire [3-1:0] node2904;
	wire [3-1:0] node2907;
	wire [3-1:0] node2910;
	wire [3-1:0] node2911;
	wire [3-1:0] node2912;
	wire [3-1:0] node2913;
	wire [3-1:0] node2914;
	wire [3-1:0] node2915;
	wire [3-1:0] node2916;
	wire [3-1:0] node2917;
	wire [3-1:0] node2919;
	wire [3-1:0] node2922;
	wire [3-1:0] node2925;
	wire [3-1:0] node2926;
	wire [3-1:0] node2928;
	wire [3-1:0] node2931;
	wire [3-1:0] node2934;
	wire [3-1:0] node2935;
	wire [3-1:0] node2936;
	wire [3-1:0] node2938;
	wire [3-1:0] node2941;
	wire [3-1:0] node2944;
	wire [3-1:0] node2945;
	wire [3-1:0] node2949;
	wire [3-1:0] node2950;
	wire [3-1:0] node2951;
	wire [3-1:0] node2952;
	wire [3-1:0] node2953;
	wire [3-1:0] node2957;
	wire [3-1:0] node2960;
	wire [3-1:0] node2961;
	wire [3-1:0] node2962;
	wire [3-1:0] node2966;
	wire [3-1:0] node2969;
	wire [3-1:0] node2970;
	wire [3-1:0] node2971;
	wire [3-1:0] node2972;
	wire [3-1:0] node2976;
	wire [3-1:0] node2979;
	wire [3-1:0] node2980;
	wire [3-1:0] node2983;
	wire [3-1:0] node2984;
	wire [3-1:0] node2988;
	wire [3-1:0] node2989;
	wire [3-1:0] node2990;
	wire [3-1:0] node2991;
	wire [3-1:0] node2993;
	wire [3-1:0] node2994;
	wire [3-1:0] node2997;
	wire [3-1:0] node3001;
	wire [3-1:0] node3002;
	wire [3-1:0] node3003;
	wire [3-1:0] node3004;
	wire [3-1:0] node3009;
	wire [3-1:0] node3010;
	wire [3-1:0] node3013;
	wire [3-1:0] node3015;
	wire [3-1:0] node3018;
	wire [3-1:0] node3019;
	wire [3-1:0] node3020;
	wire [3-1:0] node3022;
	wire [3-1:0] node3024;
	wire [3-1:0] node3027;
	wire [3-1:0] node3028;
	wire [3-1:0] node3029;
	wire [3-1:0] node3032;
	wire [3-1:0] node3035;
	wire [3-1:0] node3036;
	wire [3-1:0] node3040;
	wire [3-1:0] node3041;
	wire [3-1:0] node3043;
	wire [3-1:0] node3045;
	wire [3-1:0] node3048;
	wire [3-1:0] node3049;
	wire [3-1:0] node3050;
	wire [3-1:0] node3054;
	wire [3-1:0] node3055;
	wire [3-1:0] node3059;
	wire [3-1:0] node3060;
	wire [3-1:0] node3061;
	wire [3-1:0] node3062;
	wire [3-1:0] node3063;
	wire [3-1:0] node3064;
	wire [3-1:0] node3066;
	wire [3-1:0] node3069;
	wire [3-1:0] node3070;
	wire [3-1:0] node3073;
	wire [3-1:0] node3076;
	wire [3-1:0] node3078;
	wire [3-1:0] node3081;
	wire [3-1:0] node3082;
	wire [3-1:0] node3084;
	wire [3-1:0] node3086;
	wire [3-1:0] node3089;
	wire [3-1:0] node3090;
	wire [3-1:0] node3091;
	wire [3-1:0] node3096;
	wire [3-1:0] node3097;
	wire [3-1:0] node3098;
	wire [3-1:0] node3099;
	wire [3-1:0] node3103;
	wire [3-1:0] node3104;
	wire [3-1:0] node3107;
	wire [3-1:0] node3110;
	wire [3-1:0] node3111;
	wire [3-1:0] node3113;
	wire [3-1:0] node3117;
	wire [3-1:0] node3118;
	wire [3-1:0] node3119;
	wire [3-1:0] node3120;
	wire [3-1:0] node3121;
	wire [3-1:0] node3126;
	wire [3-1:0] node3127;
	wire [3-1:0] node3128;
	wire [3-1:0] node3131;
	wire [3-1:0] node3134;
	wire [3-1:0] node3135;
	wire [3-1:0] node3136;
	wire [3-1:0] node3139;
	wire [3-1:0] node3142;
	wire [3-1:0] node3143;
	wire [3-1:0] node3147;
	wire [3-1:0] node3148;
	wire [3-1:0] node3149;
	wire [3-1:0] node3151;
	wire [3-1:0] node3152;
	wire [3-1:0] node3155;
	wire [3-1:0] node3158;
	wire [3-1:0] node3160;
	wire [3-1:0] node3163;
	wire [3-1:0] node3164;
	wire [3-1:0] node3166;
	wire [3-1:0] node3168;
	wire [3-1:0] node3171;
	wire [3-1:0] node3172;
	wire [3-1:0] node3173;
	wire [3-1:0] node3177;
	wire [3-1:0] node3180;
	wire [3-1:0] node3181;
	wire [3-1:0] node3182;
	wire [3-1:0] node3183;
	wire [3-1:0] node3184;
	wire [3-1:0] node3185;
	wire [3-1:0] node3186;
	wire [3-1:0] node3187;
	wire [3-1:0] node3191;
	wire [3-1:0] node3192;
	wire [3-1:0] node3196;
	wire [3-1:0] node3197;
	wire [3-1:0] node3200;
	wire [3-1:0] node3203;
	wire [3-1:0] node3204;
	wire [3-1:0] node3205;
	wire [3-1:0] node3209;
	wire [3-1:0] node3210;
	wire [3-1:0] node3211;
	wire [3-1:0] node3215;
	wire [3-1:0] node3218;
	wire [3-1:0] node3219;
	wire [3-1:0] node3220;
	wire [3-1:0] node3221;
	wire [3-1:0] node3225;
	wire [3-1:0] node3227;
	wire [3-1:0] node3229;
	wire [3-1:0] node3234;
	wire [3-1:0] node3235;
	wire [3-1:0] node3236;
	wire [3-1:0] node3237;
	wire [3-1:0] node3238;
	wire [3-1:0] node3239;
	wire [3-1:0] node3240;
	wire [3-1:0] node3244;
	wire [3-1:0] node3245;
	wire [3-1:0] node3248;
	wire [3-1:0] node3251;
	wire [3-1:0] node3253;
	wire [3-1:0] node3256;
	wire [3-1:0] node3257;
	wire [3-1:0] node3258;
	wire [3-1:0] node3262;
	wire [3-1:0] node3265;
	wire [3-1:0] node3266;
	wire [3-1:0] node3267;
	wire [3-1:0] node3268;
	wire [3-1:0] node3270;
	wire [3-1:0] node3274;
	wire [3-1:0] node3275;
	wire [3-1:0] node3277;
	wire [3-1:0] node3281;
	wire [3-1:0] node3282;
	wire [3-1:0] node3283;
	wire [3-1:0] node3286;
	wire [3-1:0] node3289;
	wire [3-1:0] node3290;
	wire [3-1:0] node3291;
	wire [3-1:0] node3294;
	wire [3-1:0] node3297;
	wire [3-1:0] node3298;
	wire [3-1:0] node3302;
	wire [3-1:0] node3303;
	wire [3-1:0] node3304;
	wire [3-1:0] node3305;
	wire [3-1:0] node3306;
	wire [3-1:0] node3309;
	wire [3-1:0] node3310;
	wire [3-1:0] node3314;
	wire [3-1:0] node3315;
	wire [3-1:0] node3316;
	wire [3-1:0] node3319;
	wire [3-1:0] node3323;
	wire [3-1:0] node3324;
	wire [3-1:0] node3325;
	wire [3-1:0] node3327;
	wire [3-1:0] node3330;
	wire [3-1:0] node3332;
	wire [3-1:0] node3335;
	wire [3-1:0] node3336;
	wire [3-1:0] node3340;
	wire [3-1:0] node3341;
	wire [3-1:0] node3342;
	wire [3-1:0] node3344;
	wire [3-1:0] node3347;
	wire [3-1:0] node3349;
	wire [3-1:0] node3351;

	assign outp = (inp[6]) ? node1360 : node1;
		assign node1 = (inp[3]) ? node1001 : node2;
			assign node2 = (inp[9]) ? node566 : node3;
				assign node3 = (inp[0]) ? node277 : node4;
					assign node4 = (inp[4]) ? node142 : node5;
						assign node5 = (inp[1]) ? node63 : node6;
							assign node6 = (inp[7]) ? node50 : node7;
								assign node7 = (inp[10]) ? node31 : node8;
									assign node8 = (inp[5]) ? node18 : node9;
										assign node9 = (inp[11]) ? node15 : node10;
											assign node10 = (inp[8]) ? node12 : 3'b011;
												assign node12 = (inp[2]) ? 3'b011 : 3'b111;
											assign node15 = (inp[8]) ? 3'b011 : 3'b101;
										assign node18 = (inp[2]) ? node24 : node19;
											assign node19 = (inp[11]) ? 3'b001 : node20;
												assign node20 = (inp[8]) ? 3'b011 : 3'b111;
											assign node24 = (inp[11]) ? node28 : node25;
												assign node25 = (inp[8]) ? 3'b001 : 3'b101;
												assign node28 = (inp[8]) ? 3'b101 : 3'b001;
									assign node31 = (inp[5]) ? node41 : node32;
										assign node32 = (inp[2]) ? node36 : node33;
											assign node33 = (inp[8]) ? 3'b001 : 3'b101;
											assign node36 = (inp[11]) ? node38 : 3'b101;
												assign node38 = (inp[8]) ? 3'b101 : 3'b001;
										assign node41 = (inp[11]) ? node45 : node42;
											assign node42 = (inp[8]) ? 3'b101 : 3'b001;
											assign node45 = (inp[2]) ? node47 : 3'b001;
												assign node47 = (inp[8]) ? 3'b000 : 3'b110;
								assign node50 = (inp[10]) ? node58 : node51;
									assign node51 = (inp[8]) ? node53 : 3'b001;
										assign node53 = (inp[5]) ? 3'b001 : node54;
											assign node54 = (inp[2]) ? 3'b001 : 3'b000;
									assign node58 = (inp[8]) ? 3'b001 : node59;
										assign node59 = (inp[5]) ? 3'b000 : 3'b001;
							assign node63 = (inp[7]) ? node99 : node64;
								assign node64 = (inp[10]) ? node80 : node65;
									assign node65 = (inp[11]) ? node73 : node66;
										assign node66 = (inp[8]) ? node68 : 3'b001;
											assign node68 = (inp[2]) ? node70 : 3'b011;
												assign node70 = (inp[5]) ? 3'b001 : 3'b101;
										assign node73 = (inp[8]) ? node77 : node74;
											assign node74 = (inp[5]) ? 3'b110 : 3'b001;
											assign node77 = (inp[5]) ? 3'b001 : 3'b101;
									assign node80 = (inp[8]) ? node88 : node81;
										assign node81 = (inp[2]) ? node83 : 3'b110;
											assign node83 = (inp[11]) ? node85 : 3'b110;
												assign node85 = (inp[5]) ? 3'b010 : 3'b110;
										assign node88 = (inp[5]) ? node94 : node89;
											assign node89 = (inp[11]) ? 3'b001 : node90;
												assign node90 = (inp[2]) ? 3'b001 : 3'b101;
											assign node94 = (inp[2]) ? 3'b110 : node95;
												assign node95 = (inp[11]) ? 3'b110 : 3'b001;
								assign node99 = (inp[8]) ? node121 : node100;
									assign node100 = (inp[11]) ? node112 : node101;
										assign node101 = (inp[5]) ? node107 : node102;
											assign node102 = (inp[10]) ? 3'b101 : node103;
												assign node103 = (inp[2]) ? 3'b011 : 3'b111;
											assign node107 = (inp[10]) ? node109 : 3'b101;
												assign node109 = (inp[2]) ? 3'b001 : 3'b101;
										assign node112 = (inp[10]) ? node116 : node113;
											assign node113 = (inp[5]) ? 3'b101 : 3'b001;
											assign node116 = (inp[5]) ? 3'b001 : node117;
												assign node117 = (inp[2]) ? 3'b001 : 3'b101;
									assign node121 = (inp[10]) ? node131 : node122;
										assign node122 = (inp[5]) ? node126 : node123;
											assign node123 = (inp[2]) ? 3'b011 : 3'b111;
											assign node126 = (inp[11]) ? node128 : 3'b011;
												assign node128 = (inp[2]) ? 3'b101 : 3'b011;
										assign node131 = (inp[11]) ? node135 : node132;
											assign node132 = (inp[5]) ? 3'b101 : 3'b011;
											assign node135 = (inp[5]) ? node139 : node136;
												assign node136 = (inp[2]) ? 3'b101 : 3'b001;
												assign node139 = (inp[2]) ? 3'b001 : 3'b101;
						assign node142 = (inp[7]) ? node206 : node143;
							assign node143 = (inp[1]) ? node179 : node144;
								assign node144 = (inp[8]) ? node166 : node145;
									assign node145 = (inp[11]) ? node159 : node146;
										assign node146 = (inp[2]) ? node152 : node147;
											assign node147 = (inp[5]) ? 3'b110 : node148;
												assign node148 = (inp[10]) ? 3'b110 : 3'b100;
											assign node152 = (inp[10]) ? node156 : node153;
												assign node153 = (inp[5]) ? 3'b110 : 3'b000;
												assign node156 = (inp[5]) ? 3'b000 : 3'b110;
										assign node159 = (inp[10]) ? node163 : node160;
											assign node160 = (inp[5]) ? 3'b110 : 3'b010;
											assign node163 = (inp[5]) ? 3'b010 : 3'b110;
									assign node166 = (inp[2]) ? node174 : node167;
										assign node167 = (inp[10]) ? node171 : node168;
											assign node168 = (inp[5]) ? 3'b000 : 3'b100;
											assign node171 = (inp[5]) ? 3'b110 : 3'b000;
										assign node174 = (inp[10]) ? 3'b110 : node175;
											assign node175 = (inp[5]) ? 3'b010 : 3'b000;
								assign node179 = (inp[8]) ? node191 : node180;
									assign node180 = (inp[10]) ? node184 : node181;
										assign node181 = (inp[5]) ? 3'b010 : 3'b110;
										assign node184 = (inp[5]) ? node186 : 3'b010;
											assign node186 = (inp[2]) ? 3'b100 : node187;
												assign node187 = (inp[11]) ? 3'b100 : 3'b000;
									assign node191 = (inp[10]) ? node199 : node192;
										assign node192 = (inp[5]) ? 3'b110 : node193;
											assign node193 = (inp[2]) ? node195 : 3'b000;
												assign node195 = (inp[11]) ? 3'b110 : 3'b001;
										assign node199 = (inp[5]) ? 3'b010 : node200;
											assign node200 = (inp[11]) ? node202 : 3'b110;
												assign node202 = (inp[2]) ? 3'b010 : 3'b110;
							assign node206 = (inp[1]) ? node248 : node207;
								assign node207 = (inp[10]) ? node229 : node208;
									assign node208 = (inp[5]) ? node220 : node209;
										assign node209 = (inp[8]) ? node215 : node210;
											assign node210 = (inp[2]) ? node212 : 3'b001;
												assign node212 = (inp[11]) ? 3'b101 : 3'b111;
											assign node215 = (inp[2]) ? 3'b011 : node216;
												assign node216 = (inp[11]) ? 3'b011 : 3'b111;
										assign node220 = (inp[2]) ? node224 : node221;
											assign node221 = (inp[11]) ? 3'b101 : 3'b111;
											assign node224 = (inp[8]) ? 3'b101 : node225;
												assign node225 = (inp[11]) ? 3'b001 : 3'b101;
									assign node229 = (inp[8]) ? node237 : node230;
										assign node230 = (inp[11]) ? node232 : 3'b001;
											assign node232 = (inp[2]) ? node234 : 3'b001;
												assign node234 = (inp[5]) ? 3'b110 : 3'b001;
										assign node237 = (inp[5]) ? node243 : node238;
											assign node238 = (inp[11]) ? 3'b101 : node239;
												assign node239 = (inp[2]) ? 3'b101 : 3'b001;
											assign node243 = (inp[11]) ? 3'b001 : node244;
												assign node244 = (inp[2]) ? 3'b001 : 3'b101;
								assign node248 = (inp[8]) ? node262 : node249;
									assign node249 = (inp[10]) ? node257 : node250;
										assign node250 = (inp[11]) ? node252 : 3'b001;
											assign node252 = (inp[5]) ? 3'b110 : node253;
												assign node253 = (inp[2]) ? 3'b001 : 3'b101;
										assign node257 = (inp[11]) ? node259 : 3'b110;
											assign node259 = (inp[2]) ? 3'b010 : 3'b110;
									assign node262 = (inp[5]) ? node270 : node263;
										assign node263 = (inp[10]) ? node265 : 3'b101;
											assign node265 = (inp[11]) ? 3'b001 : node266;
												assign node266 = (inp[2]) ? 3'b001 : 3'b101;
										assign node270 = (inp[10]) ? node274 : node271;
											assign node271 = (inp[11]) ? 3'b001 : 3'b101;
											assign node274 = (inp[11]) ? 3'b110 : 3'b001;
					assign node277 = (inp[4]) ? node417 : node278;
						assign node278 = (inp[7]) ? node364 : node279;
							assign node279 = (inp[10]) ? node327 : node280;
								assign node280 = (inp[1]) ? node306 : node281;
									assign node281 = (inp[11]) ? node291 : node282;
										assign node282 = (inp[5]) ? node288 : node283;
											assign node283 = (inp[2]) ? 3'b001 : node284;
												assign node284 = (inp[8]) ? 3'b101 : 3'b001;
											assign node288 = (inp[8]) ? 3'b001 : 3'b110;
										assign node291 = (inp[8]) ? node299 : node292;
											assign node292 = (inp[5]) ? node296 : node293;
												assign node293 = (inp[2]) ? 3'b110 : 3'b010;
												assign node296 = (inp[2]) ? 3'b010 : 3'b110;
											assign node299 = (inp[5]) ? node303 : node300;
												assign node300 = (inp[2]) ? 3'b001 : 3'b000;
												assign node303 = (inp[2]) ? 3'b110 : 3'b010;
									assign node306 = (inp[5]) ? node320 : node307;
										assign node307 = (inp[2]) ? node315 : node308;
											assign node308 = (inp[11]) ? node312 : node309;
												assign node309 = (inp[8]) ? 3'b001 : 3'b111;
												assign node312 = (inp[8]) ? 3'b110 : 3'b000;
											assign node315 = (inp[8]) ? 3'b110 : node316;
												assign node316 = (inp[11]) ? 3'b010 : 3'b110;
										assign node320 = (inp[8]) ? node324 : node321;
											assign node321 = (inp[11]) ? 3'b110 : 3'b010;
											assign node324 = (inp[11]) ? 3'b010 : 3'b110;
								assign node327 = (inp[5]) ? node351 : node328;
									assign node328 = (inp[1]) ? node338 : node329;
										assign node329 = (inp[2]) ? node333 : node330;
											assign node330 = (inp[8]) ? 3'b010 : 3'b110;
											assign node333 = (inp[11]) ? node335 : 3'b110;
												assign node335 = (inp[8]) ? 3'b110 : 3'b010;
										assign node338 = (inp[2]) ? node346 : node339;
											assign node339 = (inp[11]) ? node343 : node340;
												assign node340 = (inp[8]) ? 3'b110 : 3'b010;
												assign node343 = (inp[8]) ? 3'b010 : 3'b110;
											assign node346 = (inp[8]) ? 3'b010 : node347;
												assign node347 = (inp[11]) ? 3'b100 : 3'b010;
									assign node351 = (inp[1]) ? node359 : node352;
										assign node352 = (inp[11]) ? node356 : node353;
											assign node353 = (inp[8]) ? 3'b110 : 3'b010;
											assign node356 = (inp[8]) ? 3'b010 : 3'b000;
										assign node359 = (inp[11]) ? 3'b100 : node360;
											assign node360 = (inp[8]) ? 3'b010 : 3'b100;
							assign node364 = (inp[1]) ? node392 : node365;
								assign node365 = (inp[8]) ? node373 : node366;
									assign node366 = (inp[10]) ? node370 : node367;
										assign node367 = (inp[5]) ? 3'b001 : 3'b101;
										assign node370 = (inp[5]) ? 3'b110 : 3'b001;
									assign node373 = (inp[5]) ? node385 : node374;
										assign node374 = (inp[10]) ? node380 : node375;
											assign node375 = (inp[2]) ? node377 : 3'b010;
												assign node377 = (inp[11]) ? 3'b101 : 3'b011;
											assign node380 = (inp[11]) ? node382 : 3'b101;
												assign node382 = (inp[2]) ? 3'b001 : 3'b101;
										assign node385 = (inp[10]) ? 3'b001 : node386;
											assign node386 = (inp[2]) ? node388 : 3'b101;
												assign node388 = (inp[11]) ? 3'b001 : 3'b101;
								assign node392 = (inp[10]) ? node404 : node393;
									assign node393 = (inp[8]) ? node401 : node394;
										assign node394 = (inp[5]) ? 3'b110 : node395;
											assign node395 = (inp[2]) ? 3'b001 : node396;
												assign node396 = (inp[11]) ? 3'b001 : 3'b101;
										assign node401 = (inp[5]) ? 3'b001 : 3'b101;
									assign node404 = (inp[8]) ? node412 : node405;
										assign node405 = (inp[5]) ? node407 : 3'b110;
											assign node407 = (inp[11]) ? 3'b010 : node408;
												assign node408 = (inp[2]) ? 3'b010 : 3'b110;
										assign node412 = (inp[5]) ? 3'b110 : node413;
											assign node413 = (inp[11]) ? 3'b010 : 3'b001;
						assign node417 = (inp[7]) ? node479 : node418;
							assign node418 = (inp[10]) ? node452 : node419;
								assign node419 = (inp[1]) ? node435 : node420;
									assign node420 = (inp[8]) ? node428 : node421;
										assign node421 = (inp[5]) ? 3'b100 : node422;
											assign node422 = (inp[11]) ? 3'b010 : node423;
												assign node423 = (inp[2]) ? 3'b010 : 3'b110;
										assign node428 = (inp[5]) ? 3'b010 : node429;
											assign node429 = (inp[11]) ? node431 : 3'b110;
												assign node431 = (inp[2]) ? 3'b010 : 3'b110;
									assign node435 = (inp[5]) ? node443 : node436;
										assign node436 = (inp[2]) ? node438 : 3'b100;
											assign node438 = (inp[11]) ? 3'b100 : node439;
												assign node439 = (inp[8]) ? 3'b010 : 3'b100;
										assign node443 = (inp[11]) ? node449 : node444;
											assign node444 = (inp[2]) ? 3'b100 : node445;
												assign node445 = (inp[8]) ? 3'b000 : 3'b100;
											assign node449 = (inp[8]) ? 3'b100 : 3'b000;
								assign node452 = (inp[1]) ? node468 : node453;
									assign node453 = (inp[8]) ? node461 : node454;
										assign node454 = (inp[5]) ? node456 : 3'b100;
											assign node456 = (inp[2]) ? 3'b000 : node457;
												assign node457 = (inp[11]) ? 3'b000 : 3'b100;
										assign node461 = (inp[5]) ? 3'b100 : node462;
											assign node462 = (inp[11]) ? node464 : 3'b010;
												assign node464 = (inp[2]) ? 3'b100 : 3'b000;
									assign node468 = (inp[8]) ? node470 : 3'b000;
										assign node470 = (inp[11]) ? 3'b000 : node471;
											assign node471 = (inp[2]) ? node475 : node472;
												assign node472 = (inp[5]) ? 3'b100 : 3'b000;
												assign node475 = (inp[5]) ? 3'b000 : 3'b100;
							assign node479 = (inp[10]) ? node527 : node480;
								assign node480 = (inp[11]) ? node498 : node481;
									assign node481 = (inp[5]) ? node491 : node482;
										assign node482 = (inp[1]) ? node488 : node483;
											assign node483 = (inp[2]) ? 3'b001 : node484;
												assign node484 = (inp[8]) ? 3'b101 : 3'b001;
											assign node488 = (inp[8]) ? 3'b001 : 3'b110;
										assign node491 = (inp[8]) ? node495 : node492;
											assign node492 = (inp[1]) ? 3'b010 : 3'b110;
											assign node495 = (inp[1]) ? 3'b110 : 3'b001;
									assign node498 = (inp[5]) ? node512 : node499;
										assign node499 = (inp[8]) ? node507 : node500;
											assign node500 = (inp[2]) ? node504 : node501;
												assign node501 = (inp[1]) ? 3'b100 : 3'b010;
												assign node504 = (inp[1]) ? 3'b010 : 3'b110;
											assign node507 = (inp[1]) ? 3'b110 : node508;
												assign node508 = (inp[2]) ? 3'b001 : 3'b000;
										assign node512 = (inp[8]) ? node520 : node513;
											assign node513 = (inp[2]) ? node517 : node514;
												assign node514 = (inp[1]) ? 3'b010 : 3'b110;
												assign node517 = (inp[1]) ? 3'b100 : 3'b010;
											assign node520 = (inp[1]) ? node524 : node521;
												assign node521 = (inp[2]) ? 3'b110 : 3'b010;
												assign node524 = (inp[2]) ? 3'b010 : 3'b110;
								assign node527 = (inp[5]) ? node547 : node528;
									assign node528 = (inp[1]) ? node538 : node529;
										assign node529 = (inp[8]) ? node535 : node530;
											assign node530 = (inp[2]) ? node532 : 3'b110;
												assign node532 = (inp[11]) ? 3'b010 : 3'b110;
											assign node535 = (inp[2]) ? 3'b110 : 3'b010;
										assign node538 = (inp[8]) ? node544 : node539;
											assign node539 = (inp[11]) ? node541 : 3'b010;
												assign node541 = (inp[2]) ? 3'b100 : 3'b010;
											assign node544 = (inp[2]) ? 3'b010 : 3'b110;
									assign node547 = (inp[11]) ? node555 : node548;
										assign node548 = (inp[1]) ? node552 : node549;
											assign node549 = (inp[8]) ? 3'b110 : 3'b010;
											assign node552 = (inp[8]) ? 3'b010 : 3'b100;
										assign node555 = (inp[1]) ? node561 : node556;
											assign node556 = (inp[8]) ? 3'b010 : node557;
												assign node557 = (inp[2]) ? 3'b100 : 3'b000;
											assign node561 = (inp[8]) ? 3'b100 : node562;
												assign node562 = (inp[2]) ? 3'b000 : 3'b100;
				assign node566 = (inp[7]) ? node724 : node567;
					assign node567 = (inp[0]) ? node663 : node568;
						assign node568 = (inp[10]) ? node616 : node569;
							assign node569 = (inp[1]) ? node585 : node570;
								assign node570 = (inp[4]) ? 3'b010 : node571;
									assign node571 = (inp[11]) ? node577 : node572;
										assign node572 = (inp[5]) ? node574 : 3'b010;
											assign node574 = (inp[8]) ? 3'b010 : 3'b100;
										assign node577 = (inp[2]) ? 3'b100 : node578;
											assign node578 = (inp[5]) ? node580 : 3'b000;
												assign node580 = (inp[8]) ? 3'b000 : 3'b100;
								assign node585 = (inp[4]) ? node605 : node586;
									assign node586 = (inp[5]) ? node600 : node587;
										assign node587 = (inp[8]) ? node595 : node588;
											assign node588 = (inp[11]) ? node592 : node589;
												assign node589 = (inp[2]) ? 3'b010 : 3'b011;
												assign node592 = (inp[2]) ? 3'b010 : 3'b110;
											assign node595 = (inp[11]) ? 3'b110 : node596;
												assign node596 = (inp[2]) ? 3'b110 : 3'b111;
										assign node600 = (inp[8]) ? 3'b010 : node601;
											assign node601 = (inp[11]) ? 3'b100 : 3'b010;
									assign node605 = (inp[5]) ? node613 : node606;
										assign node606 = (inp[8]) ? node608 : 3'b100;
											assign node608 = (inp[2]) ? node610 : 3'b000;
												assign node610 = (inp[11]) ? 3'b000 : 3'b010;
										assign node613 = (inp[8]) ? 3'b100 : 3'b000;
							assign node616 = (inp[4]) ? node656 : node617;
								assign node617 = (inp[1]) ? node641 : node618;
									assign node618 = (inp[2]) ? node628 : node619;
										assign node619 = (inp[5]) ? node625 : node620;
											assign node620 = (inp[8]) ? node622 : 3'b100;
												assign node622 = (inp[11]) ? 3'b100 : 3'b000;
											assign node625 = (inp[8]) ? 3'b100 : 3'b000;
										assign node628 = (inp[11]) ? node636 : node629;
											assign node629 = (inp[5]) ? node633 : node630;
												assign node630 = (inp[8]) ? 3'b000 : 3'b100;
												assign node633 = (inp[8]) ? 3'b100 : 3'b000;
											assign node636 = (inp[5]) ? 3'b000 : node637;
												assign node637 = (inp[8]) ? 3'b100 : 3'b000;
									assign node641 = (inp[5]) ? node647 : node642;
										assign node642 = (inp[8]) ? 3'b010 : node643;
											assign node643 = (inp[11]) ? 3'b100 : 3'b010;
										assign node647 = (inp[2]) ? node651 : node648;
											assign node648 = (inp[11]) ? 3'b100 : 3'b110;
											assign node651 = (inp[11]) ? node653 : 3'b100;
												assign node653 = (inp[8]) ? 3'b100 : 3'b000;
								assign node656 = (inp[5]) ? 3'b000 : node657;
									assign node657 = (inp[1]) ? node659 : 3'b010;
										assign node659 = (inp[8]) ? 3'b100 : 3'b000;
						assign node663 = (inp[4]) ? node713 : node664;
							assign node664 = (inp[1]) ? node698 : node665;
								assign node665 = (inp[10]) ? node683 : node666;
									assign node666 = (inp[5]) ? node672 : node667;
										assign node667 = (inp[11]) ? node669 : 3'b010;
											assign node669 = (inp[2]) ? 3'b010 : 3'b000;
										assign node672 = (inp[2]) ? node678 : node673;
											assign node673 = (inp[8]) ? node675 : 3'b100;
												assign node675 = (inp[11]) ? 3'b000 : 3'b010;
											assign node678 = (inp[8]) ? 3'b100 : node679;
												assign node679 = (inp[11]) ? 3'b000 : 3'b100;
									assign node683 = (inp[5]) ? node693 : node684;
										assign node684 = (inp[2]) ? node686 : 3'b100;
											assign node686 = (inp[11]) ? node690 : node687;
												assign node687 = (inp[8]) ? 3'b000 : 3'b100;
												assign node690 = (inp[8]) ? 3'b100 : 3'b000;
										assign node693 = (inp[8]) ? node695 : 3'b000;
											assign node695 = (inp[11]) ? 3'b000 : 3'b100;
								assign node698 = (inp[10]) ? 3'b000 : node699;
									assign node699 = (inp[11]) ? node705 : node700;
										assign node700 = (inp[8]) ? 3'b100 : node701;
											assign node701 = (inp[5]) ? 3'b000 : 3'b100;
										assign node705 = (inp[2]) ? node707 : 3'b000;
											assign node707 = (inp[5]) ? 3'b000 : node708;
												assign node708 = (inp[8]) ? 3'b100 : 3'b000;
							assign node713 = (inp[5]) ? 3'b000 : node714;
								assign node714 = (inp[8]) ? node716 : 3'b000;
									assign node716 = (inp[10]) ? 3'b000 : node717;
										assign node717 = (inp[1]) ? 3'b000 : node718;
											assign node718 = (inp[2]) ? 3'b100 : 3'b000;
					assign node724 = (inp[10]) ? node884 : node725;
						assign node725 = (inp[0]) ? node809 : node726;
							assign node726 = (inp[4]) ? node764 : node727;
								assign node727 = (inp[8]) ? node743 : node728;
									assign node728 = (inp[1]) ? node734 : node729;
										assign node729 = (inp[5]) ? 3'b000 : node730;
											assign node730 = (inp[11]) ? 3'b000 : 3'b101;
										assign node734 = (inp[5]) ? 3'b110 : node735;
											assign node735 = (inp[11]) ? node739 : node736;
												assign node736 = (inp[2]) ? 3'b001 : 3'b101;
												assign node739 = (inp[2]) ? 3'b110 : 3'b010;
									assign node743 = (inp[1]) ? node753 : node744;
										assign node744 = (inp[5]) ? node748 : node745;
											assign node745 = (inp[11]) ? 3'b100 : 3'b000;
											assign node748 = (inp[11]) ? node750 : 3'b101;
												assign node750 = (inp[2]) ? 3'b000 : 3'b101;
										assign node753 = (inp[5]) ? node759 : node754;
											assign node754 = (inp[11]) ? node756 : 3'b101;
												assign node756 = (inp[2]) ? 3'b001 : 3'b101;
											assign node759 = (inp[2]) ? node761 : 3'b001;
												assign node761 = (inp[11]) ? 3'b110 : 3'b001;
								assign node764 = (inp[11]) ? node790 : node765;
									assign node765 = (inp[2]) ? node781 : node766;
										assign node766 = (inp[1]) ? node774 : node767;
											assign node767 = (inp[8]) ? node771 : node768;
												assign node768 = (inp[5]) ? 3'b100 : 3'b010;
												assign node771 = (inp[5]) ? 3'b010 : 3'b110;
											assign node774 = (inp[5]) ? node778 : node775;
												assign node775 = (inp[8]) ? 3'b001 : 3'b011;
												assign node778 = (inp[8]) ? 3'b110 : 3'b010;
										assign node781 = (inp[8]) ? node783 : 3'b010;
											assign node783 = (inp[1]) ? node787 : node784;
												assign node784 = (inp[5]) ? 3'b110 : 3'b010;
												assign node787 = (inp[5]) ? 3'b010 : 3'b110;
									assign node790 = (inp[1]) ? node800 : node791;
										assign node791 = (inp[8]) ? node795 : node792;
											assign node792 = (inp[5]) ? 3'b000 : 3'b100;
											assign node795 = (inp[5]) ? 3'b100 : node796;
												assign node796 = (inp[2]) ? 3'b010 : 3'b000;
										assign node800 = (inp[5]) ? node806 : node801;
											assign node801 = (inp[2]) ? node803 : 3'b110;
												assign node803 = (inp[8]) ? 3'b110 : 3'b010;
											assign node806 = (inp[8]) ? 3'b010 : 3'b100;
							assign node809 = (inp[4]) ? node851 : node810;
								assign node810 = (inp[2]) ? node828 : node811;
									assign node811 = (inp[1]) ? node821 : node812;
										assign node812 = (inp[8]) ? node818 : node813;
											assign node813 = (inp[5]) ? 3'b010 : node814;
												assign node814 = (inp[11]) ? 3'b110 : 3'b010;
											assign node818 = (inp[5]) ? 3'b110 : 3'b000;
										assign node821 = (inp[8]) ? node825 : node822;
											assign node822 = (inp[5]) ? 3'b100 : 3'b110;
											assign node825 = (inp[5]) ? 3'b010 : 3'b110;
									assign node828 = (inp[1]) ? node842 : node829;
										assign node829 = (inp[11]) ? node837 : node830;
											assign node830 = (inp[5]) ? node834 : node831;
												assign node831 = (inp[8]) ? 3'b010 : 3'b110;
												assign node834 = (inp[8]) ? 3'b110 : 3'b010;
											assign node837 = (inp[5]) ? node839 : 3'b110;
												assign node839 = (inp[8]) ? 3'b110 : 3'b010;
										assign node842 = (inp[8]) ? node846 : node843;
											assign node843 = (inp[5]) ? 3'b100 : 3'b010;
											assign node846 = (inp[11]) ? 3'b010 : node847;
												assign node847 = (inp[5]) ? 3'b010 : 3'b110;
								assign node851 = (inp[1]) ? node871 : node852;
									assign node852 = (inp[11]) ? node862 : node853;
										assign node853 = (inp[5]) ? node859 : node854;
											assign node854 = (inp[8]) ? node856 : 3'b010;
												assign node856 = (inp[2]) ? 3'b010 : 3'b110;
											assign node859 = (inp[8]) ? 3'b010 : 3'b100;
										assign node862 = (inp[5]) ? node868 : node863;
											assign node863 = (inp[8]) ? node865 : 3'b100;
												assign node865 = (inp[2]) ? 3'b010 : 3'b000;
											assign node868 = (inp[8]) ? 3'b100 : 3'b000;
									assign node871 = (inp[11]) ? node877 : node872;
										assign node872 = (inp[8]) ? 3'b100 : node873;
											assign node873 = (inp[5]) ? 3'b000 : 3'b100;
										assign node877 = (inp[5]) ? 3'b000 : node878;
											assign node878 = (inp[8]) ? node880 : 3'b000;
												assign node880 = (inp[2]) ? 3'b100 : 3'b000;
						assign node884 = (inp[4]) ? node946 : node885;
							assign node885 = (inp[5]) ? node921 : node886;
								assign node886 = (inp[0]) ? node906 : node887;
									assign node887 = (inp[1]) ? node897 : node888;
										assign node888 = (inp[8]) ? node892 : node889;
											assign node889 = (inp[11]) ? 3'b100 : 3'b000;
											assign node892 = (inp[11]) ? node894 : 3'b101;
												assign node894 = (inp[2]) ? 3'b000 : 3'b001;
										assign node897 = (inp[2]) ? node901 : node898;
											assign node898 = (inp[8]) ? 3'b001 : 3'b110;
											assign node901 = (inp[11]) ? node903 : 3'b110;
												assign node903 = (inp[8]) ? 3'b110 : 3'b010;
									assign node906 = (inp[1]) ? node914 : node907;
										assign node907 = (inp[8]) ? node909 : 3'b010;
											assign node909 = (inp[11]) ? node911 : 3'b110;
												assign node911 = (inp[2]) ? 3'b010 : 3'b110;
										assign node914 = (inp[8]) ? node916 : 3'b100;
											assign node916 = (inp[11]) ? node918 : 3'b010;
												assign node918 = (inp[2]) ? 3'b100 : 3'b000;
								assign node921 = (inp[8]) ? node935 : node922;
									assign node922 = (inp[1]) ? node928 : node923;
										assign node923 = (inp[2]) ? 3'b100 : node924;
											assign node924 = (inp[11]) ? 3'b100 : 3'b000;
										assign node928 = (inp[0]) ? node930 : 3'b001;
											assign node930 = (inp[2]) ? 3'b000 : node931;
												assign node931 = (inp[11]) ? 3'b000 : 3'b100;
									assign node935 = (inp[1]) ? node941 : node936;
										assign node936 = (inp[0]) ? 3'b010 : node937;
											assign node937 = (inp[2]) ? 3'b100 : 3'b000;
										assign node941 = (inp[0]) ? 3'b100 : node942;
											assign node942 = (inp[2]) ? 3'b010 : 3'b110;
							assign node946 = (inp[0]) ? node980 : node947;
								assign node947 = (inp[1]) ? node963 : node948;
									assign node948 = (inp[11]) ? node958 : node949;
										assign node949 = (inp[8]) ? node953 : node950;
											assign node950 = (inp[5]) ? 3'b000 : 3'b100;
											assign node953 = (inp[5]) ? 3'b100 : node954;
												assign node954 = (inp[2]) ? 3'b100 : 3'b000;
										assign node958 = (inp[8]) ? node960 : 3'b000;
											assign node960 = (inp[5]) ? 3'b000 : 3'b100;
									assign node963 = (inp[8]) ? node969 : node964;
										assign node964 = (inp[2]) ? node966 : 3'b100;
											assign node966 = (inp[11]) ? 3'b000 : 3'b100;
										assign node969 = (inp[2]) ? node977 : node970;
											assign node970 = (inp[5]) ? node974 : node971;
												assign node971 = (inp[11]) ? 3'b010 : 3'b110;
												assign node974 = (inp[11]) ? 3'b100 : 3'b010;
											assign node977 = (inp[5]) ? 3'b100 : 3'b000;
								assign node980 = (inp[1]) ? 3'b000 : node981;
									assign node981 = (inp[5]) ? node995 : node982;
										assign node982 = (inp[2]) ? node990 : node983;
											assign node983 = (inp[11]) ? node987 : node984;
												assign node984 = (inp[8]) ? 3'b000 : 3'b100;
												assign node987 = (inp[8]) ? 3'b100 : 3'b000;
											assign node990 = (inp[11]) ? node992 : 3'b100;
												assign node992 = (inp[8]) ? 3'b100 : 3'b000;
										assign node995 = (inp[11]) ? 3'b000 : node996;
											assign node996 = (inp[8]) ? 3'b100 : 3'b000;
			assign node1001 = (inp[9]) ? node1315 : node1002;
				assign node1002 = (inp[7]) ? node1082 : node1003;
					assign node1003 = (inp[4]) ? node1067 : node1004;
						assign node1004 = (inp[10]) ? node1048 : node1005;
							assign node1005 = (inp[11]) ? node1027 : node1006;
								assign node1006 = (inp[1]) ? node1012 : node1007;
									assign node1007 = (inp[8]) ? 3'b100 : node1008;
										assign node1008 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1012 = (inp[0]) ? node1022 : node1013;
										assign node1013 = (inp[5]) ? node1019 : node1014;
											assign node1014 = (inp[8]) ? node1016 : 3'b010;
												assign node1016 = (inp[2]) ? 3'b010 : 3'b110;
											assign node1019 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1022 = (inp[5]) ? 3'b000 : node1023;
											assign node1023 = (inp[2]) ? 3'b100 : 3'b000;
								assign node1027 = (inp[0]) ? node1039 : node1028;
									assign node1028 = (inp[1]) ? node1030 : 3'b000;
										assign node1030 = (inp[2]) ? node1032 : 3'b100;
											assign node1032 = (inp[8]) ? node1036 : node1033;
												assign node1033 = (inp[5]) ? 3'b000 : 3'b100;
												assign node1036 = (inp[5]) ? 3'b100 : 3'b010;
									assign node1039 = (inp[1]) ? 3'b000 : node1040;
										assign node1040 = (inp[5]) ? 3'b000 : node1041;
											assign node1041 = (inp[8]) ? node1043 : 3'b000;
												assign node1043 = (inp[2]) ? 3'b100 : 3'b000;
							assign node1048 = (inp[0]) ? 3'b000 : node1049;
								assign node1049 = (inp[1]) ? node1051 : 3'b000;
									assign node1051 = (inp[5]) ? node1061 : node1052;
										assign node1052 = (inp[2]) ? 3'b100 : node1053;
											assign node1053 = (inp[8]) ? node1057 : node1054;
												assign node1054 = (inp[11]) ? 3'b000 : 3'b100;
												assign node1057 = (inp[11]) ? 3'b100 : 3'b000;
										assign node1061 = (inp[11]) ? 3'b000 : node1062;
											assign node1062 = (inp[8]) ? 3'b100 : 3'b000;
						assign node1067 = (inp[8]) ? node1069 : 3'b000;
							assign node1069 = (inp[5]) ? 3'b000 : node1070;
								assign node1070 = (inp[11]) ? 3'b000 : node1071;
									assign node1071 = (inp[2]) ? node1073 : 3'b000;
										assign node1073 = (inp[0]) ? 3'b000 : node1074;
											assign node1074 = (inp[10]) ? 3'b000 : node1075;
												assign node1075 = (inp[1]) ? 3'b100 : 3'b000;
					assign node1082 = (inp[4]) ? node1250 : node1083;
						assign node1083 = (inp[0]) ? node1187 : node1084;
							assign node1084 = (inp[1]) ? node1142 : node1085;
								assign node1085 = (inp[11]) ? node1115 : node1086;
									assign node1086 = (inp[2]) ? node1100 : node1087;
										assign node1087 = (inp[5]) ? node1095 : node1088;
											assign node1088 = (inp[8]) ? node1092 : node1089;
												assign node1089 = (inp[10]) ? 3'b110 : 3'b100;
												assign node1092 = (inp[10]) ? 3'b000 : 3'b100;
											assign node1095 = (inp[8]) ? 3'b110 : node1096;
												assign node1096 = (inp[10]) ? 3'b100 : 3'b110;
										assign node1100 = (inp[10]) ? node1108 : node1101;
											assign node1101 = (inp[8]) ? node1105 : node1102;
												assign node1102 = (inp[5]) ? 3'b110 : 3'b000;
												assign node1105 = (inp[5]) ? 3'b000 : 3'b100;
											assign node1108 = (inp[5]) ? node1112 : node1109;
												assign node1109 = (inp[8]) ? 3'b000 : 3'b110;
												assign node1112 = (inp[8]) ? 3'b110 : 3'b000;
									assign node1115 = (inp[8]) ? node1129 : node1116;
										assign node1116 = (inp[2]) ? node1122 : node1117;
											assign node1117 = (inp[5]) ? node1119 : 3'b010;
												assign node1119 = (inp[10]) ? 3'b010 : 3'b110;
											assign node1122 = (inp[5]) ? node1126 : node1123;
												assign node1123 = (inp[10]) ? 3'b110 : 3'b010;
												assign node1126 = (inp[10]) ? 3'b010 : 3'b110;
										assign node1129 = (inp[10]) ? node1137 : node1130;
											assign node1130 = (inp[5]) ? node1134 : node1131;
												assign node1131 = (inp[2]) ? 3'b000 : 3'b100;
												assign node1134 = (inp[2]) ? 3'b010 : 3'b000;
											assign node1137 = (inp[5]) ? 3'b110 : node1138;
												assign node1138 = (inp[2]) ? 3'b110 : 3'b000;
								assign node1142 = (inp[11]) ? node1172 : node1143;
									assign node1143 = (inp[2]) ? node1157 : node1144;
										assign node1144 = (inp[8]) ? node1150 : node1145;
											assign node1145 = (inp[5]) ? node1147 : 3'b010;
												assign node1147 = (inp[10]) ? 3'b000 : 3'b010;
											assign node1150 = (inp[10]) ? node1154 : node1151;
												assign node1151 = (inp[5]) ? 3'b110 : 3'b000;
												assign node1154 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1157 = (inp[8]) ? node1165 : node1158;
											assign node1158 = (inp[10]) ? node1162 : node1159;
												assign node1159 = (inp[5]) ? 3'b010 : 3'b110;
												assign node1162 = (inp[5]) ? 3'b100 : 3'b010;
											assign node1165 = (inp[5]) ? node1169 : node1166;
												assign node1166 = (inp[10]) ? 3'b110 : 3'b001;
												assign node1169 = (inp[10]) ? 3'b010 : 3'b110;
									assign node1172 = (inp[10]) ? node1180 : node1173;
										assign node1173 = (inp[2]) ? node1175 : 3'b100;
											assign node1175 = (inp[5]) ? 3'b010 : node1176;
												assign node1176 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1180 = (inp[2]) ? 3'b100 : node1181;
											assign node1181 = (inp[8]) ? 3'b010 : node1182;
												assign node1182 = (inp[5]) ? 3'b100 : 3'b110;
							assign node1187 = (inp[10]) ? node1215 : node1188;
								assign node1188 = (inp[5]) ? node1202 : node1189;
									assign node1189 = (inp[1]) ? node1197 : node1190;
										assign node1190 = (inp[11]) ? node1192 : 3'b110;
											assign node1192 = (inp[8]) ? node1194 : 3'b010;
												assign node1194 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1197 = (inp[11]) ? 3'b100 : node1198;
											assign node1198 = (inp[8]) ? 3'b010 : 3'b000;
									assign node1202 = (inp[8]) ? node1210 : node1203;
										assign node1203 = (inp[1]) ? node1205 : 3'b100;
											assign node1205 = (inp[11]) ? 3'b000 : node1206;
												assign node1206 = (inp[2]) ? 3'b000 : 3'b100;
										assign node1210 = (inp[2]) ? 3'b100 : node1211;
											assign node1211 = (inp[11]) ? 3'b100 : 3'b010;
								assign node1215 = (inp[11]) ? node1239 : node1216;
									assign node1216 = (inp[2]) ? node1228 : node1217;
										assign node1217 = (inp[1]) ? node1223 : node1218;
											assign node1218 = (inp[5]) ? 3'b100 : node1219;
												assign node1219 = (inp[8]) ? 3'b010 : 3'b100;
											assign node1223 = (inp[5]) ? node1225 : 3'b100;
												assign node1225 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1228 = (inp[8]) ? node1234 : node1229;
											assign node1229 = (inp[5]) ? 3'b000 : node1230;
												assign node1230 = (inp[1]) ? 3'b000 : 3'b100;
											assign node1234 = (inp[1]) ? node1236 : 3'b100;
												assign node1236 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1239 = (inp[1]) ? 3'b000 : node1240;
										assign node1240 = (inp[5]) ? node1246 : node1241;
											assign node1241 = (inp[2]) ? 3'b100 : node1242;
												assign node1242 = (inp[8]) ? 3'b000 : 3'b100;
											assign node1246 = (inp[8]) ? 3'b100 : 3'b000;
						assign node1250 = (inp[0]) ? node1302 : node1251;
							assign node1251 = (inp[1]) ? node1267 : node1252;
								assign node1252 = (inp[10]) ? 3'b000 : node1253;
									assign node1253 = (inp[11]) ? node1259 : node1254;
										assign node1254 = (inp[5]) ? node1256 : 3'b100;
											assign node1256 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1259 = (inp[5]) ? 3'b000 : node1260;
											assign node1260 = (inp[2]) ? node1262 : 3'b000;
												assign node1262 = (inp[8]) ? 3'b100 : 3'b000;
								assign node1267 = (inp[10]) ? node1287 : node1268;
									assign node1268 = (inp[11]) ? node1278 : node1269;
										assign node1269 = (inp[8]) ? node1273 : node1270;
											assign node1270 = (inp[5]) ? 3'b100 : 3'b010;
											assign node1273 = (inp[2]) ? 3'b010 : node1274;
												assign node1274 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1278 = (inp[2]) ? node1280 : 3'b100;
											assign node1280 = (inp[8]) ? node1284 : node1281;
												assign node1281 = (inp[5]) ? 3'b000 : 3'b100;
												assign node1284 = (inp[5]) ? 3'b100 : 3'b010;
									assign node1287 = (inp[8]) ? node1293 : node1288;
										assign node1288 = (inp[5]) ? 3'b000 : node1289;
											assign node1289 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1293 = (inp[5]) ? node1299 : node1294;
											assign node1294 = (inp[11]) ? 3'b100 : node1295;
												assign node1295 = (inp[2]) ? 3'b100 : 3'b000;
											assign node1299 = (inp[11]) ? 3'b000 : 3'b100;
							assign node1302 = (inp[1]) ? 3'b000 : node1303;
								assign node1303 = (inp[10]) ? 3'b000 : node1304;
									assign node1304 = (inp[11]) ? node1306 : 3'b100;
										assign node1306 = (inp[5]) ? 3'b000 : node1307;
											assign node1307 = (inp[2]) ? node1309 : 3'b000;
												assign node1309 = (inp[8]) ? 3'b100 : 3'b000;
				assign node1315 = (inp[7]) ? node1317 : 3'b000;
					assign node1317 = (inp[4]) ? 3'b000 : node1318;
						assign node1318 = (inp[0]) ? node1346 : node1319;
							assign node1319 = (inp[1]) ? node1325 : node1320;
								assign node1320 = (inp[10]) ? node1322 : 3'b010;
									assign node1322 = (inp[5]) ? 3'b000 : 3'b010;
								assign node1325 = (inp[10]) ? node1339 : node1326;
									assign node1326 = (inp[5]) ? node1334 : node1327;
										assign node1327 = (inp[8]) ? node1329 : 3'b100;
											assign node1329 = (inp[11]) ? 3'b100 : node1330;
												assign node1330 = (inp[2]) ? 3'b010 : 3'b000;
										assign node1334 = (inp[8]) ? node1336 : 3'b000;
											assign node1336 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1339 = (inp[8]) ? node1341 : 3'b000;
										assign node1341 = (inp[11]) ? 3'b000 : node1342;
											assign node1342 = (inp[5]) ? 3'b000 : 3'b100;
							assign node1346 = (inp[10]) ? 3'b000 : node1347;
								assign node1347 = (inp[5]) ? 3'b000 : node1348;
									assign node1348 = (inp[2]) ? node1350 : 3'b000;
										assign node1350 = (inp[8]) ? node1352 : 3'b000;
											assign node1352 = (inp[11]) ? 3'b000 : node1353;
												assign node1353 = (inp[1]) ? 3'b000 : 3'b100;
		assign node1360 = (inp[3]) ? node2372 : node1361;
			assign node1361 = (inp[9]) ? node1777 : node1362;
				assign node1362 = (inp[0]) ? node1496 : node1363;
					assign node1363 = (inp[1]) ? node1393 : node1364;
						assign node1364 = (inp[7]) ? 3'b111 : node1365;
							assign node1365 = (inp[4]) ? node1367 : 3'b111;
								assign node1367 = (inp[10]) ? node1375 : node1368;
									assign node1368 = (inp[2]) ? node1370 : 3'b111;
										assign node1370 = (inp[5]) ? node1372 : 3'b111;
											assign node1372 = (inp[11]) ? 3'b011 : 3'b111;
									assign node1375 = (inp[2]) ? node1381 : node1376;
										assign node1376 = (inp[11]) ? 3'b011 : node1377;
											assign node1377 = (inp[5]) ? 3'b011 : 3'b111;
										assign node1381 = (inp[8]) ? node1387 : node1382;
											assign node1382 = (inp[5]) ? node1384 : 3'b111;
												assign node1384 = (inp[11]) ? 3'b111 : 3'b011;
											assign node1387 = (inp[11]) ? node1389 : 3'b011;
												assign node1389 = (inp[5]) ? 3'b111 : 3'b011;
						assign node1393 = (inp[7]) ? node1469 : node1394;
							assign node1394 = (inp[4]) ? node1438 : node1395;
								assign node1395 = (inp[2]) ? node1417 : node1396;
									assign node1396 = (inp[8]) ? node1404 : node1397;
										assign node1397 = (inp[5]) ? node1399 : 3'b011;
											assign node1399 = (inp[11]) ? node1401 : 3'b011;
												assign node1401 = (inp[10]) ? 3'b010 : 3'b011;
										assign node1404 = (inp[10]) ? node1410 : node1405;
											assign node1405 = (inp[5]) ? node1407 : 3'b010;
												assign node1407 = (inp[11]) ? 3'b111 : 3'b011;
											assign node1410 = (inp[11]) ? node1414 : node1411;
												assign node1411 = (inp[5]) ? 3'b111 : 3'b011;
												assign node1414 = (inp[5]) ? 3'b011 : 3'b111;
									assign node1417 = (inp[10]) ? node1427 : node1418;
										assign node1418 = (inp[5]) ? node1422 : node1419;
											assign node1419 = (inp[8]) ? 3'b011 : 3'b111;
											assign node1422 = (inp[11]) ? node1424 : 3'b111;
												assign node1424 = (inp[8]) ? 3'b111 : 3'b011;
										assign node1427 = (inp[11]) ? node1433 : node1428;
											assign node1428 = (inp[8]) ? node1430 : 3'b011;
												assign node1430 = (inp[5]) ? 3'b011 : 3'b111;
											assign node1433 = (inp[8]) ? node1435 : 3'b110;
												assign node1435 = (inp[5]) ? 3'b011 : 3'b111;
								assign node1438 = (inp[8]) ? node1454 : node1439;
									assign node1439 = (inp[10]) ? node1447 : node1440;
										assign node1440 = (inp[11]) ? 3'b101 : node1441;
											assign node1441 = (inp[5]) ? 3'b101 : node1442;
												assign node1442 = (inp[2]) ? 3'b011 : 3'b111;
										assign node1447 = (inp[11]) ? 3'b001 : node1448;
											assign node1448 = (inp[5]) ? node1450 : 3'b101;
												assign node1450 = (inp[2]) ? 3'b001 : 3'b101;
									assign node1454 = (inp[10]) ? node1460 : node1455;
										assign node1455 = (inp[11]) ? 3'b011 : node1456;
											assign node1456 = (inp[5]) ? 3'b011 : 3'b111;
										assign node1460 = (inp[11]) ? node1464 : node1461;
											assign node1461 = (inp[5]) ? 3'b101 : 3'b011;
											assign node1464 = (inp[5]) ? node1466 : 3'b101;
												assign node1466 = (inp[2]) ? 3'b001 : 3'b101;
							assign node1469 = (inp[4]) ? node1471 : 3'b111;
								assign node1471 = (inp[10]) ? node1483 : node1472;
									assign node1472 = (inp[5]) ? node1478 : node1473;
										assign node1473 = (inp[8]) ? 3'b111 : node1474;
											assign node1474 = (inp[11]) ? 3'b101 : 3'b111;
										assign node1478 = (inp[11]) ? node1480 : 3'b111;
											assign node1480 = (inp[8]) ? 3'b111 : 3'b011;
									assign node1483 = (inp[11]) ? node1491 : node1484;
										assign node1484 = (inp[8]) ? node1486 : 3'b011;
											assign node1486 = (inp[5]) ? node1488 : 3'b111;
												assign node1488 = (inp[2]) ? 3'b011 : 3'b111;
										assign node1491 = (inp[8]) ? 3'b011 : node1492;
											assign node1492 = (inp[5]) ? 3'b101 : 3'b011;
					assign node1496 = (inp[4]) ? node1634 : node1497;
						assign node1497 = (inp[7]) ? node1579 : node1498;
							assign node1498 = (inp[1]) ? node1536 : node1499;
								assign node1499 = (inp[10]) ? node1517 : node1500;
									assign node1500 = (inp[11]) ? node1508 : node1501;
										assign node1501 = (inp[8]) ? node1503 : 3'b011;
											assign node1503 = (inp[2]) ? node1505 : 3'b111;
												assign node1505 = (inp[5]) ? 3'b011 : 3'b111;
										assign node1508 = (inp[5]) ? node1514 : node1509;
											assign node1509 = (inp[8]) ? 3'b111 : node1510;
												assign node1510 = (inp[2]) ? 3'b011 : 3'b111;
											assign node1514 = (inp[8]) ? 3'b011 : 3'b101;
									assign node1517 = (inp[11]) ? node1527 : node1518;
										assign node1518 = (inp[5]) ? node1524 : node1519;
											assign node1519 = (inp[8]) ? node1521 : 3'b111;
												assign node1521 = (inp[2]) ? 3'b011 : 3'b111;
											assign node1524 = (inp[2]) ? 3'b101 : 3'b111;
										assign node1527 = (inp[5]) ? node1531 : node1528;
											assign node1528 = (inp[8]) ? 3'b011 : 3'b101;
											assign node1531 = (inp[2]) ? node1533 : 3'b101;
												assign node1533 = (inp[8]) ? 3'b101 : 3'b001;
								assign node1536 = (inp[10]) ? node1560 : node1537;
									assign node1537 = (inp[5]) ? node1549 : node1538;
										assign node1538 = (inp[8]) ? node1544 : node1539;
											assign node1539 = (inp[11]) ? node1541 : 3'b011;
												assign node1541 = (inp[2]) ? 3'b101 : 3'b001;
											assign node1544 = (inp[2]) ? 3'b011 : node1545;
												assign node1545 = (inp[11]) ? 3'b010 : 3'b111;
										assign node1549 = (inp[8]) ? node1555 : node1550;
											assign node1550 = (inp[2]) ? node1552 : 3'b101;
												assign node1552 = (inp[11]) ? 3'b001 : 3'b101;
											assign node1555 = (inp[11]) ? node1557 : 3'b011;
												assign node1557 = (inp[2]) ? 3'b101 : 3'b001;
									assign node1560 = (inp[11]) ? node1570 : node1561;
										assign node1561 = (inp[5]) ? node1567 : node1562;
											assign node1562 = (inp[8]) ? node1564 : 3'b101;
												assign node1564 = (inp[2]) ? 3'b101 : 3'b001;
											assign node1567 = (inp[8]) ? 3'b101 : 3'b001;
										assign node1570 = (inp[5]) ? node1576 : node1571;
											assign node1571 = (inp[2]) ? node1573 : 3'b001;
												assign node1573 = (inp[8]) ? 3'b101 : 3'b001;
											assign node1576 = (inp[2]) ? 3'b110 : 3'b010;
							assign node1579 = (inp[1]) ? node1591 : node1580;
								assign node1580 = (inp[11]) ? node1582 : 3'b111;
									assign node1582 = (inp[10]) ? node1584 : 3'b111;
										assign node1584 = (inp[8]) ? node1586 : 3'b011;
											assign node1586 = (inp[2]) ? node1588 : 3'b111;
												assign node1588 = (inp[5]) ? 3'b011 : 3'b111;
								assign node1591 = (inp[5]) ? node1619 : node1592;
									assign node1592 = (inp[8]) ? node1606 : node1593;
										assign node1593 = (inp[2]) ? node1601 : node1594;
											assign node1594 = (inp[10]) ? node1598 : node1595;
												assign node1595 = (inp[11]) ? 3'b011 : 3'b111;
												assign node1598 = (inp[11]) ? 3'b111 : 3'b011;
											assign node1601 = (inp[11]) ? 3'b011 : node1602;
												assign node1602 = (inp[10]) ? 3'b011 : 3'b111;
										assign node1606 = (inp[11]) ? node1612 : node1607;
											assign node1607 = (inp[10]) ? 3'b111 : node1608;
												assign node1608 = (inp[2]) ? 3'b111 : 3'b101;
											assign node1612 = (inp[10]) ? node1616 : node1613;
												assign node1613 = (inp[2]) ? 3'b111 : 3'b011;
												assign node1616 = (inp[2]) ? 3'b011 : 3'b111;
									assign node1619 = (inp[10]) ? node1627 : node1620;
										assign node1620 = (inp[8]) ? node1622 : 3'b011;
											assign node1622 = (inp[11]) ? node1624 : 3'b111;
												assign node1624 = (inp[2]) ? 3'b011 : 3'b111;
										assign node1627 = (inp[8]) ? node1629 : 3'b101;
											assign node1629 = (inp[11]) ? node1631 : 3'b011;
												assign node1631 = (inp[2]) ? 3'b101 : 3'b001;
						assign node1634 = (inp[7]) ? node1706 : node1635;
							assign node1635 = (inp[10]) ? node1669 : node1636;
								assign node1636 = (inp[1]) ? node1656 : node1637;
									assign node1637 = (inp[8]) ? node1645 : node1638;
										assign node1638 = (inp[5]) ? 3'b001 : node1639;
											assign node1639 = (inp[2]) ? node1641 : 3'b001;
												assign node1641 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1645 = (inp[5]) ? node1651 : node1646;
											assign node1646 = (inp[11]) ? node1648 : 3'b011;
												assign node1648 = (inp[2]) ? 3'b101 : 3'b011;
											assign node1651 = (inp[2]) ? node1653 : 3'b101;
												assign node1653 = (inp[11]) ? 3'b001 : 3'b101;
									assign node1656 = (inp[8]) ? node1662 : node1657;
										assign node1657 = (inp[5]) ? 3'b110 : node1658;
											assign node1658 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1662 = (inp[5]) ? 3'b001 : node1663;
											assign node1663 = (inp[2]) ? node1665 : 3'b101;
												assign node1665 = (inp[11]) ? 3'b001 : 3'b101;
								assign node1669 = (inp[1]) ? node1691 : node1670;
									assign node1670 = (inp[8]) ? node1680 : node1671;
										assign node1671 = (inp[5]) ? node1675 : node1672;
											assign node1672 = (inp[11]) ? 3'b000 : 3'b001;
											assign node1675 = (inp[11]) ? 3'b110 : node1676;
												assign node1676 = (inp[2]) ? 3'b110 : 3'b010;
										assign node1680 = (inp[5]) ? node1686 : node1681;
											assign node1681 = (inp[2]) ? node1683 : 3'b101;
												assign node1683 = (inp[11]) ? 3'b001 : 3'b101;
											assign node1686 = (inp[2]) ? node1688 : 3'b001;
												assign node1688 = (inp[11]) ? 3'b110 : 3'b001;
									assign node1691 = (inp[11]) ? node1697 : node1692;
										assign node1692 = (inp[5]) ? 3'b110 : node1693;
											assign node1693 = (inp[2]) ? 3'b110 : 3'b001;
										assign node1697 = (inp[5]) ? node1703 : node1698;
											assign node1698 = (inp[2]) ? 3'b110 : node1699;
												assign node1699 = (inp[8]) ? 3'b010 : 3'b110;
											assign node1703 = (inp[8]) ? 3'b110 : 3'b010;
							assign node1706 = (inp[1]) ? node1746 : node1707;
								assign node1707 = (inp[10]) ? node1725 : node1708;
									assign node1708 = (inp[11]) ? node1716 : node1709;
										assign node1709 = (inp[8]) ? node1711 : 3'b011;
											assign node1711 = (inp[5]) ? node1713 : 3'b111;
												assign node1713 = (inp[2]) ? 3'b011 : 3'b111;
										assign node1716 = (inp[5]) ? node1722 : node1717;
											assign node1717 = (inp[8]) ? 3'b111 : node1718;
												assign node1718 = (inp[2]) ? 3'b011 : 3'b111;
											assign node1722 = (inp[8]) ? 3'b011 : 3'b101;
									assign node1725 = (inp[5]) ? node1735 : node1726;
										assign node1726 = (inp[8]) ? node1730 : node1727;
											assign node1727 = (inp[11]) ? 3'b101 : 3'b111;
											assign node1730 = (inp[11]) ? 3'b011 : node1731;
												assign node1731 = (inp[2]) ? 3'b011 : 3'b111;
										assign node1735 = (inp[2]) ? node1741 : node1736;
											assign node1736 = (inp[11]) ? 3'b101 : node1737;
												assign node1737 = (inp[8]) ? 3'b011 : 3'b111;
											assign node1741 = (inp[11]) ? node1743 : 3'b101;
												assign node1743 = (inp[8]) ? 3'b101 : 3'b001;
								assign node1746 = (inp[11]) ? node1756 : node1747;
									assign node1747 = (inp[10]) ? node1753 : node1748;
										assign node1748 = (inp[5]) ? 3'b101 : node1749;
											assign node1749 = (inp[8]) ? 3'b011 : 3'b101;
										assign node1753 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1756 = (inp[8]) ? node1768 : node1757;
										assign node1757 = (inp[10]) ? node1763 : node1758;
											assign node1758 = (inp[2]) ? node1760 : 3'b001;
												assign node1760 = (inp[5]) ? 3'b001 : 3'b101;
											assign node1763 = (inp[5]) ? node1765 : 3'b001;
												assign node1765 = (inp[2]) ? 3'b110 : 3'b010;
										assign node1768 = (inp[5]) ? node1774 : node1769;
											assign node1769 = (inp[10]) ? 3'b101 : node1770;
												assign node1770 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1774 = (inp[10]) ? 3'b001 : 3'b101;
				assign node1777 = (inp[0]) ? node2057 : node1778;
					assign node1778 = (inp[4]) ? node1922 : node1779;
						assign node1779 = (inp[7]) ? node1863 : node1780;
							assign node1780 = (inp[10]) ? node1822 : node1781;
								assign node1781 = (inp[8]) ? node1803 : node1782;
									assign node1782 = (inp[11]) ? node1794 : node1783;
										assign node1783 = (inp[2]) ? node1789 : node1784;
											assign node1784 = (inp[1]) ? node1786 : 3'b011;
												assign node1786 = (inp[5]) ? 3'b111 : 3'b011;
											assign node1789 = (inp[5]) ? 3'b101 : node1790;
												assign node1790 = (inp[1]) ? 3'b111 : 3'b011;
										assign node1794 = (inp[1]) ? node1798 : node1795;
											assign node1795 = (inp[5]) ? 3'b101 : 3'b011;
											assign node1798 = (inp[2]) ? node1800 : 3'b001;
												assign node1800 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1803 = (inp[1]) ? node1815 : node1804;
										assign node1804 = (inp[5]) ? node1810 : node1805;
											assign node1805 = (inp[11]) ? node1807 : 3'b111;
												assign node1807 = (inp[2]) ? 3'b011 : 3'b111;
											assign node1810 = (inp[2]) ? 3'b011 : node1811;
												assign node1811 = (inp[11]) ? 3'b011 : 3'b111;
										assign node1815 = (inp[5]) ? node1817 : 3'b011;
											assign node1817 = (inp[11]) ? 3'b101 : node1818;
												assign node1818 = (inp[2]) ? 3'b101 : 3'b011;
								assign node1822 = (inp[1]) ? node1842 : node1823;
									assign node1823 = (inp[8]) ? node1831 : node1824;
										assign node1824 = (inp[5]) ? node1826 : 3'b101;
											assign node1826 = (inp[11]) ? 3'b001 : node1827;
												assign node1827 = (inp[2]) ? 3'b111 : 3'b101;
										assign node1831 = (inp[11]) ? node1837 : node1832;
											assign node1832 = (inp[2]) ? node1834 : 3'b011;
												assign node1834 = (inp[5]) ? 3'b111 : 3'b011;
											assign node1837 = (inp[5]) ? 3'b101 : node1838;
												assign node1838 = (inp[2]) ? 3'b111 : 3'b011;
									assign node1842 = (inp[8]) ? node1854 : node1843;
										assign node1843 = (inp[2]) ? node1849 : node1844;
											assign node1844 = (inp[5]) ? 3'b001 : node1845;
												assign node1845 = (inp[11]) ? 3'b001 : 3'b101;
											assign node1849 = (inp[5]) ? node1851 : 3'b001;
												assign node1851 = (inp[11]) ? 3'b111 : 3'b001;
										assign node1854 = (inp[2]) ? 3'b101 : node1855;
											assign node1855 = (inp[5]) ? node1859 : node1856;
												assign node1856 = (inp[11]) ? 3'b101 : 3'b001;
												assign node1859 = (inp[11]) ? 3'b001 : 3'b101;
							assign node1863 = (inp[10]) ? node1891 : node1864;
								assign node1864 = (inp[8]) ? node1882 : node1865;
									assign node1865 = (inp[11]) ? node1871 : node1866;
										assign node1866 = (inp[5]) ? node1868 : 3'b111;
											assign node1868 = (inp[1]) ? 3'b011 : 3'b111;
										assign node1871 = (inp[5]) ? node1877 : node1872;
											assign node1872 = (inp[1]) ? node1874 : 3'b011;
												assign node1874 = (inp[2]) ? 3'b011 : 3'b111;
											assign node1877 = (inp[1]) ? node1879 : 3'b111;
												assign node1879 = (inp[2]) ? 3'b111 : 3'b011;
									assign node1882 = (inp[1]) ? node1884 : 3'b111;
										assign node1884 = (inp[2]) ? node1886 : 3'b111;
											assign node1886 = (inp[5]) ? node1888 : 3'b111;
												assign node1888 = (inp[11]) ? 3'b011 : 3'b111;
								assign node1891 = (inp[1]) ? node1907 : node1892;
									assign node1892 = (inp[8]) ? node1900 : node1893;
										assign node1893 = (inp[2]) ? 3'b011 : node1894;
											assign node1894 = (inp[5]) ? 3'b011 : node1895;
												assign node1895 = (inp[11]) ? 3'b111 : 3'b011;
										assign node1900 = (inp[2]) ? node1902 : 3'b111;
											assign node1902 = (inp[11]) ? 3'b111 : node1903;
												assign node1903 = (inp[5]) ? 3'b011 : 3'b111;
									assign node1907 = (inp[8]) ? node1915 : node1908;
										assign node1908 = (inp[5]) ? 3'b101 : node1909;
											assign node1909 = (inp[11]) ? node1911 : 3'b001;
												assign node1911 = (inp[2]) ? 3'b111 : 3'b011;
										assign node1915 = (inp[5]) ? node1919 : node1916;
											assign node1916 = (inp[11]) ? 3'b011 : 3'b111;
											assign node1919 = (inp[2]) ? 3'b001 : 3'b011;
						assign node1922 = (inp[7]) ? node1988 : node1923;
							assign node1923 = (inp[10]) ? node1949 : node1924;
								assign node1924 = (inp[1]) ? node1934 : node1925;
									assign node1925 = (inp[11]) ? 3'b101 : node1926;
										assign node1926 = (inp[8]) ? node1928 : 3'b001;
											assign node1928 = (inp[5]) ? 3'b101 : node1929;
												assign node1929 = (inp[2]) ? 3'b101 : 3'b011;
									assign node1934 = (inp[8]) ? node1942 : node1935;
										assign node1935 = (inp[5]) ? 3'b110 : node1936;
											assign node1936 = (inp[11]) ? 3'b010 : node1937;
												assign node1937 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1942 = (inp[11]) ? node1946 : node1943;
											assign node1943 = (inp[5]) ? 3'b001 : 3'b101;
											assign node1946 = (inp[5]) ? 3'b110 : 3'b001;
								assign node1949 = (inp[11]) ? node1969 : node1950;
									assign node1950 = (inp[8]) ? node1958 : node1951;
										assign node1951 = (inp[5]) ? node1953 : 3'b110;
											assign node1953 = (inp[1]) ? node1955 : 3'b110;
												assign node1955 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1958 = (inp[5]) ? node1964 : node1959;
											assign node1959 = (inp[2]) ? 3'b011 : node1960;
												assign node1960 = (inp[1]) ? 3'b001 : 3'b101;
											assign node1964 = (inp[1]) ? 3'b110 : node1965;
												assign node1965 = (inp[2]) ? 3'b110 : 3'b001;
									assign node1969 = (inp[1]) ? node1977 : node1970;
										assign node1970 = (inp[8]) ? node1972 : 3'b000;
											assign node1972 = (inp[2]) ? node1974 : 3'b001;
												assign node1974 = (inp[5]) ? 3'b000 : 3'b001;
										assign node1977 = (inp[8]) ? node1983 : node1978;
											assign node1978 = (inp[5]) ? 3'b010 : node1979;
												assign node1979 = (inp[2]) ? 3'b010 : 3'b110;
											assign node1983 = (inp[5]) ? 3'b110 : node1984;
												assign node1984 = (inp[2]) ? 3'b110 : 3'b001;
							assign node1988 = (inp[1]) ? node2026 : node1989;
								assign node1989 = (inp[8]) ? node2013 : node1990;
									assign node1990 = (inp[11]) ? node2006 : node1991;
										assign node1991 = (inp[5]) ? node1999 : node1992;
											assign node1992 = (inp[10]) ? node1996 : node1993;
												assign node1993 = (inp[2]) ? 3'b011 : 3'b101;
												assign node1996 = (inp[2]) ? 3'b101 : 3'b011;
											assign node1999 = (inp[10]) ? node2003 : node2000;
												assign node2000 = (inp[2]) ? 3'b101 : 3'b011;
												assign node2003 = (inp[2]) ? 3'b111 : 3'b101;
										assign node2006 = (inp[5]) ? node2010 : node2007;
											assign node2007 = (inp[2]) ? 3'b101 : 3'b011;
											assign node2010 = (inp[10]) ? 3'b001 : 3'b101;
									assign node2013 = (inp[10]) ? node2019 : node2014;
										assign node2014 = (inp[5]) ? node2016 : 3'b111;
											assign node2016 = (inp[11]) ? 3'b011 : 3'b111;
										assign node2019 = (inp[2]) ? node2021 : 3'b011;
											assign node2021 = (inp[5]) ? 3'b111 : node2022;
												assign node2022 = (inp[11]) ? 3'b111 : 3'b011;
								assign node2026 = (inp[10]) ? node2042 : node2027;
									assign node2027 = (inp[5]) ? node2035 : node2028;
										assign node2028 = (inp[11]) ? node2030 : 3'b011;
											assign node2030 = (inp[8]) ? 3'b011 : node2031;
												assign node2031 = (inp[2]) ? 3'b101 : 3'b001;
										assign node2035 = (inp[2]) ? 3'b101 : node2036;
											assign node2036 = (inp[11]) ? node2038 : 3'b111;
												assign node2038 = (inp[8]) ? 3'b101 : 3'b001;
									assign node2042 = (inp[5]) ? node2048 : node2043;
										assign node2043 = (inp[11]) ? node2045 : 3'b101;
											assign node2045 = (inp[8]) ? 3'b101 : 3'b001;
										assign node2048 = (inp[2]) ? node2054 : node2049;
											assign node2049 = (inp[8]) ? node2051 : 3'b001;
												assign node2051 = (inp[11]) ? 3'b001 : 3'b101;
											assign node2054 = (inp[11]) ? 3'b110 : 3'b001;
					assign node2057 = (inp[7]) ? node2205 : node2058;
						assign node2058 = (inp[10]) ? node2130 : node2059;
							assign node2059 = (inp[4]) ? node2097 : node2060;
								assign node2060 = (inp[1]) ? node2074 : node2061;
									assign node2061 = (inp[8]) ? node2069 : node2062;
										assign node2062 = (inp[11]) ? node2064 : 3'b001;
											assign node2064 = (inp[5]) ? 3'b110 : node2065;
												assign node2065 = (inp[2]) ? 3'b001 : 3'b101;
										assign node2069 = (inp[5]) ? node2071 : 3'b101;
											assign node2071 = (inp[2]) ? 3'b001 : 3'b101;
									assign node2074 = (inp[11]) ? node2084 : node2075;
										assign node2075 = (inp[8]) ? node2079 : node2076;
											assign node2076 = (inp[5]) ? 3'b110 : 3'b001;
											assign node2079 = (inp[5]) ? 3'b001 : node2080;
												assign node2080 = (inp[2]) ? 3'b001 : 3'b101;
										assign node2084 = (inp[5]) ? node2090 : node2085;
											assign node2085 = (inp[8]) ? 3'b001 : node2086;
												assign node2086 = (inp[2]) ? 3'b110 : 3'b010;
											assign node2090 = (inp[2]) ? node2094 : node2091;
												assign node2091 = (inp[8]) ? 3'b010 : 3'b110;
												assign node2094 = (inp[8]) ? 3'b110 : 3'b010;
								assign node2097 = (inp[5]) ? node2119 : node2098;
									assign node2098 = (inp[1]) ? node2112 : node2099;
										assign node2099 = (inp[2]) ? node2105 : node2100;
											assign node2100 = (inp[8]) ? 3'b001 : node2101;
												assign node2101 = (inp[11]) ? 3'b101 : 3'b010;
											assign node2105 = (inp[11]) ? node2109 : node2106;
												assign node2106 = (inp[8]) ? 3'b001 : 3'b110;
												assign node2109 = (inp[8]) ? 3'b110 : 3'b010;
										assign node2112 = (inp[11]) ? node2114 : 3'b110;
											assign node2114 = (inp[8]) ? node2116 : 3'b010;
												assign node2116 = (inp[2]) ? 3'b010 : 3'b110;
									assign node2119 = (inp[1]) ? node2127 : node2120;
										assign node2120 = (inp[8]) ? node2122 : 3'b010;
											assign node2122 = (inp[11]) ? node2124 : 3'b110;
												assign node2124 = (inp[2]) ? 3'b010 : 3'b110;
										assign node2127 = (inp[8]) ? 3'b010 : 3'b100;
							assign node2130 = (inp[4]) ? node2172 : node2131;
								assign node2131 = (inp[1]) ? node2149 : node2132;
									assign node2132 = (inp[8]) ? node2140 : node2133;
										assign node2133 = (inp[5]) ? node2135 : 3'b110;
											assign node2135 = (inp[11]) ? node2137 : 3'b110;
												assign node2137 = (inp[2]) ? 3'b010 : 3'b110;
										assign node2140 = (inp[5]) ? node2144 : node2141;
											assign node2141 = (inp[11]) ? 3'b001 : 3'b011;
											assign node2144 = (inp[2]) ? 3'b110 : node2145;
												assign node2145 = (inp[11]) ? 3'b110 : 3'b001;
									assign node2149 = (inp[5]) ? node2163 : node2150;
										assign node2150 = (inp[11]) ? node2156 : node2151;
											assign node2151 = (inp[2]) ? 3'b110 : node2152;
												assign node2152 = (inp[8]) ? 3'b010 : 3'b110;
											assign node2156 = (inp[8]) ? node2160 : node2157;
												assign node2157 = (inp[2]) ? 3'b010 : 3'b110;
												assign node2160 = (inp[2]) ? 3'b110 : 3'b010;
										assign node2163 = (inp[8]) ? node2169 : node2164;
											assign node2164 = (inp[11]) ? node2166 : 3'b010;
												assign node2166 = (inp[2]) ? 3'b100 : 3'b000;
											assign node2169 = (inp[11]) ? 3'b010 : 3'b110;
								assign node2172 = (inp[1]) ? node2192 : node2173;
									assign node2173 = (inp[5]) ? node2185 : node2174;
										assign node2174 = (inp[8]) ? node2180 : node2175;
											assign node2175 = (inp[2]) ? node2177 : 3'b010;
												assign node2177 = (inp[11]) ? 3'b100 : 3'b010;
											assign node2180 = (inp[2]) ? node2182 : 3'b110;
												assign node2182 = (inp[11]) ? 3'b010 : 3'b110;
										assign node2185 = (inp[11]) ? 3'b100 : node2186;
											assign node2186 = (inp[8]) ? 3'b010 : node2187;
												assign node2187 = (inp[2]) ? 3'b100 : 3'b000;
									assign node2192 = (inp[8]) ? node2200 : node2193;
										assign node2193 = (inp[5]) ? node2195 : 3'b100;
											assign node2195 = (inp[11]) ? 3'b000 : node2196;
												assign node2196 = (inp[2]) ? 3'b000 : 3'b100;
										assign node2200 = (inp[5]) ? 3'b100 : node2201;
											assign node2201 = (inp[11]) ? 3'b100 : 3'b010;
						assign node2205 = (inp[4]) ? node2293 : node2206;
							assign node2206 = (inp[1]) ? node2248 : node2207;
								assign node2207 = (inp[5]) ? node2229 : node2208;
									assign node2208 = (inp[8]) ? node2218 : node2209;
										assign node2209 = (inp[10]) ? 3'b101 : node2210;
											assign node2210 = (inp[11]) ? node2214 : node2211;
												assign node2211 = (inp[2]) ? 3'b011 : 3'b111;
												assign node2214 = (inp[2]) ? 3'b101 : 3'b001;
										assign node2218 = (inp[10]) ? node2224 : node2219;
											assign node2219 = (inp[2]) ? node2221 : 3'b111;
												assign node2221 = (inp[11]) ? 3'b011 : 3'b111;
											assign node2224 = (inp[2]) ? node2226 : 3'b011;
												assign node2226 = (inp[11]) ? 3'b101 : 3'b011;
									assign node2229 = (inp[11]) ? node2243 : node2230;
										assign node2230 = (inp[2]) ? node2236 : node2231;
											assign node2231 = (inp[10]) ? node2233 : 3'b101;
												assign node2233 = (inp[8]) ? 3'b101 : 3'b111;
											assign node2236 = (inp[10]) ? node2240 : node2237;
												assign node2237 = (inp[8]) ? 3'b011 : 3'b101;
												assign node2240 = (inp[8]) ? 3'b101 : 3'b011;
										assign node2243 = (inp[10]) ? node2245 : 3'b101;
											assign node2245 = (inp[8]) ? 3'b101 : 3'b001;
								assign node2248 = (inp[10]) ? node2272 : node2249;
									assign node2249 = (inp[8]) ? node2261 : node2250;
										assign node2250 = (inp[2]) ? node2256 : node2251;
											assign node2251 = (inp[5]) ? 3'b001 : node2252;
												assign node2252 = (inp[11]) ? 3'b011 : 3'b001;
											assign node2256 = (inp[11]) ? 3'b001 : node2257;
												assign node2257 = (inp[5]) ? 3'b001 : 3'b101;
										assign node2261 = (inp[5]) ? node2267 : node2262;
											assign node2262 = (inp[11]) ? node2264 : 3'b011;
												assign node2264 = (inp[2]) ? 3'b101 : 3'b111;
											assign node2267 = (inp[2]) ? node2269 : 3'b101;
												assign node2269 = (inp[11]) ? 3'b001 : 3'b101;
									assign node2272 = (inp[8]) ? node2282 : node2273;
										assign node2273 = (inp[5]) ? node2279 : node2274;
											assign node2274 = (inp[11]) ? node2276 : 3'b001;
												assign node2276 = (inp[2]) ? 3'b110 : 3'b100;
											assign node2279 = (inp[2]) ? 3'b110 : 3'b010;
										assign node2282 = (inp[2]) ? node2288 : node2283;
											assign node2283 = (inp[5]) ? 3'b001 : node2284;
												assign node2284 = (inp[11]) ? 3'b001 : 3'b101;
											assign node2288 = (inp[11]) ? 3'b110 : node2289;
												assign node2289 = (inp[5]) ? 3'b001 : 3'b101;
							assign node2293 = (inp[10]) ? node2333 : node2294;
								assign node2294 = (inp[11]) ? node2314 : node2295;
									assign node2295 = (inp[2]) ? node2307 : node2296;
										assign node2296 = (inp[1]) ? node2302 : node2297;
											assign node2297 = (inp[8]) ? node2299 : 3'b001;
												assign node2299 = (inp[5]) ? 3'b101 : 3'b011;
											assign node2302 = (inp[8]) ? node2304 : 3'b110;
												assign node2304 = (inp[5]) ? 3'b001 : 3'b101;
										assign node2307 = (inp[1]) ? 3'b001 : node2308;
											assign node2308 = (inp[5]) ? 3'b001 : node2309;
												assign node2309 = (inp[8]) ? 3'b101 : 3'b001;
									assign node2314 = (inp[5]) ? node2324 : node2315;
										assign node2315 = (inp[1]) ? node2319 : node2316;
											assign node2316 = (inp[2]) ? 3'b001 : 3'b101;
											assign node2319 = (inp[8]) ? node2321 : 3'b110;
												assign node2321 = (inp[2]) ? 3'b001 : 3'b000;
										assign node2324 = (inp[1]) ? node2328 : node2325;
											assign node2325 = (inp[8]) ? 3'b001 : 3'b110;
											assign node2328 = (inp[8]) ? node2330 : 3'b010;
												assign node2330 = (inp[2]) ? 3'b110 : 3'b010;
								assign node2333 = (inp[1]) ? node2353 : node2334;
									assign node2334 = (inp[8]) ? node2340 : node2335;
										assign node2335 = (inp[5]) ? node2337 : 3'b110;
											assign node2337 = (inp[11]) ? 3'b010 : 3'b110;
										assign node2340 = (inp[5]) ? node2348 : node2341;
											assign node2341 = (inp[2]) ? node2345 : node2342;
												assign node2342 = (inp[11]) ? 3'b001 : 3'b101;
												assign node2345 = (inp[11]) ? 3'b001 : 3'b011;
											assign node2348 = (inp[2]) ? 3'b110 : node2349;
												assign node2349 = (inp[11]) ? 3'b110 : 3'b001;
									assign node2353 = (inp[5]) ? node2363 : node2354;
										assign node2354 = (inp[8]) ? node2360 : node2355;
											assign node2355 = (inp[11]) ? node2357 : 3'b110;
												assign node2357 = (inp[2]) ? 3'b010 : 3'b110;
											assign node2360 = (inp[2]) ? 3'b110 : 3'b010;
										assign node2363 = (inp[8]) ? node2369 : node2364;
											assign node2364 = (inp[11]) ? node2366 : 3'b010;
												assign node2366 = (inp[2]) ? 3'b100 : 3'b000;
											assign node2369 = (inp[11]) ? 3'b010 : 3'b110;
			assign node2372 = (inp[9]) ? node2910 : node2373;
				assign node2373 = (inp[7]) ? node2643 : node2374;
					assign node2374 = (inp[4]) ? node2506 : node2375;
						assign node2375 = (inp[10]) ? node2439 : node2376;
							assign node2376 = (inp[5]) ? node2412 : node2377;
								assign node2377 = (inp[0]) ? node2393 : node2378;
									assign node2378 = (inp[2]) ? node2388 : node2379;
										assign node2379 = (inp[11]) ? node2383 : node2380;
											assign node2380 = (inp[1]) ? 3'b011 : 3'b111;
											assign node2383 = (inp[1]) ? 3'b101 : node2384;
												assign node2384 = (inp[8]) ? 3'b111 : 3'b101;
										assign node2388 = (inp[1]) ? node2390 : 3'b101;
											assign node2390 = (inp[8]) ? 3'b101 : 3'b001;
									assign node2393 = (inp[1]) ? node2403 : node2394;
										assign node2394 = (inp[8]) ? node2400 : node2395;
											assign node2395 = (inp[2]) ? node2397 : 3'b001;
												assign node2397 = (inp[11]) ? 3'b101 : 3'b001;
											assign node2400 = (inp[2]) ? 3'b001 : 3'b011;
										assign node2403 = (inp[2]) ? 3'b110 : node2404;
											assign node2404 = (inp[11]) ? node2408 : node2405;
												assign node2405 = (inp[8]) ? 3'b001 : 3'b111;
												assign node2408 = (inp[8]) ? 3'b110 : 3'b100;
								assign node2412 = (inp[1]) ? node2420 : node2413;
									assign node2413 = (inp[8]) ? node2417 : node2414;
										assign node2414 = (inp[0]) ? 3'b010 : 3'b110;
										assign node2417 = (inp[2]) ? 3'b110 : 3'b100;
									assign node2420 = (inp[0]) ? node2430 : node2421;
										assign node2421 = (inp[11]) ? node2427 : node2422;
											assign node2422 = (inp[8]) ? node2424 : 3'b001;
												assign node2424 = (inp[2]) ? 3'b001 : 3'b101;
											assign node2427 = (inp[8]) ? 3'b001 : 3'b110;
										assign node2430 = (inp[8]) ? node2436 : node2431;
											assign node2431 = (inp[2]) ? node2433 : 3'b010;
												assign node2433 = (inp[11]) ? 3'b100 : 3'b010;
											assign node2436 = (inp[11]) ? 3'b010 : 3'b110;
							assign node2439 = (inp[0]) ? node2471 : node2440;
								assign node2440 = (inp[1]) ? node2454 : node2441;
									assign node2441 = (inp[2]) ? node2449 : node2442;
										assign node2442 = (inp[5]) ? node2446 : node2443;
											assign node2443 = (inp[8]) ? 3'b100 : 3'b110;
											assign node2446 = (inp[8]) ? 3'b110 : 3'b100;
										assign node2449 = (inp[8]) ? 3'b110 : node2450;
											assign node2450 = (inp[5]) ? 3'b100 : 3'b110;
									assign node2454 = (inp[8]) ? node2462 : node2455;
										assign node2455 = (inp[5]) ? node2457 : 3'b110;
											assign node2457 = (inp[11]) ? node2459 : 3'b110;
												assign node2459 = (inp[2]) ? 3'b010 : 3'b110;
										assign node2462 = (inp[5]) ? node2468 : node2463;
											assign node2463 = (inp[11]) ? 3'b001 : node2464;
												assign node2464 = (inp[2]) ? 3'b001 : 3'b101;
											assign node2468 = (inp[2]) ? 3'b110 : 3'b001;
								assign node2471 = (inp[5]) ? node2489 : node2472;
									assign node2472 = (inp[8]) ? node2482 : node2473;
										assign node2473 = (inp[11]) ? node2477 : node2474;
											assign node2474 = (inp[1]) ? 3'b010 : 3'b110;
											assign node2477 = (inp[1]) ? node2479 : 3'b010;
												assign node2479 = (inp[2]) ? 3'b100 : 3'b010;
										assign node2482 = (inp[1]) ? node2486 : node2483;
											assign node2483 = (inp[2]) ? 3'b110 : 3'b100;
											assign node2486 = (inp[2]) ? 3'b010 : 3'b110;
									assign node2489 = (inp[8]) ? node2499 : node2490;
										assign node2490 = (inp[11]) ? node2492 : 3'b100;
											assign node2492 = (inp[1]) ? node2496 : node2493;
												assign node2493 = (inp[2]) ? 3'b100 : 3'b000;
												assign node2496 = (inp[2]) ? 3'b000 : 3'b100;
										assign node2499 = (inp[11]) ? node2503 : node2500;
											assign node2500 = (inp[1]) ? 3'b010 : 3'b110;
											assign node2503 = (inp[1]) ? 3'b100 : 3'b010;
						assign node2506 = (inp[0]) ? node2584 : node2507;
							assign node2507 = (inp[5]) ? node2551 : node2508;
								assign node2508 = (inp[8]) ? node2528 : node2509;
									assign node2509 = (inp[1]) ? node2521 : node2510;
										assign node2510 = (inp[2]) ? node2516 : node2511;
											assign node2511 = (inp[11]) ? node2513 : 3'b110;
												assign node2513 = (inp[10]) ? 3'b010 : 3'b110;
											assign node2516 = (inp[10]) ? 3'b110 : node2517;
												assign node2517 = (inp[11]) ? 3'b110 : 3'b000;
										assign node2521 = (inp[11]) ? node2523 : 3'b110;
											assign node2523 = (inp[10]) ? node2525 : 3'b000;
												assign node2525 = (inp[2]) ? 3'b100 : 3'b110;
									assign node2528 = (inp[10]) ? node2542 : node2529;
										assign node2529 = (inp[2]) ? node2537 : node2530;
											assign node2530 = (inp[11]) ? node2534 : node2531;
												assign node2531 = (inp[1]) ? 3'b000 : 3'b100;
												assign node2534 = (inp[1]) ? 3'b100 : 3'b000;
											assign node2537 = (inp[11]) ? node2539 : 3'b001;
												assign node2539 = (inp[1]) ? 3'b110 : 3'b000;
										assign node2542 = (inp[1]) ? node2548 : node2543;
											assign node2543 = (inp[11]) ? node2545 : 3'b000;
												assign node2545 = (inp[2]) ? 3'b110 : 3'b100;
											assign node2548 = (inp[11]) ? 3'b010 : 3'b110;
								assign node2551 = (inp[10]) ? node2563 : node2552;
									assign node2552 = (inp[1]) ? node2560 : node2553;
										assign node2553 = (inp[8]) ? node2555 : 3'b110;
											assign node2555 = (inp[11]) ? node2557 : 3'b000;
												assign node2557 = (inp[2]) ? 3'b110 : 3'b000;
										assign node2560 = (inp[8]) ? 3'b110 : 3'b010;
									assign node2563 = (inp[8]) ? node2573 : node2564;
										assign node2564 = (inp[1]) ? node2570 : node2565;
											assign node2565 = (inp[11]) ? 3'b010 : node2566;
												assign node2566 = (inp[2]) ? 3'b000 : 3'b100;
											assign node2570 = (inp[11]) ? 3'b100 : 3'b000;
										assign node2573 = (inp[1]) ? node2579 : node2574;
											assign node2574 = (inp[2]) ? node2576 : 3'b110;
												assign node2576 = (inp[11]) ? 3'b010 : 3'b110;
											assign node2579 = (inp[11]) ? node2581 : 3'b010;
												assign node2581 = (inp[2]) ? 3'b100 : 3'b010;
							assign node2584 = (inp[10]) ? node2616 : node2585;
								assign node2585 = (inp[1]) ? node2597 : node2586;
									assign node2586 = (inp[5]) ? node2594 : node2587;
										assign node2587 = (inp[8]) ? 3'b110 : node2588;
											assign node2588 = (inp[11]) ? 3'b010 : node2589;
												assign node2589 = (inp[2]) ? 3'b010 : 3'b110;
										assign node2594 = (inp[8]) ? 3'b010 : 3'b100;
									assign node2597 = (inp[11]) ? node2611 : node2598;
										assign node2598 = (inp[8]) ? node2606 : node2599;
											assign node2599 = (inp[5]) ? node2603 : node2600;
												assign node2600 = (inp[2]) ? 3'b100 : 3'b000;
												assign node2603 = (inp[2]) ? 3'b000 : 3'b100;
											assign node2606 = (inp[2]) ? node2608 : 3'b010;
												assign node2608 = (inp[5]) ? 3'b100 : 3'b010;
										assign node2611 = (inp[8]) ? 3'b100 : node2612;
											assign node2612 = (inp[5]) ? 3'b000 : 3'b100;
								assign node2616 = (inp[1]) ? node2636 : node2617;
									assign node2617 = (inp[11]) ? node2627 : node2618;
										assign node2618 = (inp[5]) ? node2622 : node2619;
											assign node2619 = (inp[8]) ? 3'b010 : 3'b100;
											assign node2622 = (inp[8]) ? 3'b100 : node2623;
												assign node2623 = (inp[2]) ? 3'b000 : 3'b100;
										assign node2627 = (inp[5]) ? node2633 : node2628;
											assign node2628 = (inp[8]) ? node2630 : 3'b100;
												assign node2630 = (inp[2]) ? 3'b100 : 3'b000;
											assign node2633 = (inp[8]) ? 3'b100 : 3'b000;
									assign node2636 = (inp[11]) ? 3'b000 : node2637;
										assign node2637 = (inp[5]) ? node2639 : 3'b100;
											assign node2639 = (inp[8]) ? 3'b100 : 3'b000;
					assign node2643 = (inp[0]) ? node2761 : node2644;
						assign node2644 = (inp[4]) ? node2694 : node2645;
							assign node2645 = (inp[1]) ? node2667 : node2646;
								assign node2646 = (inp[10]) ? node2654 : node2647;
									assign node2647 = (inp[5]) ? node2649 : 3'b111;
										assign node2649 = (inp[11]) ? node2651 : 3'b111;
											assign node2651 = (inp[2]) ? 3'b011 : 3'b111;
									assign node2654 = (inp[2]) ? node2660 : node2655;
										assign node2655 = (inp[11]) ? 3'b011 : node2656;
											assign node2656 = (inp[5]) ? 3'b011 : 3'b111;
										assign node2660 = (inp[11]) ? node2664 : node2661;
											assign node2661 = (inp[5]) ? 3'b011 : 3'b111;
											assign node2664 = (inp[5]) ? 3'b111 : 3'b011;
								assign node2667 = (inp[8]) ? node2683 : node2668;
									assign node2668 = (inp[10]) ? node2676 : node2669;
										assign node2669 = (inp[5]) ? 3'b101 : node2670;
											assign node2670 = (inp[11]) ? 3'b101 : node2671;
												assign node2671 = (inp[2]) ? 3'b011 : 3'b111;
										assign node2676 = (inp[11]) ? 3'b001 : node2677;
											assign node2677 = (inp[5]) ? node2679 : 3'b101;
												assign node2679 = (inp[2]) ? 3'b001 : 3'b101;
									assign node2683 = (inp[10]) ? node2689 : node2684;
										assign node2684 = (inp[5]) ? 3'b011 : node2685;
											assign node2685 = (inp[11]) ? 3'b011 : 3'b111;
										assign node2689 = (inp[11]) ? 3'b101 : node2690;
											assign node2690 = (inp[5]) ? 3'b101 : 3'b011;
							assign node2694 = (inp[8]) ? node2720 : node2695;
								assign node2695 = (inp[10]) ? node2711 : node2696;
									assign node2696 = (inp[11]) ? node2702 : node2697;
										assign node2697 = (inp[1]) ? 3'b001 : node2698;
											assign node2698 = (inp[5]) ? 3'b101 : 3'b011;
										assign node2702 = (inp[1]) ? node2706 : node2703;
											assign node2703 = (inp[5]) ? 3'b001 : 3'b100;
											assign node2706 = (inp[5]) ? 3'b110 : node2707;
												assign node2707 = (inp[2]) ? 3'b001 : 3'b101;
									assign node2711 = (inp[1]) ? 3'b110 : node2712;
										assign node2712 = (inp[11]) ? node2716 : node2713;
											assign node2713 = (inp[5]) ? 3'b001 : 3'b101;
											assign node2716 = (inp[5]) ? 3'b110 : 3'b001;
								assign node2720 = (inp[10]) ? node2740 : node2721;
									assign node2721 = (inp[5]) ? node2729 : node2722;
										assign node2722 = (inp[1]) ? node2724 : 3'b011;
											assign node2724 = (inp[2]) ? 3'b101 : node2725;
												assign node2725 = (inp[11]) ? 3'b101 : 3'b011;
										assign node2729 = (inp[1]) ? node2735 : node2730;
											assign node2730 = (inp[11]) ? 3'b101 : node2731;
												assign node2731 = (inp[2]) ? 3'b101 : 3'b011;
											assign node2735 = (inp[11]) ? 3'b001 : node2736;
												assign node2736 = (inp[2]) ? 3'b001 : 3'b101;
									assign node2740 = (inp[1]) ? node2752 : node2741;
										assign node2741 = (inp[11]) ? node2747 : node2742;
											assign node2742 = (inp[2]) ? node2744 : 3'b101;
												assign node2744 = (inp[5]) ? 3'b001 : 3'b101;
											assign node2747 = (inp[2]) ? 3'b001 : node2748;
												assign node2748 = (inp[5]) ? 3'b001 : 3'b101;
										assign node2752 = (inp[5]) ? node2756 : node2753;
											assign node2753 = (inp[2]) ? 3'b001 : 3'b101;
											assign node2756 = (inp[11]) ? 3'b110 : node2757;
												assign node2757 = (inp[2]) ? 3'b110 : 3'b001;
						assign node2761 = (inp[4]) ? node2829 : node2762;
							assign node2762 = (inp[10]) ? node2792 : node2763;
								assign node2763 = (inp[11]) ? node2779 : node2764;
									assign node2764 = (inp[8]) ? node2772 : node2765;
										assign node2765 = (inp[5]) ? node2769 : node2766;
											assign node2766 = (inp[1]) ? 3'b001 : 3'b101;
											assign node2769 = (inp[1]) ? 3'b110 : 3'b001;
										assign node2772 = (inp[1]) ? node2776 : node2773;
											assign node2773 = (inp[5]) ? 3'b101 : 3'b011;
											assign node2776 = (inp[5]) ? 3'b001 : 3'b101;
									assign node2779 = (inp[8]) ? node2781 : 3'b001;
										assign node2781 = (inp[5]) ? node2787 : node2782;
											assign node2782 = (inp[1]) ? 3'b101 : node2783;
												assign node2783 = (inp[2]) ? 3'b101 : 3'b011;
											assign node2787 = (inp[1]) ? 3'b001 : node2788;
												assign node2788 = (inp[2]) ? 3'b001 : 3'b101;
								assign node2792 = (inp[1]) ? node2816 : node2793;
									assign node2793 = (inp[8]) ? node2805 : node2794;
										assign node2794 = (inp[5]) ? node2800 : node2795;
											assign node2795 = (inp[11]) ? node2797 : 3'b001;
												assign node2797 = (inp[2]) ? 3'b110 : 3'b000;
											assign node2800 = (inp[2]) ? 3'b110 : node2801;
												assign node2801 = (inp[11]) ? 3'b110 : 3'b010;
										assign node2805 = (inp[5]) ? node2811 : node2806;
											assign node2806 = (inp[11]) ? node2808 : 3'b101;
												assign node2808 = (inp[2]) ? 3'b001 : 3'b101;
											assign node2811 = (inp[11]) ? node2813 : 3'b001;
												assign node2813 = (inp[2]) ? 3'b110 : 3'b001;
									assign node2816 = (inp[5]) ? node2822 : node2817;
										assign node2817 = (inp[8]) ? node2819 : 3'b110;
											assign node2819 = (inp[2]) ? 3'b110 : 3'b010;
										assign node2822 = (inp[8]) ? 3'b110 : node2823;
											assign node2823 = (inp[11]) ? 3'b010 : node2824;
												assign node2824 = (inp[2]) ? 3'b010 : 3'b110;
							assign node2829 = (inp[10]) ? node2869 : node2830;
								assign node2830 = (inp[5]) ? node2852 : node2831;
									assign node2831 = (inp[8]) ? node2843 : node2832;
										assign node2832 = (inp[2]) ? node2838 : node2833;
											assign node2833 = (inp[11]) ? 3'b100 : node2834;
												assign node2834 = (inp[1]) ? 3'b111 : 3'b110;
											assign node2838 = (inp[11]) ? node2840 : 3'b110;
												assign node2840 = (inp[1]) ? 3'b010 : 3'b110;
										assign node2843 = (inp[1]) ? node2847 : node2844;
											assign node2844 = (inp[2]) ? 3'b001 : 3'b101;
											assign node2847 = (inp[2]) ? 3'b110 : node2848;
												assign node2848 = (inp[11]) ? 3'b110 : 3'b001;
									assign node2852 = (inp[8]) ? node2858 : node2853;
										assign node2853 = (inp[11]) ? 3'b010 : node2854;
											assign node2854 = (inp[1]) ? 3'b010 : 3'b110;
										assign node2858 = (inp[1]) ? node2864 : node2859;
											assign node2859 = (inp[2]) ? 3'b110 : node2860;
												assign node2860 = (inp[11]) ? 3'b110 : 3'b001;
											assign node2864 = (inp[2]) ? node2866 : 3'b110;
												assign node2866 = (inp[11]) ? 3'b010 : 3'b110;
								assign node2869 = (inp[11]) ? node2887 : node2870;
									assign node2870 = (inp[1]) ? node2878 : node2871;
										assign node2871 = (inp[8]) ? node2873 : 3'b010;
											assign node2873 = (inp[5]) ? node2875 : 3'b001;
												assign node2875 = (inp[2]) ? 3'b010 : 3'b110;
										assign node2878 = (inp[8]) ? node2882 : node2879;
											assign node2879 = (inp[5]) ? 3'b100 : 3'b010;
											assign node2882 = (inp[2]) ? 3'b010 : node2883;
												assign node2883 = (inp[5]) ? 3'b010 : 3'b110;
									assign node2887 = (inp[8]) ? node2903 : node2888;
										assign node2888 = (inp[5]) ? node2896 : node2889;
											assign node2889 = (inp[2]) ? node2893 : node2890;
												assign node2890 = (inp[1]) ? 3'b010 : 3'b000;
												assign node2893 = (inp[1]) ? 3'b100 : 3'b000;
											assign node2896 = (inp[2]) ? node2900 : node2897;
												assign node2897 = (inp[1]) ? 3'b100 : 3'b000;
												assign node2900 = (inp[1]) ? 3'b000 : 3'b100;
										assign node2903 = (inp[1]) ? node2907 : node2904;
											assign node2904 = (inp[5]) ? 3'b010 : 3'b110;
											assign node2907 = (inp[5]) ? 3'b100 : 3'b010;
				assign node2910 = (inp[0]) ? node3180 : node2911;
					assign node2911 = (inp[4]) ? node3059 : node2912;
						assign node2912 = (inp[7]) ? node2988 : node2913;
							assign node2913 = (inp[1]) ? node2949 : node2914;
								assign node2914 = (inp[10]) ? node2934 : node2915;
									assign node2915 = (inp[5]) ? node2925 : node2916;
										assign node2916 = (inp[11]) ? node2922 : node2917;
											assign node2917 = (inp[8]) ? node2919 : 3'b001;
												assign node2919 = (inp[2]) ? 3'b000 : 3'b100;
											assign node2922 = (inp[8]) ? 3'b001 : 3'b111;
										assign node2925 = (inp[11]) ? node2931 : node2926;
											assign node2926 = (inp[8]) ? node2928 : 3'b110;
												assign node2928 = (inp[2]) ? 3'b111 : 3'b001;
											assign node2931 = (inp[8]) ? 3'b110 : 3'b010;
									assign node2934 = (inp[5]) ? node2944 : node2935;
										assign node2935 = (inp[11]) ? node2941 : node2936;
											assign node2936 = (inp[8]) ? node2938 : 3'b110;
												assign node2938 = (inp[2]) ? 3'b111 : 3'b011;
											assign node2941 = (inp[8]) ? 3'b110 : 3'b010;
										assign node2944 = (inp[11]) ? 3'b010 : node2945;
											assign node2945 = (inp[8]) ? 3'b110 : 3'b010;
								assign node2949 = (inp[11]) ? node2969 : node2950;
									assign node2950 = (inp[10]) ? node2960 : node2951;
										assign node2951 = (inp[5]) ? node2957 : node2952;
											assign node2952 = (inp[2]) ? 3'b100 : node2953;
												assign node2953 = (inp[8]) ? 3'b111 : 3'b101;
											assign node2957 = (inp[8]) ? 3'b000 : 3'b010;
										assign node2960 = (inp[5]) ? node2966 : node2961;
											assign node2961 = (inp[2]) ? 3'b010 : node2962;
												assign node2962 = (inp[8]) ? 3'b000 : 3'b010;
											assign node2966 = (inp[8]) ? 3'b110 : 3'b100;
									assign node2969 = (inp[10]) ? node2979 : node2970;
										assign node2970 = (inp[5]) ? node2976 : node2971;
											assign node2971 = (inp[8]) ? 3'b100 : node2972;
												assign node2972 = (inp[2]) ? 3'b010 : 3'b110;
											assign node2976 = (inp[8]) ? 3'b010 : 3'b100;
										assign node2979 = (inp[5]) ? node2983 : node2980;
											assign node2980 = (inp[8]) ? 3'b010 : 3'b100;
											assign node2983 = (inp[8]) ? 3'b100 : node2984;
												assign node2984 = (inp[2]) ? 3'b000 : 3'b100;
							assign node2988 = (inp[10]) ? node3018 : node2989;
								assign node2989 = (inp[1]) ? node3001 : node2990;
									assign node2990 = (inp[11]) ? 3'b101 : node2991;
										assign node2991 = (inp[8]) ? node2993 : 3'b001;
											assign node2993 = (inp[2]) ? node2997 : node2994;
												assign node2994 = (inp[5]) ? 3'b101 : 3'b011;
												assign node2997 = (inp[5]) ? 3'b001 : 3'b101;
									assign node3001 = (inp[8]) ? node3009 : node3002;
										assign node3002 = (inp[5]) ? 3'b110 : node3003;
											assign node3003 = (inp[11]) ? 3'b110 : node3004;
												assign node3004 = (inp[2]) ? 3'b001 : 3'b101;
										assign node3009 = (inp[5]) ? node3013 : node3010;
											assign node3010 = (inp[11]) ? 3'b001 : 3'b101;
											assign node3013 = (inp[2]) ? node3015 : 3'b001;
												assign node3015 = (inp[11]) ? 3'b110 : 3'b001;
								assign node3018 = (inp[11]) ? node3040 : node3019;
									assign node3019 = (inp[8]) ? node3027 : node3020;
										assign node3020 = (inp[5]) ? node3022 : 3'b110;
											assign node3022 = (inp[1]) ? node3024 : 3'b110;
												assign node3024 = (inp[2]) ? 3'b001 : 3'b101;
										assign node3027 = (inp[5]) ? node3035 : node3028;
											assign node3028 = (inp[2]) ? node3032 : node3029;
												assign node3029 = (inp[1]) ? 3'b001 : 3'b101;
												assign node3032 = (inp[1]) ? 3'b001 : 3'b011;
											assign node3035 = (inp[2]) ? 3'b110 : node3036;
												assign node3036 = (inp[1]) ? 3'b110 : 3'b001;
									assign node3040 = (inp[1]) ? node3048 : node3041;
										assign node3041 = (inp[8]) ? node3043 : 3'b000;
											assign node3043 = (inp[5]) ? node3045 : 3'b001;
												assign node3045 = (inp[2]) ? 3'b000 : 3'b001;
										assign node3048 = (inp[8]) ? node3054 : node3049;
											assign node3049 = (inp[2]) ? 3'b010 : node3050;
												assign node3050 = (inp[5]) ? 3'b010 : 3'b110;
											assign node3054 = (inp[5]) ? 3'b110 : node3055;
												assign node3055 = (inp[2]) ? 3'b110 : 3'b001;
						assign node3059 = (inp[1]) ? node3117 : node3060;
							assign node3060 = (inp[7]) ? node3096 : node3061;
								assign node3061 = (inp[10]) ? node3081 : node3062;
									assign node3062 = (inp[2]) ? node3076 : node3063;
										assign node3063 = (inp[11]) ? node3069 : node3064;
											assign node3064 = (inp[5]) ? node3066 : 3'b110;
												assign node3066 = (inp[8]) ? 3'b010 : 3'b110;
											assign node3069 = (inp[8]) ? node3073 : node3070;
												assign node3070 = (inp[5]) ? 3'b110 : 3'b010;
												assign node3073 = (inp[5]) ? 3'b010 : 3'b110;
										assign node3076 = (inp[5]) ? node3078 : 3'b010;
											assign node3078 = (inp[8]) ? 3'b010 : 3'b110;
									assign node3081 = (inp[5]) ? node3089 : node3082;
										assign node3082 = (inp[8]) ? node3084 : 3'b110;
											assign node3084 = (inp[2]) ? node3086 : 3'b010;
												assign node3086 = (inp[11]) ? 3'b110 : 3'b010;
										assign node3089 = (inp[8]) ? 3'b100 : node3090;
											assign node3090 = (inp[11]) ? 3'b000 : node3091;
												assign node3091 = (inp[2]) ? 3'b000 : 3'b100;
								assign node3096 = (inp[10]) ? node3110 : node3097;
									assign node3097 = (inp[5]) ? node3103 : node3098;
										assign node3098 = (inp[8]) ? 3'b001 : node3099;
											assign node3099 = (inp[11]) ? 3'b110 : 3'b001;
										assign node3103 = (inp[8]) ? node3107 : node3104;
											assign node3104 = (inp[11]) ? 3'b010 : 3'b110;
											assign node3107 = (inp[11]) ? 3'b110 : 3'b001;
									assign node3110 = (inp[5]) ? 3'b010 : node3111;
										assign node3111 = (inp[11]) ? node3113 : 3'b110;
											assign node3113 = (inp[8]) ? 3'b110 : 3'b010;
							assign node3117 = (inp[7]) ? node3147 : node3118;
								assign node3118 = (inp[8]) ? node3126 : node3119;
									assign node3119 = (inp[5]) ? 3'b000 : node3120;
										assign node3120 = (inp[10]) ? 3'b000 : node3121;
											assign node3121 = (inp[11]) ? 3'b000 : 3'b100;
									assign node3126 = (inp[11]) ? node3134 : node3127;
										assign node3127 = (inp[10]) ? node3131 : node3128;
											assign node3128 = (inp[5]) ? 3'b100 : 3'b000;
											assign node3131 = (inp[5]) ? 3'b000 : 3'b100;
										assign node3134 = (inp[2]) ? node3142 : node3135;
											assign node3135 = (inp[10]) ? node3139 : node3136;
												assign node3136 = (inp[5]) ? 3'b100 : 3'b000;
												assign node3139 = (inp[5]) ? 3'b000 : 3'b100;
											assign node3142 = (inp[10]) ? 3'b000 : node3143;
												assign node3143 = (inp[5]) ? 3'b000 : 3'b100;
								assign node3147 = (inp[10]) ? node3163 : node3148;
									assign node3148 = (inp[2]) ? node3158 : node3149;
										assign node3149 = (inp[5]) ? node3151 : 3'b110;
											assign node3151 = (inp[11]) ? node3155 : node3152;
												assign node3152 = (inp[8]) ? 3'b110 : 3'b010;
												assign node3155 = (inp[8]) ? 3'b010 : 3'b100;
										assign node3158 = (inp[8]) ? node3160 : 3'b010;
											assign node3160 = (inp[5]) ? 3'b010 : 3'b110;
									assign node3163 = (inp[8]) ? node3171 : node3164;
										assign node3164 = (inp[11]) ? node3166 : 3'b100;
											assign node3166 = (inp[2]) ? node3168 : 3'b100;
												assign node3168 = (inp[5]) ? 3'b000 : 3'b100;
										assign node3171 = (inp[2]) ? node3177 : node3172;
											assign node3172 = (inp[5]) ? 3'b010 : node3173;
												assign node3173 = (inp[11]) ? 3'b010 : 3'b110;
											assign node3177 = (inp[5]) ? 3'b100 : 3'b010;
					assign node3180 = (inp[7]) ? node3234 : node3181;
						assign node3181 = (inp[4]) ? 3'b000 : node3182;
							assign node3182 = (inp[1]) ? node3218 : node3183;
								assign node3183 = (inp[5]) ? node3203 : node3184;
									assign node3184 = (inp[11]) ? node3196 : node3185;
										assign node3185 = (inp[10]) ? node3191 : node3186;
											assign node3186 = (inp[2]) ? 3'b010 : node3187;
												assign node3187 = (inp[8]) ? 3'b110 : 3'b010;
											assign node3191 = (inp[8]) ? 3'b010 : node3192;
												assign node3192 = (inp[2]) ? 3'b100 : 3'b110;
										assign node3196 = (inp[10]) ? node3200 : node3197;
											assign node3197 = (inp[8]) ? 3'b010 : 3'b100;
											assign node3200 = (inp[8]) ? 3'b100 : 3'b000;
									assign node3203 = (inp[8]) ? node3209 : node3204;
										assign node3204 = (inp[11]) ? 3'b000 : node3205;
											assign node3205 = (inp[2]) ? 3'b100 : 3'b000;
										assign node3209 = (inp[11]) ? node3215 : node3210;
											assign node3210 = (inp[10]) ? 3'b100 : node3211;
												assign node3211 = (inp[2]) ? 3'b100 : 3'b010;
											assign node3215 = (inp[10]) ? 3'b000 : 3'b100;
								assign node3218 = (inp[10]) ? 3'b000 : node3219;
									assign node3219 = (inp[11]) ? node3225 : node3220;
										assign node3220 = (inp[8]) ? 3'b100 : node3221;
											assign node3221 = (inp[5]) ? 3'b000 : 3'b100;
										assign node3225 = (inp[2]) ? node3227 : 3'b000;
											assign node3227 = (inp[8]) ? node3229 : 3'b000;
												assign node3229 = (inp[5]) ? 3'b000 : 3'b100;
						assign node3234 = (inp[4]) ? node3302 : node3235;
							assign node3235 = (inp[10]) ? node3265 : node3236;
								assign node3236 = (inp[1]) ? node3256 : node3237;
									assign node3237 = (inp[5]) ? node3251 : node3238;
										assign node3238 = (inp[2]) ? node3244 : node3239;
											assign node3239 = (inp[8]) ? 3'b001 : node3240;
												assign node3240 = (inp[11]) ? 3'b101 : 3'b010;
											assign node3244 = (inp[11]) ? node3248 : node3245;
												assign node3245 = (inp[8]) ? 3'b001 : 3'b110;
												assign node3248 = (inp[8]) ? 3'b110 : 3'b010;
										assign node3251 = (inp[8]) ? node3253 : 3'b010;
											assign node3253 = (inp[2]) ? 3'b010 : 3'b110;
									assign node3256 = (inp[8]) ? node3262 : node3257;
										assign node3257 = (inp[5]) ? 3'b100 : node3258;
											assign node3258 = (inp[11]) ? 3'b010 : 3'b110;
										assign node3262 = (inp[5]) ? 3'b010 : 3'b110;
								assign node3265 = (inp[1]) ? node3281 : node3266;
									assign node3266 = (inp[8]) ? node3274 : node3267;
										assign node3267 = (inp[2]) ? 3'b100 : node3268;
											assign node3268 = (inp[5]) ? node3270 : 3'b010;
												assign node3270 = (inp[11]) ? 3'b100 : 3'b000;
										assign node3274 = (inp[5]) ? 3'b010 : node3275;
											assign node3275 = (inp[11]) ? node3277 : 3'b110;
												assign node3277 = (inp[2]) ? 3'b010 : 3'b110;
									assign node3281 = (inp[11]) ? node3289 : node3282;
										assign node3282 = (inp[5]) ? node3286 : node3283;
											assign node3283 = (inp[8]) ? 3'b010 : 3'b100;
											assign node3286 = (inp[8]) ? 3'b100 : 3'b000;
										assign node3289 = (inp[2]) ? node3297 : node3290;
											assign node3290 = (inp[8]) ? node3294 : node3291;
												assign node3291 = (inp[5]) ? 3'b000 : 3'b100;
												assign node3294 = (inp[5]) ? 3'b100 : 3'b000;
											assign node3297 = (inp[8]) ? 3'b100 : node3298;
												assign node3298 = (inp[5]) ? 3'b000 : 3'b100;
							assign node3302 = (inp[1]) ? node3340 : node3303;
								assign node3303 = (inp[5]) ? node3323 : node3304;
									assign node3304 = (inp[10]) ? node3314 : node3305;
										assign node3305 = (inp[8]) ? node3309 : node3306;
											assign node3306 = (inp[11]) ? 3'b100 : 3'b010;
											assign node3309 = (inp[2]) ? 3'b010 : node3310;
												assign node3310 = (inp[11]) ? 3'b010 : 3'b110;
										assign node3314 = (inp[2]) ? 3'b100 : node3315;
											assign node3315 = (inp[11]) ? node3319 : node3316;
												assign node3316 = (inp[8]) ? 3'b010 : 3'b110;
												assign node3319 = (inp[8]) ? 3'b100 : 3'b000;
									assign node3323 = (inp[10]) ? node3335 : node3324;
										assign node3324 = (inp[2]) ? node3330 : node3325;
											assign node3325 = (inp[11]) ? node3327 : 3'b010;
												assign node3327 = (inp[8]) ? 3'b100 : 3'b000;
											assign node3330 = (inp[11]) ? node3332 : 3'b100;
												assign node3332 = (inp[8]) ? 3'b100 : 3'b000;
										assign node3335 = (inp[11]) ? 3'b000 : node3336;
											assign node3336 = (inp[8]) ? 3'b100 : 3'b000;
								assign node3340 = (inp[10]) ? 3'b000 : node3341;
									assign node3341 = (inp[11]) ? node3347 : node3342;
										assign node3342 = (inp[5]) ? node3344 : 3'b100;
											assign node3344 = (inp[8]) ? 3'b100 : 3'b000;
										assign node3347 = (inp[2]) ? node3349 : 3'b000;
											assign node3349 = (inp[8]) ? node3351 : 3'b000;
												assign node3351 = (inp[5]) ? 3'b000 : 3'b100;

endmodule