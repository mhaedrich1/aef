module dtc_split875_bm57 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node287;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node302;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node331;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node341;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node368;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node399;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node420;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node427;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node457;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node463;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node474;
	wire [3-1:0] node476;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node496;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node505;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node512;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node519;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node537;
	wire [3-1:0] node539;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node548;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node560;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node572;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node586;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node594;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node601;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node620;
	wire [3-1:0] node622;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node646;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node662;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node682;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node691;
	wire [3-1:0] node694;
	wire [3-1:0] node695;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node711;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node720;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node725;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node732;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node743;
	wire [3-1:0] node746;
	wire [3-1:0] node748;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node758;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node765;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node773;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node780;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node786;
	wire [3-1:0] node789;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node804;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node811;
	wire [3-1:0] node814;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node828;
	wire [3-1:0] node831;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node838;
	wire [3-1:0] node841;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node847;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node863;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node868;
	wire [3-1:0] node871;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node879;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node886;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node900;
	wire [3-1:0] node903;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node916;
	wire [3-1:0] node918;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node926;
	wire [3-1:0] node929;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node937;
	wire [3-1:0] node938;
	wire [3-1:0] node942;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node947;
	wire [3-1:0] node950;
	wire [3-1:0] node951;
	wire [3-1:0] node954;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node969;
	wire [3-1:0] node970;
	wire [3-1:0] node971;
	wire [3-1:0] node974;
	wire [3-1:0] node977;
	wire [3-1:0] node978;
	wire [3-1:0] node981;
	wire [3-1:0] node984;
	wire [3-1:0] node985;
	wire [3-1:0] node987;
	wire [3-1:0] node989;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node994;
	wire [3-1:0] node997;
	wire [3-1:0] node1000;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1008;
	wire [3-1:0] node1011;
	wire [3-1:0] node1012;
	wire [3-1:0] node1015;
	wire [3-1:0] node1018;
	wire [3-1:0] node1019;
	wire [3-1:0] node1021;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1031;
	wire [3-1:0] node1032;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1046;
	wire [3-1:0] node1047;
	wire [3-1:0] node1048;
	wire [3-1:0] node1049;
	wire [3-1:0] node1050;
	wire [3-1:0] node1053;
	wire [3-1:0] node1055;
	wire [3-1:0] node1058;
	wire [3-1:0] node1059;
	wire [3-1:0] node1061;
	wire [3-1:0] node1064;
	wire [3-1:0] node1065;
	wire [3-1:0] node1069;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1074;
	wire [3-1:0] node1076;
	wire [3-1:0] node1079;
	wire [3-1:0] node1080;
	wire [3-1:0] node1081;
	wire [3-1:0] node1084;
	wire [3-1:0] node1087;
	wire [3-1:0] node1088;
	wire [3-1:0] node1092;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1095;
	wire [3-1:0] node1098;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1106;
	wire [3-1:0] node1108;
	wire [3-1:0] node1109;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1115;
	wire [3-1:0] node1116;
	wire [3-1:0] node1117;
	wire [3-1:0] node1118;
	wire [3-1:0] node1122;
	wire [3-1:0] node1123;
	wire [3-1:0] node1126;
	wire [3-1:0] node1129;
	wire [3-1:0] node1131;
	wire [3-1:0] node1132;
	wire [3-1:0] node1136;
	wire [3-1:0] node1137;
	wire [3-1:0] node1138;
	wire [3-1:0] node1141;
	wire [3-1:0] node1142;
	wire [3-1:0] node1145;
	wire [3-1:0] node1148;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1154;
	wire [3-1:0] node1155;
	wire [3-1:0] node1158;
	wire [3-1:0] node1161;
	wire [3-1:0] node1162;
	wire [3-1:0] node1163;
	wire [3-1:0] node1164;
	wire [3-1:0] node1167;
	wire [3-1:0] node1170;
	wire [3-1:0] node1171;
	wire [3-1:0] node1174;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1183;
	wire [3-1:0] node1186;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1191;
	wire [3-1:0] node1192;
	wire [3-1:0] node1195;
	wire [3-1:0] node1198;
	wire [3-1:0] node1199;
	wire [3-1:0] node1202;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1208;
	wire [3-1:0] node1211;
	wire [3-1:0] node1212;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1220;
	wire [3-1:0] node1223;
	wire [3-1:0] node1225;
	wire [3-1:0] node1228;
	wire [3-1:0] node1229;
	wire [3-1:0] node1230;
	wire [3-1:0] node1233;
	wire [3-1:0] node1236;
	wire [3-1:0] node1239;
	wire [3-1:0] node1240;
	wire [3-1:0] node1241;
	wire [3-1:0] node1242;
	wire [3-1:0] node1245;
	wire [3-1:0] node1248;
	wire [3-1:0] node1249;
	wire [3-1:0] node1252;
	wire [3-1:0] node1255;
	wire [3-1:0] node1256;
	wire [3-1:0] node1257;
	wire [3-1:0] node1260;
	wire [3-1:0] node1263;
	wire [3-1:0] node1264;
	wire [3-1:0] node1267;
	wire [3-1:0] node1270;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1274;
	wire [3-1:0] node1275;
	wire [3-1:0] node1278;
	wire [3-1:0] node1281;
	wire [3-1:0] node1282;
	wire [3-1:0] node1286;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1291;
	wire [3-1:0] node1294;
	wire [3-1:0] node1297;
	wire [3-1:0] node1298;
	wire [3-1:0] node1299;
	wire [3-1:0] node1302;
	wire [3-1:0] node1303;
	wire [3-1:0] node1306;
	wire [3-1:0] node1309;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1314;
	wire [3-1:0] node1317;
	wire [3-1:0] node1318;
	wire [3-1:0] node1322;
	wire [3-1:0] node1323;
	wire [3-1:0] node1324;
	wire [3-1:0] node1325;
	wire [3-1:0] node1328;
	wire [3-1:0] node1331;
	wire [3-1:0] node1332;
	wire [3-1:0] node1336;
	wire [3-1:0] node1339;
	wire [3-1:0] node1340;
	wire [3-1:0] node1341;
	wire [3-1:0] node1342;
	wire [3-1:0] node1343;
	wire [3-1:0] node1344;
	wire [3-1:0] node1345;
	wire [3-1:0] node1348;
	wire [3-1:0] node1349;
	wire [3-1:0] node1351;
	wire [3-1:0] node1354;
	wire [3-1:0] node1355;
	wire [3-1:0] node1359;
	wire [3-1:0] node1360;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1365;
	wire [3-1:0] node1368;
	wire [3-1:0] node1369;
	wire [3-1:0] node1370;
	wire [3-1:0] node1373;
	wire [3-1:0] node1376;
	wire [3-1:0] node1377;
	wire [3-1:0] node1380;
	wire [3-1:0] node1383;
	wire [3-1:0] node1384;
	wire [3-1:0] node1385;
	wire [3-1:0] node1390;
	wire [3-1:0] node1391;
	wire [3-1:0] node1392;
	wire [3-1:0] node1395;
	wire [3-1:0] node1396;
	wire [3-1:0] node1398;
	wire [3-1:0] node1401;
	wire [3-1:0] node1402;
	wire [3-1:0] node1406;
	wire [3-1:0] node1407;
	wire [3-1:0] node1408;
	wire [3-1:0] node1409;
	wire [3-1:0] node1412;
	wire [3-1:0] node1415;
	wire [3-1:0] node1416;
	wire [3-1:0] node1419;
	wire [3-1:0] node1422;
	wire [3-1:0] node1423;
	wire [3-1:0] node1424;
	wire [3-1:0] node1428;
	wire [3-1:0] node1429;
	wire [3-1:0] node1433;
	wire [3-1:0] node1434;
	wire [3-1:0] node1435;
	wire [3-1:0] node1436;
	wire [3-1:0] node1439;
	wire [3-1:0] node1440;
	wire [3-1:0] node1442;
	wire [3-1:0] node1445;
	wire [3-1:0] node1446;
	wire [3-1:0] node1450;
	wire [3-1:0] node1451;
	wire [3-1:0] node1452;
	wire [3-1:0] node1453;
	wire [3-1:0] node1456;
	wire [3-1:0] node1459;
	wire [3-1:0] node1460;
	wire [3-1:0] node1461;
	wire [3-1:0] node1464;
	wire [3-1:0] node1467;
	wire [3-1:0] node1468;
	wire [3-1:0] node1471;
	wire [3-1:0] node1474;
	wire [3-1:0] node1475;
	wire [3-1:0] node1477;
	wire [3-1:0] node1480;
	wire [3-1:0] node1481;
	wire [3-1:0] node1485;
	wire [3-1:0] node1486;
	wire [3-1:0] node1487;
	wire [3-1:0] node1490;
	wire [3-1:0] node1491;
	wire [3-1:0] node1494;
	wire [3-1:0] node1495;
	wire [3-1:0] node1499;
	wire [3-1:0] node1500;
	wire [3-1:0] node1501;
	wire [3-1:0] node1502;
	wire [3-1:0] node1503;
	wire [3-1:0] node1506;
	wire [3-1:0] node1509;
	wire [3-1:0] node1510;
	wire [3-1:0] node1513;
	wire [3-1:0] node1516;
	wire [3-1:0] node1517;
	wire [3-1:0] node1518;
	wire [3-1:0] node1522;
	wire [3-1:0] node1523;
	wire [3-1:0] node1526;
	wire [3-1:0] node1529;
	wire [3-1:0] node1530;
	wire [3-1:0] node1531;
	wire [3-1:0] node1535;
	wire [3-1:0] node1537;
	wire [3-1:0] node1540;
	wire [3-1:0] node1541;
	wire [3-1:0] node1542;
	wire [3-1:0] node1543;
	wire [3-1:0] node1544;
	wire [3-1:0] node1545;
	wire [3-1:0] node1546;
	wire [3-1:0] node1549;
	wire [3-1:0] node1552;
	wire [3-1:0] node1553;
	wire [3-1:0] node1554;
	wire [3-1:0] node1557;
	wire [3-1:0] node1560;
	wire [3-1:0] node1561;
	wire [3-1:0] node1564;
	wire [3-1:0] node1567;
	wire [3-1:0] node1568;
	wire [3-1:0] node1571;
	wire [3-1:0] node1574;
	wire [3-1:0] node1575;
	wire [3-1:0] node1576;
	wire [3-1:0] node1579;
	wire [3-1:0] node1582;
	wire [3-1:0] node1583;
	wire [3-1:0] node1586;
	wire [3-1:0] node1589;
	wire [3-1:0] node1590;
	wire [3-1:0] node1591;
	wire [3-1:0] node1594;
	wire [3-1:0] node1597;
	wire [3-1:0] node1598;
	wire [3-1:0] node1599;
	wire [3-1:0] node1600;
	wire [3-1:0] node1601;
	wire [3-1:0] node1604;
	wire [3-1:0] node1607;
	wire [3-1:0] node1608;
	wire [3-1:0] node1611;
	wire [3-1:0] node1614;
	wire [3-1:0] node1615;
	wire [3-1:0] node1618;
	wire [3-1:0] node1621;
	wire [3-1:0] node1622;
	wire [3-1:0] node1623;
	wire [3-1:0] node1624;
	wire [3-1:0] node1627;
	wire [3-1:0] node1630;
	wire [3-1:0] node1631;
	wire [3-1:0] node1635;
	wire [3-1:0] node1636;
	wire [3-1:0] node1637;
	wire [3-1:0] node1640;
	wire [3-1:0] node1643;
	wire [3-1:0] node1644;
	wire [3-1:0] node1647;
	wire [3-1:0] node1650;
	wire [3-1:0] node1651;
	wire [3-1:0] node1652;
	wire [3-1:0] node1653;
	wire [3-1:0] node1654;
	wire [3-1:0] node1655;
	wire [3-1:0] node1658;
	wire [3-1:0] node1661;
	wire [3-1:0] node1662;
	wire [3-1:0] node1665;
	wire [3-1:0] node1668;
	wire [3-1:0] node1669;
	wire [3-1:0] node1670;
	wire [3-1:0] node1673;
	wire [3-1:0] node1676;
	wire [3-1:0] node1677;
	wire [3-1:0] node1680;
	wire [3-1:0] node1683;
	wire [3-1:0] node1684;
	wire [3-1:0] node1685;
	wire [3-1:0] node1688;
	wire [3-1:0] node1691;
	wire [3-1:0] node1692;
	wire [3-1:0] node1695;
	wire [3-1:0] node1698;
	wire [3-1:0] node1699;
	wire [3-1:0] node1702;
	wire [3-1:0] node1705;
	wire [3-1:0] node1706;
	wire [3-1:0] node1707;
	wire [3-1:0] node1708;
	wire [3-1:0] node1709;
	wire [3-1:0] node1710;
	wire [3-1:0] node1712;
	wire [3-1:0] node1715;
	wire [3-1:0] node1717;
	wire [3-1:0] node1720;
	wire [3-1:0] node1721;
	wire [3-1:0] node1723;
	wire [3-1:0] node1726;
	wire [3-1:0] node1728;
	wire [3-1:0] node1731;
	wire [3-1:0] node1732;
	wire [3-1:0] node1733;
	wire [3-1:0] node1734;
	wire [3-1:0] node1735;
	wire [3-1:0] node1736;
	wire [3-1:0] node1739;
	wire [3-1:0] node1742;
	wire [3-1:0] node1744;
	wire [3-1:0] node1747;
	wire [3-1:0] node1748;
	wire [3-1:0] node1749;
	wire [3-1:0] node1752;
	wire [3-1:0] node1755;
	wire [3-1:0] node1756;
	wire [3-1:0] node1759;
	wire [3-1:0] node1762;
	wire [3-1:0] node1763;
	wire [3-1:0] node1764;
	wire [3-1:0] node1767;
	wire [3-1:0] node1770;
	wire [3-1:0] node1772;
	wire [3-1:0] node1773;
	wire [3-1:0] node1776;
	wire [3-1:0] node1779;
	wire [3-1:0] node1780;
	wire [3-1:0] node1781;
	wire [3-1:0] node1782;
	wire [3-1:0] node1785;
	wire [3-1:0] node1788;
	wire [3-1:0] node1789;
	wire [3-1:0] node1791;
	wire [3-1:0] node1794;
	wire [3-1:0] node1795;
	wire [3-1:0] node1799;
	wire [3-1:0] node1800;
	wire [3-1:0] node1801;
	wire [3-1:0] node1804;
	wire [3-1:0] node1807;
	wire [3-1:0] node1808;
	wire [3-1:0] node1811;
	wire [3-1:0] node1814;
	wire [3-1:0] node1815;
	wire [3-1:0] node1816;
	wire [3-1:0] node1817;
	wire [3-1:0] node1818;
	wire [3-1:0] node1820;
	wire [3-1:0] node1823;
	wire [3-1:0] node1826;
	wire [3-1:0] node1827;
	wire [3-1:0] node1829;
	wire [3-1:0] node1832;
	wire [3-1:0] node1833;
	wire [3-1:0] node1836;
	wire [3-1:0] node1839;
	wire [3-1:0] node1840;
	wire [3-1:0] node1841;
	wire [3-1:0] node1842;
	wire [3-1:0] node1847;
	wire [3-1:0] node1848;
	wire [3-1:0] node1849;
	wire [3-1:0] node1854;
	wire [3-1:0] node1855;
	wire [3-1:0] node1856;
	wire [3-1:0] node1857;
	wire [3-1:0] node1858;
	wire [3-1:0] node1859;
	wire [3-1:0] node1862;
	wire [3-1:0] node1865;
	wire [3-1:0] node1866;
	wire [3-1:0] node1869;
	wire [3-1:0] node1873;
	wire [3-1:0] node1874;
	wire [3-1:0] node1878;
	wire [3-1:0] node1879;
	wire [3-1:0] node1880;
	wire [3-1:0] node1881;
	wire [3-1:0] node1884;
	wire [3-1:0] node1888;
	wire [3-1:0] node1889;
	wire [3-1:0] node1893;
	wire [3-1:0] node1894;
	wire [3-1:0] node1895;
	wire [3-1:0] node1896;
	wire [3-1:0] node1897;
	wire [3-1:0] node1898;
	wire [3-1:0] node1900;
	wire [3-1:0] node1903;
	wire [3-1:0] node1904;
	wire [3-1:0] node1908;
	wire [3-1:0] node1909;
	wire [3-1:0] node1911;
	wire [3-1:0] node1914;
	wire [3-1:0] node1916;
	wire [3-1:0] node1919;
	wire [3-1:0] node1920;
	wire [3-1:0] node1921;
	wire [3-1:0] node1923;
	wire [3-1:0] node1926;
	wire [3-1:0] node1928;
	wire [3-1:0] node1931;
	wire [3-1:0] node1932;
	wire [3-1:0] node1933;
	wire [3-1:0] node1937;
	wire [3-1:0] node1939;
	wire [3-1:0] node1942;
	wire [3-1:0] node1943;
	wire [3-1:0] node1944;
	wire [3-1:0] node1945;
	wire [3-1:0] node1946;
	wire [3-1:0] node1947;
	wire [3-1:0] node1950;
	wire [3-1:0] node1954;
	wire [3-1:0] node1955;
	wire [3-1:0] node1956;
	wire [3-1:0] node1959;
	wire [3-1:0] node1962;
	wire [3-1:0] node1963;
	wire [3-1:0] node1966;
	wire [3-1:0] node1969;
	wire [3-1:0] node1970;
	wire [3-1:0] node1972;
	wire [3-1:0] node1975;
	wire [3-1:0] node1976;
	wire [3-1:0] node1977;
	wire [3-1:0] node1981;
	wire [3-1:0] node1982;
	wire [3-1:0] node1985;
	wire [3-1:0] node1988;
	wire [3-1:0] node1989;
	wire [3-1:0] node1990;
	wire [3-1:0] node1993;
	wire [3-1:0] node1996;
	wire [3-1:0] node1997;
	wire [3-1:0] node2000;
	wire [3-1:0] node2003;
	wire [3-1:0] node2004;
	wire [3-1:0] node2005;
	wire [3-1:0] node2009;
	wire [3-1:0] node2010;
	wire [3-1:0] node2014;
	wire [3-1:0] node2015;
	wire [3-1:0] node2016;
	wire [3-1:0] node2017;
	wire [3-1:0] node2018;
	wire [3-1:0] node2019;
	wire [3-1:0] node2020;
	wire [3-1:0] node2021;
	wire [3-1:0] node2022;
	wire [3-1:0] node2023;
	wire [3-1:0] node2024;
	wire [3-1:0] node2027;
	wire [3-1:0] node2030;
	wire [3-1:0] node2031;
	wire [3-1:0] node2034;
	wire [3-1:0] node2037;
	wire [3-1:0] node2038;
	wire [3-1:0] node2039;
	wire [3-1:0] node2042;
	wire [3-1:0] node2045;
	wire [3-1:0] node2046;
	wire [3-1:0] node2049;
	wire [3-1:0] node2052;
	wire [3-1:0] node2053;
	wire [3-1:0] node2054;
	wire [3-1:0] node2055;
	wire [3-1:0] node2058;
	wire [3-1:0] node2061;
	wire [3-1:0] node2064;
	wire [3-1:0] node2065;
	wire [3-1:0] node2068;
	wire [3-1:0] node2071;
	wire [3-1:0] node2072;
	wire [3-1:0] node2073;
	wire [3-1:0] node2074;
	wire [3-1:0] node2077;
	wire [3-1:0] node2078;
	wire [3-1:0] node2081;
	wire [3-1:0] node2084;
	wire [3-1:0] node2085;
	wire [3-1:0] node2087;
	wire [3-1:0] node2090;
	wire [3-1:0] node2091;
	wire [3-1:0] node2094;
	wire [3-1:0] node2097;
	wire [3-1:0] node2098;
	wire [3-1:0] node2099;
	wire [3-1:0] node2100;
	wire [3-1:0] node2104;
	wire [3-1:0] node2105;
	wire [3-1:0] node2108;
	wire [3-1:0] node2111;
	wire [3-1:0] node2112;
	wire [3-1:0] node2114;
	wire [3-1:0] node2117;
	wire [3-1:0] node2119;
	wire [3-1:0] node2122;
	wire [3-1:0] node2123;
	wire [3-1:0] node2124;
	wire [3-1:0] node2125;
	wire [3-1:0] node2127;
	wire [3-1:0] node2130;
	wire [3-1:0] node2131;
	wire [3-1:0] node2135;
	wire [3-1:0] node2136;
	wire [3-1:0] node2138;
	wire [3-1:0] node2139;
	wire [3-1:0] node2142;
	wire [3-1:0] node2145;
	wire [3-1:0] node2146;
	wire [3-1:0] node2149;
	wire [3-1:0] node2152;
	wire [3-1:0] node2153;
	wire [3-1:0] node2154;
	wire [3-1:0] node2156;
	wire [3-1:0] node2159;
	wire [3-1:0] node2160;
	wire [3-1:0] node2164;
	wire [3-1:0] node2167;
	wire [3-1:0] node2168;
	wire [3-1:0] node2169;
	wire [3-1:0] node2170;
	wire [3-1:0] node2171;
	wire [3-1:0] node2172;
	wire [3-1:0] node2175;
	wire [3-1:0] node2176;
	wire [3-1:0] node2179;
	wire [3-1:0] node2182;
	wire [3-1:0] node2183;
	wire [3-1:0] node2184;
	wire [3-1:0] node2187;
	wire [3-1:0] node2190;
	wire [3-1:0] node2192;
	wire [3-1:0] node2195;
	wire [3-1:0] node2196;
	wire [3-1:0] node2197;
	wire [3-1:0] node2200;
	wire [3-1:0] node2202;
	wire [3-1:0] node2205;
	wire [3-1:0] node2206;
	wire [3-1:0] node2207;
	wire [3-1:0] node2210;
	wire [3-1:0] node2213;
	wire [3-1:0] node2214;
	wire [3-1:0] node2218;
	wire [3-1:0] node2219;
	wire [3-1:0] node2220;
	wire [3-1:0] node2221;
	wire [3-1:0] node2224;
	wire [3-1:0] node2227;
	wire [3-1:0] node2228;
	wire [3-1:0] node2231;
	wire [3-1:0] node2232;
	wire [3-1:0] node2235;
	wire [3-1:0] node2238;
	wire [3-1:0] node2239;
	wire [3-1:0] node2240;
	wire [3-1:0] node2241;
	wire [3-1:0] node2244;
	wire [3-1:0] node2247;
	wire [3-1:0] node2248;
	wire [3-1:0] node2251;
	wire [3-1:0] node2254;
	wire [3-1:0] node2255;
	wire [3-1:0] node2256;
	wire [3-1:0] node2259;
	wire [3-1:0] node2262;
	wire [3-1:0] node2263;
	wire [3-1:0] node2266;
	wire [3-1:0] node2269;
	wire [3-1:0] node2270;
	wire [3-1:0] node2271;
	wire [3-1:0] node2272;
	wire [3-1:0] node2274;
	wire [3-1:0] node2277;
	wire [3-1:0] node2279;
	wire [3-1:0] node2282;
	wire [3-1:0] node2283;
	wire [3-1:0] node2284;
	wire [3-1:0] node2288;
	wire [3-1:0] node2289;
	wire [3-1:0] node2292;
	wire [3-1:0] node2295;
	wire [3-1:0] node2296;
	wire [3-1:0] node2297;
	wire [3-1:0] node2299;
	wire [3-1:0] node2302;
	wire [3-1:0] node2303;
	wire [3-1:0] node2307;
	wire [3-1:0] node2310;
	wire [3-1:0] node2311;
	wire [3-1:0] node2312;
	wire [3-1:0] node2313;
	wire [3-1:0] node2314;
	wire [3-1:0] node2315;
	wire [3-1:0] node2316;
	wire [3-1:0] node2319;
	wire [3-1:0] node2322;
	wire [3-1:0] node2323;
	wire [3-1:0] node2324;
	wire [3-1:0] node2327;
	wire [3-1:0] node2330;
	wire [3-1:0] node2331;
	wire [3-1:0] node2335;
	wire [3-1:0] node2336;
	wire [3-1:0] node2337;
	wire [3-1:0] node2338;
	wire [3-1:0] node2343;
	wire [3-1:0] node2344;
	wire [3-1:0] node2348;
	wire [3-1:0] node2349;
	wire [3-1:0] node2350;
	wire [3-1:0] node2351;
	wire [3-1:0] node2354;
	wire [3-1:0] node2357;
	wire [3-1:0] node2358;
	wire [3-1:0] node2359;
	wire [3-1:0] node2362;
	wire [3-1:0] node2365;
	wire [3-1:0] node2368;
	wire [3-1:0] node2369;
	wire [3-1:0] node2370;
	wire [3-1:0] node2372;
	wire [3-1:0] node2376;
	wire [3-1:0] node2377;
	wire [3-1:0] node2380;
	wire [3-1:0] node2383;
	wire [3-1:0] node2384;
	wire [3-1:0] node2385;
	wire [3-1:0] node2386;
	wire [3-1:0] node2387;
	wire [3-1:0] node2391;
	wire [3-1:0] node2392;
	wire [3-1:0] node2396;
	wire [3-1:0] node2397;
	wire [3-1:0] node2398;
	wire [3-1:0] node2401;
	wire [3-1:0] node2404;
	wire [3-1:0] node2405;
	wire [3-1:0] node2406;
	wire [3-1:0] node2409;
	wire [3-1:0] node2412;
	wire [3-1:0] node2413;
	wire [3-1:0] node2417;
	wire [3-1:0] node2418;
	wire [3-1:0] node2419;
	wire [3-1:0] node2421;
	wire [3-1:0] node2424;
	wire [3-1:0] node2425;
	wire [3-1:0] node2429;
	wire [3-1:0] node2432;
	wire [3-1:0] node2433;
	wire [3-1:0] node2434;
	wire [3-1:0] node2435;
	wire [3-1:0] node2436;
	wire [3-1:0] node2438;
	wire [3-1:0] node2441;
	wire [3-1:0] node2443;
	wire [3-1:0] node2444;
	wire [3-1:0] node2448;
	wire [3-1:0] node2449;
	wire [3-1:0] node2450;
	wire [3-1:0] node2451;
	wire [3-1:0] node2454;
	wire [3-1:0] node2457;
	wire [3-1:0] node2460;
	wire [3-1:0] node2461;
	wire [3-1:0] node2464;
	wire [3-1:0] node2467;
	wire [3-1:0] node2468;
	wire [3-1:0] node2469;
	wire [3-1:0] node2471;
	wire [3-1:0] node2474;
	wire [3-1:0] node2475;
	wire [3-1:0] node2478;
	wire [3-1:0] node2480;
	wire [3-1:0] node2483;
	wire [3-1:0] node2484;
	wire [3-1:0] node2485;
	wire [3-1:0] node2486;
	wire [3-1:0] node2490;
	wire [3-1:0] node2492;
	wire [3-1:0] node2495;
	wire [3-1:0] node2498;
	wire [3-1:0] node2499;
	wire [3-1:0] node2500;
	wire [3-1:0] node2501;
	wire [3-1:0] node2503;
	wire [3-1:0] node2506;
	wire [3-1:0] node2507;
	wire [3-1:0] node2511;
	wire [3-1:0] node2512;
	wire [3-1:0] node2513;
	wire [3-1:0] node2516;
	wire [3-1:0] node2519;
	wire [3-1:0] node2520;
	wire [3-1:0] node2521;
	wire [3-1:0] node2524;
	wire [3-1:0] node2527;
	wire [3-1:0] node2528;
	wire [3-1:0] node2532;
	wire [3-1:0] node2533;
	wire [3-1:0] node2536;
	wire [3-1:0] node2537;
	wire [3-1:0] node2538;
	wire [3-1:0] node2543;
	wire [3-1:0] node2544;
	wire [3-1:0] node2545;
	wire [3-1:0] node2546;
	wire [3-1:0] node2547;
	wire [3-1:0] node2548;
	wire [3-1:0] node2549;
	wire [3-1:0] node2550;
	wire [3-1:0] node2551;
	wire [3-1:0] node2555;
	wire [3-1:0] node2556;
	wire [3-1:0] node2559;
	wire [3-1:0] node2562;
	wire [3-1:0] node2563;
	wire [3-1:0] node2566;
	wire [3-1:0] node2569;
	wire [3-1:0] node2570;
	wire [3-1:0] node2572;
	wire [3-1:0] node2574;
	wire [3-1:0] node2577;
	wire [3-1:0] node2579;
	wire [3-1:0] node2581;
	wire [3-1:0] node2584;
	wire [3-1:0] node2585;
	wire [3-1:0] node2586;
	wire [3-1:0] node2587;
	wire [3-1:0] node2589;
	wire [3-1:0] node2592;
	wire [3-1:0] node2594;
	wire [3-1:0] node2597;
	wire [3-1:0] node2598;
	wire [3-1:0] node2600;
	wire [3-1:0] node2603;
	wire [3-1:0] node2605;
	wire [3-1:0] node2608;
	wire [3-1:0] node2609;
	wire [3-1:0] node2610;
	wire [3-1:0] node2613;
	wire [3-1:0] node2616;
	wire [3-1:0] node2617;
	wire [3-1:0] node2618;
	wire [3-1:0] node2621;
	wire [3-1:0] node2625;
	wire [3-1:0] node2626;
	wire [3-1:0] node2627;
	wire [3-1:0] node2628;
	wire [3-1:0] node2629;
	wire [3-1:0] node2630;
	wire [3-1:0] node2634;
	wire [3-1:0] node2635;
	wire [3-1:0] node2639;
	wire [3-1:0] node2640;
	wire [3-1:0] node2642;
	wire [3-1:0] node2646;
	wire [3-1:0] node2647;
	wire [3-1:0] node2648;
	wire [3-1:0] node2649;
	wire [3-1:0] node2653;
	wire [3-1:0] node2656;
	wire [3-1:0] node2657;
	wire [3-1:0] node2658;
	wire [3-1:0] node2662;
	wire [3-1:0] node2665;
	wire [3-1:0] node2666;
	wire [3-1:0] node2667;
	wire [3-1:0] node2668;
	wire [3-1:0] node2669;
	wire [3-1:0] node2672;
	wire [3-1:0] node2676;
	wire [3-1:0] node2677;
	wire [3-1:0] node2678;
	wire [3-1:0] node2682;
	wire [3-1:0] node2683;
	wire [3-1:0] node2687;
	wire [3-1:0] node2688;
	wire [3-1:0] node2689;
	wire [3-1:0] node2690;
	wire [3-1:0] node2694;
	wire [3-1:0] node2695;
	wire [3-1:0] node2699;
	wire [3-1:0] node2700;
	wire [3-1:0] node2701;
	wire [3-1:0] node2705;
	wire [3-1:0] node2706;
	wire [3-1:0] node2710;
	wire [3-1:0] node2711;
	wire [3-1:0] node2712;
	wire [3-1:0] node2713;
	wire [3-1:0] node2714;
	wire [3-1:0] node2717;
	wire [3-1:0] node2721;
	wire [3-1:0] node2722;
	wire [3-1:0] node2726;
	wire [3-1:0] node2727;
	wire [3-1:0] node2728;
	wire [3-1:0] node2729;
	wire [3-1:0] node2730;
	wire [3-1:0] node2733;
	wire [3-1:0] node2736;
	wire [3-1:0] node2737;
	wire [3-1:0] node2740;
	wire [3-1:0] node2744;
	wire [3-1:0] node2745;
	wire [3-1:0] node2749;
	wire [3-1:0] node2750;
	wire [3-1:0] node2751;
	wire [3-1:0] node2752;
	wire [3-1:0] node2753;
	wire [3-1:0] node2754;
	wire [3-1:0] node2755;
	wire [3-1:0] node2757;
	wire [3-1:0] node2760;
	wire [3-1:0] node2761;
	wire [3-1:0] node2764;
	wire [3-1:0] node2767;
	wire [3-1:0] node2768;
	wire [3-1:0] node2769;
	wire [3-1:0] node2772;
	wire [3-1:0] node2775;
	wire [3-1:0] node2776;
	wire [3-1:0] node2780;
	wire [3-1:0] node2781;
	wire [3-1:0] node2782;
	wire [3-1:0] node2783;
	wire [3-1:0] node2786;
	wire [3-1:0] node2790;
	wire [3-1:0] node2791;
	wire [3-1:0] node2794;
	wire [3-1:0] node2795;
	wire [3-1:0] node2799;
	wire [3-1:0] node2800;
	wire [3-1:0] node2801;
	wire [3-1:0] node2802;
	wire [3-1:0] node2803;
	wire [3-1:0] node2806;
	wire [3-1:0] node2809;
	wire [3-1:0] node2810;
	wire [3-1:0] node2813;
	wire [3-1:0] node2816;
	wire [3-1:0] node2817;
	wire [3-1:0] node2818;
	wire [3-1:0] node2821;
	wire [3-1:0] node2824;
	wire [3-1:0] node2825;
	wire [3-1:0] node2828;
	wire [3-1:0] node2831;
	wire [3-1:0] node2832;
	wire [3-1:0] node2833;
	wire [3-1:0] node2837;
	wire [3-1:0] node2838;
	wire [3-1:0] node2839;
	wire [3-1:0] node2843;
	wire [3-1:0] node2845;
	wire [3-1:0] node2848;
	wire [3-1:0] node2849;
	wire [3-1:0] node2850;
	wire [3-1:0] node2851;
	wire [3-1:0] node2852;
	wire [3-1:0] node2855;
	wire [3-1:0] node2858;
	wire [3-1:0] node2859;
	wire [3-1:0] node2860;
	wire [3-1:0] node2863;
	wire [3-1:0] node2866;
	wire [3-1:0] node2867;
	wire [3-1:0] node2870;
	wire [3-1:0] node2873;
	wire [3-1:0] node2874;
	wire [3-1:0] node2875;
	wire [3-1:0] node2876;
	wire [3-1:0] node2880;
	wire [3-1:0] node2881;
	wire [3-1:0] node2885;
	wire [3-1:0] node2886;
	wire [3-1:0] node2887;
	wire [3-1:0] node2892;
	wire [3-1:0] node2893;
	wire [3-1:0] node2894;
	wire [3-1:0] node2895;
	wire [3-1:0] node2899;
	wire [3-1:0] node2900;
	wire [3-1:0] node2904;
	wire [3-1:0] node2905;
	wire [3-1:0] node2906;
	wire [3-1:0] node2910;
	wire [3-1:0] node2911;
	wire [3-1:0] node2915;
	wire [3-1:0] node2916;
	wire [3-1:0] node2917;
	wire [3-1:0] node2918;
	wire [3-1:0] node2919;
	wire [3-1:0] node2923;
	wire [3-1:0] node2924;
	wire [3-1:0] node2929;
	wire [3-1:0] node2930;
	wire [3-1:0] node2931;
	wire [3-1:0] node2932;
	wire [3-1:0] node2936;
	wire [3-1:0] node2937;
	wire [3-1:0] node2942;
	wire [3-1:0] node2943;
	wire [3-1:0] node2944;
	wire [3-1:0] node2945;
	wire [3-1:0] node2946;
	wire [3-1:0] node2947;
	wire [3-1:0] node2948;
	wire [3-1:0] node2949;
	wire [3-1:0] node2950;
	wire [3-1:0] node2953;
	wire [3-1:0] node2956;
	wire [3-1:0] node2957;
	wire [3-1:0] node2960;
	wire [3-1:0] node2963;
	wire [3-1:0] node2964;
	wire [3-1:0] node2966;
	wire [3-1:0] node2967;
	wire [3-1:0] node2970;
	wire [3-1:0] node2973;
	wire [3-1:0] node2974;
	wire [3-1:0] node2975;
	wire [3-1:0] node2978;
	wire [3-1:0] node2981;
	wire [3-1:0] node2983;
	wire [3-1:0] node2986;
	wire [3-1:0] node2987;
	wire [3-1:0] node2988;
	wire [3-1:0] node2991;
	wire [3-1:0] node2994;
	wire [3-1:0] node2995;
	wire [3-1:0] node2996;
	wire [3-1:0] node2999;
	wire [3-1:0] node3002;
	wire [3-1:0] node3003;
	wire [3-1:0] node3006;
	wire [3-1:0] node3009;
	wire [3-1:0] node3010;
	wire [3-1:0] node3011;
	wire [3-1:0] node3012;
	wire [3-1:0] node3016;
	wire [3-1:0] node3018;
	wire [3-1:0] node3021;
	wire [3-1:0] node3022;
	wire [3-1:0] node3023;
	wire [3-1:0] node3027;
	wire [3-1:0] node3028;
	wire [3-1:0] node3032;
	wire [3-1:0] node3033;
	wire [3-1:0] node3034;
	wire [3-1:0] node3035;
	wire [3-1:0] node3036;
	wire [3-1:0] node3037;
	wire [3-1:0] node3040;
	wire [3-1:0] node3043;
	wire [3-1:0] node3044;
	wire [3-1:0] node3047;
	wire [3-1:0] node3050;
	wire [3-1:0] node3051;
	wire [3-1:0] node3052;
	wire [3-1:0] node3055;
	wire [3-1:0] node3058;
	wire [3-1:0] node3060;
	wire [3-1:0] node3061;
	wire [3-1:0] node3064;
	wire [3-1:0] node3067;
	wire [3-1:0] node3068;
	wire [3-1:0] node3069;
	wire [3-1:0] node3072;
	wire [3-1:0] node3075;
	wire [3-1:0] node3076;
	wire [3-1:0] node3079;
	wire [3-1:0] node3082;
	wire [3-1:0] node3083;
	wire [3-1:0] node3084;
	wire [3-1:0] node3085;
	wire [3-1:0] node3086;
	wire [3-1:0] node3087;
	wire [3-1:0] node3090;
	wire [3-1:0] node3093;
	wire [3-1:0] node3094;
	wire [3-1:0] node3097;
	wire [3-1:0] node3100;
	wire [3-1:0] node3101;
	wire [3-1:0] node3104;
	wire [3-1:0] node3107;
	wire [3-1:0] node3108;
	wire [3-1:0] node3109;
	wire [3-1:0] node3110;
	wire [3-1:0] node3113;
	wire [3-1:0] node3116;
	wire [3-1:0] node3117;
	wire [3-1:0] node3120;
	wire [3-1:0] node3123;
	wire [3-1:0] node3124;
	wire [3-1:0] node3127;
	wire [3-1:0] node3130;
	wire [3-1:0] node3131;
	wire [3-1:0] node3134;
	wire [3-1:0] node3137;
	wire [3-1:0] node3138;
	wire [3-1:0] node3139;
	wire [3-1:0] node3140;
	wire [3-1:0] node3141;
	wire [3-1:0] node3142;
	wire [3-1:0] node3143;
	wire [3-1:0] node3147;
	wire [3-1:0] node3149;
	wire [3-1:0] node3152;
	wire [3-1:0] node3153;
	wire [3-1:0] node3155;
	wire [3-1:0] node3158;
	wire [3-1:0] node3160;
	wire [3-1:0] node3163;
	wire [3-1:0] node3164;
	wire [3-1:0] node3165;
	wire [3-1:0] node3166;
	wire [3-1:0] node3170;
	wire [3-1:0] node3172;
	wire [3-1:0] node3175;
	wire [3-1:0] node3176;
	wire [3-1:0] node3178;
	wire [3-1:0] node3181;
	wire [3-1:0] node3182;
	wire [3-1:0] node3186;
	wire [3-1:0] node3187;
	wire [3-1:0] node3190;
	wire [3-1:0] node3193;
	wire [3-1:0] node3194;
	wire [3-1:0] node3195;
	wire [3-1:0] node3196;
	wire [3-1:0] node3197;
	wire [3-1:0] node3201;
	wire [3-1:0] node3202;
	wire [3-1:0] node3207;
	wire [3-1:0] node3208;
	wire [3-1:0] node3209;
	wire [3-1:0] node3210;
	wire [3-1:0] node3214;
	wire [3-1:0] node3215;
	wire [3-1:0] node3220;
	wire [3-1:0] node3221;
	wire [3-1:0] node3222;
	wire [3-1:0] node3223;
	wire [3-1:0] node3224;
	wire [3-1:0] node3225;
	wire [3-1:0] node3226;
	wire [3-1:0] node3227;
	wire [3-1:0] node3230;
	wire [3-1:0] node3233;
	wire [3-1:0] node3234;
	wire [3-1:0] node3237;
	wire [3-1:0] node3240;
	wire [3-1:0] node3241;
	wire [3-1:0] node3242;
	wire [3-1:0] node3246;
	wire [3-1:0] node3247;
	wire [3-1:0] node3248;
	wire [3-1:0] node3251;
	wire [3-1:0] node3254;
	wire [3-1:0] node3256;
	wire [3-1:0] node3259;
	wire [3-1:0] node3260;
	wire [3-1:0] node3261;
	wire [3-1:0] node3264;
	wire [3-1:0] node3267;
	wire [3-1:0] node3268;
	wire [3-1:0] node3269;
	wire [3-1:0] node3272;
	wire [3-1:0] node3275;
	wire [3-1:0] node3276;
	wire [3-1:0] node3277;
	wire [3-1:0] node3280;
	wire [3-1:0] node3283;
	wire [3-1:0] node3285;
	wire [3-1:0] node3288;
	wire [3-1:0] node3289;
	wire [3-1:0] node3290;
	wire [3-1:0] node3293;
	wire [3-1:0] node3296;
	wire [3-1:0] node3297;
	wire [3-1:0] node3300;
	wire [3-1:0] node3303;
	wire [3-1:0] node3304;
	wire [3-1:0] node3305;
	wire [3-1:0] node3309;
	wire [3-1:0] node3310;
	wire [3-1:0] node3314;
	wire [3-1:0] node3315;
	wire [3-1:0] node3316;
	wire [3-1:0] node3317;
	wire [3-1:0] node3321;
	wire [3-1:0] node3322;
	wire [3-1:0] node3326;
	wire [3-1:0] node3327;

	assign outp = (inp[5]) ? node2014 : node1;
		assign node1 = (inp[8]) ? node1339 : node2;
			assign node2 = (inp[6]) ? node714 : node3;
				assign node3 = (inp[4]) ? node389 : node4;
					assign node4 = (inp[1]) ? node196 : node5;
						assign node5 = (inp[7]) ? node113 : node6;
							assign node6 = (inp[11]) ? node56 : node7;
								assign node7 = (inp[2]) ? node27 : node8;
									assign node8 = (inp[9]) ? node18 : node9;
										assign node9 = (inp[0]) ? node11 : 3'b010;
											assign node11 = (inp[3]) ? node15 : node12;
												assign node12 = (inp[10]) ? 3'b011 : 3'b001;
												assign node15 = (inp[10]) ? 3'b001 : 3'b011;
										assign node18 = (inp[0]) ? 3'b000 : node19;
											assign node19 = (inp[10]) ? node23 : node20;
												assign node20 = (inp[3]) ? 3'b011 : 3'b001;
												assign node23 = (inp[3]) ? 3'b001 : 3'b011;
									assign node27 = (inp[0]) ? node41 : node28;
										assign node28 = (inp[9]) ? node34 : node29;
											assign node29 = (inp[3]) ? 3'b001 : node30;
												assign node30 = (inp[10]) ? 3'b010 : 3'b000;
											assign node34 = (inp[10]) ? node38 : node35;
												assign node35 = (inp[3]) ? 3'b011 : 3'b001;
												assign node38 = (inp[3]) ? 3'b000 : 3'b011;
										assign node41 = (inp[9]) ? node49 : node42;
											assign node42 = (inp[3]) ? node46 : node43;
												assign node43 = (inp[10]) ? 3'b011 : 3'b001;
												assign node46 = (inp[10]) ? 3'b000 : 3'b011;
											assign node49 = (inp[3]) ? node53 : node50;
												assign node50 = (inp[10]) ? 3'b010 : 3'b000;
												assign node53 = (inp[10]) ? 3'b001 : 3'b010;
								assign node56 = (inp[2]) ? node86 : node57;
									assign node57 = (inp[0]) ? node71 : node58;
										assign node58 = (inp[9]) ? node64 : node59;
											assign node59 = (inp[10]) ? 3'b001 : node60;
												assign node60 = (inp[3]) ? 3'b010 : 3'b000;
											assign node64 = (inp[10]) ? node68 : node65;
												assign node65 = (inp[3]) ? 3'b011 : 3'b001;
												assign node68 = (inp[3]) ? 3'b000 : 3'b010;
										assign node71 = (inp[3]) ? node79 : node72;
											assign node72 = (inp[10]) ? node76 : node73;
												assign node73 = (inp[9]) ? 3'b000 : 3'b001;
												assign node76 = (inp[9]) ? 3'b011 : 3'b010;
											assign node79 = (inp[10]) ? node83 : node80;
												assign node80 = (inp[9]) ? 3'b010 : 3'b011;
												assign node83 = (inp[9]) ? 3'b001 : 3'b000;
									assign node86 = (inp[10]) ? node98 : node87;
										assign node87 = (inp[3]) ? node93 : node88;
											assign node88 = (inp[0]) ? node90 : 3'b001;
												assign node90 = (inp[9]) ? 3'b000 : 3'b001;
											assign node93 = (inp[9]) ? 3'b011 : node94;
												assign node94 = (inp[0]) ? 3'b011 : 3'b010;
										assign node98 = (inp[3]) ? node106 : node99;
											assign node99 = (inp[9]) ? node103 : node100;
												assign node100 = (inp[0]) ? 3'b010 : 3'b011;
												assign node103 = (inp[0]) ? 3'b011 : 3'b010;
											assign node106 = (inp[9]) ? node110 : node107;
												assign node107 = (inp[0]) ? 3'b001 : 3'b000;
												assign node110 = (inp[0]) ? 3'b000 : 3'b001;
							assign node113 = (inp[9]) ? node151 : node114;
								assign node114 = (inp[0]) ? node132 : node115;
									assign node115 = (inp[3]) ? node123 : node116;
										assign node116 = (inp[11]) ? node120 : node117;
											assign node117 = (inp[10]) ? 3'b010 : 3'b000;
											assign node120 = (inp[10]) ? 3'b000 : 3'b010;
										assign node123 = (inp[10]) ? node127 : node124;
											assign node124 = (inp[11]) ? 3'b000 : 3'b011;
											assign node127 = (inp[11]) ? 3'b011 : node128;
												assign node128 = (inp[2]) ? 3'b000 : 3'b001;
									assign node132 = (inp[3]) ? node142 : node133;
										assign node133 = (inp[10]) ? node139 : node134;
											assign node134 = (inp[11]) ? node136 : 3'b001;
												assign node136 = (inp[2]) ? 3'b010 : 3'b011;
											assign node139 = (inp[11]) ? 3'b001 : 3'b011;
										assign node142 = (inp[11]) ? node148 : node143;
											assign node143 = (inp[10]) ? node145 : 3'b010;
												assign node145 = (inp[2]) ? 3'b001 : 3'b000;
											assign node148 = (inp[10]) ? 3'b010 : 3'b001;
								assign node151 = (inp[0]) ? node171 : node152;
									assign node152 = (inp[3]) ? node162 : node153;
										assign node153 = (inp[10]) ? node159 : node154;
											assign node154 = (inp[11]) ? node156 : 3'b001;
												assign node156 = (inp[2]) ? 3'b010 : 3'b011;
											assign node159 = (inp[11]) ? 3'b001 : 3'b011;
										assign node162 = (inp[10]) ? node166 : node163;
											assign node163 = (inp[11]) ? 3'b001 : 3'b010;
											assign node166 = (inp[11]) ? 3'b010 : node167;
												assign node167 = (inp[2]) ? 3'b001 : 3'b000;
									assign node171 = (inp[3]) ? node181 : node172;
										assign node172 = (inp[11]) ? node176 : node173;
											assign node173 = (inp[10]) ? 3'b010 : 3'b000;
											assign node176 = (inp[10]) ? 3'b000 : node177;
												assign node177 = (inp[2]) ? 3'b011 : 3'b010;
										assign node181 = (inp[2]) ? node189 : node182;
											assign node182 = (inp[10]) ? node186 : node183;
												assign node183 = (inp[11]) ? 3'b000 : 3'b011;
												assign node186 = (inp[11]) ? 3'b011 : 3'b001;
											assign node189 = (inp[11]) ? node193 : node190;
												assign node190 = (inp[10]) ? 3'b000 : 3'b011;
												assign node193 = (inp[10]) ? 3'b011 : 3'b000;
						assign node196 = (inp[2]) ? node282 : node197;
							assign node197 = (inp[0]) ? node241 : node198;
								assign node198 = (inp[9]) ? node222 : node199;
									assign node199 = (inp[3]) ? node207 : node200;
										assign node200 = (inp[10]) ? node202 : 3'b000;
											assign node202 = (inp[11]) ? node204 : 3'b010;
												assign node204 = (inp[7]) ? 3'b000 : 3'b011;
										assign node207 = (inp[10]) ? node215 : node208;
											assign node208 = (inp[11]) ? node212 : node209;
												assign node209 = (inp[7]) ? 3'b011 : 3'b010;
												assign node212 = (inp[7]) ? 3'b000 : 3'b010;
											assign node215 = (inp[11]) ? node219 : node216;
												assign node216 = (inp[7]) ? 3'b000 : 3'b001;
												assign node219 = (inp[7]) ? 3'b011 : 3'b000;
									assign node222 = (inp[10]) ? node234 : node223;
										assign node223 = (inp[3]) ? node229 : node224;
											assign node224 = (inp[7]) ? node226 : 3'b001;
												assign node226 = (inp[11]) ? 3'b010 : 3'b001;
											assign node229 = (inp[7]) ? node231 : 3'b011;
												assign node231 = (inp[11]) ? 3'b001 : 3'b010;
										assign node234 = (inp[11]) ? 3'b010 : node235;
											assign node235 = (inp[3]) ? node237 : 3'b011;
												assign node237 = (inp[7]) ? 3'b001 : 3'b000;
								assign node241 = (inp[9]) ? node265 : node242;
									assign node242 = (inp[3]) ? node250 : node243;
										assign node243 = (inp[10]) ? node247 : node244;
											assign node244 = (inp[11]) ? 3'b010 : 3'b001;
											assign node247 = (inp[11]) ? 3'b001 : 3'b011;
										assign node250 = (inp[10]) ? node258 : node251;
											assign node251 = (inp[11]) ? node255 : node252;
												assign node252 = (inp[7]) ? 3'b010 : 3'b011;
												assign node255 = (inp[7]) ? 3'b001 : 3'b011;
											assign node258 = (inp[11]) ? node262 : node259;
												assign node259 = (inp[7]) ? 3'b001 : 3'b000;
												assign node262 = (inp[7]) ? 3'b010 : 3'b001;
									assign node265 = (inp[11]) ? node275 : node266;
										assign node266 = (inp[3]) ? node270 : node267;
											assign node267 = (inp[10]) ? 3'b010 : 3'b000;
											assign node270 = (inp[10]) ? node272 : 3'b010;
												assign node272 = (inp[7]) ? 3'b000 : 3'b001;
										assign node275 = (inp[7]) ? 3'b011 : node276;
											assign node276 = (inp[3]) ? 3'b000 : node277;
												assign node277 = (inp[10]) ? 3'b011 : 3'b000;
							assign node282 = (inp[11]) ? node334 : node283;
								assign node283 = (inp[3]) ? node305 : node284;
									assign node284 = (inp[10]) ? node290 : node285;
										assign node285 = (inp[0]) ? node287 : 3'b001;
											assign node287 = (inp[9]) ? 3'b001 : 3'b000;
										assign node290 = (inp[7]) ? node298 : node291;
											assign node291 = (inp[0]) ? node295 : node292;
												assign node292 = (inp[9]) ? 3'b010 : 3'b011;
												assign node295 = (inp[9]) ? 3'b011 : 3'b010;
											assign node298 = (inp[9]) ? node302 : node299;
												assign node299 = (inp[0]) ? 3'b010 : 3'b011;
												assign node302 = (inp[0]) ? 3'b011 : 3'b010;
									assign node305 = (inp[10]) ? node321 : node306;
										assign node306 = (inp[7]) ? node314 : node307;
											assign node307 = (inp[9]) ? node311 : node308;
												assign node308 = (inp[0]) ? 3'b010 : 3'b011;
												assign node311 = (inp[0]) ? 3'b011 : 3'b010;
											assign node314 = (inp[9]) ? node318 : node315;
												assign node315 = (inp[0]) ? 3'b011 : 3'b010;
												assign node318 = (inp[0]) ? 3'b010 : 3'b011;
										assign node321 = (inp[0]) ? node329 : node322;
											assign node322 = (inp[7]) ? node326 : node323;
												assign node323 = (inp[9]) ? 3'b000 : 3'b001;
												assign node326 = (inp[9]) ? 3'b001 : 3'b000;
											assign node329 = (inp[9]) ? node331 : 3'b001;
												assign node331 = (inp[7]) ? 3'b000 : 3'b001;
								assign node334 = (inp[10]) ? node364 : node335;
									assign node335 = (inp[7]) ? node351 : node336;
										assign node336 = (inp[3]) ? node344 : node337;
											assign node337 = (inp[0]) ? node341 : node338;
												assign node338 = (inp[9]) ? 3'b000 : 3'b001;
												assign node341 = (inp[9]) ? 3'b001 : 3'b000;
											assign node344 = (inp[9]) ? node348 : node345;
												assign node345 = (inp[0]) ? 3'b010 : 3'b011;
												assign node348 = (inp[0]) ? 3'b011 : 3'b010;
										assign node351 = (inp[3]) ? node357 : node352;
											assign node352 = (inp[9]) ? 3'b010 : node353;
												assign node353 = (inp[0]) ? 3'b010 : 3'b011;
											assign node357 = (inp[0]) ? node361 : node358;
												assign node358 = (inp[9]) ? 3'b000 : 3'b001;
												assign node361 = (inp[9]) ? 3'b001 : 3'b000;
									assign node364 = (inp[9]) ? node378 : node365;
										assign node365 = (inp[0]) ? node371 : node366;
											assign node366 = (inp[7]) ? node368 : 3'b010;
												assign node368 = (inp[3]) ? 3'b010 : 3'b001;
											assign node371 = (inp[3]) ? node375 : node372;
												assign node372 = (inp[7]) ? 3'b000 : 3'b011;
												assign node375 = (inp[7]) ? 3'b011 : 3'b001;
										assign node378 = (inp[0]) ? node384 : node379;
											assign node379 = (inp[7]) ? node381 : 3'b011;
												assign node381 = (inp[3]) ? 3'b011 : 3'b000;
											assign node384 = (inp[7]) ? 3'b010 : node385;
												assign node385 = (inp[3]) ? 3'b000 : 3'b010;
					assign node389 = (inp[3]) ? node563 : node390;
						assign node390 = (inp[1]) ? node490 : node391;
							assign node391 = (inp[9]) ? node443 : node392;
								assign node392 = (inp[11]) ? node414 : node393;
									assign node393 = (inp[10]) ? node407 : node394;
										assign node394 = (inp[7]) ? node402 : node395;
											assign node395 = (inp[0]) ? node399 : node396;
												assign node396 = (inp[2]) ? 3'b101 : 3'b100;
												assign node399 = (inp[2]) ? 3'b100 : 3'b101;
											assign node402 = (inp[0]) ? 3'b100 : node403;
												assign node403 = (inp[2]) ? 3'b101 : 3'b100;
										assign node407 = (inp[2]) ? node411 : node408;
											assign node408 = (inp[0]) ? 3'b111 : 3'b110;
											assign node411 = (inp[0]) ? 3'b110 : 3'b111;
									assign node414 = (inp[10]) ? node430 : node415;
										assign node415 = (inp[7]) ? node423 : node416;
											assign node416 = (inp[0]) ? node420 : node417;
												assign node417 = (inp[2]) ? 3'b111 : 3'b110;
												assign node420 = (inp[2]) ? 3'b110 : 3'b111;
											assign node423 = (inp[0]) ? node427 : node424;
												assign node424 = (inp[2]) ? 3'b111 : 3'b110;
												assign node427 = (inp[2]) ? 3'b110 : 3'b111;
										assign node430 = (inp[2]) ? node436 : node431;
											assign node431 = (inp[7]) ? 3'b101 : node432;
												assign node432 = (inp[0]) ? 3'b100 : 3'b101;
											assign node436 = (inp[0]) ? node440 : node437;
												assign node437 = (inp[7]) ? 3'b101 : 3'b100;
												assign node440 = (inp[7]) ? 3'b100 : 3'b101;
								assign node443 = (inp[7]) ? node467 : node444;
									assign node444 = (inp[2]) ? node460 : node445;
										assign node445 = (inp[0]) ? node453 : node446;
											assign node446 = (inp[11]) ? node450 : node447;
												assign node447 = (inp[10]) ? 3'b110 : 3'b100;
												assign node450 = (inp[10]) ? 3'b101 : 3'b110;
											assign node453 = (inp[10]) ? node457 : node454;
												assign node454 = (inp[11]) ? 3'b111 : 3'b101;
												assign node457 = (inp[11]) ? 3'b100 : 3'b111;
										assign node460 = (inp[0]) ? 3'b110 : node461;
											assign node461 = (inp[10]) ? node463 : 3'b111;
												assign node463 = (inp[11]) ? 3'b100 : 3'b111;
									assign node467 = (inp[11]) ? node479 : node468;
										assign node468 = (inp[10]) ? node474 : node469;
											assign node469 = (inp[2]) ? 3'b100 : node470;
												assign node470 = (inp[0]) ? 3'b101 : 3'b100;
											assign node474 = (inp[2]) ? node476 : 3'b110;
												assign node476 = (inp[0]) ? 3'b110 : 3'b111;
										assign node479 = (inp[10]) ? node485 : node480;
											assign node480 = (inp[2]) ? 3'b110 : node481;
												assign node481 = (inp[0]) ? 3'b111 : 3'b110;
											assign node485 = (inp[0]) ? 3'b100 : node486;
												assign node486 = (inp[2]) ? 3'b101 : 3'b100;
							assign node490 = (inp[11]) ? node522 : node491;
								assign node491 = (inp[10]) ? node499 : node492;
									assign node492 = (inp[2]) ? node496 : node493;
										assign node493 = (inp[0]) ? 3'b101 : 3'b100;
										assign node496 = (inp[0]) ? 3'b100 : 3'b101;
									assign node499 = (inp[9]) ? node515 : node500;
										assign node500 = (inp[7]) ? node508 : node501;
											assign node501 = (inp[0]) ? node505 : node502;
												assign node502 = (inp[2]) ? 3'b111 : 3'b110;
												assign node505 = (inp[2]) ? 3'b110 : 3'b111;
											assign node508 = (inp[0]) ? node512 : node509;
												assign node509 = (inp[2]) ? 3'b111 : 3'b110;
												assign node512 = (inp[2]) ? 3'b110 : 3'b111;
										assign node515 = (inp[0]) ? node519 : node516;
											assign node516 = (inp[2]) ? 3'b111 : 3'b110;
											assign node519 = (inp[2]) ? 3'b110 : 3'b111;
								assign node522 = (inp[10]) ? node542 : node523;
									assign node523 = (inp[2]) ? node531 : node524;
										assign node524 = (inp[7]) ? node528 : node525;
											assign node525 = (inp[0]) ? 3'b111 : 3'b110;
											assign node528 = (inp[0]) ? 3'b110 : 3'b111;
										assign node531 = (inp[9]) ? node537 : node532;
											assign node532 = (inp[7]) ? 3'b110 : node533;
												assign node533 = (inp[0]) ? 3'b110 : 3'b111;
											assign node537 = (inp[7]) ? node539 : 3'b110;
												assign node539 = (inp[0]) ? 3'b111 : 3'b110;
									assign node542 = (inp[9]) ? node556 : node543;
										assign node543 = (inp[7]) ? node551 : node544;
											assign node544 = (inp[2]) ? node548 : node545;
												assign node545 = (inp[0]) ? 3'b101 : 3'b100;
												assign node548 = (inp[0]) ? 3'b100 : 3'b101;
											assign node551 = (inp[2]) ? 3'b100 : node552;
												assign node552 = (inp[0]) ? 3'b101 : 3'b100;
										assign node556 = (inp[2]) ? node560 : node557;
											assign node557 = (inp[0]) ? 3'b101 : 3'b100;
											assign node560 = (inp[0]) ? 3'b100 : 3'b101;
						assign node563 = (inp[10]) ? node625 : node564;
							assign node564 = (inp[11]) ? node604 : node565;
								assign node565 = (inp[1]) ? node589 : node566;
									assign node566 = (inp[2]) ? node582 : node567;
										assign node567 = (inp[9]) ? node575 : node568;
											assign node568 = (inp[7]) ? node572 : node569;
												assign node569 = (inp[0]) ? 3'b101 : 3'b100;
												assign node572 = (inp[0]) ? 3'b100 : 3'b101;
											assign node575 = (inp[0]) ? node579 : node576;
												assign node576 = (inp[7]) ? 3'b101 : 3'b100;
												assign node579 = (inp[7]) ? 3'b100 : 3'b101;
										assign node582 = (inp[0]) ? node586 : node583;
											assign node583 = (inp[7]) ? 3'b100 : 3'b101;
											assign node586 = (inp[7]) ? 3'b101 : 3'b100;
									assign node589 = (inp[7]) ? node597 : node590;
										assign node590 = (inp[2]) ? node594 : node591;
											assign node591 = (inp[0]) ? 3'b100 : 3'b101;
											assign node594 = (inp[0]) ? 3'b101 : 3'b100;
										assign node597 = (inp[0]) ? node601 : node598;
											assign node598 = (inp[2]) ? 3'b101 : 3'b100;
											assign node601 = (inp[2]) ? 3'b100 : 3'b101;
								assign node604 = (inp[0]) ? node614 : node605;
									assign node605 = (inp[2]) ? node609 : node606;
										assign node606 = (inp[7]) ? 3'b110 : 3'b111;
										assign node609 = (inp[7]) ? 3'b111 : node610;
											assign node610 = (inp[1]) ? 3'b110 : 3'b111;
									assign node614 = (inp[2]) ? node620 : node615;
										assign node615 = (inp[7]) ? 3'b111 : node616;
											assign node616 = (inp[1]) ? 3'b110 : 3'b111;
										assign node620 = (inp[1]) ? node622 : 3'b110;
											assign node622 = (inp[7]) ? 3'b110 : 3'b111;
							assign node625 = (inp[11]) ? node685 : node626;
								assign node626 = (inp[9]) ? node656 : node627;
									assign node627 = (inp[7]) ? node641 : node628;
										assign node628 = (inp[0]) ? node636 : node629;
											assign node629 = (inp[1]) ? node633 : node630;
												assign node630 = (inp[2]) ? 3'b111 : 3'b110;
												assign node633 = (inp[2]) ? 3'b110 : 3'b111;
											assign node636 = (inp[2]) ? 3'b110 : node637;
												assign node637 = (inp[1]) ? 3'b110 : 3'b111;
										assign node641 = (inp[2]) ? node649 : node642;
											assign node642 = (inp[0]) ? node646 : node643;
												assign node643 = (inp[1]) ? 3'b110 : 3'b111;
												assign node646 = (inp[1]) ? 3'b111 : 3'b110;
											assign node649 = (inp[1]) ? node653 : node650;
												assign node650 = (inp[0]) ? 3'b111 : 3'b110;
												assign node653 = (inp[0]) ? 3'b110 : 3'b111;
									assign node656 = (inp[7]) ? node670 : node657;
										assign node657 = (inp[2]) ? node665 : node658;
											assign node658 = (inp[1]) ? node662 : node659;
												assign node659 = (inp[0]) ? 3'b111 : 3'b110;
												assign node662 = (inp[0]) ? 3'b110 : 3'b111;
											assign node665 = (inp[1]) ? 3'b111 : node666;
												assign node666 = (inp[0]) ? 3'b110 : 3'b111;
										assign node670 = (inp[1]) ? node678 : node671;
											assign node671 = (inp[2]) ? node675 : node672;
												assign node672 = (inp[0]) ? 3'b110 : 3'b111;
												assign node675 = (inp[0]) ? 3'b111 : 3'b110;
											assign node678 = (inp[2]) ? node682 : node679;
												assign node679 = (inp[0]) ? 3'b111 : 3'b110;
												assign node682 = (inp[0]) ? 3'b110 : 3'b111;
								assign node685 = (inp[7]) ? node699 : node686;
									assign node686 = (inp[1]) ? node694 : node687;
										assign node687 = (inp[0]) ? node691 : node688;
											assign node688 = (inp[2]) ? 3'b101 : 3'b100;
											assign node691 = (inp[2]) ? 3'b100 : 3'b101;
										assign node694 = (inp[0]) ? 3'b101 : node695;
											assign node695 = (inp[2]) ? 3'b101 : 3'b100;
									assign node699 = (inp[1]) ? node707 : node700;
										assign node700 = (inp[0]) ? node704 : node701;
											assign node701 = (inp[2]) ? 3'b100 : 3'b101;
											assign node704 = (inp[2]) ? 3'b101 : 3'b100;
										assign node707 = (inp[2]) ? node711 : node708;
											assign node708 = (inp[0]) ? 3'b101 : 3'b100;
											assign node711 = (inp[0]) ? 3'b100 : 3'b101;
				assign node714 = (inp[1]) ? node1044 : node715;
					assign node715 = (inp[0]) ? node889 : node716;
						assign node716 = (inp[2]) ? node798 : node717;
							assign node717 = (inp[10]) ? node751 : node718;
								assign node718 = (inp[11]) ? node736 : node719;
									assign node719 = (inp[4]) ? 3'b100 : node720;
										assign node720 = (inp[9]) ? node728 : node721;
											assign node721 = (inp[3]) ? node725 : node722;
												assign node722 = (inp[7]) ? 3'b110 : 3'b100;
												assign node725 = (inp[7]) ? 3'b101 : 3'b110;
											assign node728 = (inp[7]) ? node732 : node729;
												assign node729 = (inp[3]) ? 3'b111 : 3'b101;
												assign node732 = (inp[3]) ? 3'b100 : 3'b111;
									assign node736 = (inp[3]) ? node746 : node737;
										assign node737 = (inp[4]) ? node743 : node738;
											assign node738 = (inp[9]) ? 3'b100 : node739;
												assign node739 = (inp[7]) ? 3'b101 : 3'b100;
											assign node743 = (inp[7]) ? 3'b111 : 3'b110;
										assign node746 = (inp[9]) ? node748 : 3'b110;
											assign node748 = (inp[4]) ? 3'b110 : 3'b111;
								assign node751 = (inp[11]) ? node783 : node752;
									assign node752 = (inp[4]) ? node768 : node753;
										assign node753 = (inp[9]) ? node761 : node754;
											assign node754 = (inp[7]) ? node758 : node755;
												assign node755 = (inp[3]) ? 3'b101 : 3'b110;
												assign node758 = (inp[3]) ? 3'b110 : 3'b101;
											assign node761 = (inp[3]) ? node765 : node762;
												assign node762 = (inp[7]) ? 3'b100 : 3'b111;
												assign node765 = (inp[7]) ? 3'b111 : 3'b100;
										assign node768 = (inp[9]) ? node776 : node769;
											assign node769 = (inp[3]) ? node773 : node770;
												assign node770 = (inp[7]) ? 3'b111 : 3'b110;
												assign node773 = (inp[7]) ? 3'b110 : 3'b111;
											assign node776 = (inp[7]) ? node780 : node777;
												assign node777 = (inp[3]) ? 3'b111 : 3'b110;
												assign node780 = (inp[3]) ? 3'b110 : 3'b111;
									assign node783 = (inp[3]) ? node793 : node784;
										assign node784 = (inp[4]) ? 3'b101 : node785;
											assign node785 = (inp[9]) ? node789 : node786;
												assign node786 = (inp[7]) ? 3'b110 : 3'b111;
												assign node789 = (inp[7]) ? 3'b111 : 3'b110;
										assign node793 = (inp[4]) ? 3'b100 : node794;
											assign node794 = (inp[7]) ? 3'b101 : 3'b100;
							assign node798 = (inp[4]) ? node850 : node799;
								assign node799 = (inp[9]) ? node825 : node800;
									assign node800 = (inp[3]) ? node814 : node801;
										assign node801 = (inp[10]) ? node807 : node802;
											assign node802 = (inp[11]) ? node804 : 3'b110;
												assign node804 = (inp[7]) ? 3'b101 : 3'b100;
											assign node807 = (inp[11]) ? node811 : node808;
												assign node808 = (inp[7]) ? 3'b101 : 3'b111;
												assign node811 = (inp[7]) ? 3'b111 : 3'b110;
										assign node814 = (inp[10]) ? node820 : node815;
											assign node815 = (inp[11]) ? 3'b110 : node816;
												assign node816 = (inp[7]) ? 3'b100 : 3'b110;
											assign node820 = (inp[11]) ? 3'b100 : node821;
												assign node821 = (inp[7]) ? 3'b110 : 3'b101;
									assign node825 = (inp[3]) ? node841 : node826;
										assign node826 = (inp[10]) ? node834 : node827;
											assign node827 = (inp[11]) ? node831 : node828;
												assign node828 = (inp[7]) ? 3'b111 : 3'b101;
												assign node831 = (inp[7]) ? 3'b100 : 3'b101;
											assign node834 = (inp[7]) ? node838 : node835;
												assign node835 = (inp[11]) ? 3'b111 : 3'b110;
												assign node838 = (inp[11]) ? 3'b110 : 3'b100;
										assign node841 = (inp[7]) ? node843 : 3'b111;
											assign node843 = (inp[10]) ? node847 : node844;
												assign node844 = (inp[11]) ? 3'b111 : 3'b101;
												assign node847 = (inp[11]) ? 3'b101 : 3'b111;
								assign node850 = (inp[3]) ? node866 : node851;
									assign node851 = (inp[7]) ? node859 : node852;
										assign node852 = (inp[11]) ? node856 : node853;
											assign node853 = (inp[10]) ? 3'b111 : 3'b101;
											assign node856 = (inp[10]) ? 3'b101 : 3'b111;
										assign node859 = (inp[11]) ? node863 : node860;
											assign node860 = (inp[10]) ? 3'b110 : 3'b101;
											assign node863 = (inp[10]) ? 3'b100 : 3'b110;
									assign node866 = (inp[7]) ? node874 : node867;
										assign node867 = (inp[11]) ? node871 : node868;
											assign node868 = (inp[10]) ? 3'b110 : 3'b101;
											assign node871 = (inp[10]) ? 3'b101 : 3'b111;
										assign node874 = (inp[9]) ? node882 : node875;
											assign node875 = (inp[10]) ? node879 : node876;
												assign node876 = (inp[11]) ? 3'b111 : 3'b101;
												assign node879 = (inp[11]) ? 3'b101 : 3'b111;
											assign node882 = (inp[10]) ? node886 : node883;
												assign node883 = (inp[11]) ? 3'b111 : 3'b101;
												assign node886 = (inp[11]) ? 3'b101 : 3'b111;
						assign node889 = (inp[2]) ? node957 : node890;
							assign node890 = (inp[4]) ? node932 : node891;
								assign node891 = (inp[9]) ? node911 : node892;
									assign node892 = (inp[10]) ? node898 : node893;
										assign node893 = (inp[3]) ? 3'b111 : node894;
											assign node894 = (inp[7]) ? 3'b111 : 3'b101;
										assign node898 = (inp[3]) ? node906 : node899;
											assign node899 = (inp[7]) ? node903 : node900;
												assign node900 = (inp[11]) ? 3'b110 : 3'b111;
												assign node903 = (inp[11]) ? 3'b111 : 3'b100;
											assign node906 = (inp[11]) ? 3'b101 : node907;
												assign node907 = (inp[7]) ? 3'b111 : 3'b100;
									assign node911 = (inp[10]) ? node921 : node912;
										assign node912 = (inp[3]) ? node916 : node913;
											assign node913 = (inp[7]) ? 3'b101 : 3'b100;
											assign node916 = (inp[7]) ? node918 : 3'b110;
												assign node918 = (inp[11]) ? 3'b110 : 3'b101;
										assign node921 = (inp[11]) ? node929 : node922;
											assign node922 = (inp[7]) ? node926 : node923;
												assign node923 = (inp[3]) ? 3'b101 : 3'b110;
												assign node926 = (inp[3]) ? 3'b110 : 3'b101;
											assign node929 = (inp[7]) ? 3'b110 : 3'b111;
								assign node932 = (inp[7]) ? node942 : node933;
									assign node933 = (inp[10]) ? node937 : node934;
										assign node934 = (inp[11]) ? 3'b111 : 3'b101;
										assign node937 = (inp[11]) ? 3'b101 : node938;
											assign node938 = (inp[3]) ? 3'b110 : 3'b111;
									assign node942 = (inp[3]) ? node950 : node943;
										assign node943 = (inp[10]) ? node947 : node944;
											assign node944 = (inp[11]) ? 3'b110 : 3'b101;
											assign node947 = (inp[11]) ? 3'b100 : 3'b110;
										assign node950 = (inp[10]) ? node954 : node951;
											assign node951 = (inp[11]) ? 3'b111 : 3'b101;
											assign node954 = (inp[11]) ? 3'b101 : 3'b111;
							assign node957 = (inp[9]) ? node1003 : node958;
								assign node958 = (inp[4]) ? node984 : node959;
									assign node959 = (inp[10]) ? node969 : node960;
										assign node960 = (inp[3]) ? node964 : node961;
											assign node961 = (inp[7]) ? 3'b111 : 3'b101;
											assign node964 = (inp[11]) ? 3'b111 : node965;
												assign node965 = (inp[7]) ? 3'b101 : 3'b111;
										assign node969 = (inp[3]) ? node977 : node970;
											assign node970 = (inp[11]) ? node974 : node971;
												assign node971 = (inp[7]) ? 3'b100 : 3'b110;
												assign node974 = (inp[7]) ? 3'b110 : 3'b111;
											assign node977 = (inp[7]) ? node981 : node978;
												assign node978 = (inp[11]) ? 3'b101 : 3'b100;
												assign node981 = (inp[11]) ? 3'b101 : 3'b111;
									assign node984 = (inp[10]) ? node992 : node985;
										assign node985 = (inp[11]) ? node987 : 3'b100;
											assign node987 = (inp[7]) ? node989 : 3'b110;
												assign node989 = (inp[3]) ? 3'b110 : 3'b111;
										assign node992 = (inp[11]) ? node1000 : node993;
											assign node993 = (inp[7]) ? node997 : node994;
												assign node994 = (inp[3]) ? 3'b111 : 3'b110;
												assign node997 = (inp[3]) ? 3'b110 : 3'b111;
											assign node1000 = (inp[3]) ? 3'b100 : 3'b101;
								assign node1003 = (inp[3]) ? node1029 : node1004;
									assign node1004 = (inp[7]) ? node1018 : node1005;
										assign node1005 = (inp[10]) ? node1011 : node1006;
											assign node1006 = (inp[11]) ? node1008 : 3'b100;
												assign node1008 = (inp[4]) ? 3'b110 : 3'b100;
											assign node1011 = (inp[4]) ? node1015 : node1012;
												assign node1012 = (inp[11]) ? 3'b110 : 3'b111;
												assign node1015 = (inp[11]) ? 3'b100 : 3'b110;
										assign node1018 = (inp[10]) ? node1024 : node1019;
											assign node1019 = (inp[11]) ? node1021 : 3'b100;
												assign node1021 = (inp[4]) ? 3'b111 : 3'b101;
											assign node1024 = (inp[4]) ? 3'b111 : node1025;
												assign node1025 = (inp[11]) ? 3'b111 : 3'b101;
									assign node1029 = (inp[10]) ? node1037 : node1030;
										assign node1030 = (inp[11]) ? 3'b110 : node1031;
											assign node1031 = (inp[7]) ? 3'b100 : node1032;
												assign node1032 = (inp[4]) ? 3'b100 : 3'b110;
										assign node1037 = (inp[11]) ? 3'b100 : node1038;
											assign node1038 = (inp[7]) ? 3'b110 : node1039;
												assign node1039 = (inp[4]) ? 3'b111 : 3'b101;
					assign node1044 = (inp[0]) ? node1186 : node1045;
						assign node1045 = (inp[2]) ? node1113 : node1046;
							assign node1046 = (inp[4]) ? node1092 : node1047;
								assign node1047 = (inp[9]) ? node1069 : node1048;
									assign node1048 = (inp[10]) ? node1058 : node1049;
										assign node1049 = (inp[3]) ? node1053 : node1050;
											assign node1050 = (inp[7]) ? 3'b111 : 3'b101;
											assign node1053 = (inp[7]) ? node1055 : 3'b111;
												assign node1055 = (inp[11]) ? 3'b111 : 3'b101;
										assign node1058 = (inp[3]) ? node1064 : node1059;
											assign node1059 = (inp[11]) ? node1061 : 3'b110;
												assign node1061 = (inp[7]) ? 3'b110 : 3'b111;
											assign node1064 = (inp[11]) ? 3'b101 : node1065;
												assign node1065 = (inp[7]) ? 3'b111 : 3'b100;
									assign node1069 = (inp[7]) ? node1079 : node1070;
										assign node1070 = (inp[10]) ? node1074 : node1071;
											assign node1071 = (inp[3]) ? 3'b110 : 3'b100;
											assign node1074 = (inp[3]) ? node1076 : 3'b110;
												assign node1076 = (inp[11]) ? 3'b100 : 3'b101;
										assign node1079 = (inp[3]) ? node1087 : node1080;
											assign node1080 = (inp[11]) ? node1084 : node1081;
												assign node1081 = (inp[10]) ? 3'b101 : 3'b110;
												assign node1084 = (inp[10]) ? 3'b111 : 3'b101;
											assign node1087 = (inp[11]) ? 3'b100 : node1088;
												assign node1088 = (inp[10]) ? 3'b110 : 3'b100;
								assign node1092 = (inp[10]) ? node1106 : node1093;
									assign node1093 = (inp[11]) ? node1101 : node1094;
										assign node1094 = (inp[7]) ? node1098 : node1095;
											assign node1095 = (inp[3]) ? 3'b100 : 3'b101;
											assign node1098 = (inp[3]) ? 3'b101 : 3'b100;
										assign node1101 = (inp[7]) ? 3'b110 : node1102;
											assign node1102 = (inp[3]) ? 3'b110 : 3'b111;
									assign node1106 = (inp[11]) ? node1108 : 3'b110;
										assign node1108 = (inp[7]) ? 3'b100 : node1109;
											assign node1109 = (inp[3]) ? 3'b100 : 3'b101;
							assign node1113 = (inp[4]) ? node1161 : node1114;
								assign node1114 = (inp[9]) ? node1136 : node1115;
									assign node1115 = (inp[3]) ? node1129 : node1116;
										assign node1116 = (inp[10]) ? node1122 : node1117;
											assign node1117 = (inp[11]) ? 3'b101 : node1118;
												assign node1118 = (inp[7]) ? 3'b110 : 3'b100;
											assign node1122 = (inp[7]) ? node1126 : node1123;
												assign node1123 = (inp[11]) ? 3'b111 : 3'b110;
												assign node1126 = (inp[11]) ? 3'b110 : 3'b101;
										assign node1129 = (inp[10]) ? node1131 : 3'b110;
											assign node1131 = (inp[11]) ? 3'b100 : node1132;
												assign node1132 = (inp[7]) ? 3'b110 : 3'b101;
									assign node1136 = (inp[7]) ? node1148 : node1137;
										assign node1137 = (inp[10]) ? node1141 : node1138;
											assign node1138 = (inp[3]) ? 3'b111 : 3'b101;
											assign node1141 = (inp[3]) ? node1145 : node1142;
												assign node1142 = (inp[11]) ? 3'b110 : 3'b111;
												assign node1145 = (inp[11]) ? 3'b101 : 3'b100;
										assign node1148 = (inp[10]) ? node1154 : node1149;
											assign node1149 = (inp[3]) ? 3'b100 : node1150;
												assign node1150 = (inp[11]) ? 3'b100 : 3'b111;
											assign node1154 = (inp[11]) ? node1158 : node1155;
												assign node1155 = (inp[3]) ? 3'b111 : 3'b100;
												assign node1158 = (inp[3]) ? 3'b101 : 3'b111;
								assign node1161 = (inp[3]) ? node1177 : node1162;
									assign node1162 = (inp[7]) ? node1170 : node1163;
										assign node1163 = (inp[10]) ? node1167 : node1164;
											assign node1164 = (inp[11]) ? 3'b110 : 3'b100;
											assign node1167 = (inp[11]) ? 3'b100 : 3'b111;
										assign node1170 = (inp[10]) ? node1174 : node1171;
											assign node1171 = (inp[11]) ? 3'b111 : 3'b101;
											assign node1174 = (inp[11]) ? 3'b101 : 3'b111;
									assign node1177 = (inp[11]) ? node1183 : node1178;
										assign node1178 = (inp[10]) ? 3'b111 : node1179;
											assign node1179 = (inp[7]) ? 3'b100 : 3'b101;
										assign node1183 = (inp[10]) ? 3'b101 : 3'b111;
						assign node1186 = (inp[2]) ? node1270 : node1187;
							assign node1187 = (inp[4]) ? node1239 : node1188;
								assign node1188 = (inp[9]) ? node1216 : node1189;
									assign node1189 = (inp[3]) ? node1205 : node1190;
										assign node1190 = (inp[10]) ? node1198 : node1191;
											assign node1191 = (inp[11]) ? node1195 : node1192;
												assign node1192 = (inp[7]) ? 3'b110 : 3'b100;
												assign node1195 = (inp[7]) ? 3'b101 : 3'b100;
											assign node1198 = (inp[11]) ? node1202 : node1199;
												assign node1199 = (inp[7]) ? 3'b101 : 3'b111;
												assign node1202 = (inp[7]) ? 3'b111 : 3'b110;
										assign node1205 = (inp[10]) ? node1211 : node1206;
											assign node1206 = (inp[7]) ? node1208 : 3'b110;
												assign node1208 = (inp[11]) ? 3'b110 : 3'b100;
											assign node1211 = (inp[11]) ? 3'b100 : node1212;
												assign node1212 = (inp[7]) ? 3'b110 : 3'b101;
									assign node1216 = (inp[10]) ? node1228 : node1217;
										assign node1217 = (inp[3]) ? node1223 : node1218;
											assign node1218 = (inp[11]) ? node1220 : 3'b111;
												assign node1220 = (inp[7]) ? 3'b100 : 3'b101;
											assign node1223 = (inp[7]) ? node1225 : 3'b111;
												assign node1225 = (inp[11]) ? 3'b111 : 3'b101;
										assign node1228 = (inp[3]) ? node1236 : node1229;
											assign node1229 = (inp[11]) ? node1233 : node1230;
												assign node1230 = (inp[7]) ? 3'b100 : 3'b110;
												assign node1233 = (inp[7]) ? 3'b110 : 3'b111;
											assign node1236 = (inp[11]) ? 3'b101 : 3'b100;
								assign node1239 = (inp[7]) ? node1255 : node1240;
									assign node1240 = (inp[3]) ? node1248 : node1241;
										assign node1241 = (inp[11]) ? node1245 : node1242;
											assign node1242 = (inp[10]) ? 3'b111 : 3'b100;
											assign node1245 = (inp[10]) ? 3'b100 : 3'b110;
										assign node1248 = (inp[11]) ? node1252 : node1249;
											assign node1249 = (inp[10]) ? 3'b111 : 3'b101;
											assign node1252 = (inp[10]) ? 3'b101 : 3'b111;
									assign node1255 = (inp[3]) ? node1263 : node1256;
										assign node1256 = (inp[10]) ? node1260 : node1257;
											assign node1257 = (inp[11]) ? 3'b111 : 3'b101;
											assign node1260 = (inp[11]) ? 3'b101 : 3'b111;
										assign node1263 = (inp[10]) ? node1267 : node1264;
											assign node1264 = (inp[11]) ? 3'b111 : 3'b100;
											assign node1267 = (inp[11]) ? 3'b101 : 3'b111;
							assign node1270 = (inp[4]) ? node1322 : node1271;
								assign node1271 = (inp[9]) ? node1297 : node1272;
									assign node1272 = (inp[10]) ? node1286 : node1273;
										assign node1273 = (inp[3]) ? node1281 : node1274;
											assign node1274 = (inp[11]) ? node1278 : node1275;
												assign node1275 = (inp[7]) ? 3'b111 : 3'b101;
												assign node1278 = (inp[7]) ? 3'b100 : 3'b101;
											assign node1281 = (inp[11]) ? 3'b111 : node1282;
												assign node1282 = (inp[7]) ? 3'b100 : 3'b111;
										assign node1286 = (inp[3]) ? node1294 : node1287;
											assign node1287 = (inp[11]) ? node1291 : node1288;
												assign node1288 = (inp[7]) ? 3'b100 : 3'b111;
												assign node1291 = (inp[7]) ? 3'b111 : 3'b110;
											assign node1294 = (inp[11]) ? 3'b101 : 3'b100;
									assign node1297 = (inp[10]) ? node1309 : node1298;
										assign node1298 = (inp[7]) ? node1302 : node1299;
											assign node1299 = (inp[3]) ? 3'b110 : 3'b100;
											assign node1302 = (inp[3]) ? node1306 : node1303;
												assign node1303 = (inp[11]) ? 3'b101 : 3'b110;
												assign node1306 = (inp[11]) ? 3'b110 : 3'b101;
										assign node1309 = (inp[3]) ? node1317 : node1310;
											assign node1310 = (inp[7]) ? node1314 : node1311;
												assign node1311 = (inp[11]) ? 3'b111 : 3'b110;
												assign node1314 = (inp[11]) ? 3'b110 : 3'b101;
											assign node1317 = (inp[11]) ? 3'b100 : node1318;
												assign node1318 = (inp[7]) ? 3'b110 : 3'b101;
								assign node1322 = (inp[10]) ? node1336 : node1323;
									assign node1323 = (inp[11]) ? node1331 : node1324;
										assign node1324 = (inp[7]) ? node1328 : node1325;
											assign node1325 = (inp[3]) ? 3'b100 : 3'b101;
											assign node1328 = (inp[3]) ? 3'b101 : 3'b100;
										assign node1331 = (inp[3]) ? 3'b110 : node1332;
											assign node1332 = (inp[7]) ? 3'b110 : 3'b111;
									assign node1336 = (inp[11]) ? 3'b100 : 3'b110;
			assign node1339 = (inp[4]) ? node1705 : node1340;
				assign node1340 = (inp[6]) ? node1540 : node1341;
					assign node1341 = (inp[1]) ? node1433 : node1342;
						assign node1342 = (inp[9]) ? node1390 : node1343;
							assign node1343 = (inp[10]) ? node1359 : node1344;
								assign node1344 = (inp[7]) ? node1348 : node1345;
									assign node1345 = (inp[3]) ? 3'b110 : 3'b100;
									assign node1348 = (inp[3]) ? node1354 : node1349;
										assign node1349 = (inp[11]) ? node1351 : 3'b110;
											assign node1351 = (inp[2]) ? 3'b111 : 3'b110;
										assign node1354 = (inp[11]) ? 3'b100 : node1355;
											assign node1355 = (inp[2]) ? 3'b100 : 3'b101;
								assign node1359 = (inp[7]) ? node1383 : node1360;
									assign node1360 = (inp[3]) ? node1368 : node1361;
										assign node1361 = (inp[2]) ? node1365 : node1362;
											assign node1362 = (inp[11]) ? 3'b101 : 3'b100;
											assign node1365 = (inp[11]) ? 3'b100 : 3'b101;
										assign node1368 = (inp[0]) ? node1376 : node1369;
											assign node1369 = (inp[2]) ? node1373 : node1370;
												assign node1370 = (inp[11]) ? 3'b111 : 3'b110;
												assign node1373 = (inp[11]) ? 3'b110 : 3'b111;
											assign node1376 = (inp[11]) ? node1380 : node1377;
												assign node1377 = (inp[2]) ? 3'b111 : 3'b110;
												assign node1380 = (inp[2]) ? 3'b110 : 3'b111;
									assign node1383 = (inp[3]) ? 3'b100 : node1384;
										assign node1384 = (inp[11]) ? 3'b110 : node1385;
											assign node1385 = (inp[2]) ? 3'b111 : 3'b110;
							assign node1390 = (inp[10]) ? node1406 : node1391;
								assign node1391 = (inp[7]) ? node1395 : node1392;
									assign node1392 = (inp[3]) ? 3'b111 : 3'b101;
									assign node1395 = (inp[3]) ? node1401 : node1396;
										assign node1396 = (inp[2]) ? node1398 : 3'b111;
											assign node1398 = (inp[11]) ? 3'b110 : 3'b111;
										assign node1401 = (inp[11]) ? 3'b101 : node1402;
											assign node1402 = (inp[2]) ? 3'b101 : 3'b100;
								assign node1406 = (inp[7]) ? node1422 : node1407;
									assign node1407 = (inp[3]) ? node1415 : node1408;
										assign node1408 = (inp[11]) ? node1412 : node1409;
											assign node1409 = (inp[2]) ? 3'b100 : 3'b101;
											assign node1412 = (inp[2]) ? 3'b101 : 3'b100;
										assign node1415 = (inp[11]) ? node1419 : node1416;
											assign node1416 = (inp[2]) ? 3'b110 : 3'b111;
											assign node1419 = (inp[2]) ? 3'b111 : 3'b110;
									assign node1422 = (inp[3]) ? node1428 : node1423;
										assign node1423 = (inp[11]) ? 3'b111 : node1424;
											assign node1424 = (inp[2]) ? 3'b110 : 3'b111;
										assign node1428 = (inp[2]) ? 3'b101 : node1429;
											assign node1429 = (inp[11]) ? 3'b100 : 3'b101;
						assign node1433 = (inp[9]) ? node1485 : node1434;
							assign node1434 = (inp[10]) ? node1450 : node1435;
								assign node1435 = (inp[7]) ? node1439 : node1436;
									assign node1436 = (inp[3]) ? 3'b111 : 3'b101;
									assign node1439 = (inp[3]) ? node1445 : node1440;
										assign node1440 = (inp[11]) ? node1442 : 3'b111;
											assign node1442 = (inp[2]) ? 3'b110 : 3'b111;
										assign node1445 = (inp[2]) ? 3'b101 : node1446;
											assign node1446 = (inp[11]) ? 3'b101 : 3'b100;
								assign node1450 = (inp[7]) ? node1474 : node1451;
									assign node1451 = (inp[3]) ? node1459 : node1452;
										assign node1452 = (inp[11]) ? node1456 : node1453;
											assign node1453 = (inp[2]) ? 3'b100 : 3'b101;
											assign node1456 = (inp[2]) ? 3'b101 : 3'b100;
										assign node1459 = (inp[0]) ? node1467 : node1460;
											assign node1460 = (inp[2]) ? node1464 : node1461;
												assign node1461 = (inp[11]) ? 3'b110 : 3'b111;
												assign node1464 = (inp[11]) ? 3'b111 : 3'b110;
											assign node1467 = (inp[2]) ? node1471 : node1468;
												assign node1468 = (inp[11]) ? 3'b110 : 3'b111;
												assign node1471 = (inp[11]) ? 3'b111 : 3'b110;
									assign node1474 = (inp[3]) ? node1480 : node1475;
										assign node1475 = (inp[2]) ? node1477 : 3'b111;
											assign node1477 = (inp[11]) ? 3'b111 : 3'b110;
										assign node1480 = (inp[2]) ? 3'b101 : node1481;
											assign node1481 = (inp[11]) ? 3'b100 : 3'b101;
							assign node1485 = (inp[10]) ? node1499 : node1486;
								assign node1486 = (inp[7]) ? node1490 : node1487;
									assign node1487 = (inp[3]) ? 3'b110 : 3'b100;
									assign node1490 = (inp[3]) ? node1494 : node1491;
										assign node1491 = (inp[11]) ? 3'b111 : 3'b110;
										assign node1494 = (inp[2]) ? 3'b100 : node1495;
											assign node1495 = (inp[11]) ? 3'b100 : 3'b101;
								assign node1499 = (inp[7]) ? node1529 : node1500;
									assign node1500 = (inp[3]) ? node1516 : node1501;
										assign node1501 = (inp[0]) ? node1509 : node1502;
											assign node1502 = (inp[11]) ? node1506 : node1503;
												assign node1503 = (inp[2]) ? 3'b101 : 3'b100;
												assign node1506 = (inp[2]) ? 3'b100 : 3'b101;
											assign node1509 = (inp[2]) ? node1513 : node1510;
												assign node1510 = (inp[11]) ? 3'b101 : 3'b100;
												assign node1513 = (inp[11]) ? 3'b100 : 3'b101;
										assign node1516 = (inp[0]) ? node1522 : node1517;
											assign node1517 = (inp[2]) ? 3'b111 : node1518;
												assign node1518 = (inp[11]) ? 3'b111 : 3'b110;
											assign node1522 = (inp[11]) ? node1526 : node1523;
												assign node1523 = (inp[2]) ? 3'b111 : 3'b110;
												assign node1526 = (inp[2]) ? 3'b110 : 3'b111;
									assign node1529 = (inp[3]) ? node1535 : node1530;
										assign node1530 = (inp[11]) ? 3'b110 : node1531;
											assign node1531 = (inp[2]) ? 3'b111 : 3'b110;
										assign node1535 = (inp[11]) ? node1537 : 3'b100;
											assign node1537 = (inp[2]) ? 3'b100 : 3'b101;
					assign node1540 = (inp[11]) ? node1650 : node1541;
						assign node1541 = (inp[3]) ? node1589 : node1542;
							assign node1542 = (inp[2]) ? node1574 : node1543;
								assign node1543 = (inp[7]) ? node1567 : node1544;
									assign node1544 = (inp[1]) ? node1552 : node1545;
										assign node1545 = (inp[10]) ? node1549 : node1546;
											assign node1546 = (inp[9]) ? 3'b001 : 3'b000;
											assign node1549 = (inp[9]) ? 3'b000 : 3'b001;
										assign node1552 = (inp[0]) ? node1560 : node1553;
											assign node1553 = (inp[10]) ? node1557 : node1554;
												assign node1554 = (inp[9]) ? 3'b001 : 3'b000;
												assign node1557 = (inp[9]) ? 3'b000 : 3'b001;
											assign node1560 = (inp[9]) ? node1564 : node1561;
												assign node1561 = (inp[10]) ? 3'b001 : 3'b000;
												assign node1564 = (inp[10]) ? 3'b000 : 3'b001;
									assign node1567 = (inp[10]) ? node1571 : node1568;
										assign node1568 = (inp[9]) ? 3'b001 : 3'b000;
										assign node1571 = (inp[9]) ? 3'b000 : 3'b001;
								assign node1574 = (inp[9]) ? node1582 : node1575;
									assign node1575 = (inp[10]) ? node1579 : node1576;
										assign node1576 = (inp[7]) ? 3'b001 : 3'b000;
										assign node1579 = (inp[7]) ? 3'b000 : 3'b001;
									assign node1582 = (inp[7]) ? node1586 : node1583;
										assign node1583 = (inp[10]) ? 3'b000 : 3'b001;
										assign node1586 = (inp[10]) ? 3'b001 : 3'b000;
							assign node1589 = (inp[7]) ? node1597 : node1590;
								assign node1590 = (inp[9]) ? node1594 : node1591;
									assign node1591 = (inp[10]) ? 3'b011 : 3'b010;
									assign node1594 = (inp[10]) ? 3'b010 : 3'b011;
								assign node1597 = (inp[1]) ? node1621 : node1598;
									assign node1598 = (inp[9]) ? node1614 : node1599;
										assign node1599 = (inp[0]) ? node1607 : node1600;
											assign node1600 = (inp[10]) ? node1604 : node1601;
												assign node1601 = (inp[2]) ? 3'b010 : 3'b011;
												assign node1604 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1607 = (inp[2]) ? node1611 : node1608;
												assign node1608 = (inp[10]) ? 3'b010 : 3'b011;
												assign node1611 = (inp[10]) ? 3'b011 : 3'b010;
										assign node1614 = (inp[2]) ? node1618 : node1615;
											assign node1615 = (inp[10]) ? 3'b011 : 3'b010;
											assign node1618 = (inp[10]) ? 3'b010 : 3'b011;
									assign node1621 = (inp[9]) ? node1635 : node1622;
										assign node1622 = (inp[0]) ? node1630 : node1623;
											assign node1623 = (inp[10]) ? node1627 : node1624;
												assign node1624 = (inp[2]) ? 3'b010 : 3'b011;
												assign node1627 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1630 = (inp[10]) ? 3'b010 : node1631;
												assign node1631 = (inp[2]) ? 3'b010 : 3'b011;
										assign node1635 = (inp[0]) ? node1643 : node1636;
											assign node1636 = (inp[10]) ? node1640 : node1637;
												assign node1637 = (inp[2]) ? 3'b011 : 3'b010;
												assign node1640 = (inp[2]) ? 3'b010 : 3'b011;
											assign node1643 = (inp[10]) ? node1647 : node1644;
												assign node1644 = (inp[2]) ? 3'b011 : 3'b010;
												assign node1647 = (inp[2]) ? 3'b010 : 3'b011;
						assign node1650 = (inp[3]) ? node1698 : node1651;
							assign node1651 = (inp[10]) ? node1683 : node1652;
								assign node1652 = (inp[0]) ? node1668 : node1653;
									assign node1653 = (inp[1]) ? node1661 : node1654;
										assign node1654 = (inp[9]) ? node1658 : node1655;
											assign node1655 = (inp[7]) ? 3'b011 : 3'b010;
											assign node1658 = (inp[7]) ? 3'b010 : 3'b011;
										assign node1661 = (inp[9]) ? node1665 : node1662;
											assign node1662 = (inp[7]) ? 3'b011 : 3'b010;
											assign node1665 = (inp[7]) ? 3'b010 : 3'b011;
									assign node1668 = (inp[2]) ? node1676 : node1669;
										assign node1669 = (inp[9]) ? node1673 : node1670;
											assign node1670 = (inp[7]) ? 3'b011 : 3'b010;
											assign node1673 = (inp[7]) ? 3'b010 : 3'b011;
										assign node1676 = (inp[9]) ? node1680 : node1677;
											assign node1677 = (inp[7]) ? 3'b011 : 3'b010;
											assign node1680 = (inp[7]) ? 3'b010 : 3'b011;
								assign node1683 = (inp[2]) ? node1691 : node1684;
									assign node1684 = (inp[9]) ? node1688 : node1685;
										assign node1685 = (inp[7]) ? 3'b011 : 3'b010;
										assign node1688 = (inp[7]) ? 3'b010 : 3'b011;
									assign node1691 = (inp[7]) ? node1695 : node1692;
										assign node1692 = (inp[9]) ? 3'b011 : 3'b010;
										assign node1695 = (inp[9]) ? 3'b010 : 3'b011;
							assign node1698 = (inp[9]) ? node1702 : node1699;
								assign node1699 = (inp[2]) ? 3'b001 : 3'b000;
								assign node1702 = (inp[2]) ? 3'b000 : 3'b001;
				assign node1705 = (inp[11]) ? node1893 : node1706;
					assign node1706 = (inp[7]) ? node1814 : node1707;
						assign node1707 = (inp[6]) ? node1731 : node1708;
							assign node1708 = (inp[1]) ? node1720 : node1709;
								assign node1709 = (inp[2]) ? node1715 : node1710;
									assign node1710 = (inp[10]) ? node1712 : 3'b000;
										assign node1712 = (inp[3]) ? 3'b001 : 3'b000;
									assign node1715 = (inp[3]) ? node1717 : 3'b001;
										assign node1717 = (inp[10]) ? 3'b000 : 3'b001;
								assign node1720 = (inp[2]) ? node1726 : node1721;
									assign node1721 = (inp[3]) ? node1723 : 3'b001;
										assign node1723 = (inp[10]) ? 3'b000 : 3'b001;
									assign node1726 = (inp[3]) ? node1728 : 3'b000;
										assign node1728 = (inp[10]) ? 3'b001 : 3'b000;
							assign node1731 = (inp[1]) ? node1779 : node1732;
								assign node1732 = (inp[9]) ? node1762 : node1733;
									assign node1733 = (inp[0]) ? node1747 : node1734;
										assign node1734 = (inp[3]) ? node1742 : node1735;
											assign node1735 = (inp[2]) ? node1739 : node1736;
												assign node1736 = (inp[10]) ? 3'b011 : 3'b010;
												assign node1739 = (inp[10]) ? 3'b010 : 3'b011;
											assign node1742 = (inp[10]) ? node1744 : 3'b010;
												assign node1744 = (inp[2]) ? 3'b010 : 3'b011;
										assign node1747 = (inp[3]) ? node1755 : node1748;
											assign node1748 = (inp[2]) ? node1752 : node1749;
												assign node1749 = (inp[10]) ? 3'b011 : 3'b010;
												assign node1752 = (inp[10]) ? 3'b010 : 3'b011;
											assign node1755 = (inp[2]) ? node1759 : node1756;
												assign node1756 = (inp[10]) ? 3'b011 : 3'b010;
												assign node1759 = (inp[10]) ? 3'b010 : 3'b011;
									assign node1762 = (inp[0]) ? node1770 : node1763;
										assign node1763 = (inp[10]) ? node1767 : node1764;
											assign node1764 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1767 = (inp[2]) ? 3'b010 : 3'b011;
										assign node1770 = (inp[3]) ? node1772 : 3'b010;
											assign node1772 = (inp[10]) ? node1776 : node1773;
												assign node1773 = (inp[2]) ? 3'b011 : 3'b010;
												assign node1776 = (inp[2]) ? 3'b010 : 3'b011;
								assign node1779 = (inp[3]) ? node1799 : node1780;
									assign node1780 = (inp[0]) ? node1788 : node1781;
										assign node1781 = (inp[10]) ? node1785 : node1782;
											assign node1782 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1785 = (inp[2]) ? 3'b010 : 3'b011;
										assign node1788 = (inp[9]) ? node1794 : node1789;
											assign node1789 = (inp[2]) ? node1791 : 3'b011;
												assign node1791 = (inp[10]) ? 3'b010 : 3'b011;
											assign node1794 = (inp[2]) ? 3'b011 : node1795;
												assign node1795 = (inp[10]) ? 3'b011 : 3'b010;
									assign node1799 = (inp[0]) ? node1807 : node1800;
										assign node1800 = (inp[10]) ? node1804 : node1801;
											assign node1801 = (inp[2]) ? 3'b011 : 3'b010;
											assign node1804 = (inp[2]) ? 3'b010 : 3'b011;
										assign node1807 = (inp[2]) ? node1811 : node1808;
											assign node1808 = (inp[10]) ? 3'b011 : 3'b010;
											assign node1811 = (inp[10]) ? 3'b010 : 3'b011;
						assign node1814 = (inp[0]) ? node1854 : node1815;
							assign node1815 = (inp[1]) ? node1839 : node1816;
								assign node1816 = (inp[2]) ? node1826 : node1817;
									assign node1817 = (inp[6]) ? node1823 : node1818;
										assign node1818 = (inp[3]) ? node1820 : 3'b010;
											assign node1820 = (inp[10]) ? 3'b010 : 3'b011;
										assign node1823 = (inp[10]) ? 3'b011 : 3'b010;
									assign node1826 = (inp[3]) ? node1832 : node1827;
										assign node1827 = (inp[10]) ? node1829 : 3'b011;
											assign node1829 = (inp[6]) ? 3'b010 : 3'b011;
										assign node1832 = (inp[6]) ? node1836 : node1833;
											assign node1833 = (inp[10]) ? 3'b011 : 3'b010;
											assign node1836 = (inp[10]) ? 3'b010 : 3'b011;
								assign node1839 = (inp[2]) ? node1847 : node1840;
									assign node1840 = (inp[10]) ? 3'b011 : node1841;
										assign node1841 = (inp[6]) ? 3'b010 : node1842;
											assign node1842 = (inp[3]) ? 3'b010 : 3'b011;
									assign node1847 = (inp[10]) ? 3'b010 : node1848;
										assign node1848 = (inp[6]) ? 3'b011 : node1849;
											assign node1849 = (inp[3]) ? 3'b011 : 3'b010;
							assign node1854 = (inp[2]) ? node1878 : node1855;
								assign node1855 = (inp[10]) ? node1873 : node1856;
									assign node1856 = (inp[6]) ? 3'b010 : node1857;
										assign node1857 = (inp[9]) ? node1865 : node1858;
											assign node1858 = (inp[1]) ? node1862 : node1859;
												assign node1859 = (inp[3]) ? 3'b011 : 3'b010;
												assign node1862 = (inp[3]) ? 3'b010 : 3'b011;
											assign node1865 = (inp[3]) ? node1869 : node1866;
												assign node1866 = (inp[1]) ? 3'b011 : 3'b010;
												assign node1869 = (inp[1]) ? 3'b010 : 3'b011;
									assign node1873 = (inp[6]) ? 3'b011 : node1874;
										assign node1874 = (inp[1]) ? 3'b011 : 3'b010;
								assign node1878 = (inp[10]) ? node1888 : node1879;
									assign node1879 = (inp[6]) ? 3'b011 : node1880;
										assign node1880 = (inp[3]) ? node1884 : node1881;
											assign node1881 = (inp[1]) ? 3'b010 : 3'b011;
											assign node1884 = (inp[1]) ? 3'b011 : 3'b010;
									assign node1888 = (inp[1]) ? 3'b010 : node1889;
										assign node1889 = (inp[6]) ? 3'b010 : 3'b011;
					assign node1893 = (inp[6]) ? node2003 : node1894;
						assign node1894 = (inp[7]) ? node1942 : node1895;
							assign node1895 = (inp[0]) ? node1919 : node1896;
								assign node1896 = (inp[2]) ? node1908 : node1897;
									assign node1897 = (inp[1]) ? node1903 : node1898;
										assign node1898 = (inp[10]) ? node1900 : 3'b010;
											assign node1900 = (inp[3]) ? 3'b010 : 3'b011;
										assign node1903 = (inp[3]) ? 3'b011 : node1904;
											assign node1904 = (inp[10]) ? 3'b010 : 3'b011;
									assign node1908 = (inp[1]) ? node1914 : node1909;
										assign node1909 = (inp[10]) ? node1911 : 3'b011;
											assign node1911 = (inp[3]) ? 3'b011 : 3'b010;
										assign node1914 = (inp[10]) ? node1916 : 3'b010;
											assign node1916 = (inp[3]) ? 3'b010 : 3'b011;
								assign node1919 = (inp[1]) ? node1931 : node1920;
									assign node1920 = (inp[2]) ? node1926 : node1921;
										assign node1921 = (inp[10]) ? node1923 : 3'b010;
											assign node1923 = (inp[3]) ? 3'b010 : 3'b011;
										assign node1926 = (inp[10]) ? node1928 : 3'b011;
											assign node1928 = (inp[3]) ? 3'b011 : 3'b010;
									assign node1931 = (inp[2]) ? node1937 : node1932;
										assign node1932 = (inp[3]) ? 3'b011 : node1933;
											assign node1933 = (inp[10]) ? 3'b010 : 3'b011;
										assign node1937 = (inp[10]) ? node1939 : 3'b010;
											assign node1939 = (inp[3]) ? 3'b010 : 3'b011;
							assign node1942 = (inp[10]) ? node1988 : node1943;
								assign node1943 = (inp[9]) ? node1969 : node1944;
									assign node1944 = (inp[1]) ? node1954 : node1945;
										assign node1945 = (inp[0]) ? 3'b000 : node1946;
											assign node1946 = (inp[3]) ? node1950 : node1947;
												assign node1947 = (inp[2]) ? 3'b000 : 3'b001;
												assign node1950 = (inp[2]) ? 3'b001 : 3'b000;
										assign node1954 = (inp[0]) ? node1962 : node1955;
											assign node1955 = (inp[2]) ? node1959 : node1956;
												assign node1956 = (inp[3]) ? 3'b001 : 3'b000;
												assign node1959 = (inp[3]) ? 3'b000 : 3'b001;
											assign node1962 = (inp[2]) ? node1966 : node1963;
												assign node1963 = (inp[3]) ? 3'b001 : 3'b000;
												assign node1966 = (inp[3]) ? 3'b000 : 3'b001;
									assign node1969 = (inp[1]) ? node1975 : node1970;
										assign node1970 = (inp[3]) ? node1972 : 3'b001;
											assign node1972 = (inp[2]) ? 3'b001 : 3'b000;
										assign node1975 = (inp[0]) ? node1981 : node1976;
											assign node1976 = (inp[2]) ? 3'b000 : node1977;
												assign node1977 = (inp[3]) ? 3'b001 : 3'b000;
											assign node1981 = (inp[3]) ? node1985 : node1982;
												assign node1982 = (inp[2]) ? 3'b001 : 3'b000;
												assign node1985 = (inp[2]) ? 3'b000 : 3'b001;
								assign node1988 = (inp[3]) ? node1996 : node1989;
									assign node1989 = (inp[2]) ? node1993 : node1990;
										assign node1990 = (inp[1]) ? 3'b001 : 3'b000;
										assign node1993 = (inp[1]) ? 3'b000 : 3'b001;
									assign node1996 = (inp[2]) ? node2000 : node1997;
										assign node1997 = (inp[1]) ? 3'b001 : 3'b000;
										assign node2000 = (inp[1]) ? 3'b000 : 3'b001;
						assign node2003 = (inp[2]) ? node2009 : node2004;
							assign node2004 = (inp[7]) ? 3'b001 : node2005;
								assign node2005 = (inp[3]) ? 3'b001 : 3'b000;
							assign node2009 = (inp[3]) ? 3'b000 : node2010;
								assign node2010 = (inp[7]) ? 3'b000 : 3'b001;
		assign node2014 = (inp[4]) ? node2942 : node2015;
			assign node2015 = (inp[6]) ? node2543 : node2016;
				assign node2016 = (inp[1]) ? node2310 : node2017;
					assign node2017 = (inp[9]) ? node2167 : node2018;
						assign node2018 = (inp[8]) ? node2122 : node2019;
							assign node2019 = (inp[3]) ? node2071 : node2020;
								assign node2020 = (inp[10]) ? node2052 : node2021;
									assign node2021 = (inp[7]) ? node2037 : node2022;
										assign node2022 = (inp[11]) ? node2030 : node2023;
											assign node2023 = (inp[2]) ? node2027 : node2024;
												assign node2024 = (inp[0]) ? 3'b101 : 3'b100;
												assign node2027 = (inp[0]) ? 3'b100 : 3'b101;
											assign node2030 = (inp[2]) ? node2034 : node2031;
												assign node2031 = (inp[0]) ? 3'b111 : 3'b110;
												assign node2034 = (inp[0]) ? 3'b110 : 3'b111;
										assign node2037 = (inp[11]) ? node2045 : node2038;
											assign node2038 = (inp[2]) ? node2042 : node2039;
												assign node2039 = (inp[0]) ? 3'b101 : 3'b100;
												assign node2042 = (inp[0]) ? 3'b100 : 3'b101;
											assign node2045 = (inp[0]) ? node2049 : node2046;
												assign node2046 = (inp[2]) ? 3'b100 : 3'b101;
												assign node2049 = (inp[2]) ? 3'b101 : 3'b100;
									assign node2052 = (inp[7]) ? node2064 : node2053;
										assign node2053 = (inp[11]) ? node2061 : node2054;
											assign node2054 = (inp[2]) ? node2058 : node2055;
												assign node2055 = (inp[0]) ? 3'b111 : 3'b110;
												assign node2058 = (inp[0]) ? 3'b110 : 3'b111;
											assign node2061 = (inp[0]) ? 3'b100 : 3'b101;
										assign node2064 = (inp[0]) ? node2068 : node2065;
											assign node2065 = (inp[2]) ? 3'b111 : 3'b110;
											assign node2068 = (inp[2]) ? 3'b110 : 3'b111;
								assign node2071 = (inp[10]) ? node2097 : node2072;
									assign node2072 = (inp[7]) ? node2084 : node2073;
										assign node2073 = (inp[11]) ? node2077 : node2074;
											assign node2074 = (inp[0]) ? 3'b111 : 3'b110;
											assign node2077 = (inp[2]) ? node2081 : node2078;
												assign node2078 = (inp[0]) ? 3'b100 : 3'b101;
												assign node2081 = (inp[0]) ? 3'b101 : 3'b100;
										assign node2084 = (inp[2]) ? node2090 : node2085;
											assign node2085 = (inp[11]) ? node2087 : 3'b110;
												assign node2087 = (inp[0]) ? 3'b111 : 3'b110;
											assign node2090 = (inp[11]) ? node2094 : node2091;
												assign node2091 = (inp[0]) ? 3'b110 : 3'b111;
												assign node2094 = (inp[0]) ? 3'b111 : 3'b110;
									assign node2097 = (inp[11]) ? node2111 : node2098;
										assign node2098 = (inp[2]) ? node2104 : node2099;
											assign node2099 = (inp[7]) ? 3'b100 : node2100;
												assign node2100 = (inp[0]) ? 3'b100 : 3'b101;
											assign node2104 = (inp[7]) ? node2108 : node2105;
												assign node2105 = (inp[0]) ? 3'b101 : 3'b100;
												assign node2108 = (inp[0]) ? 3'b100 : 3'b101;
										assign node2111 = (inp[7]) ? node2117 : node2112;
											assign node2112 = (inp[0]) ? node2114 : 3'b110;
												assign node2114 = (inp[2]) ? 3'b110 : 3'b111;
											assign node2117 = (inp[0]) ? node2119 : 3'b100;
												assign node2119 = (inp[2]) ? 3'b100 : 3'b101;
							assign node2122 = (inp[10]) ? node2152 : node2123;
								assign node2123 = (inp[7]) ? node2135 : node2124;
									assign node2124 = (inp[3]) ? node2130 : node2125;
										assign node2125 = (inp[2]) ? node2127 : 3'b100;
											assign node2127 = (inp[11]) ? 3'b100 : 3'b101;
										assign node2130 = (inp[2]) ? 3'b110 : node2131;
											assign node2131 = (inp[11]) ? 3'b111 : 3'b110;
									assign node2135 = (inp[3]) ? node2145 : node2136;
										assign node2136 = (inp[0]) ? node2138 : 3'b111;
											assign node2138 = (inp[2]) ? node2142 : node2139;
												assign node2139 = (inp[11]) ? 3'b111 : 3'b110;
												assign node2142 = (inp[11]) ? 3'b110 : 3'b111;
										assign node2145 = (inp[11]) ? node2149 : node2146;
											assign node2146 = (inp[2]) ? 3'b101 : 3'b100;
											assign node2149 = (inp[2]) ? 3'b100 : 3'b101;
								assign node2152 = (inp[7]) ? node2164 : node2153;
									assign node2153 = (inp[3]) ? node2159 : node2154;
										assign node2154 = (inp[11]) ? node2156 : 3'b100;
											assign node2156 = (inp[2]) ? 3'b101 : 3'b100;
										assign node2159 = (inp[2]) ? 3'b110 : node2160;
											assign node2160 = (inp[11]) ? 3'b110 : 3'b111;
									assign node2164 = (inp[3]) ? 3'b100 : 3'b110;
						assign node2167 = (inp[8]) ? node2269 : node2168;
							assign node2168 = (inp[10]) ? node2218 : node2169;
								assign node2169 = (inp[3]) ? node2195 : node2170;
									assign node2170 = (inp[7]) ? node2182 : node2171;
										assign node2171 = (inp[11]) ? node2175 : node2172;
											assign node2172 = (inp[0]) ? 3'b101 : 3'b100;
											assign node2175 = (inp[0]) ? node2179 : node2176;
												assign node2176 = (inp[2]) ? 3'b110 : 3'b111;
												assign node2179 = (inp[2]) ? 3'b111 : 3'b110;
										assign node2182 = (inp[11]) ? node2190 : node2183;
											assign node2183 = (inp[0]) ? node2187 : node2184;
												assign node2184 = (inp[2]) ? 3'b100 : 3'b101;
												assign node2187 = (inp[2]) ? 3'b101 : 3'b100;
											assign node2190 = (inp[2]) ? node2192 : 3'b100;
												assign node2192 = (inp[0]) ? 3'b100 : 3'b101;
									assign node2195 = (inp[7]) ? node2205 : node2196;
										assign node2196 = (inp[11]) ? node2200 : node2197;
											assign node2197 = (inp[0]) ? 3'b110 : 3'b111;
											assign node2200 = (inp[2]) ? node2202 : 3'b100;
												assign node2202 = (inp[0]) ? 3'b100 : 3'b101;
										assign node2205 = (inp[2]) ? node2213 : node2206;
											assign node2206 = (inp[0]) ? node2210 : node2207;
												assign node2207 = (inp[11]) ? 3'b111 : 3'b110;
												assign node2210 = (inp[11]) ? 3'b110 : 3'b111;
											assign node2213 = (inp[0]) ? 3'b110 : node2214;
												assign node2214 = (inp[11]) ? 3'b111 : 3'b110;
								assign node2218 = (inp[3]) ? node2238 : node2219;
									assign node2219 = (inp[11]) ? node2227 : node2220;
										assign node2220 = (inp[2]) ? node2224 : node2221;
											assign node2221 = (inp[0]) ? 3'b110 : 3'b111;
											assign node2224 = (inp[0]) ? 3'b111 : 3'b110;
										assign node2227 = (inp[7]) ? node2231 : node2228;
											assign node2228 = (inp[0]) ? 3'b101 : 3'b100;
											assign node2231 = (inp[0]) ? node2235 : node2232;
												assign node2232 = (inp[2]) ? 3'b110 : 3'b111;
												assign node2235 = (inp[2]) ? 3'b111 : 3'b110;
									assign node2238 = (inp[7]) ? node2254 : node2239;
										assign node2239 = (inp[11]) ? node2247 : node2240;
											assign node2240 = (inp[0]) ? node2244 : node2241;
												assign node2241 = (inp[2]) ? 3'b101 : 3'b100;
												assign node2244 = (inp[2]) ? 3'b100 : 3'b101;
											assign node2247 = (inp[0]) ? node2251 : node2248;
												assign node2248 = (inp[2]) ? 3'b110 : 3'b111;
												assign node2251 = (inp[2]) ? 3'b111 : 3'b110;
										assign node2254 = (inp[11]) ? node2262 : node2255;
											assign node2255 = (inp[0]) ? node2259 : node2256;
												assign node2256 = (inp[2]) ? 3'b100 : 3'b101;
												assign node2259 = (inp[2]) ? 3'b101 : 3'b100;
											assign node2262 = (inp[2]) ? node2266 : node2263;
												assign node2263 = (inp[0]) ? 3'b100 : 3'b101;
												assign node2266 = (inp[0]) ? 3'b101 : 3'b100;
							assign node2269 = (inp[10]) ? node2295 : node2270;
								assign node2270 = (inp[7]) ? node2282 : node2271;
									assign node2271 = (inp[3]) ? node2277 : node2272;
										assign node2272 = (inp[2]) ? node2274 : 3'b101;
											assign node2274 = (inp[11]) ? 3'b101 : 3'b100;
										assign node2277 = (inp[11]) ? node2279 : 3'b111;
											assign node2279 = (inp[2]) ? 3'b111 : 3'b110;
									assign node2282 = (inp[3]) ? node2288 : node2283;
										assign node2283 = (inp[11]) ? 3'b110 : node2284;
											assign node2284 = (inp[2]) ? 3'b110 : 3'b111;
										assign node2288 = (inp[11]) ? node2292 : node2289;
											assign node2289 = (inp[2]) ? 3'b100 : 3'b101;
											assign node2292 = (inp[2]) ? 3'b101 : 3'b100;
								assign node2295 = (inp[7]) ? node2307 : node2296;
									assign node2296 = (inp[3]) ? node2302 : node2297;
										assign node2297 = (inp[11]) ? node2299 : 3'b101;
											assign node2299 = (inp[2]) ? 3'b100 : 3'b101;
										assign node2302 = (inp[2]) ? 3'b111 : node2303;
											assign node2303 = (inp[11]) ? 3'b111 : 3'b110;
									assign node2307 = (inp[3]) ? 3'b101 : 3'b111;
					assign node2310 = (inp[9]) ? node2432 : node2311;
						assign node2311 = (inp[8]) ? node2383 : node2312;
							assign node2312 = (inp[0]) ? node2348 : node2313;
								assign node2313 = (inp[10]) ? node2335 : node2314;
									assign node2314 = (inp[3]) ? node2322 : node2315;
										assign node2315 = (inp[7]) ? node2319 : node2316;
											assign node2316 = (inp[11]) ? 3'b110 : 3'b100;
											assign node2319 = (inp[11]) ? 3'b101 : 3'b100;
										assign node2322 = (inp[2]) ? node2330 : node2323;
											assign node2323 = (inp[11]) ? node2327 : node2324;
												assign node2324 = (inp[7]) ? 3'b110 : 3'b111;
												assign node2327 = (inp[7]) ? 3'b111 : 3'b101;
											assign node2330 = (inp[11]) ? 3'b110 : node2331;
												assign node2331 = (inp[7]) ? 3'b111 : 3'b110;
									assign node2335 = (inp[3]) ? node2343 : node2336;
										assign node2336 = (inp[7]) ? 3'b110 : node2337;
											assign node2337 = (inp[2]) ? 3'b101 : node2338;
												assign node2338 = (inp[11]) ? 3'b100 : 3'b110;
										assign node2343 = (inp[7]) ? 3'b100 : node2344;
											assign node2344 = (inp[11]) ? 3'b110 : 3'b101;
								assign node2348 = (inp[10]) ? node2368 : node2349;
									assign node2349 = (inp[3]) ? node2357 : node2350;
										assign node2350 = (inp[7]) ? node2354 : node2351;
											assign node2351 = (inp[11]) ? 3'b111 : 3'b101;
											assign node2354 = (inp[11]) ? 3'b100 : 3'b101;
										assign node2357 = (inp[11]) ? node2365 : node2358;
											assign node2358 = (inp[2]) ? node2362 : node2359;
												assign node2359 = (inp[7]) ? 3'b111 : 3'b110;
												assign node2362 = (inp[7]) ? 3'b110 : 3'b111;
											assign node2365 = (inp[7]) ? 3'b111 : 3'b100;
									assign node2368 = (inp[3]) ? node2376 : node2369;
										assign node2369 = (inp[7]) ? 3'b111 : node2370;
											assign node2370 = (inp[11]) ? node2372 : 3'b111;
												assign node2372 = (inp[2]) ? 3'b100 : 3'b101;
										assign node2376 = (inp[11]) ? node2380 : node2377;
											assign node2377 = (inp[7]) ? 3'b101 : 3'b100;
											assign node2380 = (inp[7]) ? 3'b101 : 3'b111;
							assign node2383 = (inp[10]) ? node2417 : node2384;
								assign node2384 = (inp[7]) ? node2396 : node2385;
									assign node2385 = (inp[3]) ? node2391 : node2386;
										assign node2386 = (inp[11]) ? 3'b101 : node2387;
											assign node2387 = (inp[2]) ? 3'b100 : 3'b101;
										assign node2391 = (inp[2]) ? 3'b111 : node2392;
											assign node2392 = (inp[11]) ? 3'b110 : 3'b111;
									assign node2396 = (inp[3]) ? node2404 : node2397;
										assign node2397 = (inp[2]) ? node2401 : node2398;
											assign node2398 = (inp[11]) ? 3'b110 : 3'b111;
											assign node2401 = (inp[11]) ? 3'b111 : 3'b110;
										assign node2404 = (inp[0]) ? node2412 : node2405;
											assign node2405 = (inp[11]) ? node2409 : node2406;
												assign node2406 = (inp[2]) ? 3'b100 : 3'b101;
												assign node2409 = (inp[2]) ? 3'b101 : 3'b100;
											assign node2412 = (inp[2]) ? 3'b100 : node2413;
												assign node2413 = (inp[11]) ? 3'b100 : 3'b101;
								assign node2417 = (inp[7]) ? node2429 : node2418;
									assign node2418 = (inp[3]) ? node2424 : node2419;
										assign node2419 = (inp[2]) ? node2421 : 3'b101;
											assign node2421 = (inp[11]) ? 3'b100 : 3'b101;
										assign node2424 = (inp[2]) ? 3'b111 : node2425;
											assign node2425 = (inp[11]) ? 3'b111 : 3'b110;
									assign node2429 = (inp[3]) ? 3'b101 : 3'b111;
						assign node2432 = (inp[8]) ? node2498 : node2433;
							assign node2433 = (inp[0]) ? node2467 : node2434;
								assign node2434 = (inp[3]) ? node2448 : node2435;
									assign node2435 = (inp[10]) ? node2441 : node2436;
										assign node2436 = (inp[11]) ? node2438 : 3'b101;
											assign node2438 = (inp[7]) ? 3'b100 : 3'b111;
										assign node2441 = (inp[11]) ? node2443 : 3'b111;
											assign node2443 = (inp[7]) ? 3'b111 : node2444;
												assign node2444 = (inp[2]) ? 3'b100 : 3'b101;
									assign node2448 = (inp[10]) ? node2460 : node2449;
										assign node2449 = (inp[11]) ? node2457 : node2450;
											assign node2450 = (inp[7]) ? node2454 : node2451;
												assign node2451 = (inp[2]) ? 3'b111 : 3'b110;
												assign node2454 = (inp[2]) ? 3'b110 : 3'b111;
											assign node2457 = (inp[7]) ? 3'b110 : 3'b100;
										assign node2460 = (inp[11]) ? node2464 : node2461;
											assign node2461 = (inp[7]) ? 3'b101 : 3'b100;
											assign node2464 = (inp[7]) ? 3'b101 : 3'b111;
								assign node2467 = (inp[10]) ? node2483 : node2468;
									assign node2468 = (inp[3]) ? node2474 : node2469;
										assign node2469 = (inp[11]) ? node2471 : 3'b100;
											assign node2471 = (inp[7]) ? 3'b101 : 3'b110;
										assign node2474 = (inp[7]) ? node2478 : node2475;
											assign node2475 = (inp[11]) ? 3'b101 : 3'b111;
											assign node2478 = (inp[11]) ? node2480 : 3'b110;
												assign node2480 = (inp[2]) ? 3'b110 : 3'b111;
									assign node2483 = (inp[7]) ? node2495 : node2484;
										assign node2484 = (inp[2]) ? node2490 : node2485;
											assign node2485 = (inp[3]) ? 3'b101 : node2486;
												assign node2486 = (inp[11]) ? 3'b100 : 3'b110;
											assign node2490 = (inp[3]) ? node2492 : 3'b101;
												assign node2492 = (inp[11]) ? 3'b110 : 3'b101;
										assign node2495 = (inp[3]) ? 3'b100 : 3'b110;
							assign node2498 = (inp[10]) ? node2532 : node2499;
								assign node2499 = (inp[7]) ? node2511 : node2500;
									assign node2500 = (inp[3]) ? node2506 : node2501;
										assign node2501 = (inp[2]) ? node2503 : 3'b100;
											assign node2503 = (inp[11]) ? 3'b100 : 3'b101;
										assign node2506 = (inp[2]) ? 3'b110 : node2507;
											assign node2507 = (inp[11]) ? 3'b111 : 3'b110;
									assign node2511 = (inp[3]) ? node2519 : node2512;
										assign node2512 = (inp[11]) ? node2516 : node2513;
											assign node2513 = (inp[2]) ? 3'b111 : 3'b110;
											assign node2516 = (inp[2]) ? 3'b110 : 3'b111;
										assign node2519 = (inp[0]) ? node2527 : node2520;
											assign node2520 = (inp[11]) ? node2524 : node2521;
												assign node2521 = (inp[2]) ? 3'b101 : 3'b100;
												assign node2524 = (inp[2]) ? 3'b100 : 3'b101;
											assign node2527 = (inp[2]) ? 3'b101 : node2528;
												assign node2528 = (inp[11]) ? 3'b101 : 3'b100;
								assign node2532 = (inp[3]) ? node2536 : node2533;
									assign node2533 = (inp[7]) ? 3'b110 : 3'b100;
									assign node2536 = (inp[7]) ? 3'b100 : node2537;
										assign node2537 = (inp[11]) ? 3'b110 : node2538;
											assign node2538 = (inp[2]) ? 3'b110 : 3'b111;
				assign node2543 = (inp[3]) ? node2749 : node2544;
					assign node2544 = (inp[8]) ? node2710 : node2545;
						assign node2545 = (inp[10]) ? node2625 : node2546;
							assign node2546 = (inp[11]) ? node2584 : node2547;
								assign node2547 = (inp[7]) ? node2569 : node2548;
									assign node2548 = (inp[1]) ? node2562 : node2549;
										assign node2549 = (inp[2]) ? node2555 : node2550;
											assign node2550 = (inp[0]) ? 3'b011 : node2551;
												assign node2551 = (inp[9]) ? 3'b011 : 3'b010;
											assign node2555 = (inp[0]) ? node2559 : node2556;
												assign node2556 = (inp[9]) ? 3'b010 : 3'b011;
												assign node2559 = (inp[9]) ? 3'b011 : 3'b010;
										assign node2562 = (inp[9]) ? node2566 : node2563;
											assign node2563 = (inp[0]) ? 3'b010 : 3'b011;
											assign node2566 = (inp[0]) ? 3'b011 : 3'b010;
									assign node2569 = (inp[0]) ? node2577 : node2570;
										assign node2570 = (inp[9]) ? node2572 : 3'b000;
											assign node2572 = (inp[1]) ? node2574 : 3'b001;
												assign node2574 = (inp[2]) ? 3'b000 : 3'b001;
										assign node2577 = (inp[9]) ? node2579 : 3'b001;
											assign node2579 = (inp[1]) ? node2581 : 3'b000;
												assign node2581 = (inp[2]) ? 3'b001 : 3'b000;
								assign node2584 = (inp[7]) ? node2608 : node2585;
									assign node2585 = (inp[9]) ? node2597 : node2586;
										assign node2586 = (inp[0]) ? node2592 : node2587;
											assign node2587 = (inp[1]) ? node2589 : 3'b000;
												assign node2589 = (inp[2]) ? 3'b001 : 3'b000;
											assign node2592 = (inp[2]) ? node2594 : 3'b001;
												assign node2594 = (inp[1]) ? 3'b000 : 3'b001;
										assign node2597 = (inp[0]) ? node2603 : node2598;
											assign node2598 = (inp[1]) ? node2600 : 3'b001;
												assign node2600 = (inp[2]) ? 3'b000 : 3'b001;
											assign node2603 = (inp[1]) ? node2605 : 3'b000;
												assign node2605 = (inp[2]) ? 3'b001 : 3'b000;
									assign node2608 = (inp[2]) ? node2616 : node2609;
										assign node2609 = (inp[9]) ? node2613 : node2610;
											assign node2610 = (inp[0]) ? 3'b000 : 3'b001;
											assign node2613 = (inp[0]) ? 3'b001 : 3'b000;
										assign node2616 = (inp[9]) ? 3'b000 : node2617;
											assign node2617 = (inp[0]) ? node2621 : node2618;
												assign node2618 = (inp[1]) ? 3'b000 : 3'b001;
												assign node2621 = (inp[1]) ? 3'b001 : 3'b000;
							assign node2625 = (inp[11]) ? node2665 : node2626;
								assign node2626 = (inp[7]) ? node2646 : node2627;
									assign node2627 = (inp[9]) ? node2639 : node2628;
										assign node2628 = (inp[0]) ? node2634 : node2629;
											assign node2629 = (inp[2]) ? 3'b000 : node2630;
												assign node2630 = (inp[1]) ? 3'b000 : 3'b001;
											assign node2634 = (inp[2]) ? 3'b001 : node2635;
												assign node2635 = (inp[1]) ? 3'b001 : 3'b000;
										assign node2639 = (inp[1]) ? 3'b000 : node2640;
											assign node2640 = (inp[0]) ? node2642 : 3'b000;
												assign node2642 = (inp[2]) ? 3'b000 : 3'b001;
									assign node2646 = (inp[9]) ? node2656 : node2647;
										assign node2647 = (inp[0]) ? node2653 : node2648;
											assign node2648 = (inp[2]) ? 3'b010 : node2649;
												assign node2649 = (inp[1]) ? 3'b010 : 3'b011;
											assign node2653 = (inp[2]) ? 3'b011 : 3'b010;
										assign node2656 = (inp[0]) ? node2662 : node2657;
											assign node2657 = (inp[2]) ? 3'b011 : node2658;
												assign node2658 = (inp[1]) ? 3'b011 : 3'b010;
											assign node2662 = (inp[2]) ? 3'b010 : 3'b011;
								assign node2665 = (inp[7]) ? node2687 : node2666;
									assign node2666 = (inp[0]) ? node2676 : node2667;
										assign node2667 = (inp[2]) ? 3'b011 : node2668;
											assign node2668 = (inp[9]) ? node2672 : node2669;
												assign node2669 = (inp[1]) ? 3'b011 : 3'b010;
												assign node2672 = (inp[1]) ? 3'b010 : 3'b011;
										assign node2676 = (inp[9]) ? node2682 : node2677;
											assign node2677 = (inp[2]) ? 3'b010 : node2678;
												assign node2678 = (inp[1]) ? 3'b010 : 3'b011;
											assign node2682 = (inp[2]) ? 3'b011 : node2683;
												assign node2683 = (inp[1]) ? 3'b011 : 3'b010;
									assign node2687 = (inp[0]) ? node2699 : node2688;
										assign node2688 = (inp[9]) ? node2694 : node2689;
											assign node2689 = (inp[2]) ? 3'b010 : node2690;
												assign node2690 = (inp[1]) ? 3'b010 : 3'b011;
											assign node2694 = (inp[1]) ? 3'b011 : node2695;
												assign node2695 = (inp[2]) ? 3'b011 : 3'b010;
										assign node2699 = (inp[9]) ? node2705 : node2700;
											assign node2700 = (inp[1]) ? 3'b011 : node2701;
												assign node2701 = (inp[2]) ? 3'b011 : 3'b010;
											assign node2705 = (inp[2]) ? 3'b010 : node2706;
												assign node2706 = (inp[1]) ? 3'b010 : 3'b011;
						assign node2710 = (inp[9]) ? node2726 : node2711;
							assign node2711 = (inp[7]) ? node2721 : node2712;
								assign node2712 = (inp[11]) ? 3'b010 : node2713;
									assign node2713 = (inp[10]) ? node2717 : node2714;
										assign node2714 = (inp[2]) ? 3'b011 : 3'b010;
										assign node2717 = (inp[2]) ? 3'b010 : 3'b011;
								assign node2721 = (inp[11]) ? 3'b011 : node2722;
									assign node2722 = (inp[10]) ? 3'b011 : 3'b010;
							assign node2726 = (inp[7]) ? node2744 : node2727;
								assign node2727 = (inp[11]) ? 3'b011 : node2728;
									assign node2728 = (inp[1]) ? node2736 : node2729;
										assign node2729 = (inp[10]) ? node2733 : node2730;
											assign node2730 = (inp[2]) ? 3'b010 : 3'b011;
											assign node2733 = (inp[2]) ? 3'b011 : 3'b010;
										assign node2736 = (inp[10]) ? node2740 : node2737;
											assign node2737 = (inp[2]) ? 3'b010 : 3'b011;
											assign node2740 = (inp[2]) ? 3'b011 : 3'b010;
								assign node2744 = (inp[10]) ? 3'b010 : node2745;
									assign node2745 = (inp[11]) ? 3'b010 : 3'b011;
					assign node2749 = (inp[8]) ? node2915 : node2750;
						assign node2750 = (inp[10]) ? node2848 : node2751;
							assign node2751 = (inp[7]) ? node2799 : node2752;
								assign node2752 = (inp[11]) ? node2780 : node2753;
									assign node2753 = (inp[1]) ? node2767 : node2754;
										assign node2754 = (inp[2]) ? node2760 : node2755;
											assign node2755 = (inp[9]) ? node2757 : 3'b001;
												assign node2757 = (inp[0]) ? 3'b001 : 3'b000;
											assign node2760 = (inp[0]) ? node2764 : node2761;
												assign node2761 = (inp[9]) ? 3'b001 : 3'b000;
												assign node2764 = (inp[9]) ? 3'b000 : 3'b001;
										assign node2767 = (inp[2]) ? node2775 : node2768;
											assign node2768 = (inp[9]) ? node2772 : node2769;
												assign node2769 = (inp[0]) ? 3'b001 : 3'b000;
												assign node2772 = (inp[0]) ? 3'b000 : 3'b001;
											assign node2775 = (inp[9]) ? 3'b000 : node2776;
												assign node2776 = (inp[0]) ? 3'b001 : 3'b000;
									assign node2780 = (inp[9]) ? node2790 : node2781;
										assign node2781 = (inp[2]) ? 3'b011 : node2782;
											assign node2782 = (inp[1]) ? node2786 : node2783;
												assign node2783 = (inp[0]) ? 3'b010 : 3'b011;
												assign node2786 = (inp[0]) ? 3'b011 : 3'b010;
										assign node2790 = (inp[0]) ? node2794 : node2791;
											assign node2791 = (inp[1]) ? 3'b011 : 3'b010;
											assign node2794 = (inp[1]) ? 3'b010 : node2795;
												assign node2795 = (inp[2]) ? 3'b010 : 3'b011;
								assign node2799 = (inp[1]) ? node2831 : node2800;
									assign node2800 = (inp[0]) ? node2816 : node2801;
										assign node2801 = (inp[9]) ? node2809 : node2802;
											assign node2802 = (inp[11]) ? node2806 : node2803;
												assign node2803 = (inp[2]) ? 3'b011 : 3'b010;
												assign node2806 = (inp[2]) ? 3'b010 : 3'b011;
											assign node2809 = (inp[2]) ? node2813 : node2810;
												assign node2810 = (inp[11]) ? 3'b010 : 3'b011;
												assign node2813 = (inp[11]) ? 3'b011 : 3'b010;
										assign node2816 = (inp[2]) ? node2824 : node2817;
											assign node2817 = (inp[9]) ? node2821 : node2818;
												assign node2818 = (inp[11]) ? 3'b010 : 3'b011;
												assign node2821 = (inp[11]) ? 3'b011 : 3'b010;
											assign node2824 = (inp[11]) ? node2828 : node2825;
												assign node2825 = (inp[9]) ? 3'b011 : 3'b010;
												assign node2828 = (inp[9]) ? 3'b010 : 3'b011;
									assign node2831 = (inp[0]) ? node2837 : node2832;
										assign node2832 = (inp[11]) ? 3'b010 : node2833;
											assign node2833 = (inp[9]) ? 3'b010 : 3'b011;
										assign node2837 = (inp[2]) ? node2843 : node2838;
											assign node2838 = (inp[9]) ? 3'b010 : node2839;
												assign node2839 = (inp[11]) ? 3'b011 : 3'b010;
											assign node2843 = (inp[9]) ? node2845 : 3'b011;
												assign node2845 = (inp[11]) ? 3'b010 : 3'b011;
							assign node2848 = (inp[11]) ? node2892 : node2849;
								assign node2849 = (inp[7]) ? node2873 : node2850;
									assign node2850 = (inp[2]) ? node2858 : node2851;
										assign node2851 = (inp[9]) ? node2855 : node2852;
											assign node2852 = (inp[0]) ? 3'b010 : 3'b011;
											assign node2855 = (inp[0]) ? 3'b011 : 3'b010;
										assign node2858 = (inp[0]) ? node2866 : node2859;
											assign node2859 = (inp[1]) ? node2863 : node2860;
												assign node2860 = (inp[9]) ? 3'b010 : 3'b011;
												assign node2863 = (inp[9]) ? 3'b011 : 3'b010;
											assign node2866 = (inp[1]) ? node2870 : node2867;
												assign node2867 = (inp[9]) ? 3'b011 : 3'b010;
												assign node2870 = (inp[9]) ? 3'b010 : 3'b011;
									assign node2873 = (inp[9]) ? node2885 : node2874;
										assign node2874 = (inp[0]) ? node2880 : node2875;
											assign node2875 = (inp[2]) ? 3'b000 : node2876;
												assign node2876 = (inp[1]) ? 3'b000 : 3'b001;
											assign node2880 = (inp[1]) ? 3'b001 : node2881;
												assign node2881 = (inp[2]) ? 3'b001 : 3'b000;
										assign node2885 = (inp[0]) ? 3'b000 : node2886;
											assign node2886 = (inp[2]) ? 3'b001 : node2887;
												assign node2887 = (inp[1]) ? 3'b001 : 3'b000;
								assign node2892 = (inp[9]) ? node2904 : node2893;
									assign node2893 = (inp[0]) ? node2899 : node2894;
										assign node2894 = (inp[1]) ? 3'b000 : node2895;
											assign node2895 = (inp[2]) ? 3'b000 : 3'b001;
										assign node2899 = (inp[2]) ? 3'b001 : node2900;
											assign node2900 = (inp[1]) ? 3'b001 : 3'b000;
									assign node2904 = (inp[0]) ? node2910 : node2905;
										assign node2905 = (inp[1]) ? 3'b001 : node2906;
											assign node2906 = (inp[2]) ? 3'b001 : 3'b000;
										assign node2910 = (inp[2]) ? 3'b000 : node2911;
											assign node2911 = (inp[1]) ? 3'b000 : 3'b001;
						assign node2915 = (inp[9]) ? node2929 : node2916;
							assign node2916 = (inp[11]) ? 3'b001 : node2917;
								assign node2917 = (inp[10]) ? node2923 : node2918;
									assign node2918 = (inp[7]) ? 3'b000 : node2919;
										assign node2919 = (inp[2]) ? 3'b000 : 3'b001;
									assign node2923 = (inp[7]) ? 3'b001 : node2924;
										assign node2924 = (inp[2]) ? 3'b001 : 3'b000;
							assign node2929 = (inp[11]) ? 3'b000 : node2930;
								assign node2930 = (inp[10]) ? node2936 : node2931;
									assign node2931 = (inp[2]) ? 3'b001 : node2932;
										assign node2932 = (inp[7]) ? 3'b001 : 3'b000;
									assign node2936 = (inp[2]) ? 3'b000 : node2937;
										assign node2937 = (inp[7]) ? 3'b000 : 3'b001;
			assign node2942 = (inp[7]) ? node3220 : node2943;
				assign node2943 = (inp[6]) ? node3137 : node2944;
					assign node2944 = (inp[8]) ? node3032 : node2945;
						assign node2945 = (inp[10]) ? node3009 : node2946;
							assign node2946 = (inp[2]) ? node2986 : node2947;
								assign node2947 = (inp[1]) ? node2963 : node2948;
									assign node2948 = (inp[11]) ? node2956 : node2949;
										assign node2949 = (inp[3]) ? node2953 : node2950;
											assign node2950 = (inp[0]) ? 3'b001 : 3'b000;
											assign node2953 = (inp[0]) ? 3'b000 : 3'b001;
										assign node2956 = (inp[3]) ? node2960 : node2957;
											assign node2957 = (inp[0]) ? 3'b001 : 3'b000;
											assign node2960 = (inp[0]) ? 3'b000 : 3'b001;
									assign node2963 = (inp[9]) ? node2973 : node2964;
										assign node2964 = (inp[11]) ? node2966 : 3'b001;
											assign node2966 = (inp[3]) ? node2970 : node2967;
												assign node2967 = (inp[0]) ? 3'b000 : 3'b001;
												assign node2970 = (inp[0]) ? 3'b001 : 3'b000;
										assign node2973 = (inp[0]) ? node2981 : node2974;
											assign node2974 = (inp[3]) ? node2978 : node2975;
												assign node2975 = (inp[11]) ? 3'b001 : 3'b000;
												assign node2978 = (inp[11]) ? 3'b000 : 3'b001;
											assign node2981 = (inp[3]) ? node2983 : 3'b001;
												assign node2983 = (inp[11]) ? 3'b001 : 3'b000;
								assign node2986 = (inp[11]) ? node2994 : node2987;
									assign node2987 = (inp[0]) ? node2991 : node2988;
										assign node2988 = (inp[3]) ? 3'b001 : 3'b000;
										assign node2991 = (inp[3]) ? 3'b000 : 3'b001;
									assign node2994 = (inp[3]) ? node3002 : node2995;
										assign node2995 = (inp[1]) ? node2999 : node2996;
											assign node2996 = (inp[0]) ? 3'b001 : 3'b000;
											assign node2999 = (inp[0]) ? 3'b000 : 3'b001;
										assign node3002 = (inp[0]) ? node3006 : node3003;
											assign node3003 = (inp[1]) ? 3'b000 : 3'b001;
											assign node3006 = (inp[1]) ? 3'b001 : 3'b000;
							assign node3009 = (inp[0]) ? node3021 : node3010;
								assign node3010 = (inp[3]) ? node3016 : node3011;
									assign node3011 = (inp[1]) ? 3'b010 : node3012;
										assign node3012 = (inp[11]) ? 3'b011 : 3'b010;
									assign node3016 = (inp[11]) ? node3018 : 3'b011;
										assign node3018 = (inp[1]) ? 3'b011 : 3'b010;
								assign node3021 = (inp[3]) ? node3027 : node3022;
									assign node3022 = (inp[1]) ? 3'b011 : node3023;
										assign node3023 = (inp[11]) ? 3'b010 : 3'b011;
									assign node3027 = (inp[1]) ? 3'b010 : node3028;
										assign node3028 = (inp[11]) ? 3'b011 : 3'b010;
						assign node3032 = (inp[2]) ? node3082 : node3033;
							assign node3033 = (inp[9]) ? node3067 : node3034;
								assign node3034 = (inp[11]) ? node3050 : node3035;
									assign node3035 = (inp[10]) ? node3043 : node3036;
										assign node3036 = (inp[3]) ? node3040 : node3037;
											assign node3037 = (inp[1]) ? 3'b011 : 3'b010;
											assign node3040 = (inp[1]) ? 3'b010 : 3'b011;
										assign node3043 = (inp[1]) ? node3047 : node3044;
											assign node3044 = (inp[3]) ? 3'b011 : 3'b010;
											assign node3047 = (inp[3]) ? 3'b010 : 3'b011;
									assign node3050 = (inp[0]) ? node3058 : node3051;
										assign node3051 = (inp[3]) ? node3055 : node3052;
											assign node3052 = (inp[1]) ? 3'b011 : 3'b010;
											assign node3055 = (inp[1]) ? 3'b010 : 3'b011;
										assign node3058 = (inp[10]) ? node3060 : 3'b011;
											assign node3060 = (inp[1]) ? node3064 : node3061;
												assign node3061 = (inp[3]) ? 3'b011 : 3'b010;
												assign node3064 = (inp[3]) ? 3'b010 : 3'b011;
								assign node3067 = (inp[11]) ? node3075 : node3068;
									assign node3068 = (inp[1]) ? node3072 : node3069;
										assign node3069 = (inp[3]) ? 3'b011 : 3'b010;
										assign node3072 = (inp[3]) ? 3'b010 : 3'b011;
									assign node3075 = (inp[1]) ? node3079 : node3076;
										assign node3076 = (inp[3]) ? 3'b011 : 3'b010;
										assign node3079 = (inp[3]) ? 3'b010 : 3'b011;
							assign node3082 = (inp[9]) ? node3130 : node3083;
								assign node3083 = (inp[0]) ? node3107 : node3084;
									assign node3084 = (inp[10]) ? node3100 : node3085;
										assign node3085 = (inp[11]) ? node3093 : node3086;
											assign node3086 = (inp[3]) ? node3090 : node3087;
												assign node3087 = (inp[1]) ? 3'b011 : 3'b010;
												assign node3090 = (inp[1]) ? 3'b010 : 3'b011;
											assign node3093 = (inp[3]) ? node3097 : node3094;
												assign node3094 = (inp[1]) ? 3'b011 : 3'b010;
												assign node3097 = (inp[1]) ? 3'b010 : 3'b011;
										assign node3100 = (inp[1]) ? node3104 : node3101;
											assign node3101 = (inp[3]) ? 3'b011 : 3'b010;
											assign node3104 = (inp[3]) ? 3'b010 : 3'b011;
									assign node3107 = (inp[10]) ? node3123 : node3108;
										assign node3108 = (inp[11]) ? node3116 : node3109;
											assign node3109 = (inp[1]) ? node3113 : node3110;
												assign node3110 = (inp[3]) ? 3'b011 : 3'b010;
												assign node3113 = (inp[3]) ? 3'b010 : 3'b011;
											assign node3116 = (inp[1]) ? node3120 : node3117;
												assign node3117 = (inp[3]) ? 3'b011 : 3'b010;
												assign node3120 = (inp[3]) ? 3'b010 : 3'b011;
										assign node3123 = (inp[1]) ? node3127 : node3124;
											assign node3124 = (inp[3]) ? 3'b011 : 3'b010;
											assign node3127 = (inp[3]) ? 3'b010 : 3'b011;
								assign node3130 = (inp[1]) ? node3134 : node3131;
									assign node3131 = (inp[3]) ? 3'b011 : 3'b010;
									assign node3134 = (inp[3]) ? 3'b010 : 3'b011;
					assign node3137 = (inp[10]) ? node3193 : node3138;
						assign node3138 = (inp[8]) ? node3186 : node3139;
							assign node3139 = (inp[9]) ? node3163 : node3140;
								assign node3140 = (inp[3]) ? node3152 : node3141;
									assign node3141 = (inp[0]) ? node3147 : node3142;
										assign node3142 = (inp[11]) ? 3'b010 : node3143;
											assign node3143 = (inp[1]) ? 3'b011 : 3'b010;
										assign node3147 = (inp[1]) ? node3149 : 3'b011;
											assign node3149 = (inp[11]) ? 3'b011 : 3'b010;
									assign node3152 = (inp[0]) ? node3158 : node3153;
										assign node3153 = (inp[1]) ? node3155 : 3'b011;
											assign node3155 = (inp[11]) ? 3'b011 : 3'b010;
										assign node3158 = (inp[1]) ? node3160 : 3'b010;
											assign node3160 = (inp[11]) ? 3'b010 : 3'b011;
								assign node3163 = (inp[3]) ? node3175 : node3164;
									assign node3164 = (inp[0]) ? node3170 : node3165;
										assign node3165 = (inp[11]) ? 3'b010 : node3166;
											assign node3166 = (inp[1]) ? 3'b011 : 3'b010;
										assign node3170 = (inp[1]) ? node3172 : 3'b011;
											assign node3172 = (inp[11]) ? 3'b011 : 3'b010;
									assign node3175 = (inp[0]) ? node3181 : node3176;
										assign node3176 = (inp[1]) ? node3178 : 3'b011;
											assign node3178 = (inp[11]) ? 3'b011 : 3'b010;
										assign node3181 = (inp[11]) ? 3'b010 : node3182;
											assign node3182 = (inp[1]) ? 3'b011 : 3'b010;
							assign node3186 = (inp[11]) ? node3190 : node3187;
								assign node3187 = (inp[3]) ? 3'b001 : 3'b000;
								assign node3190 = (inp[3]) ? 3'b000 : 3'b001;
						assign node3193 = (inp[3]) ? node3207 : node3194;
							assign node3194 = (inp[8]) ? 3'b001 : node3195;
								assign node3195 = (inp[0]) ? node3201 : node3196;
									assign node3196 = (inp[1]) ? 3'b000 : node3197;
										assign node3197 = (inp[11]) ? 3'b000 : 3'b001;
									assign node3201 = (inp[11]) ? 3'b001 : node3202;
										assign node3202 = (inp[1]) ? 3'b001 : 3'b000;
							assign node3207 = (inp[8]) ? 3'b000 : node3208;
								assign node3208 = (inp[0]) ? node3214 : node3209;
									assign node3209 = (inp[11]) ? 3'b001 : node3210;
										assign node3210 = (inp[1]) ? 3'b001 : 3'b000;
									assign node3214 = (inp[1]) ? 3'b000 : node3215;
										assign node3215 = (inp[11]) ? 3'b000 : 3'b001;
				assign node3220 = (inp[10]) ? node3314 : node3221;
					assign node3221 = (inp[8]) ? node3303 : node3222;
						assign node3222 = (inp[6]) ? node3288 : node3223;
							assign node3223 = (inp[9]) ? node3259 : node3224;
								assign node3224 = (inp[2]) ? node3240 : node3225;
									assign node3225 = (inp[1]) ? node3233 : node3226;
										assign node3226 = (inp[11]) ? node3230 : node3227;
											assign node3227 = (inp[0]) ? 3'b011 : 3'b010;
											assign node3230 = (inp[0]) ? 3'b010 : 3'b011;
										assign node3233 = (inp[11]) ? node3237 : node3234;
											assign node3234 = (inp[0]) ? 3'b011 : 3'b010;
											assign node3237 = (inp[0]) ? 3'b010 : 3'b011;
									assign node3240 = (inp[1]) ? node3246 : node3241;
										assign node3241 = (inp[11]) ? 3'b010 : node3242;
											assign node3242 = (inp[0]) ? 3'b011 : 3'b010;
										assign node3246 = (inp[3]) ? node3254 : node3247;
											assign node3247 = (inp[0]) ? node3251 : node3248;
												assign node3248 = (inp[11]) ? 3'b011 : 3'b010;
												assign node3251 = (inp[11]) ? 3'b010 : 3'b011;
											assign node3254 = (inp[11]) ? node3256 : 3'b010;
												assign node3256 = (inp[0]) ? 3'b010 : 3'b011;
								assign node3259 = (inp[3]) ? node3267 : node3260;
									assign node3260 = (inp[11]) ? node3264 : node3261;
										assign node3261 = (inp[0]) ? 3'b011 : 3'b010;
										assign node3264 = (inp[0]) ? 3'b010 : 3'b011;
									assign node3267 = (inp[1]) ? node3275 : node3268;
										assign node3268 = (inp[11]) ? node3272 : node3269;
											assign node3269 = (inp[0]) ? 3'b011 : 3'b010;
											assign node3272 = (inp[0]) ? 3'b010 : 3'b011;
										assign node3275 = (inp[2]) ? node3283 : node3276;
											assign node3276 = (inp[11]) ? node3280 : node3277;
												assign node3277 = (inp[0]) ? 3'b011 : 3'b010;
												assign node3280 = (inp[0]) ? 3'b010 : 3'b011;
											assign node3283 = (inp[0]) ? node3285 : 3'b011;
												assign node3285 = (inp[11]) ? 3'b010 : 3'b011;
							assign node3288 = (inp[3]) ? node3296 : node3289;
								assign node3289 = (inp[0]) ? node3293 : node3290;
									assign node3290 = (inp[11]) ? 3'b011 : 3'b010;
									assign node3293 = (inp[11]) ? 3'b010 : 3'b011;
								assign node3296 = (inp[11]) ? node3300 : node3297;
									assign node3297 = (inp[0]) ? 3'b011 : 3'b010;
									assign node3300 = (inp[0]) ? 3'b010 : 3'b011;
						assign node3303 = (inp[11]) ? node3309 : node3304;
							assign node3304 = (inp[6]) ? 3'b001 : node3305;
								assign node3305 = (inp[1]) ? 3'b001 : 3'b000;
							assign node3309 = (inp[1]) ? 3'b000 : node3310;
								assign node3310 = (inp[6]) ? 3'b000 : 3'b001;
					assign node3314 = (inp[0]) ? node3326 : node3315;
						assign node3315 = (inp[8]) ? node3321 : node3316;
							assign node3316 = (inp[1]) ? 3'b001 : node3317;
								assign node3317 = (inp[6]) ? 3'b001 : 3'b000;
							assign node3321 = (inp[1]) ? 3'b000 : node3322;
								assign node3322 = (inp[6]) ? 3'b000 : 3'b001;
						assign node3326 = (inp[1]) ? 3'b000 : node3327;
							assign node3327 = (inp[6]) ? 3'b000 : 3'b001;

endmodule