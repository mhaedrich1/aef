module dtc_split05_bm84 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;

	assign outp = (inp[9]) ? node84 : node1;
		assign node1 = (inp[6]) ? node43 : node2;
			assign node2 = (inp[10]) ? node18 : node3;
				assign node3 = (inp[0]) ? node11 : node4;
					assign node4 = (inp[11]) ? node6 : 3'b111;
						assign node6 = (inp[4]) ? node8 : 3'b101;
							assign node8 = (inp[2]) ? 3'b111 : 3'b011;
					assign node11 = (inp[2]) ? node13 : 3'b111;
						assign node13 = (inp[11]) ? 3'b011 : node14;
							assign node14 = (inp[3]) ? 3'b011 : 3'b111;
				assign node18 = (inp[2]) ? node32 : node19;
					assign node19 = (inp[0]) ? node25 : node20;
						assign node20 = (inp[7]) ? node22 : 3'b101;
							assign node22 = (inp[1]) ? 3'b001 : 3'b101;
						assign node25 = (inp[8]) ? node29 : node26;
							assign node26 = (inp[7]) ? 3'b101 : 3'b011;
							assign node29 = (inp[11]) ? 3'b101 : 3'b001;
					assign node32 = (inp[11]) ? node36 : node33;
						assign node33 = (inp[3]) ? 3'b011 : 3'b001;
						assign node36 = (inp[8]) ? node40 : node37;
							assign node37 = (inp[0]) ? 3'b101 : 3'b011;
							assign node40 = (inp[4]) ? 3'b010 : 3'b110;
			assign node43 = (inp[10]) ? node73 : node44;
				assign node44 = (inp[11]) ? node60 : node45;
					assign node45 = (inp[7]) ? node53 : node46;
						assign node46 = (inp[4]) ? node50 : node47;
							assign node47 = (inp[5]) ? 3'b001 : 3'b011;
							assign node50 = (inp[2]) ? 3'b001 : 3'b101;
						assign node53 = (inp[5]) ? node57 : node54;
							assign node54 = (inp[8]) ? 3'b000 : 3'b001;
							assign node57 = (inp[4]) ? 3'b110 : 3'b001;
					assign node60 = (inp[4]) ? node66 : node61;
						assign node61 = (inp[1]) ? 3'b110 : node62;
							assign node62 = (inp[7]) ? 3'b010 : 3'b110;
						assign node66 = (inp[7]) ? node70 : node67;
							assign node67 = (inp[3]) ? 3'b110 : 3'b001;
							assign node70 = (inp[0]) ? 3'b000 : 3'b010;
				assign node73 = (inp[7]) ? node81 : node74;
					assign node74 = (inp[11]) ? node78 : node75;
						assign node75 = (inp[8]) ? 3'b010 : 3'b110;
						assign node78 = (inp[8]) ? 3'b100 : 3'b010;
					assign node81 = (inp[11]) ? 3'b000 : 3'b100;
		assign node84 = (inp[6]) ? node116 : node85;
			assign node85 = (inp[7]) ? node103 : node86;
				assign node86 = (inp[10]) ? node96 : node87;
					assign node87 = (inp[8]) ? node93 : node88;
						assign node88 = (inp[4]) ? node90 : 3'b001;
							assign node90 = (inp[3]) ? 3'b110 : 3'b101;
						assign node93 = (inp[11]) ? 3'b010 : 3'b000;
					assign node96 = (inp[8]) ? node100 : node97;
						assign node97 = (inp[11]) ? 3'b100 : 3'b010;
						assign node100 = (inp[11]) ? 3'b000 : 3'b100;
				assign node103 = (inp[10]) ? 3'b000 : node104;
					assign node104 = (inp[11]) ? node110 : node105;
						assign node105 = (inp[5]) ? node107 : 3'b010;
							assign node107 = (inp[2]) ? 3'b100 : 3'b010;
						assign node110 = (inp[4]) ? node112 : 3'b100;
							assign node112 = (inp[2]) ? 3'b100 : 3'b000;
			assign node116 = (inp[7]) ? 3'b000 : node117;
				assign node117 = (inp[10]) ? 3'b000 : node118;
					assign node118 = (inp[8]) ? 3'b000 : node119;
						assign node119 = (inp[11]) ? 3'b000 : 3'b100;

endmodule