module dtc_split5_bm15 (
	input  wire [15-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node6;
	wire [1-1:0] node8;
	wire [1-1:0] node10;
	wire [1-1:0] node12;
	wire [1-1:0] node14;
	wire [1-1:0] node16;
	wire [1-1:0] node19;
	wire [1-1:0] node20;
	wire [1-1:0] node22;
	wire [1-1:0] node24;
	wire [1-1:0] node26;
	wire [1-1:0] node28;
	wire [1-1:0] node30;
	wire [1-1:0] node33;
	wire [1-1:0] node34;
	wire [1-1:0] node36;
	wire [1-1:0] node38;
	wire [1-1:0] node40;
	wire [1-1:0] node41;
	wire [1-1:0] node45;
	wire [1-1:0] node46;
	wire [1-1:0] node48;
	wire [1-1:0] node50;
	wire [1-1:0] node52;
	wire [1-1:0] node55;
	wire [1-1:0] node56;
	wire [1-1:0] node58;
	wire [1-1:0] node60;
	wire [1-1:0] node63;
	wire [1-1:0] node64;
	wire [1-1:0] node66;
	wire [1-1:0] node70;
	wire [1-1:0] node71;
	wire [1-1:0] node72;
	wire [1-1:0] node74;
	wire [1-1:0] node76;
	wire [1-1:0] node78;
	wire [1-1:0] node80;
	wire [1-1:0] node83;
	wire [1-1:0] node84;
	wire [1-1:0] node86;
	wire [1-1:0] node88;
	wire [1-1:0] node90;
	wire [1-1:0] node92;
	wire [1-1:0] node95;
	wire [1-1:0] node96;
	wire [1-1:0] node98;
	wire [1-1:0] node100;
	wire [1-1:0] node102;
	wire [1-1:0] node105;
	wire [1-1:0] node106;
	wire [1-1:0] node108;
	wire [1-1:0] node110;
	wire [1-1:0] node113;
	wire [1-1:0] node114;
	wire [1-1:0] node116;
	wire [1-1:0] node119;
	wire [1-1:0] node120;
	wire [1-1:0] node124;
	wire [1-1:0] node125;
	wire [1-1:0] node126;
	wire [1-1:0] node128;
	wire [1-1:0] node130;
	wire [1-1:0] node132;
	wire [1-1:0] node133;
	wire [1-1:0] node137;
	wire [1-1:0] node138;
	wire [1-1:0] node140;
	wire [1-1:0] node142;
	wire [1-1:0] node144;
	wire [1-1:0] node147;
	wire [1-1:0] node148;
	wire [1-1:0] node150;
	wire [1-1:0] node152;
	wire [1-1:0] node155;
	wire [1-1:0] node156;
	wire [1-1:0] node158;
	wire [1-1:0] node161;
	wire [1-1:0] node162;
	wire [1-1:0] node166;
	wire [1-1:0] node167;
	wire [1-1:0] node168;
	wire [1-1:0] node170;
	wire [1-1:0] node172;
	wire [1-1:0] node174;
	wire [1-1:0] node177;
	wire [1-1:0] node178;
	wire [1-1:0] node180;
	wire [1-1:0] node181;
	wire [1-1:0] node184;
	wire [1-1:0] node187;
	wire [1-1:0] node189;
	wire [1-1:0] node190;
	wire [1-1:0] node194;
	wire [1-1:0] node195;
	wire [1-1:0] node197;
	wire [1-1:0] node198;
	wire [1-1:0] node200;
	wire [1-1:0] node203;
	wire [1-1:0] node204;
	wire [1-1:0] node208;
	wire [1-1:0] node209;
	wire [1-1:0] node210;
	wire [1-1:0] node212;
	wire [1-1:0] node215;
	wire [1-1:0] node216;
	wire [1-1:0] node220;
	wire [1-1:0] node221;
	wire [1-1:0] node222;
	wire [1-1:0] node227;
	wire [1-1:0] node228;
	wire [1-1:0] node229;
	wire [1-1:0] node230;
	wire [1-1:0] node232;
	wire [1-1:0] node234;
	wire [1-1:0] node236;
	wire [1-1:0] node238;
	wire [1-1:0] node240;
	wire [1-1:0] node243;
	wire [1-1:0] node244;
	wire [1-1:0] node246;
	wire [1-1:0] node248;
	wire [1-1:0] node250;
	wire [1-1:0] node251;
	wire [1-1:0] node254;
	wire [1-1:0] node257;
	wire [1-1:0] node258;
	wire [1-1:0] node260;
	wire [1-1:0] node262;
	wire [1-1:0] node264;
	wire [1-1:0] node267;
	wire [1-1:0] node268;
	wire [1-1:0] node270;
	wire [1-1:0] node272;
	wire [1-1:0] node275;
	wire [1-1:0] node276;
	wire [1-1:0] node278;
	wire [1-1:0] node282;
	wire [1-1:0] node283;
	wire [1-1:0] node284;
	wire [1-1:0] node286;
	wire [1-1:0] node288;
	wire [1-1:0] node290;
	wire [1-1:0] node293;
	wire [1-1:0] node294;
	wire [1-1:0] node296;
	wire [1-1:0] node298;
	wire [1-1:0] node300;
	wire [1-1:0] node303;
	wire [1-1:0] node304;
	wire [1-1:0] node306;
	wire [1-1:0] node309;
	wire [1-1:0] node310;
	wire [1-1:0] node312;
	wire [1-1:0] node315;
	wire [1-1:0] node316;
	wire [1-1:0] node320;
	wire [1-1:0] node321;
	wire [1-1:0] node322;
	wire [1-1:0] node324;
	wire [1-1:0] node326;
	wire [1-1:0] node328;
	wire [1-1:0] node331;
	wire [1-1:0] node332;
	wire [1-1:0] node334;
	wire [1-1:0] node336;
	wire [1-1:0] node339;
	wire [1-1:0] node340;
	wire [1-1:0] node343;
	wire [1-1:0] node344;
	wire [1-1:0] node348;
	wire [1-1:0] node349;
	wire [1-1:0] node350;
	wire [1-1:0] node352;
	wire [1-1:0] node354;
	wire [1-1:0] node357;
	wire [1-1:0] node358;
	wire [1-1:0] node360;
	wire [1-1:0] node364;
	wire [1-1:0] node365;
	wire [1-1:0] node366;
	wire [1-1:0] node368;
	wire [1-1:0] node371;
	wire [1-1:0] node372;
	wire [1-1:0] node377;
	wire [1-1:0] node378;
	wire [1-1:0] node379;
	wire [1-1:0] node380;
	wire [1-1:0] node382;
	wire [1-1:0] node384;
	wire [1-1:0] node386;
	wire [1-1:0] node389;
	wire [1-1:0] node390;
	wire [1-1:0] node392;
	wire [1-1:0] node394;
	wire [1-1:0] node396;
	wire [1-1:0] node399;
	wire [1-1:0] node400;
	wire [1-1:0] node402;
	wire [1-1:0] node404;
	wire [1-1:0] node407;
	wire [1-1:0] node408;
	wire [1-1:0] node409;
	wire [1-1:0] node414;
	wire [1-1:0] node415;
	wire [1-1:0] node416;
	wire [1-1:0] node418;
	wire [1-1:0] node420;
	wire [1-1:0] node422;
	wire [1-1:0] node425;
	wire [1-1:0] node426;
	wire [1-1:0] node428;
	wire [1-1:0] node430;
	wire [1-1:0] node433;
	wire [1-1:0] node434;
	wire [1-1:0] node436;
	wire [1-1:0] node440;
	wire [1-1:0] node441;
	wire [1-1:0] node442;
	wire [1-1:0] node444;
	wire [1-1:0] node446;
	wire [1-1:0] node449;
	wire [1-1:0] node450;
	wire [1-1:0] node452;
	wire [1-1:0] node455;
	wire [1-1:0] node456;
	wire [1-1:0] node460;
	wire [1-1:0] node461;
	wire [1-1:0] node462;
	wire [1-1:0] node464;
	wire [1-1:0] node467;
	wire [1-1:0] node468;
	wire [1-1:0] node472;
	wire [1-1:0] node473;
	wire [1-1:0] node474;
	wire [1-1:0] node479;
	wire [1-1:0] node480;
	wire [1-1:0] node481;
	wire [1-1:0] node482;
	wire [1-1:0] node484;
	wire [1-1:0] node486;
	wire [1-1:0] node488;
	wire [1-1:0] node491;
	wire [1-1:0] node492;
	wire [1-1:0] node494;
	wire [1-1:0] node495;
	wire [1-1:0] node498;
	wire [1-1:0] node501;
	wire [1-1:0] node502;
	wire [1-1:0] node504;
	wire [1-1:0] node508;
	wire [1-1:0] node509;
	wire [1-1:0] node510;
	wire [1-1:0] node512;
	wire [1-1:0] node514;
	wire [1-1:0] node517;
	wire [1-1:0] node518;
	wire [1-1:0] node520;
	wire [1-1:0] node523;
	wire [1-1:0] node524;
	wire [1-1:0] node528;
	wire [1-1:0] node529;
	wire [1-1:0] node530;
	wire [1-1:0] node532;
	wire [1-1:0] node535;
	wire [1-1:0] node536;
	wire [1-1:0] node540;
	wire [1-1:0] node541;
	wire [1-1:0] node542;
	wire [1-1:0] node547;
	wire [1-1:0] node548;
	wire [1-1:0] node549;
	wire [1-1:0] node550;
	wire [1-1:0] node552;
	wire [1-1:0] node554;
	wire [1-1:0] node557;
	wire [1-1:0] node558;
	wire [1-1:0] node560;
	wire [1-1:0] node563;
	wire [1-1:0] node564;
	wire [1-1:0] node568;
	wire [1-1:0] node569;
	wire [1-1:0] node570;
	wire [1-1:0] node572;
	wire [1-1:0] node575;
	wire [1-1:0] node576;
	wire [1-1:0] node581;
	wire [1-1:0] node582;
	wire [1-1:0] node583;
	wire [1-1:0] node584;
	wire [1-1:0] node586;
	wire [1-1:0] node589;
	wire [1-1:0] node590;
	wire [1-1:0] node594;
	wire [1-1:0] node595;
	wire [1-1:0] node596;
	wire [1-1:0] node602;
	wire [1-1:0] node603;
	wire [1-1:0] node604;
	wire [1-1:0] node605;
	wire [1-1:0] node607;
	wire [1-1:0] node608;
	wire [1-1:0] node610;
	wire [1-1:0] node612;
	wire [1-1:0] node614;
	wire [1-1:0] node616;
	wire [1-1:0] node619;
	wire [1-1:0] node620;
	wire [1-1:0] node622;
	wire [1-1:0] node624;
	wire [1-1:0] node626;
	wire [1-1:0] node629;
	wire [1-1:0] node630;
	wire [1-1:0] node632;
	wire [1-1:0] node634;
	wire [1-1:0] node637;
	wire [1-1:0] node638;
	wire [1-1:0] node639;
	wire [1-1:0] node642;
	wire [1-1:0] node645;
	wire [1-1:0] node646;
	wire [1-1:0] node650;
	wire [1-1:0] node651;
	wire [1-1:0] node652;
	wire [1-1:0] node654;
	wire [1-1:0] node656;
	wire [1-1:0] node658;
	wire [1-1:0] node661;
	wire [1-1:0] node662;
	wire [1-1:0] node664;
	wire [1-1:0] node666;
	wire [1-1:0] node668;
	wire [1-1:0] node671;
	wire [1-1:0] node672;
	wire [1-1:0] node674;
	wire [1-1:0] node676;
	wire [1-1:0] node679;
	wire [1-1:0] node680;
	wire [1-1:0] node682;
	wire [1-1:0] node686;
	wire [1-1:0] node687;
	wire [1-1:0] node689;
	wire [1-1:0] node690;
	wire [1-1:0] node692;
	wire [1-1:0] node693;
	wire [1-1:0] node696;
	wire [1-1:0] node699;
	wire [1-1:0] node700;
	wire [1-1:0] node702;
	wire [1-1:0] node705;
	wire [1-1:0] node706;
	wire [1-1:0] node710;
	wire [1-1:0] node711;
	wire [1-1:0] node712;
	wire [1-1:0] node714;
	wire [1-1:0] node716;
	wire [1-1:0] node719;
	wire [1-1:0] node720;
	wire [1-1:0] node722;
	wire [1-1:0] node726;
	wire [1-1:0] node727;
	wire [1-1:0] node728;
	wire [1-1:0] node730;
	wire [1-1:0] node733;
	wire [1-1:0] node734;
	wire [1-1:0] node739;
	wire [1-1:0] node740;
	wire [1-1:0] node741;
	wire [1-1:0] node742;
	wire [1-1:0] node744;
	wire [1-1:0] node746;
	wire [1-1:0] node748;
	wire [1-1:0] node750;
	wire [1-1:0] node753;
	wire [1-1:0] node754;
	wire [1-1:0] node756;
	wire [1-1:0] node758;
	wire [1-1:0] node760;
	wire [1-1:0] node763;
	wire [1-1:0] node764;
	wire [1-1:0] node766;
	wire [1-1:0] node768;
	wire [1-1:0] node771;
	wire [1-1:0] node772;
	wire [1-1:0] node774;
	wire [1-1:0] node777;
	wire [1-1:0] node778;
	wire [1-1:0] node782;
	wire [1-1:0] node783;
	wire [1-1:0] node784;
	wire [1-1:0] node786;
	wire [1-1:0] node788;
	wire [1-1:0] node790;
	wire [1-1:0] node793;
	wire [1-1:0] node794;
	wire [1-1:0] node796;
	wire [1-1:0] node797;
	wire [1-1:0] node801;
	wire [1-1:0] node802;
	wire [1-1:0] node804;
	wire [1-1:0] node808;
	wire [1-1:0] node809;
	wire [1-1:0] node810;
	wire [1-1:0] node812;
	wire [1-1:0] node814;
	wire [1-1:0] node817;
	wire [1-1:0] node818;
	wire [1-1:0] node820;
	wire [1-1:0] node823;
	wire [1-1:0] node824;
	wire [1-1:0] node828;
	wire [1-1:0] node829;
	wire [1-1:0] node830;
	wire [1-1:0] node832;
	wire [1-1:0] node835;
	wire [1-1:0] node836;
	wire [1-1:0] node840;
	wire [1-1:0] node841;
	wire [1-1:0] node842;
	wire [1-1:0] node847;
	wire [1-1:0] node848;
	wire [1-1:0] node849;
	wire [1-1:0] node850;
	wire [1-1:0] node852;
	wire [1-1:0] node854;
	wire [1-1:0] node856;
	wire [1-1:0] node859;
	wire [1-1:0] node860;
	wire [1-1:0] node862;
	wire [1-1:0] node864;
	wire [1-1:0] node867;
	wire [1-1:0] node868;
	wire [1-1:0] node870;
	wire [1-1:0] node873;
	wire [1-1:0] node874;
	wire [1-1:0] node877;
	wire [1-1:0] node880;
	wire [1-1:0] node881;
	wire [1-1:0] node882;
	wire [1-1:0] node884;
	wire [1-1:0] node886;
	wire [1-1:0] node889;
	wire [1-1:0] node890;
	wire [1-1:0] node892;
	wire [1-1:0] node895;
	wire [1-1:0] node896;
	wire [1-1:0] node900;
	wire [1-1:0] node901;
	wire [1-1:0] node902;
	wire [1-1:0] node905;
	wire [1-1:0] node906;
	wire [1-1:0] node910;
	wire [1-1:0] node911;
	wire [1-1:0] node912;
	wire [1-1:0] node917;
	wire [1-1:0] node918;
	wire [1-1:0] node919;
	wire [1-1:0] node920;
	wire [1-1:0] node922;
	wire [1-1:0] node924;
	wire [1-1:0] node927;
	wire [1-1:0] node928;
	wire [1-1:0] node929;
	wire [1-1:0] node932;
	wire [1-1:0] node935;
	wire [1-1:0] node936;
	wire [1-1:0] node940;
	wire [1-1:0] node941;
	wire [1-1:0] node942;
	wire [1-1:0] node944;
	wire [1-1:0] node947;
	wire [1-1:0] node948;
	wire [1-1:0] node952;
	wire [1-1:0] node953;
	wire [1-1:0] node954;
	wire [1-1:0] node959;
	wire [1-1:0] node960;
	wire [1-1:0] node961;
	wire [1-1:0] node962;
	wire [1-1:0] node964;
	wire [1-1:0] node967;
	wire [1-1:0] node968;
	wire [1-1:0] node972;
	wire [1-1:0] node973;
	wire [1-1:0] node974;
	wire [1-1:0] node979;
	wire [1-1:0] node980;
	wire [1-1:0] node981;
	wire [1-1:0] node982;
	wire [1-1:0] node988;
	wire [1-1:0] node989;
	wire [1-1:0] node990;
	wire [1-1:0] node991;
	wire [1-1:0] node992;
	wire [1-1:0] node994;
	wire [1-1:0] node996;
	wire [1-1:0] node998;
	wire [1-1:0] node1000;
	wire [1-1:0] node1003;
	wire [1-1:0] node1004;
	wire [1-1:0] node1006;
	wire [1-1:0] node1008;
	wire [1-1:0] node1010;
	wire [1-1:0] node1013;
	wire [1-1:0] node1014;
	wire [1-1:0] node1016;
	wire [1-1:0] node1018;
	wire [1-1:0] node1021;
	wire [1-1:0] node1022;
	wire [1-1:0] node1024;
	wire [1-1:0] node1027;
	wire [1-1:0] node1028;
	wire [1-1:0] node1032;
	wire [1-1:0] node1033;
	wire [1-1:0] node1034;
	wire [1-1:0] node1036;
	wire [1-1:0] node1038;
	wire [1-1:0] node1040;
	wire [1-1:0] node1043;
	wire [1-1:0] node1044;
	wire [1-1:0] node1046;
	wire [1-1:0] node1048;
	wire [1-1:0] node1051;
	wire [1-1:0] node1052;
	wire [1-1:0] node1053;
	wire [1-1:0] node1056;
	wire [1-1:0] node1059;
	wire [1-1:0] node1060;
	wire [1-1:0] node1064;
	wire [1-1:0] node1065;
	wire [1-1:0] node1067;
	wire [1-1:0] node1068;
	wire [1-1:0] node1070;
	wire [1-1:0] node1073;
	wire [1-1:0] node1074;
	wire [1-1:0] node1078;
	wire [1-1:0] node1079;
	wire [1-1:0] node1080;
	wire [1-1:0] node1082;
	wire [1-1:0] node1085;
	wire [1-1:0] node1086;
	wire [1-1:0] node1090;
	wire [1-1:0] node1091;
	wire [1-1:0] node1092;
	wire [1-1:0] node1097;
	wire [1-1:0] node1098;
	wire [1-1:0] node1099;
	wire [1-1:0] node1100;
	wire [1-1:0] node1102;
	wire [1-1:0] node1104;
	wire [1-1:0] node1106;
	wire [1-1:0] node1109;
	wire [1-1:0] node1110;
	wire [1-1:0] node1112;
	wire [1-1:0] node1115;
	wire [1-1:0] node1116;
	wire [1-1:0] node1118;
	wire [1-1:0] node1122;
	wire [1-1:0] node1123;
	wire [1-1:0] node1124;
	wire [1-1:0] node1126;
	wire [1-1:0] node1128;
	wire [1-1:0] node1131;
	wire [1-1:0] node1132;
	wire [1-1:0] node1134;
	wire [1-1:0] node1137;
	wire [1-1:0] node1138;
	wire [1-1:0] node1142;
	wire [1-1:0] node1143;
	wire [1-1:0] node1144;
	wire [1-1:0] node1146;
	wire [1-1:0] node1149;
	wire [1-1:0] node1150;
	wire [1-1:0] node1154;
	wire [1-1:0] node1155;
	wire [1-1:0] node1156;
	wire [1-1:0] node1161;
	wire [1-1:0] node1162;
	wire [1-1:0] node1163;
	wire [1-1:0] node1165;
	wire [1-1:0] node1166;
	wire [1-1:0] node1168;
	wire [1-1:0] node1171;
	wire [1-1:0] node1172;
	wire [1-1:0] node1176;
	wire [1-1:0] node1177;
	wire [1-1:0] node1178;
	wire [1-1:0] node1180;
	wire [1-1:0] node1183;
	wire [1-1:0] node1184;
	wire [1-1:0] node1188;
	wire [1-1:0] node1189;
	wire [1-1:0] node1190;
	wire [1-1:0] node1195;
	wire [1-1:0] node1196;
	wire [1-1:0] node1197;
	wire [1-1:0] node1198;
	wire [1-1:0] node1200;
	wire [1-1:0] node1203;
	wire [1-1:0] node1204;
	wire [1-1:0] node1208;
	wire [1-1:0] node1209;
	wire [1-1:0] node1210;
	wire [1-1:0] node1215;
	wire [1-1:0] node1216;
	wire [1-1:0] node1217;
	wire [1-1:0] node1218;
	wire [1-1:0] node1224;
	wire [1-1:0] node1225;
	wire [1-1:0] node1226;
	wire [1-1:0] node1227;
	wire [1-1:0] node1228;
	wire [1-1:0] node1230;
	wire [1-1:0] node1232;
	wire [1-1:0] node1234;
	wire [1-1:0] node1237;
	wire [1-1:0] node1238;
	wire [1-1:0] node1240;
	wire [1-1:0] node1242;
	wire [1-1:0] node1245;
	wire [1-1:0] node1246;
	wire [1-1:0] node1248;
	wire [1-1:0] node1251;
	wire [1-1:0] node1252;
	wire [1-1:0] node1256;
	wire [1-1:0] node1257;
	wire [1-1:0] node1258;
	wire [1-1:0] node1260;
	wire [1-1:0] node1262;
	wire [1-1:0] node1265;
	wire [1-1:0] node1266;
	wire [1-1:0] node1268;
	wire [1-1:0] node1271;
	wire [1-1:0] node1272;
	wire [1-1:0] node1276;
	wire [1-1:0] node1277;
	wire [1-1:0] node1278;
	wire [1-1:0] node1280;
	wire [1-1:0] node1283;
	wire [1-1:0] node1284;
	wire [1-1:0] node1288;
	wire [1-1:0] node1289;
	wire [1-1:0] node1290;
	wire [1-1:0] node1295;
	wire [1-1:0] node1296;
	wire [1-1:0] node1297;
	wire [1-1:0] node1298;
	wire [1-1:0] node1300;
	wire [1-1:0] node1302;
	wire [1-1:0] node1305;
	wire [1-1:0] node1306;
	wire [1-1:0] node1308;
	wire [1-1:0] node1311;
	wire [1-1:0] node1312;
	wire [1-1:0] node1316;
	wire [1-1:0] node1317;
	wire [1-1:0] node1318;
	wire [1-1:0] node1320;
	wire [1-1:0] node1323;
	wire [1-1:0] node1324;
	wire [1-1:0] node1328;
	wire [1-1:0] node1329;
	wire [1-1:0] node1330;
	wire [1-1:0] node1335;
	wire [1-1:0] node1336;
	wire [1-1:0] node1337;
	wire [1-1:0] node1338;
	wire [1-1:0] node1340;
	wire [1-1:0] node1343;
	wire [1-1:0] node1344;
	wire [1-1:0] node1348;
	wire [1-1:0] node1349;
	wire [1-1:0] node1350;
	wire [1-1:0] node1355;
	wire [1-1:0] node1356;
	wire [1-1:0] node1357;
	wire [1-1:0] node1358;
	wire [1-1:0] node1364;
	wire [1-1:0] node1365;
	wire [1-1:0] node1366;
	wire [1-1:0] node1367;
	wire [1-1:0] node1368;
	wire [1-1:0] node1370;
	wire [1-1:0] node1372;
	wire [1-1:0] node1375;
	wire [1-1:0] node1376;
	wire [1-1:0] node1378;
	wire [1-1:0] node1381;
	wire [1-1:0] node1382;
	wire [1-1:0] node1386;
	wire [1-1:0] node1387;
	wire [1-1:0] node1388;
	wire [1-1:0] node1390;
	wire [1-1:0] node1393;
	wire [1-1:0] node1394;
	wire [1-1:0] node1398;
	wire [1-1:0] node1399;
	wire [1-1:0] node1400;
	wire [1-1:0] node1405;
	wire [1-1:0] node1406;
	wire [1-1:0] node1407;
	wire [1-1:0] node1408;
	wire [1-1:0] node1410;
	wire [1-1:0] node1413;
	wire [1-1:0] node1414;
	wire [1-1:0] node1418;
	wire [1-1:0] node1419;
	wire [1-1:0] node1423;
	wire [1-1:0] node1424;
	wire [1-1:0] node1425;
	wire [1-1:0] node1426;
	wire [1-1:0] node1432;
	wire [1-1:0] node1433;
	wire [1-1:0] node1434;
	wire [1-1:0] node1435;
	wire [1-1:0] node1436;
	wire [1-1:0] node1438;
	wire [1-1:0] node1441;
	wire [1-1:0] node1442;
	wire [1-1:0] node1446;
	wire [1-1:0] node1447;
	wire [1-1:0] node1448;
	wire [1-1:0] node1453;
	wire [1-1:0] node1454;
	wire [1-1:0] node1455;
	wire [1-1:0] node1456;
	wire [1-1:0] node1462;
	wire [1-1:0] node1463;
	wire [1-1:0] node1464;
	wire [1-1:0] node1465;
	wire [1-1:0] node1466;
	wire [1-1:0] node1473;
	wire [1-1:0] node1474;
	wire [1-1:0] node1475;
	wire [1-1:0] node1476;
	wire [1-1:0] node1477;
	wire [1-1:0] node1478;
	wire [1-1:0] node1480;
	wire [1-1:0] node1482;
	wire [1-1:0] node1484;
	wire [1-1:0] node1486;
	wire [1-1:0] node1488;
	wire [1-1:0] node1491;
	wire [1-1:0] node1492;
	wire [1-1:0] node1494;
	wire [1-1:0] node1496;
	wire [1-1:0] node1498;
	wire [1-1:0] node1500;
	wire [1-1:0] node1503;
	wire [1-1:0] node1504;
	wire [1-1:0] node1506;
	wire [1-1:0] node1508;
	wire [1-1:0] node1510;
	wire [1-1:0] node1513;
	wire [1-1:0] node1514;
	wire [1-1:0] node1516;
	wire [1-1:0] node1518;
	wire [1-1:0] node1521;
	wire [1-1:0] node1522;
	wire [1-1:0] node1523;
	wire [1-1:0] node1526;
	wire [1-1:0] node1529;
	wire [1-1:0] node1530;
	wire [1-1:0] node1534;
	wire [1-1:0] node1535;
	wire [1-1:0] node1536;
	wire [1-1:0] node1538;
	wire [1-1:0] node1540;
	wire [1-1:0] node1542;
	wire [1-1:0] node1544;
	wire [1-1:0] node1547;
	wire [1-1:0] node1548;
	wire [1-1:0] node1550;
	wire [1-1:0] node1552;
	wire [1-1:0] node1554;
	wire [1-1:0] node1557;
	wire [1-1:0] node1558;
	wire [1-1:0] node1560;
	wire [1-1:0] node1562;
	wire [1-1:0] node1565;
	wire [1-1:0] node1566;
	wire [1-1:0] node1570;
	wire [1-1:0] node1571;
	wire [1-1:0] node1572;
	wire [1-1:0] node1574;
	wire [1-1:0] node1576;
	wire [1-1:0] node1578;
	wire [1-1:0] node1581;
	wire [1-1:0] node1582;
	wire [1-1:0] node1584;
	wire [1-1:0] node1586;
	wire [1-1:0] node1589;
	wire [1-1:0] node1590;
	wire [1-1:0] node1592;
	wire [1-1:0] node1595;
	wire [1-1:0] node1596;
	wire [1-1:0] node1600;
	wire [1-1:0] node1601;
	wire [1-1:0] node1602;
	wire [1-1:0] node1604;
	wire [1-1:0] node1606;
	wire [1-1:0] node1609;
	wire [1-1:0] node1610;
	wire [1-1:0] node1612;
	wire [1-1:0] node1615;
	wire [1-1:0] node1616;
	wire [1-1:0] node1620;
	wire [1-1:0] node1621;
	wire [1-1:0] node1622;
	wire [1-1:0] node1624;
	wire [1-1:0] node1627;
	wire [1-1:0] node1628;
	wire [1-1:0] node1632;
	wire [1-1:0] node1633;
	wire [1-1:0] node1634;
	wire [1-1:0] node1639;
	wire [1-1:0] node1640;
	wire [1-1:0] node1641;
	wire [1-1:0] node1642;
	wire [1-1:0] node1644;
	wire [1-1:0] node1646;
	wire [1-1:0] node1648;
	wire [1-1:0] node1650;
	wire [1-1:0] node1653;
	wire [1-1:0] node1654;
	wire [1-1:0] node1656;
	wire [1-1:0] node1658;
	wire [1-1:0] node1660;
	wire [1-1:0] node1663;
	wire [1-1:0] node1664;
	wire [1-1:0] node1666;
	wire [1-1:0] node1668;
	wire [1-1:0] node1671;
	wire [1-1:0] node1672;
	wire [1-1:0] node1674;
	wire [1-1:0] node1678;
	wire [1-1:0] node1679;
	wire [1-1:0] node1680;
	wire [1-1:0] node1682;
	wire [1-1:0] node1684;
	wire [1-1:0] node1686;
	wire [1-1:0] node1689;
	wire [1-1:0] node1690;
	wire [1-1:0] node1692;
	wire [1-1:0] node1694;
	wire [1-1:0] node1697;
	wire [1-1:0] node1698;
	wire [1-1:0] node1700;
	wire [1-1:0] node1703;
	wire [1-1:0] node1704;
	wire [1-1:0] node1708;
	wire [1-1:0] node1709;
	wire [1-1:0] node1710;
	wire [1-1:0] node1712;
	wire [1-1:0] node1714;
	wire [1-1:0] node1717;
	wire [1-1:0] node1718;
	wire [1-1:0] node1720;
	wire [1-1:0] node1723;
	wire [1-1:0] node1724;
	wire [1-1:0] node1728;
	wire [1-1:0] node1729;
	wire [1-1:0] node1730;
	wire [1-1:0] node1732;
	wire [1-1:0] node1735;
	wire [1-1:0] node1736;
	wire [1-1:0] node1740;
	wire [1-1:0] node1741;
	wire [1-1:0] node1742;
	wire [1-1:0] node1747;
	wire [1-1:0] node1748;
	wire [1-1:0] node1749;
	wire [1-1:0] node1751;
	wire [1-1:0] node1752;
	wire [1-1:0] node1754;
	wire [1-1:0] node1756;
	wire [1-1:0] node1759;
	wire [1-1:0] node1760;
	wire [1-1:0] node1762;
	wire [1-1:0] node1765;
	wire [1-1:0] node1766;
	wire [1-1:0] node1770;
	wire [1-1:0] node1771;
	wire [1-1:0] node1772;
	wire [1-1:0] node1774;
	wire [1-1:0] node1776;
	wire [1-1:0] node1779;
	wire [1-1:0] node1780;
	wire [1-1:0] node1782;
	wire [1-1:0] node1785;
	wire [1-1:0] node1786;
	wire [1-1:0] node1790;
	wire [1-1:0] node1791;
	wire [1-1:0] node1792;
	wire [1-1:0] node1794;
	wire [1-1:0] node1797;
	wire [1-1:0] node1798;
	wire [1-1:0] node1802;
	wire [1-1:0] node1803;
	wire [1-1:0] node1807;
	wire [1-1:0] node1808;
	wire [1-1:0] node1809;
	wire [1-1:0] node1810;
	wire [1-1:0] node1812;
	wire [1-1:0] node1814;
	wire [1-1:0] node1817;
	wire [1-1:0] node1818;
	wire [1-1:0] node1820;
	wire [1-1:0] node1823;
	wire [1-1:0] node1824;
	wire [1-1:0] node1828;
	wire [1-1:0] node1829;
	wire [1-1:0] node1830;
	wire [1-1:0] node1832;
	wire [1-1:0] node1835;
	wire [1-1:0] node1836;
	wire [1-1:0] node1840;
	wire [1-1:0] node1841;
	wire [1-1:0] node1842;
	wire [1-1:0] node1847;
	wire [1-1:0] node1848;
	wire [1-1:0] node1849;
	wire [1-1:0] node1850;
	wire [1-1:0] node1852;
	wire [1-1:0] node1855;
	wire [1-1:0] node1856;
	wire [1-1:0] node1860;
	wire [1-1:0] node1861;
	wire [1-1:0] node1862;
	wire [1-1:0] node1867;
	wire [1-1:0] node1868;
	wire [1-1:0] node1869;
	wire [1-1:0] node1874;
	wire [1-1:0] node1875;
	wire [1-1:0] node1876;
	wire [1-1:0] node1877;
	wire [1-1:0] node1878;
	wire [1-1:0] node1880;
	wire [1-1:0] node1882;
	wire [1-1:0] node1884;
	wire [1-1:0] node1886;
	wire [1-1:0] node1889;
	wire [1-1:0] node1890;
	wire [1-1:0] node1892;
	wire [1-1:0] node1894;
	wire [1-1:0] node1897;
	wire [1-1:0] node1898;
	wire [1-1:0] node1900;
	wire [1-1:0] node1902;
	wire [1-1:0] node1905;
	wire [1-1:0] node1906;
	wire [1-1:0] node1908;
	wire [1-1:0] node1911;
	wire [1-1:0] node1912;
	wire [1-1:0] node1916;
	wire [1-1:0] node1917;
	wire [1-1:0] node1918;
	wire [1-1:0] node1920;
	wire [1-1:0] node1922;
	wire [1-1:0] node1924;
	wire [1-1:0] node1927;
	wire [1-1:0] node1928;
	wire [1-1:0] node1930;
	wire [1-1:0] node1932;
	wire [1-1:0] node1935;
	wire [1-1:0] node1936;
	wire [1-1:0] node1937;
	wire [1-1:0] node1940;
	wire [1-1:0] node1943;
	wire [1-1:0] node1944;
	wire [1-1:0] node1948;
	wire [1-1:0] node1949;
	wire [1-1:0] node1950;
	wire [1-1:0] node1952;
	wire [1-1:0] node1954;
	wire [1-1:0] node1957;
	wire [1-1:0] node1958;
	wire [1-1:0] node1960;
	wire [1-1:0] node1963;
	wire [1-1:0] node1964;
	wire [1-1:0] node1968;
	wire [1-1:0] node1969;
	wire [1-1:0] node1970;
	wire [1-1:0] node1972;
	wire [1-1:0] node1975;
	wire [1-1:0] node1976;
	wire [1-1:0] node1981;
	wire [1-1:0] node1982;
	wire [1-1:0] node1983;
	wire [1-1:0] node1984;
	wire [1-1:0] node1986;
	wire [1-1:0] node1988;
	wire [1-1:0] node1990;
	wire [1-1:0] node1993;
	wire [1-1:0] node1994;
	wire [1-1:0] node1996;
	wire [1-1:0] node1999;
	wire [1-1:0] node2000;
	wire [1-1:0] node2002;
	wire [1-1:0] node2005;
	wire [1-1:0] node2006;
	wire [1-1:0] node2010;
	wire [1-1:0] node2011;
	wire [1-1:0] node2012;
	wire [1-1:0] node2014;
	wire [1-1:0] node2016;
	wire [1-1:0] node2019;
	wire [1-1:0] node2020;
	wire [1-1:0] node2022;
	wire [1-1:0] node2025;
	wire [1-1:0] node2026;
	wire [1-1:0] node2030;
	wire [1-1:0] node2031;
	wire [1-1:0] node2032;
	wire [1-1:0] node2034;
	wire [1-1:0] node2037;
	wire [1-1:0] node2038;
	wire [1-1:0] node2043;
	wire [1-1:0] node2044;
	wire [1-1:0] node2045;
	wire [1-1:0] node2046;
	wire [1-1:0] node2048;
	wire [1-1:0] node2049;
	wire [1-1:0] node2053;
	wire [1-1:0] node2054;
	wire [1-1:0] node2057;
	wire [1-1:0] node2058;
	wire [1-1:0] node2062;
	wire [1-1:0] node2063;
	wire [1-1:0] node2064;
	wire [1-1:0] node2066;
	wire [1-1:0] node2069;
	wire [1-1:0] node2070;
	wire [1-1:0] node2073;
	wire [1-1:0] node2076;
	wire [1-1:0] node2077;
	wire [1-1:0] node2078;
	wire [1-1:0] node2083;
	wire [1-1:0] node2084;
	wire [1-1:0] node2085;
	wire [1-1:0] node2086;
	wire [1-1:0] node2088;
	wire [1-1:0] node2091;
	wire [1-1:0] node2092;
	wire [1-1:0] node2096;
	wire [1-1:0] node2097;
	wire [1-1:0] node2098;
	wire [1-1:0] node2103;
	wire [1-1:0] node2104;
	wire [1-1:0] node2105;
	wire [1-1:0] node2106;
	wire [1-1:0] node2112;
	wire [1-1:0] node2113;
	wire [1-1:0] node2114;
	wire [1-1:0] node2115;
	wire [1-1:0] node2116;
	wire [1-1:0] node2118;
	wire [1-1:0] node2120;
	wire [1-1:0] node2122;
	wire [1-1:0] node2125;
	wire [1-1:0] node2126;
	wire [1-1:0] node2128;
	wire [1-1:0] node2130;
	wire [1-1:0] node2133;
	wire [1-1:0] node2134;
	wire [1-1:0] node2136;
	wire [1-1:0] node2139;
	wire [1-1:0] node2140;
	wire [1-1:0] node2144;
	wire [1-1:0] node2145;
	wire [1-1:0] node2146;
	wire [1-1:0] node2148;
	wire [1-1:0] node2150;
	wire [1-1:0] node2153;
	wire [1-1:0] node2154;
	wire [1-1:0] node2156;
	wire [1-1:0] node2159;
	wire [1-1:0] node2160;
	wire [1-1:0] node2164;
	wire [1-1:0] node2165;
	wire [1-1:0] node2166;
	wire [1-1:0] node2168;
	wire [1-1:0] node2171;
	wire [1-1:0] node2172;
	wire [1-1:0] node2176;
	wire [1-1:0] node2177;
	wire [1-1:0] node2178;
	wire [1-1:0] node2183;
	wire [1-1:0] node2184;
	wire [1-1:0] node2185;
	wire [1-1:0] node2186;
	wire [1-1:0] node2188;
	wire [1-1:0] node2190;
	wire [1-1:0] node2193;
	wire [1-1:0] node2194;
	wire [1-1:0] node2196;
	wire [1-1:0] node2199;
	wire [1-1:0] node2200;
	wire [1-1:0] node2204;
	wire [1-1:0] node2205;
	wire [1-1:0] node2206;
	wire [1-1:0] node2207;
	wire [1-1:0] node2210;
	wire [1-1:0] node2213;
	wire [1-1:0] node2214;
	wire [1-1:0] node2218;
	wire [1-1:0] node2219;
	wire [1-1:0] node2220;
	wire [1-1:0] node2225;
	wire [1-1:0] node2226;
	wire [1-1:0] node2227;
	wire [1-1:0] node2229;
	wire [1-1:0] node2230;
	wire [1-1:0] node2234;
	wire [1-1:0] node2235;
	wire [1-1:0] node2236;
	wire [1-1:0] node2241;
	wire [1-1:0] node2242;
	wire [1-1:0] node2243;
	wire [1-1:0] node2248;
	wire [1-1:0] node2249;
	wire [1-1:0] node2250;
	wire [1-1:0] node2251;
	wire [1-1:0] node2252;
	wire [1-1:0] node2254;
	wire [1-1:0] node2256;
	wire [1-1:0] node2259;
	wire [1-1:0] node2260;
	wire [1-1:0] node2262;
	wire [1-1:0] node2265;
	wire [1-1:0] node2266;
	wire [1-1:0] node2270;
	wire [1-1:0] node2271;
	wire [1-1:0] node2272;
	wire [1-1:0] node2274;
	wire [1-1:0] node2277;
	wire [1-1:0] node2278;
	wire [1-1:0] node2282;
	wire [1-1:0] node2283;
	wire [1-1:0] node2284;
	wire [1-1:0] node2289;
	wire [1-1:0] node2290;
	wire [1-1:0] node2291;
	wire [1-1:0] node2292;
	wire [1-1:0] node2294;
	wire [1-1:0] node2297;
	wire [1-1:0] node2298;
	wire [1-1:0] node2302;
	wire [1-1:0] node2303;
	wire [1-1:0] node2304;
	wire [1-1:0] node2309;
	wire [1-1:0] node2310;
	wire [1-1:0] node2311;
	wire [1-1:0] node2316;
	wire [1-1:0] node2317;
	wire [1-1:0] node2318;
	wire [1-1:0] node2319;
	wire [1-1:0] node2320;
	wire [1-1:0] node2322;
	wire [1-1:0] node2325;
	wire [1-1:0] node2326;
	wire [1-1:0] node2330;
	wire [1-1:0] node2331;
	wire [1-1:0] node2332;
	wire [1-1:0] node2337;
	wire [1-1:0] node2338;
	wire [1-1:0] node2339;
	wire [1-1:0] node2340;
	wire [1-1:0] node2346;
	wire [1-1:0] node2347;
	wire [1-1:0] node2348;
	wire [1-1:0] node2349;
	wire [1-1:0] node2350;
	wire [1-1:0] node2357;
	wire [1-1:0] node2358;
	wire [1-1:0] node2359;
	wire [1-1:0] node2360;
	wire [1-1:0] node2361;
	wire [1-1:0] node2362;
	wire [1-1:0] node2364;
	wire [1-1:0] node2366;
	wire [1-1:0] node2368;
	wire [1-1:0] node2370;
	wire [1-1:0] node2373;
	wire [1-1:0] node2374;
	wire [1-1:0] node2376;
	wire [1-1:0] node2378;
	wire [1-1:0] node2380;
	wire [1-1:0] node2383;
	wire [1-1:0] node2384;
	wire [1-1:0] node2386;
	wire [1-1:0] node2388;
	wire [1-1:0] node2391;
	wire [1-1:0] node2392;
	wire [1-1:0] node2394;
	wire [1-1:0] node2397;
	wire [1-1:0] node2398;
	wire [1-1:0] node2402;
	wire [1-1:0] node2403;
	wire [1-1:0] node2404;
	wire [1-1:0] node2406;
	wire [1-1:0] node2408;
	wire [1-1:0] node2410;
	wire [1-1:0] node2413;
	wire [1-1:0] node2414;
	wire [1-1:0] node2416;
	wire [1-1:0] node2418;
	wire [1-1:0] node2421;
	wire [1-1:0] node2422;
	wire [1-1:0] node2424;
	wire [1-1:0] node2427;
	wire [1-1:0] node2428;
	wire [1-1:0] node2432;
	wire [1-1:0] node2433;
	wire [1-1:0] node2434;
	wire [1-1:0] node2436;
	wire [1-1:0] node2439;
	wire [1-1:0] node2440;
	wire [1-1:0] node2442;
	wire [1-1:0] node2445;
	wire [1-1:0] node2446;
	wire [1-1:0] node2450;
	wire [1-1:0] node2451;
	wire [1-1:0] node2452;
	wire [1-1:0] node2455;
	wire [1-1:0] node2456;
	wire [1-1:0] node2460;
	wire [1-1:0] node2461;
	wire [1-1:0] node2462;
	wire [1-1:0] node2467;
	wire [1-1:0] node2468;
	wire [1-1:0] node2469;
	wire [1-1:0] node2471;
	wire [1-1:0] node2472;
	wire [1-1:0] node2474;
	wire [1-1:0] node2476;
	wire [1-1:0] node2479;
	wire [1-1:0] node2480;
	wire [1-1:0] node2482;
	wire [1-1:0] node2485;
	wire [1-1:0] node2486;
	wire [1-1:0] node2490;
	wire [1-1:0] node2491;
	wire [1-1:0] node2492;
	wire [1-1:0] node2494;
	wire [1-1:0] node2496;
	wire [1-1:0] node2499;
	wire [1-1:0] node2500;
	wire [1-1:0] node2502;
	wire [1-1:0] node2505;
	wire [1-1:0] node2506;
	wire [1-1:0] node2510;
	wire [1-1:0] node2511;
	wire [1-1:0] node2512;
	wire [1-1:0] node2514;
	wire [1-1:0] node2517;
	wire [1-1:0] node2518;
	wire [1-1:0] node2522;
	wire [1-1:0] node2523;
	wire [1-1:0] node2524;
	wire [1-1:0] node2529;
	wire [1-1:0] node2530;
	wire [1-1:0] node2531;
	wire [1-1:0] node2532;
	wire [1-1:0] node2534;
	wire [1-1:0] node2536;
	wire [1-1:0] node2539;
	wire [1-1:0] node2540;
	wire [1-1:0] node2542;
	wire [1-1:0] node2545;
	wire [1-1:0] node2546;
	wire [1-1:0] node2550;
	wire [1-1:0] node2551;
	wire [1-1:0] node2552;
	wire [1-1:0] node2554;
	wire [1-1:0] node2557;
	wire [1-1:0] node2558;
	wire [1-1:0] node2562;
	wire [1-1:0] node2563;
	wire [1-1:0] node2564;
	wire [1-1:0] node2569;
	wire [1-1:0] node2570;
	wire [1-1:0] node2571;
	wire [1-1:0] node2572;
	wire [1-1:0] node2574;
	wire [1-1:0] node2577;
	wire [1-1:0] node2578;
	wire [1-1:0] node2582;
	wire [1-1:0] node2583;
	wire [1-1:0] node2584;
	wire [1-1:0] node2589;
	wire [1-1:0] node2590;
	wire [1-1:0] node2591;
	wire [1-1:0] node2596;
	wire [1-1:0] node2597;
	wire [1-1:0] node2598;
	wire [1-1:0] node2599;
	wire [1-1:0] node2600;
	wire [1-1:0] node2602;
	wire [1-1:0] node2604;
	wire [1-1:0] node2606;
	wire [1-1:0] node2609;
	wire [1-1:0] node2610;
	wire [1-1:0] node2612;
	wire [1-1:0] node2614;
	wire [1-1:0] node2617;
	wire [1-1:0] node2618;
	wire [1-1:0] node2620;
	wire [1-1:0] node2623;
	wire [1-1:0] node2624;
	wire [1-1:0] node2628;
	wire [1-1:0] node2629;
	wire [1-1:0] node2630;
	wire [1-1:0] node2632;
	wire [1-1:0] node2634;
	wire [1-1:0] node2637;
	wire [1-1:0] node2638;
	wire [1-1:0] node2640;
	wire [1-1:0] node2643;
	wire [1-1:0] node2644;
	wire [1-1:0] node2648;
	wire [1-1:0] node2649;
	wire [1-1:0] node2650;
	wire [1-1:0] node2652;
	wire [1-1:0] node2655;
	wire [1-1:0] node2656;
	wire [1-1:0] node2660;
	wire [1-1:0] node2661;
	wire [1-1:0] node2662;
	wire [1-1:0] node2667;
	wire [1-1:0] node2668;
	wire [1-1:0] node2669;
	wire [1-1:0] node2670;
	wire [1-1:0] node2672;
	wire [1-1:0] node2674;
	wire [1-1:0] node2677;
	wire [1-1:0] node2678;
	wire [1-1:0] node2680;
	wire [1-1:0] node2683;
	wire [1-1:0] node2684;
	wire [1-1:0] node2688;
	wire [1-1:0] node2689;
	wire [1-1:0] node2690;
	wire [1-1:0] node2692;
	wire [1-1:0] node2695;
	wire [1-1:0] node2696;
	wire [1-1:0] node2701;
	wire [1-1:0] node2702;
	wire [1-1:0] node2703;
	wire [1-1:0] node2704;
	wire [1-1:0] node2706;
	wire [1-1:0] node2709;
	wire [1-1:0] node2710;
	wire [1-1:0] node2714;
	wire [1-1:0] node2715;
	wire [1-1:0] node2716;
	wire [1-1:0] node2721;
	wire [1-1:0] node2722;
	wire [1-1:0] node2723;
	wire [1-1:0] node2724;
	wire [1-1:0] node2730;
	wire [1-1:0] node2731;
	wire [1-1:0] node2732;
	wire [1-1:0] node2733;
	wire [1-1:0] node2734;
	wire [1-1:0] node2736;
	wire [1-1:0] node2738;
	wire [1-1:0] node2741;
	wire [1-1:0] node2742;
	wire [1-1:0] node2744;
	wire [1-1:0] node2748;
	wire [1-1:0] node2749;
	wire [1-1:0] node2751;
	wire [1-1:0] node2752;
	wire [1-1:0] node2755;
	wire [1-1:0] node2758;
	wire [1-1:0] node2759;
	wire [1-1:0] node2760;
	wire [1-1:0] node2765;
	wire [1-1:0] node2766;
	wire [1-1:0] node2767;
	wire [1-1:0] node2768;
	wire [1-1:0] node2770;
	wire [1-1:0] node2773;
	wire [1-1:0] node2774;
	wire [1-1:0] node2778;
	wire [1-1:0] node2779;
	wire [1-1:0] node2784;
	wire [1-1:0] node2785;
	wire [1-1:0] node2786;
	wire [1-1:0] node2787;
	wire [1-1:0] node2788;
	wire [1-1:0] node2790;
	wire [1-1:0] node2793;
	wire [1-1:0] node2794;
	wire [1-1:0] node2798;
	wire [1-1:0] node2799;
	wire [1-1:0] node2800;
	wire [1-1:0] node2805;
	wire [1-1:0] node2806;
	wire [1-1:0] node2807;
	wire [1-1:0] node2808;
	wire [1-1:0] node2815;
	wire [1-1:0] node2816;
	wire [1-1:0] node2817;
	wire [1-1:0] node2818;
	wire [1-1:0] node2819;
	wire [1-1:0] node2820;
	wire [1-1:0] node2822;
	wire [1-1:0] node2824;
	wire [1-1:0] node2826;
	wire [1-1:0] node2829;
	wire [1-1:0] node2830;
	wire [1-1:0] node2832;
	wire [1-1:0] node2834;
	wire [1-1:0] node2837;
	wire [1-1:0] node2838;
	wire [1-1:0] node2840;
	wire [1-1:0] node2843;
	wire [1-1:0] node2844;
	wire [1-1:0] node2848;
	wire [1-1:0] node2849;
	wire [1-1:0] node2850;
	wire [1-1:0] node2852;
	wire [1-1:0] node2854;
	wire [1-1:0] node2857;
	wire [1-1:0] node2858;
	wire [1-1:0] node2860;
	wire [1-1:0] node2863;
	wire [1-1:0] node2864;
	wire [1-1:0] node2868;
	wire [1-1:0] node2869;
	wire [1-1:0] node2870;
	wire [1-1:0] node2872;
	wire [1-1:0] node2875;
	wire [1-1:0] node2876;
	wire [1-1:0] node2880;
	wire [1-1:0] node2881;
	wire [1-1:0] node2882;
	wire [1-1:0] node2887;
	wire [1-1:0] node2888;
	wire [1-1:0] node2889;
	wire [1-1:0] node2890;
	wire [1-1:0] node2892;
	wire [1-1:0] node2894;
	wire [1-1:0] node2897;
	wire [1-1:0] node2898;
	wire [1-1:0] node2900;
	wire [1-1:0] node2903;
	wire [1-1:0] node2904;
	wire [1-1:0] node2908;
	wire [1-1:0] node2909;
	wire [1-1:0] node2910;
	wire [1-1:0] node2912;
	wire [1-1:0] node2915;
	wire [1-1:0] node2916;
	wire [1-1:0] node2920;
	wire [1-1:0] node2921;
	wire [1-1:0] node2922;
	wire [1-1:0] node2927;
	wire [1-1:0] node2928;
	wire [1-1:0] node2929;
	wire [1-1:0] node2930;
	wire [1-1:0] node2932;
	wire [1-1:0] node2935;
	wire [1-1:0] node2936;
	wire [1-1:0] node2940;
	wire [1-1:0] node2941;
	wire [1-1:0] node2942;
	wire [1-1:0] node2947;
	wire [1-1:0] node2948;
	wire [1-1:0] node2949;
	wire [1-1:0] node2950;
	wire [1-1:0] node2956;
	wire [1-1:0] node2957;
	wire [1-1:0] node2958;
	wire [1-1:0] node2959;
	wire [1-1:0] node2960;
	wire [1-1:0] node2962;
	wire [1-1:0] node2964;
	wire [1-1:0] node2967;
	wire [1-1:0] node2968;
	wire [1-1:0] node2971;
	wire [1-1:0] node2972;
	wire [1-1:0] node2976;
	wire [1-1:0] node2977;
	wire [1-1:0] node2978;
	wire [1-1:0] node2980;
	wire [1-1:0] node2983;
	wire [1-1:0] node2984;
	wire [1-1:0] node2988;
	wire [1-1:0] node2989;
	wire [1-1:0] node2993;
	wire [1-1:0] node2994;
	wire [1-1:0] node2995;
	wire [1-1:0] node2996;
	wire [1-1:0] node2998;
	wire [1-1:0] node3001;
	wire [1-1:0] node3002;
	wire [1-1:0] node3006;
	wire [1-1:0] node3007;
	wire [1-1:0] node3008;
	wire [1-1:0] node3013;
	wire [1-1:0] node3014;
	wire [1-1:0] node3015;
	wire [1-1:0] node3016;
	wire [1-1:0] node3022;
	wire [1-1:0] node3023;
	wire [1-1:0] node3024;
	wire [1-1:0] node3025;
	wire [1-1:0] node3026;
	wire [1-1:0] node3028;
	wire [1-1:0] node3031;
	wire [1-1:0] node3032;
	wire [1-1:0] node3036;
	wire [1-1:0] node3037;
	wire [1-1:0] node3039;
	wire [1-1:0] node3043;
	wire [1-1:0] node3044;
	wire [1-1:0] node3045;
	wire [1-1:0] node3046;
	wire [1-1:0] node3052;
	wire [1-1:0] node3053;
	wire [1-1:0] node3054;
	wire [1-1:0] node3055;
	wire [1-1:0] node3056;
	wire [1-1:0] node3063;
	wire [1-1:0] node3064;
	wire [1-1:0] node3065;
	wire [1-1:0] node3066;
	wire [1-1:0] node3067;
	wire [1-1:0] node3068;
	wire [1-1:0] node3070;
	wire [1-1:0] node3073;
	wire [1-1:0] node3074;
	wire [1-1:0] node3076;
	wire [1-1:0] node3079;
	wire [1-1:0] node3080;
	wire [1-1:0] node3084;
	wire [1-1:0] node3085;
	wire [1-1:0] node3086;
	wire [1-1:0] node3088;
	wire [1-1:0] node3091;
	wire [1-1:0] node3092;
	wire [1-1:0] node3095;
	wire [1-1:0] node3098;
	wire [1-1:0] node3099;
	wire [1-1:0] node3103;
	wire [1-1:0] node3104;
	wire [1-1:0] node3105;
	wire [1-1:0] node3106;
	wire [1-1:0] node3108;
	wire [1-1:0] node3111;
	wire [1-1:0] node3112;
	wire [1-1:0] node3116;
	wire [1-1:0] node3117;
	wire [1-1:0] node3118;
	wire [1-1:0] node3123;
	wire [1-1:0] node3124;
	wire [1-1:0] node3125;
	wire [1-1:0] node3126;
	wire [1-1:0] node3132;
	wire [1-1:0] node3133;
	wire [1-1:0] node3134;
	wire [1-1:0] node3135;
	wire [1-1:0] node3136;
	wire [1-1:0] node3138;
	wire [1-1:0] node3141;
	wire [1-1:0] node3142;
	wire [1-1:0] node3146;
	wire [1-1:0] node3147;
	wire [1-1:0] node3148;
	wire [1-1:0] node3153;
	wire [1-1:0] node3154;
	wire [1-1:0] node3155;
	wire [1-1:0] node3157;
	wire [1-1:0] node3162;
	wire [1-1:0] node3163;
	wire [1-1:0] node3164;
	wire [1-1:0] node3165;
	wire [1-1:0] node3167;
	wire [1-1:0] node3173;
	wire [1-1:0] node3174;
	wire [1-1:0] node3175;
	wire [1-1:0] node3176;
	wire [1-1:0] node3177;
	wire [1-1:0] node3178;
	wire [1-1:0] node3180;
	wire [1-1:0] node3183;
	wire [1-1:0] node3184;
	wire [1-1:0] node3188;
	wire [1-1:0] node3189;
	wire [1-1:0] node3190;
	wire [1-1:0] node3195;
	wire [1-1:0] node3196;
	wire [1-1:0] node3197;
	wire [1-1:0] node3198;
	wire [1-1:0] node3204;
	wire [1-1:0] node3205;
	wire [1-1:0] node3206;
	wire [1-1:0] node3207;
	wire [1-1:0] node3208;
	wire [1-1:0] node3215;
	wire [1-1:0] node3217;
	wire [1-1:0] node3218;
	wire [1-1:0] node3219;
	wire [1-1:0] node3220;
	wire [1-1:0] node3221;
	wire [1-1:0] node3228;
	wire [1-1:0] node3229;
	wire [1-1:0] node3230;
	wire [1-1:0] node3231;
	wire [1-1:0] node3232;
	wire [1-1:0] node3233;
	wire [1-1:0] node3234;
	wire [1-1:0] node3236;
	wire [1-1:0] node3238;
	wire [1-1:0] node3240;
	wire [1-1:0] node3242;
	wire [1-1:0] node3244;
	wire [1-1:0] node3247;
	wire [1-1:0] node3248;
	wire [1-1:0] node3250;
	wire [1-1:0] node3252;
	wire [1-1:0] node3254;
	wire [1-1:0] node3256;
	wire [1-1:0] node3259;
	wire [1-1:0] node3260;
	wire [1-1:0] node3262;
	wire [1-1:0] node3264;
	wire [1-1:0] node3266;
	wire [1-1:0] node3269;
	wire [1-1:0] node3270;
	wire [1-1:0] node3272;
	wire [1-1:0] node3274;
	wire [1-1:0] node3277;
	wire [1-1:0] node3278;
	wire [1-1:0] node3280;
	wire [1-1:0] node3283;
	wire [1-1:0] node3284;
	wire [1-1:0] node3288;
	wire [1-1:0] node3289;
	wire [1-1:0] node3290;
	wire [1-1:0] node3292;
	wire [1-1:0] node3294;
	wire [1-1:0] node3296;
	wire [1-1:0] node3298;
	wire [1-1:0] node3301;
	wire [1-1:0] node3302;
	wire [1-1:0] node3304;
	wire [1-1:0] node3306;
	wire [1-1:0] node3308;
	wire [1-1:0] node3311;
	wire [1-1:0] node3312;
	wire [1-1:0] node3314;
	wire [1-1:0] node3316;
	wire [1-1:0] node3319;
	wire [1-1:0] node3320;
	wire [1-1:0] node3322;
	wire [1-1:0] node3325;
	wire [1-1:0] node3326;
	wire [1-1:0] node3330;
	wire [1-1:0] node3331;
	wire [1-1:0] node3332;
	wire [1-1:0] node3334;
	wire [1-1:0] node3336;
	wire [1-1:0] node3338;
	wire [1-1:0] node3341;
	wire [1-1:0] node3342;
	wire [1-1:0] node3344;
	wire [1-1:0] node3346;
	wire [1-1:0] node3349;
	wire [1-1:0] node3350;
	wire [1-1:0] node3352;
	wire [1-1:0] node3356;
	wire [1-1:0] node3357;
	wire [1-1:0] node3358;
	wire [1-1:0] node3359;
	wire [1-1:0] node3361;
	wire [1-1:0] node3365;
	wire [1-1:0] node3366;
	wire [1-1:0] node3368;
	wire [1-1:0] node3371;
	wire [1-1:0] node3372;
	wire [1-1:0] node3376;
	wire [1-1:0] node3377;
	wire [1-1:0] node3379;
	wire [1-1:0] node3380;
	wire [1-1:0] node3384;
	wire [1-1:0] node3385;
	wire [1-1:0] node3386;
	wire [1-1:0] node3391;
	wire [1-1:0] node3392;
	wire [1-1:0] node3393;
	wire [1-1:0] node3394;
	wire [1-1:0] node3396;
	wire [1-1:0] node3398;
	wire [1-1:0] node3400;
	wire [1-1:0] node3402;
	wire [1-1:0] node3405;
	wire [1-1:0] node3406;
	wire [1-1:0] node3408;
	wire [1-1:0] node3410;
	wire [1-1:0] node3412;
	wire [1-1:0] node3415;
	wire [1-1:0] node3416;
	wire [1-1:0] node3418;
	wire [1-1:0] node3420;
	wire [1-1:0] node3423;
	wire [1-1:0] node3424;
	wire [1-1:0] node3426;
	wire [1-1:0] node3430;
	wire [1-1:0] node3431;
	wire [1-1:0] node3432;
	wire [1-1:0] node3434;
	wire [1-1:0] node3436;
	wire [1-1:0] node3439;
	wire [1-1:0] node3440;
	wire [1-1:0] node3442;
	wire [1-1:0] node3444;
	wire [1-1:0] node3447;
	wire [1-1:0] node3448;
	wire [1-1:0] node3450;
	wire [1-1:0] node3453;
	wire [1-1:0] node3454;
	wire [1-1:0] node3458;
	wire [1-1:0] node3459;
	wire [1-1:0] node3460;
	wire [1-1:0] node3462;
	wire [1-1:0] node3465;
	wire [1-1:0] node3466;
	wire [1-1:0] node3468;
	wire [1-1:0] node3471;
	wire [1-1:0] node3472;
	wire [1-1:0] node3476;
	wire [1-1:0] node3477;
	wire [1-1:0] node3478;
	wire [1-1:0] node3480;
	wire [1-1:0] node3483;
	wire [1-1:0] node3484;
	wire [1-1:0] node3488;
	wire [1-1:0] node3489;
	wire [1-1:0] node3493;
	wire [1-1:0] node3494;
	wire [1-1:0] node3495;
	wire [1-1:0] node3497;
	wire [1-1:0] node3498;
	wire [1-1:0] node3500;
	wire [1-1:0] node3502;
	wire [1-1:0] node3505;
	wire [1-1:0] node3506;
	wire [1-1:0] node3508;
	wire [1-1:0] node3511;
	wire [1-1:0] node3512;
	wire [1-1:0] node3516;
	wire [1-1:0] node3517;
	wire [1-1:0] node3518;
	wire [1-1:0] node3520;
	wire [1-1:0] node3521;
	wire [1-1:0] node3524;
	wire [1-1:0] node3527;
	wire [1-1:0] node3528;
	wire [1-1:0] node3530;
	wire [1-1:0] node3533;
	wire [1-1:0] node3534;
	wire [1-1:0] node3538;
	wire [1-1:0] node3539;
	wire [1-1:0] node3540;
	wire [1-1:0] node3543;
	wire [1-1:0] node3544;
	wire [1-1:0] node3548;
	wire [1-1:0] node3549;
	wire [1-1:0] node3550;
	wire [1-1:0] node3555;
	wire [1-1:0] node3556;
	wire [1-1:0] node3557;
	wire [1-1:0] node3559;
	wire [1-1:0] node3561;
	wire [1-1:0] node3562;
	wire [1-1:0] node3566;
	wire [1-1:0] node3567;
	wire [1-1:0] node3568;
	wire [1-1:0] node3570;
	wire [1-1:0] node3573;
	wire [1-1:0] node3574;
	wire [1-1:0] node3578;
	wire [1-1:0] node3579;
	wire [1-1:0] node3580;
	wire [1-1:0] node3585;
	wire [1-1:0] node3586;
	wire [1-1:0] node3587;
	wire [1-1:0] node3588;
	wire [1-1:0] node3590;
	wire [1-1:0] node3593;
	wire [1-1:0] node3594;
	wire [1-1:0] node3598;
	wire [1-1:0] node3599;
	wire [1-1:0] node3600;
	wire [1-1:0] node3606;
	wire [1-1:0] node3607;
	wire [1-1:0] node3608;
	wire [1-1:0] node3609;
	wire [1-1:0] node3610;
	wire [1-1:0] node3612;
	wire [1-1:0] node3614;
	wire [1-1:0] node3616;
	wire [1-1:0] node3618;
	wire [1-1:0] node3621;
	wire [1-1:0] node3622;
	wire [1-1:0] node3624;
	wire [1-1:0] node3626;
	wire [1-1:0] node3628;
	wire [1-1:0] node3631;
	wire [1-1:0] node3632;
	wire [1-1:0] node3634;
	wire [1-1:0] node3635;
	wire [1-1:0] node3638;
	wire [1-1:0] node3641;
	wire [1-1:0] node3642;
	wire [1-1:0] node3644;
	wire [1-1:0] node3647;
	wire [1-1:0] node3648;
	wire [1-1:0] node3652;
	wire [1-1:0] node3653;
	wire [1-1:0] node3654;
	wire [1-1:0] node3656;
	wire [1-1:0] node3658;
	wire [1-1:0] node3660;
	wire [1-1:0] node3663;
	wire [1-1:0] node3664;
	wire [1-1:0] node3666;
	wire [1-1:0] node3668;
	wire [1-1:0] node3671;
	wire [1-1:0] node3672;
	wire [1-1:0] node3674;
	wire [1-1:0] node3678;
	wire [1-1:0] node3679;
	wire [1-1:0] node3680;
	wire [1-1:0] node3682;
	wire [1-1:0] node3685;
	wire [1-1:0] node3686;
	wire [1-1:0] node3688;
	wire [1-1:0] node3691;
	wire [1-1:0] node3692;
	wire [1-1:0] node3696;
	wire [1-1:0] node3697;
	wire [1-1:0] node3698;
	wire [1-1:0] node3700;
	wire [1-1:0] node3703;
	wire [1-1:0] node3704;
	wire [1-1:0] node3707;
	wire [1-1:0] node3710;
	wire [1-1:0] node3711;
	wire [1-1:0] node3712;
	wire [1-1:0] node3717;
	wire [1-1:0] node3718;
	wire [1-1:0] node3719;
	wire [1-1:0] node3720;
	wire [1-1:0] node3722;
	wire [1-1:0] node3724;
	wire [1-1:0] node3726;
	wire [1-1:0] node3729;
	wire [1-1:0] node3730;
	wire [1-1:0] node3732;
	wire [1-1:0] node3734;
	wire [1-1:0] node3737;
	wire [1-1:0] node3738;
	wire [1-1:0] node3740;
	wire [1-1:0] node3743;
	wire [1-1:0] node3744;
	wire [1-1:0] node3748;
	wire [1-1:0] node3749;
	wire [1-1:0] node3750;
	wire [1-1:0] node3752;
	wire [1-1:0] node3754;
	wire [1-1:0] node3757;
	wire [1-1:0] node3758;
	wire [1-1:0] node3761;
	wire [1-1:0] node3762;
	wire [1-1:0] node3766;
	wire [1-1:0] node3767;
	wire [1-1:0] node3768;
	wire [1-1:0] node3770;
	wire [1-1:0] node3775;
	wire [1-1:0] node3776;
	wire [1-1:0] node3777;
	wire [1-1:0] node3778;
	wire [1-1:0] node3780;
	wire [1-1:0] node3782;
	wire [1-1:0] node3785;
	wire [1-1:0] node3786;
	wire [1-1:0] node3788;
	wire [1-1:0] node3791;
	wire [1-1:0] node3792;
	wire [1-1:0] node3796;
	wire [1-1:0] node3797;
	wire [1-1:0] node3798;
	wire [1-1:0] node3800;
	wire [1-1:0] node3803;
	wire [1-1:0] node3804;
	wire [1-1:0] node3808;
	wire [1-1:0] node3809;
	wire [1-1:0] node3811;
	wire [1-1:0] node3815;
	wire [1-1:0] node3816;
	wire [1-1:0] node3817;
	wire [1-1:0] node3818;
	wire [1-1:0] node3820;
	wire [1-1:0] node3823;
	wire [1-1:0] node3824;
	wire [1-1:0] node3828;
	wire [1-1:0] node3829;
	wire [1-1:0] node3830;
	wire [1-1:0] node3835;
	wire [1-1:0] node3836;
	wire [1-1:0] node3837;
	wire [1-1:0] node3838;
	wire [1-1:0] node3844;
	wire [1-1:0] node3845;
	wire [1-1:0] node3846;
	wire [1-1:0] node3847;
	wire [1-1:0] node3848;
	wire [1-1:0] node3850;
	wire [1-1:0] node3852;
	wire [1-1:0] node3854;
	wire [1-1:0] node3857;
	wire [1-1:0] node3858;
	wire [1-1:0] node3860;
	wire [1-1:0] node3862;
	wire [1-1:0] node3865;
	wire [1-1:0] node3866;
	wire [1-1:0] node3868;
	wire [1-1:0] node3871;
	wire [1-1:0] node3872;
	wire [1-1:0] node3876;
	wire [1-1:0] node3877;
	wire [1-1:0] node3878;
	wire [1-1:0] node3880;
	wire [1-1:0] node3882;
	wire [1-1:0] node3885;
	wire [1-1:0] node3886;
	wire [1-1:0] node3888;
	wire [1-1:0] node3892;
	wire [1-1:0] node3893;
	wire [1-1:0] node3894;
	wire [1-1:0] node3896;
	wire [1-1:0] node3899;
	wire [1-1:0] node3900;
	wire [1-1:0] node3904;
	wire [1-1:0] node3905;
	wire [1-1:0] node3906;
	wire [1-1:0] node3911;
	wire [1-1:0] node3912;
	wire [1-1:0] node3913;
	wire [1-1:0] node3914;
	wire [1-1:0] node3916;
	wire [1-1:0] node3918;
	wire [1-1:0] node3921;
	wire [1-1:0] node3922;
	wire [1-1:0] node3924;
	wire [1-1:0] node3928;
	wire [1-1:0] node3929;
	wire [1-1:0] node3930;
	wire [1-1:0] node3932;
	wire [1-1:0] node3935;
	wire [1-1:0] node3936;
	wire [1-1:0] node3940;
	wire [1-1:0] node3941;
	wire [1-1:0] node3942;
	wire [1-1:0] node3947;
	wire [1-1:0] node3948;
	wire [1-1:0] node3949;
	wire [1-1:0] node3950;
	wire [1-1:0] node3952;
	wire [1-1:0] node3955;
	wire [1-1:0] node3957;
	wire [1-1:0] node3960;
	wire [1-1:0] node3961;
	wire [1-1:0] node3962;
	wire [1-1:0] node3967;
	wire [1-1:0] node3968;
	wire [1-1:0] node3969;
	wire [1-1:0] node3970;
	wire [1-1:0] node3976;
	wire [1-1:0] node3977;
	wire [1-1:0] node3978;
	wire [1-1:0] node3979;
	wire [1-1:0] node3980;
	wire [1-1:0] node3982;
	wire [1-1:0] node3984;
	wire [1-1:0] node3987;
	wire [1-1:0] node3988;
	wire [1-1:0] node3990;
	wire [1-1:0] node3994;
	wire [1-1:0] node3995;
	wire [1-1:0] node3996;
	wire [1-1:0] node3998;
	wire [1-1:0] node4001;
	wire [1-1:0] node4002;
	wire [1-1:0] node4006;
	wire [1-1:0] node4007;
	wire [1-1:0] node4009;
	wire [1-1:0] node4013;
	wire [1-1:0] node4014;
	wire [1-1:0] node4015;
	wire [1-1:0] node4016;
	wire [1-1:0] node4018;
	wire [1-1:0] node4021;
	wire [1-1:0] node4023;
	wire [1-1:0] node4026;
	wire [1-1:0] node4027;
	wire [1-1:0] node4029;
	wire [1-1:0] node4033;
	wire [1-1:0] node4034;
	wire [1-1:0] node4035;
	wire [1-1:0] node4036;
	wire [1-1:0] node4042;
	wire [1-1:0] node4043;
	wire [1-1:0] node4044;
	wire [1-1:0] node4045;
	wire [1-1:0] node4046;
	wire [1-1:0] node4048;
	wire [1-1:0] node4051;
	wire [1-1:0] node4052;
	wire [1-1:0] node4056;
	wire [1-1:0] node4057;
	wire [1-1:0] node4058;
	wire [1-1:0] node4063;
	wire [1-1:0] node4064;
	wire [1-1:0] node4065;
	wire [1-1:0] node4070;
	wire [1-1:0] node4071;
	wire [1-1:0] node4072;
	wire [1-1:0] node4073;
	wire [1-1:0] node4074;
	wire [1-1:0] node4081;
	wire [1-1:0] node4082;
	wire [1-1:0] node4083;
	wire [1-1:0] node4084;
	wire [1-1:0] node4085;
	wire [1-1:0] node4086;
	wire [1-1:0] node4088;
	wire [1-1:0] node4090;
	wire [1-1:0] node4092;
	wire [1-1:0] node4094;
	wire [1-1:0] node4097;
	wire [1-1:0] node4098;
	wire [1-1:0] node4100;
	wire [1-1:0] node4102;
	wire [1-1:0] node4105;
	wire [1-1:0] node4106;
	wire [1-1:0] node4108;
	wire [1-1:0] node4110;
	wire [1-1:0] node4113;
	wire [1-1:0] node4114;
	wire [1-1:0] node4118;
	wire [1-1:0] node4119;
	wire [1-1:0] node4120;
	wire [1-1:0] node4122;
	wire [1-1:0] node4124;
	wire [1-1:0] node4126;
	wire [1-1:0] node4129;
	wire [1-1:0] node4130;
	wire [1-1:0] node4132;
	wire [1-1:0] node4134;
	wire [1-1:0] node4137;
	wire [1-1:0] node4138;
	wire [1-1:0] node4140;
	wire [1-1:0] node4143;
	wire [1-1:0] node4144;
	wire [1-1:0] node4148;
	wire [1-1:0] node4149;
	wire [1-1:0] node4151;
	wire [1-1:0] node4152;
	wire [1-1:0] node4154;
	wire [1-1:0] node4157;
	wire [1-1:0] node4158;
	wire [1-1:0] node4162;
	wire [1-1:0] node4163;
	wire [1-1:0] node4164;
	wire [1-1:0] node4166;
	wire [1-1:0] node4169;
	wire [1-1:0] node4170;
	wire [1-1:0] node4174;
	wire [1-1:0] node4175;
	wire [1-1:0] node4176;
	wire [1-1:0] node4181;
	wire [1-1:0] node4182;
	wire [1-1:0] node4183;
	wire [1-1:0] node4184;
	wire [1-1:0] node4186;
	wire [1-1:0] node4188;
	wire [1-1:0] node4190;
	wire [1-1:0] node4193;
	wire [1-1:0] node4194;
	wire [1-1:0] node4196;
	wire [1-1:0] node4198;
	wire [1-1:0] node4201;
	wire [1-1:0] node4202;
	wire [1-1:0] node4204;
	wire [1-1:0] node4208;
	wire [1-1:0] node4209;
	wire [1-1:0] node4210;
	wire [1-1:0] node4212;
	wire [1-1:0] node4215;
	wire [1-1:0] node4216;
	wire [1-1:0] node4218;
	wire [1-1:0] node4221;
	wire [1-1:0] node4222;
	wire [1-1:0] node4226;
	wire [1-1:0] node4227;
	wire [1-1:0] node4228;
	wire [1-1:0] node4230;
	wire [1-1:0] node4233;
	wire [1-1:0] node4234;
	wire [1-1:0] node4239;
	wire [1-1:0] node4240;
	wire [1-1:0] node4241;
	wire [1-1:0] node4243;
	wire [1-1:0] node4244;
	wire [1-1:0] node4246;
	wire [1-1:0] node4249;
	wire [1-1:0] node4250;
	wire [1-1:0] node4254;
	wire [1-1:0] node4255;
	wire [1-1:0] node4256;
	wire [1-1:0] node4258;
	wire [1-1:0] node4261;
	wire [1-1:0] node4262;
	wire [1-1:0] node4267;
	wire [1-1:0] node4268;
	wire [1-1:0] node4269;
	wire [1-1:0] node4270;
	wire [1-1:0] node4272;
	wire [1-1:0] node4275;
	wire [1-1:0] node4276;
	wire [1-1:0] node4280;
	wire [1-1:0] node4281;
	wire [1-1:0] node4282;
	wire [1-1:0] node4287;
	wire [1-1:0] node4288;
	wire [1-1:0] node4289;
	wire [1-1:0] node4290;
	wire [1-1:0] node4296;
	wire [1-1:0] node4297;
	wire [1-1:0] node4298;
	wire [1-1:0] node4299;
	wire [1-1:0] node4300;
	wire [1-1:0] node4302;
	wire [1-1:0] node4304;
	wire [1-1:0] node4307;
	wire [1-1:0] node4308;
	wire [1-1:0] node4310;
	wire [1-1:0] node4312;
	wire [1-1:0] node4315;
	wire [1-1:0] node4316;
	wire [1-1:0] node4319;
	wire [1-1:0] node4320;
	wire [1-1:0] node4324;
	wire [1-1:0] node4325;
	wire [1-1:0] node4326;
	wire [1-1:0] node4328;
	wire [1-1:0] node4330;
	wire [1-1:0] node4333;
	wire [1-1:0] node4334;
	wire [1-1:0] node4336;
	wire [1-1:0] node4339;
	wire [1-1:0] node4340;
	wire [1-1:0] node4344;
	wire [1-1:0] node4345;
	wire [1-1:0] node4346;
	wire [1-1:0] node4348;
	wire [1-1:0] node4351;
	wire [1-1:0] node4352;
	wire [1-1:0] node4357;
	wire [1-1:0] node4358;
	wire [1-1:0] node4359;
	wire [1-1:0] node4360;
	wire [1-1:0] node4362;
	wire [1-1:0] node4364;
	wire [1-1:0] node4367;
	wire [1-1:0] node4368;
	wire [1-1:0] node4370;
	wire [1-1:0] node4373;
	wire [1-1:0] node4374;
	wire [1-1:0] node4378;
	wire [1-1:0] node4379;
	wire [1-1:0] node4380;
	wire [1-1:0] node4382;
	wire [1-1:0] node4385;
	wire [1-1:0] node4386;
	wire [1-1:0] node4390;
	wire [1-1:0] node4391;
	wire [1-1:0] node4392;
	wire [1-1:0] node4397;
	wire [1-1:0] node4398;
	wire [1-1:0] node4399;
	wire [1-1:0] node4400;
	wire [1-1:0] node4402;
	wire [1-1:0] node4405;
	wire [1-1:0] node4406;
	wire [1-1:0] node4409;
	wire [1-1:0] node4412;
	wire [1-1:0] node4413;
	wire [1-1:0] node4414;
	wire [1-1:0] node4419;
	wire [1-1:0] node4420;
	wire [1-1:0] node4421;
	wire [1-1:0] node4422;
	wire [1-1:0] node4428;
	wire [1-1:0] node4429;
	wire [1-1:0] node4430;
	wire [1-1:0] node4431;
	wire [1-1:0] node4432;
	wire [1-1:0] node4434;
	wire [1-1:0] node4436;
	wire [1-1:0] node4439;
	wire [1-1:0] node4440;
	wire [1-1:0] node4442;
	wire [1-1:0] node4445;
	wire [1-1:0] node4446;
	wire [1-1:0] node4450;
	wire [1-1:0] node4451;
	wire [1-1:0] node4452;
	wire [1-1:0] node4454;
	wire [1-1:0] node4457;
	wire [1-1:0] node4458;
	wire [1-1:0] node4462;
	wire [1-1:0] node4463;
	wire [1-1:0] node4464;
	wire [1-1:0] node4469;
	wire [1-1:0] node4470;
	wire [1-1:0] node4471;
	wire [1-1:0] node4472;
	wire [1-1:0] node4474;
	wire [1-1:0] node4477;
	wire [1-1:0] node4478;
	wire [1-1:0] node4482;
	wire [1-1:0] node4483;
	wire [1-1:0] node4484;
	wire [1-1:0] node4489;
	wire [1-1:0] node4490;
	wire [1-1:0] node4491;
	wire [1-1:0] node4492;
	wire [1-1:0] node4498;
	wire [1-1:0] node4499;
	wire [1-1:0] node4500;
	wire [1-1:0] node4501;
	wire [1-1:0] node4502;
	wire [1-1:0] node4504;
	wire [1-1:0] node4507;
	wire [1-1:0] node4508;
	wire [1-1:0] node4512;
	wire [1-1:0] node4513;
	wire [1-1:0] node4514;
	wire [1-1:0] node4519;
	wire [1-1:0] node4520;
	wire [1-1:0] node4521;
	wire [1-1:0] node4522;
	wire [1-1:0] node4528;
	wire [1-1:0] node4529;
	wire [1-1:0] node4530;
	wire [1-1:0] node4531;
	wire [1-1:0] node4532;
	wire [1-1:0] node4539;
	wire [1-1:0] node4540;
	wire [1-1:0] node4541;
	wire [1-1:0] node4542;
	wire [1-1:0] node4543;
	wire [1-1:0] node4544;
	wire [1-1:0] node4546;
	wire [1-1:0] node4548;
	wire [1-1:0] node4550;
	wire [1-1:0] node4553;
	wire [1-1:0] node4554;
	wire [1-1:0] node4556;
	wire [1-1:0] node4558;
	wire [1-1:0] node4561;
	wire [1-1:0] node4562;
	wire [1-1:0] node4564;
	wire [1-1:0] node4567;
	wire [1-1:0] node4568;
	wire [1-1:0] node4572;
	wire [1-1:0] node4573;
	wire [1-1:0] node4574;
	wire [1-1:0] node4576;
	wire [1-1:0] node4578;
	wire [1-1:0] node4581;
	wire [1-1:0] node4582;
	wire [1-1:0] node4584;
	wire [1-1:0] node4587;
	wire [1-1:0] node4588;
	wire [1-1:0] node4592;
	wire [1-1:0] node4593;
	wire [1-1:0] node4594;
	wire [1-1:0] node4595;
	wire [1-1:0] node4598;
	wire [1-1:0] node4601;
	wire [1-1:0] node4604;
	wire [1-1:0] node4605;
	wire [1-1:0] node4606;
	wire [1-1:0] node4611;
	wire [1-1:0] node4612;
	wire [1-1:0] node4613;
	wire [1-1:0] node4614;
	wire [1-1:0] node4616;
	wire [1-1:0] node4618;
	wire [1-1:0] node4621;
	wire [1-1:0] node4622;
	wire [1-1:0] node4624;
	wire [1-1:0] node4627;
	wire [1-1:0] node4628;
	wire [1-1:0] node4632;
	wire [1-1:0] node4633;
	wire [1-1:0] node4634;
	wire [1-1:0] node4636;
	wire [1-1:0] node4639;
	wire [1-1:0] node4642;
	wire [1-1:0] node4643;
	wire [1-1:0] node4644;
	wire [1-1:0] node4649;
	wire [1-1:0] node4650;
	wire [1-1:0] node4651;
	wire [1-1:0] node4652;
	wire [1-1:0] node4654;
	wire [1-1:0] node4657;
	wire [1-1:0] node4658;
	wire [1-1:0] node4662;
	wire [1-1:0] node4663;
	wire [1-1:0] node4664;
	wire [1-1:0] node4669;
	wire [1-1:0] node4670;
	wire [1-1:0] node4671;
	wire [1-1:0] node4672;
	wire [1-1:0] node4678;
	wire [1-1:0] node4679;
	wire [1-1:0] node4680;
	wire [1-1:0] node4681;
	wire [1-1:0] node4682;
	wire [1-1:0] node4684;
	wire [1-1:0] node4686;
	wire [1-1:0] node4689;
	wire [1-1:0] node4690;
	wire [1-1:0] node4692;
	wire [1-1:0] node4695;
	wire [1-1:0] node4696;
	wire [1-1:0] node4700;
	wire [1-1:0] node4701;
	wire [1-1:0] node4702;
	wire [1-1:0] node4705;
	wire [1-1:0] node4706;
	wire [1-1:0] node4710;
	wire [1-1:0] node4711;
	wire [1-1:0] node4712;
	wire [1-1:0] node4717;
	wire [1-1:0] node4718;
	wire [1-1:0] node4719;
	wire [1-1:0] node4720;
	wire [1-1:0] node4722;
	wire [1-1:0] node4725;
	wire [1-1:0] node4726;
	wire [1-1:0] node4730;
	wire [1-1:0] node4731;
	wire [1-1:0] node4732;
	wire [1-1:0] node4737;
	wire [1-1:0] node4738;
	wire [1-1:0] node4739;
	wire [1-1:0] node4740;
	wire [1-1:0] node4746;
	wire [1-1:0] node4747;
	wire [1-1:0] node4748;
	wire [1-1:0] node4749;
	wire [1-1:0] node4750;
	wire [1-1:0] node4752;
	wire [1-1:0] node4755;
	wire [1-1:0] node4756;
	wire [1-1:0] node4760;
	wire [1-1:0] node4761;
	wire [1-1:0] node4765;
	wire [1-1:0] node4766;
	wire [1-1:0] node4767;
	wire [1-1:0] node4768;
	wire [1-1:0] node4774;
	wire [1-1:0] node4775;
	wire [1-1:0] node4776;
	wire [1-1:0] node4777;
	wire [1-1:0] node4778;
	wire [1-1:0] node4785;
	wire [1-1:0] node4786;
	wire [1-1:0] node4787;
	wire [1-1:0] node4788;
	wire [1-1:0] node4789;
	wire [1-1:0] node4790;
	wire [1-1:0] node4792;
	wire [1-1:0] node4794;
	wire [1-1:0] node4797;
	wire [1-1:0] node4798;
	wire [1-1:0] node4800;
	wire [1-1:0] node4803;
	wire [1-1:0] node4804;
	wire [1-1:0] node4808;
	wire [1-1:0] node4809;
	wire [1-1:0] node4810;
	wire [1-1:0] node4812;
	wire [1-1:0] node4815;
	wire [1-1:0] node4816;
	wire [1-1:0] node4820;
	wire [1-1:0] node4821;
	wire [1-1:0] node4822;
	wire [1-1:0] node4827;
	wire [1-1:0] node4828;
	wire [1-1:0] node4829;
	wire [1-1:0] node4830;
	wire [1-1:0] node4832;
	wire [1-1:0] node4835;
	wire [1-1:0] node4836;
	wire [1-1:0] node4840;
	wire [1-1:0] node4841;
	wire [1-1:0] node4842;
	wire [1-1:0] node4847;
	wire [1-1:0] node4848;
	wire [1-1:0] node4849;
	wire [1-1:0] node4850;
	wire [1-1:0] node4856;
	wire [1-1:0] node4857;
	wire [1-1:0] node4858;
	wire [1-1:0] node4859;
	wire [1-1:0] node4861;
	wire [1-1:0] node4862;
	wire [1-1:0] node4866;
	wire [1-1:0] node4867;
	wire [1-1:0] node4869;
	wire [1-1:0] node4873;
	wire [1-1:0] node4874;
	wire [1-1:0] node4875;
	wire [1-1:0] node4876;
	wire [1-1:0] node4883;
	wire [1-1:0] node4884;
	wire [1-1:0] node4885;
	wire [1-1:0] node4886;
	wire [1-1:0] node4887;
	wire [1-1:0] node4888;
	wire [1-1:0] node4890;
	wire [1-1:0] node4893;
	wire [1-1:0] node4894;
	wire [1-1:0] node4898;
	wire [1-1:0] node4899;
	wire [1-1:0] node4900;
	wire [1-1:0] node4905;
	wire [1-1:0] node4906;
	wire [1-1:0] node4907;
	wire [1-1:0] node4912;
	wire [1-1:0] node4913;
	wire [1-1:0] node4914;
	wire [1-1:0] node4915;
	wire [1-1:0] node4921;
	wire [1-1:0] node4922;
	wire [1-1:0] node4923;
	wire [1-1:0] node4924;
	wire [1-1:0] node4925;
	wire [1-1:0] node4926;
	wire [1-1:0] node4934;
	wire [1-1:0] node4935;
	wire [1-1:0] node4936;
	wire [1-1:0] node4937;
	wire [1-1:0] node4938;
	wire [1-1:0] node4939;
	wire [1-1:0] node4940;
	wire [1-1:0] node4942;
	wire [1-1:0] node4944;
	wire [1-1:0] node4946;
	wire [1-1:0] node4948;
	wire [1-1:0] node4951;
	wire [1-1:0] node4952;
	wire [1-1:0] node4954;
	wire [1-1:0] node4956;
	wire [1-1:0] node4958;
	wire [1-1:0] node4961;
	wire [1-1:0] node4962;
	wire [1-1:0] node4964;
	wire [1-1:0] node4966;
	wire [1-1:0] node4969;
	wire [1-1:0] node4970;
	wire [1-1:0] node4972;
	wire [1-1:0] node4975;
	wire [1-1:0] node4976;
	wire [1-1:0] node4980;
	wire [1-1:0] node4981;
	wire [1-1:0] node4982;
	wire [1-1:0] node4984;
	wire [1-1:0] node4986;
	wire [1-1:0] node4988;
	wire [1-1:0] node4991;
	wire [1-1:0] node4992;
	wire [1-1:0] node4994;
	wire [1-1:0] node4996;
	wire [1-1:0] node4999;
	wire [1-1:0] node5000;
	wire [1-1:0] node5001;
	wire [1-1:0] node5005;
	wire [1-1:0] node5006;
	wire [1-1:0] node5010;
	wire [1-1:0] node5011;
	wire [1-1:0] node5012;
	wire [1-1:0] node5014;
	wire [1-1:0] node5016;
	wire [1-1:0] node5019;
	wire [1-1:0] node5020;
	wire [1-1:0] node5022;
	wire [1-1:0] node5025;
	wire [1-1:0] node5026;
	wire [1-1:0] node5030;
	wire [1-1:0] node5031;
	wire [1-1:0] node5032;
	wire [1-1:0] node5034;
	wire [1-1:0] node5037;
	wire [1-1:0] node5038;
	wire [1-1:0] node5042;
	wire [1-1:0] node5043;
	wire [1-1:0] node5044;
	wire [1-1:0] node5049;
	wire [1-1:0] node5050;
	wire [1-1:0] node5051;
	wire [1-1:0] node5052;
	wire [1-1:0] node5054;
	wire [1-1:0] node5056;
	wire [1-1:0] node5058;
	wire [1-1:0] node5061;
	wire [1-1:0] node5062;
	wire [1-1:0] node5064;
	wire [1-1:0] node5066;
	wire [1-1:0] node5069;
	wire [1-1:0] node5070;
	wire [1-1:0] node5072;
	wire [1-1:0] node5075;
	wire [1-1:0] node5076;
	wire [1-1:0] node5080;
	wire [1-1:0] node5081;
	wire [1-1:0] node5082;
	wire [1-1:0] node5084;
	wire [1-1:0] node5086;
	wire [1-1:0] node5089;
	wire [1-1:0] node5090;
	wire [1-1:0] node5092;
	wire [1-1:0] node5096;
	wire [1-1:0] node5097;
	wire [1-1:0] node5098;
	wire [1-1:0] node5100;
	wire [1-1:0] node5103;
	wire [1-1:0] node5104;
	wire [1-1:0] node5108;
	wire [1-1:0] node5109;
	wire [1-1:0] node5110;
	wire [1-1:0] node5115;
	wire [1-1:0] node5116;
	wire [1-1:0] node5117;
	wire [1-1:0] node5118;
	wire [1-1:0] node5120;
	wire [1-1:0] node5122;
	wire [1-1:0] node5125;
	wire [1-1:0] node5126;
	wire [1-1:0] node5127;
	wire [1-1:0] node5130;
	wire [1-1:0] node5134;
	wire [1-1:0] node5135;
	wire [1-1:0] node5136;
	wire [1-1:0] node5138;
	wire [1-1:0] node5141;
	wire [1-1:0] node5144;
	wire [1-1:0] node5145;
	wire [1-1:0] node5146;
	wire [1-1:0] node5151;
	wire [1-1:0] node5152;
	wire [1-1:0] node5153;
	wire [1-1:0] node5154;
	wire [1-1:0] node5156;
	wire [1-1:0] node5159;
	wire [1-1:0] node5160;
	wire [1-1:0] node5164;
	wire [1-1:0] node5165;
	wire [1-1:0] node5166;
	wire [1-1:0] node5171;
	wire [1-1:0] node5172;
	wire [1-1:0] node5173;
	wire [1-1:0] node5174;
	wire [1-1:0] node5180;
	wire [1-1:0] node5181;
	wire [1-1:0] node5182;
	wire [1-1:0] node5183;
	wire [1-1:0] node5185;
	wire [1-1:0] node5186;
	wire [1-1:0] node5188;
	wire [1-1:0] node5190;
	wire [1-1:0] node5193;
	wire [1-1:0] node5194;
	wire [1-1:0] node5196;
	wire [1-1:0] node5200;
	wire [1-1:0] node5201;
	wire [1-1:0] node5202;
	wire [1-1:0] node5204;
	wire [1-1:0] node5206;
	wire [1-1:0] node5209;
	wire [1-1:0] node5210;
	wire [1-1:0] node5212;
	wire [1-1:0] node5215;
	wire [1-1:0] node5216;
	wire [1-1:0] node5220;
	wire [1-1:0] node5221;
	wire [1-1:0] node5222;
	wire [1-1:0] node5224;
	wire [1-1:0] node5227;
	wire [1-1:0] node5228;
	wire [1-1:0] node5232;
	wire [1-1:0] node5233;
	wire [1-1:0] node5234;
	wire [1-1:0] node5239;
	wire [1-1:0] node5240;
	wire [1-1:0] node5241;
	wire [1-1:0] node5243;
	wire [1-1:0] node5244;
	wire [1-1:0] node5246;
	wire [1-1:0] node5249;
	wire [1-1:0] node5250;
	wire [1-1:0] node5254;
	wire [1-1:0] node5255;
	wire [1-1:0] node5256;
	wire [1-1:0] node5258;
	wire [1-1:0] node5261;
	wire [1-1:0] node5262;
	wire [1-1:0] node5266;
	wire [1-1:0] node5267;
	wire [1-1:0] node5268;
	wire [1-1:0] node5273;
	wire [1-1:0] node5274;
	wire [1-1:0] node5275;
	wire [1-1:0] node5276;
	wire [1-1:0] node5278;
	wire [1-1:0] node5281;
	wire [1-1:0] node5282;
	wire [1-1:0] node5286;
	wire [1-1:0] node5287;
	wire [1-1:0] node5288;
	wire [1-1:0] node5293;
	wire [1-1:0] node5294;
	wire [1-1:0] node5295;
	wire [1-1:0] node5296;
	wire [1-1:0] node5302;
	wire [1-1:0] node5303;
	wire [1-1:0] node5304;
	wire [1-1:0] node5305;
	wire [1-1:0] node5306;
	wire [1-1:0] node5308;
	wire [1-1:0] node5310;
	wire [1-1:0] node5313;
	wire [1-1:0] node5314;
	wire [1-1:0] node5316;
	wire [1-1:0] node5319;
	wire [1-1:0] node5320;
	wire [1-1:0] node5324;
	wire [1-1:0] node5325;
	wire [1-1:0] node5326;
	wire [1-1:0] node5328;
	wire [1-1:0] node5331;
	wire [1-1:0] node5332;
	wire [1-1:0] node5336;
	wire [1-1:0] node5337;
	wire [1-1:0] node5338;
	wire [1-1:0] node5343;
	wire [1-1:0] node5344;
	wire [1-1:0] node5345;
	wire [1-1:0] node5346;
	wire [1-1:0] node5348;
	wire [1-1:0] node5351;
	wire [1-1:0] node5352;
	wire [1-1:0] node5356;
	wire [1-1:0] node5357;
	wire [1-1:0] node5358;
	wire [1-1:0] node5363;
	wire [1-1:0] node5364;
	wire [1-1:0] node5365;
	wire [1-1:0] node5366;
	wire [1-1:0] node5372;
	wire [1-1:0] node5373;
	wire [1-1:0] node5374;
	wire [1-1:0] node5375;
	wire [1-1:0] node5377;
	wire [1-1:0] node5378;
	wire [1-1:0] node5382;
	wire [1-1:0] node5383;
	wire [1-1:0] node5384;
	wire [1-1:0] node5389;
	wire [1-1:0] node5390;
	wire [1-1:0] node5391;
	wire [1-1:0] node5392;
	wire [1-1:0] node5398;
	wire [1-1:0] node5399;
	wire [1-1:0] node5400;
	wire [1-1:0] node5401;
	wire [1-1:0] node5402;
	wire [1-1:0] node5409;
	wire [1-1:0] node5410;
	wire [1-1:0] node5411;
	wire [1-1:0] node5412;
	wire [1-1:0] node5413;
	wire [1-1:0] node5414;
	wire [1-1:0] node5416;
	wire [1-1:0] node5418;
	wire [1-1:0] node5420;
	wire [1-1:0] node5423;
	wire [1-1:0] node5424;
	wire [1-1:0] node5426;
	wire [1-1:0] node5428;
	wire [1-1:0] node5431;
	wire [1-1:0] node5432;
	wire [1-1:0] node5434;
	wire [1-1:0] node5437;
	wire [1-1:0] node5438;
	wire [1-1:0] node5442;
	wire [1-1:0] node5443;
	wire [1-1:0] node5444;
	wire [1-1:0] node5446;
	wire [1-1:0] node5448;
	wire [1-1:0] node5451;
	wire [1-1:0] node5452;
	wire [1-1:0] node5454;
	wire [1-1:0] node5457;
	wire [1-1:0] node5458;
	wire [1-1:0] node5462;
	wire [1-1:0] node5463;
	wire [1-1:0] node5464;
	wire [1-1:0] node5466;
	wire [1-1:0] node5469;
	wire [1-1:0] node5470;
	wire [1-1:0] node5474;
	wire [1-1:0] node5475;
	wire [1-1:0] node5476;
	wire [1-1:0] node5481;
	wire [1-1:0] node5482;
	wire [1-1:0] node5483;
	wire [1-1:0] node5484;
	wire [1-1:0] node5486;
	wire [1-1:0] node5488;
	wire [1-1:0] node5491;
	wire [1-1:0] node5492;
	wire [1-1:0] node5494;
	wire [1-1:0] node5497;
	wire [1-1:0] node5498;
	wire [1-1:0] node5502;
	wire [1-1:0] node5503;
	wire [1-1:0] node5504;
	wire [1-1:0] node5506;
	wire [1-1:0] node5509;
	wire [1-1:0] node5510;
	wire [1-1:0] node5514;
	wire [1-1:0] node5515;
	wire [1-1:0] node5516;
	wire [1-1:0] node5521;
	wire [1-1:0] node5522;
	wire [1-1:0] node5523;
	wire [1-1:0] node5524;
	wire [1-1:0] node5526;
	wire [1-1:0] node5529;
	wire [1-1:0] node5530;
	wire [1-1:0] node5534;
	wire [1-1:0] node5535;
	wire [1-1:0] node5536;
	wire [1-1:0] node5541;
	wire [1-1:0] node5542;
	wire [1-1:0] node5543;
	wire [1-1:0] node5544;
	wire [1-1:0] node5550;
	wire [1-1:0] node5551;
	wire [1-1:0] node5552;
	wire [1-1:0] node5553;
	wire [1-1:0] node5554;
	wire [1-1:0] node5556;
	wire [1-1:0] node5558;
	wire [1-1:0] node5561;
	wire [1-1:0] node5563;
	wire [1-1:0] node5564;
	wire [1-1:0] node5568;
	wire [1-1:0] node5569;
	wire [1-1:0] node5570;
	wire [1-1:0] node5572;
	wire [1-1:0] node5575;
	wire [1-1:0] node5576;
	wire [1-1:0] node5580;
	wire [1-1:0] node5581;
	wire [1-1:0] node5582;
	wire [1-1:0] node5587;
	wire [1-1:0] node5588;
	wire [1-1:0] node5589;
	wire [1-1:0] node5591;
	wire [1-1:0] node5592;
	wire [1-1:0] node5596;
	wire [1-1:0] node5597;
	wire [1-1:0] node5598;
	wire [1-1:0] node5603;
	wire [1-1:0] node5604;
	wire [1-1:0] node5605;
	wire [1-1:0] node5606;
	wire [1-1:0] node5612;
	wire [1-1:0] node5613;
	wire [1-1:0] node5614;
	wire [1-1:0] node5615;
	wire [1-1:0] node5616;
	wire [1-1:0] node5618;
	wire [1-1:0] node5621;
	wire [1-1:0] node5622;
	wire [1-1:0] node5626;
	wire [1-1:0] node5627;
	wire [1-1:0] node5628;
	wire [1-1:0] node5633;
	wire [1-1:0] node5634;
	wire [1-1:0] node5635;
	wire [1-1:0] node5641;
	wire [1-1:0] node5642;
	wire [1-1:0] node5643;
	wire [1-1:0] node5644;
	wire [1-1:0] node5645;
	wire [1-1:0] node5646;
	wire [1-1:0] node5648;
	wire [1-1:0] node5650;
	wire [1-1:0] node5653;
	wire [1-1:0] node5654;
	wire [1-1:0] node5656;
	wire [1-1:0] node5659;
	wire [1-1:0] node5660;
	wire [1-1:0] node5664;
	wire [1-1:0] node5665;
	wire [1-1:0] node5666;
	wire [1-1:0] node5668;
	wire [1-1:0] node5671;
	wire [1-1:0] node5672;
	wire [1-1:0] node5677;
	wire [1-1:0] node5678;
	wire [1-1:0] node5679;
	wire [1-1:0] node5681;
	wire [1-1:0] node5682;
	wire [1-1:0] node5686;
	wire [1-1:0] node5687;
	wire [1-1:0] node5688;
	wire [1-1:0] node5693;
	wire [1-1:0] node5694;
	wire [1-1:0] node5695;
	wire [1-1:0] node5696;
	wire [1-1:0] node5702;
	wire [1-1:0] node5703;
	wire [1-1:0] node5704;
	wire [1-1:0] node5705;
	wire [1-1:0] node5706;
	wire [1-1:0] node5708;
	wire [1-1:0] node5711;
	wire [1-1:0] node5712;
	wire [1-1:0] node5716;
	wire [1-1:0] node5717;
	wire [1-1:0] node5718;
	wire [1-1:0] node5723;
	wire [1-1:0] node5724;
	wire [1-1:0] node5725;
	wire [1-1:0] node5726;
	wire [1-1:0] node5732;
	wire [1-1:0] node5733;
	wire [1-1:0] node5734;
	wire [1-1:0] node5735;
	wire [1-1:0] node5736;
	wire [1-1:0] node5743;
	wire [1-1:0] node5744;
	wire [1-1:0] node5745;
	wire [1-1:0] node5746;
	wire [1-1:0] node5747;
	wire [1-1:0] node5748;
	wire [1-1:0] node5750;
	wire [1-1:0] node5753;
	wire [1-1:0] node5754;
	wire [1-1:0] node5758;
	wire [1-1:0] node5759;
	wire [1-1:0] node5760;
	wire [1-1:0] node5765;
	wire [1-1:0] node5766;
	wire [1-1:0] node5767;
	wire [1-1:0] node5768;
	wire [1-1:0] node5774;
	wire [1-1:0] node5775;
	wire [1-1:0] node5776;
	wire [1-1:0] node5777;
	wire [1-1:0] node5778;
	wire [1-1:0] node5785;
	wire [1-1:0] node5786;
	wire [1-1:0] node5787;
	wire [1-1:0] node5788;
	wire [1-1:0] node5789;
	wire [1-1:0] node5796;
	wire [1-1:0] node5797;
	wire [1-1:0] node5798;
	wire [1-1:0] node5799;
	wire [1-1:0] node5800;
	wire [1-1:0] node5801;
	wire [1-1:0] node5802;
	wire [1-1:0] node5804;
	wire [1-1:0] node5806;
	wire [1-1:0] node5808;
	wire [1-1:0] node5811;
	wire [1-1:0] node5812;
	wire [1-1:0] node5814;
	wire [1-1:0] node5816;
	wire [1-1:0] node5819;
	wire [1-1:0] node5820;
	wire [1-1:0] node5822;
	wire [1-1:0] node5825;
	wire [1-1:0] node5826;
	wire [1-1:0] node5830;
	wire [1-1:0] node5831;
	wire [1-1:0] node5833;
	wire [1-1:0] node5834;
	wire [1-1:0] node5836;
	wire [1-1:0] node5839;
	wire [1-1:0] node5840;
	wire [1-1:0] node5844;
	wire [1-1:0] node5845;
	wire [1-1:0] node5847;
	wire [1-1:0] node5848;
	wire [1-1:0] node5852;
	wire [1-1:0] node5853;
	wire [1-1:0] node5854;
	wire [1-1:0] node5859;
	wire [1-1:0] node5860;
	wire [1-1:0] node5861;
	wire [1-1:0] node5863;
	wire [1-1:0] node5864;
	wire [1-1:0] node5866;
	wire [1-1:0] node5869;
	wire [1-1:0] node5870;
	wire [1-1:0] node5874;
	wire [1-1:0] node5875;
	wire [1-1:0] node5876;
	wire [1-1:0] node5878;
	wire [1-1:0] node5881;
	wire [1-1:0] node5882;
	wire [1-1:0] node5886;
	wire [1-1:0] node5887;
	wire [1-1:0] node5889;
	wire [1-1:0] node5893;
	wire [1-1:0] node5894;
	wire [1-1:0] node5895;
	wire [1-1:0] node5897;
	wire [1-1:0] node5898;
	wire [1-1:0] node5902;
	wire [1-1:0] node5903;
	wire [1-1:0] node5904;
	wire [1-1:0] node5907;
	wire [1-1:0] node5911;
	wire [1-1:0] node5912;
	wire [1-1:0] node5913;
	wire [1-1:0] node5914;
	wire [1-1:0] node5920;
	wire [1-1:0] node5921;
	wire [1-1:0] node5922;
	wire [1-1:0] node5923;
	wire [1-1:0] node5924;
	wire [1-1:0] node5926;
	wire [1-1:0] node5928;
	wire [1-1:0] node5931;
	wire [1-1:0] node5932;
	wire [1-1:0] node5934;
	wire [1-1:0] node5937;
	wire [1-1:0] node5938;
	wire [1-1:0] node5942;
	wire [1-1:0] node5943;
	wire [1-1:0] node5944;
	wire [1-1:0] node5946;
	wire [1-1:0] node5949;
	wire [1-1:0] node5950;
	wire [1-1:0] node5954;
	wire [1-1:0] node5955;
	wire [1-1:0] node5959;
	wire [1-1:0] node5960;
	wire [1-1:0] node5961;
	wire [1-1:0] node5963;
	wire [1-1:0] node5964;
	wire [1-1:0] node5968;
	wire [1-1:0] node5969;
	wire [1-1:0] node5970;
	wire [1-1:0] node5975;
	wire [1-1:0] node5976;
	wire [1-1:0] node5977;
	wire [1-1:0] node5978;
	wire [1-1:0] node5984;
	wire [1-1:0] node5985;
	wire [1-1:0] node5986;
	wire [1-1:0] node5987;
	wire [1-1:0] node5989;
	wire [1-1:0] node5990;
	wire [1-1:0] node5994;
	wire [1-1:0] node5995;
	wire [1-1:0] node5996;
	wire [1-1:0] node6001;
	wire [1-1:0] node6002;
	wire [1-1:0] node6003;
	wire [1-1:0] node6004;
	wire [1-1:0] node6010;
	wire [1-1:0] node6011;
	wire [1-1:0] node6012;
	wire [1-1:0] node6013;
	wire [1-1:0] node6014;
	wire [1-1:0] node6021;
	wire [1-1:0] node6022;
	wire [1-1:0] node6023;
	wire [1-1:0] node6024;
	wire [1-1:0] node6025;
	wire [1-1:0] node6026;
	wire [1-1:0] node6028;
	wire [1-1:0] node6030;
	wire [1-1:0] node6033;
	wire [1-1:0] node6034;
	wire [1-1:0] node6036;
	wire [1-1:0] node6040;
	wire [1-1:0] node6041;
	wire [1-1:0] node6042;
	wire [1-1:0] node6044;
	wire [1-1:0] node6047;
	wire [1-1:0] node6048;
	wire [1-1:0] node6052;
	wire [1-1:0] node6053;
	wire [1-1:0] node6054;
	wire [1-1:0] node6059;
	wire [1-1:0] node6060;
	wire [1-1:0] node6061;
	wire [1-1:0] node6062;
	wire [1-1:0] node6064;
	wire [1-1:0] node6067;
	wire [1-1:0] node6068;
	wire [1-1:0] node6072;
	wire [1-1:0] node6073;
	wire [1-1:0] node6074;
	wire [1-1:0] node6079;
	wire [1-1:0] node6080;
	wire [1-1:0] node6081;
	wire [1-1:0] node6086;
	wire [1-1:0] node6087;
	wire [1-1:0] node6088;
	wire [1-1:0] node6089;
	wire [1-1:0] node6090;
	wire [1-1:0] node6092;
	wire [1-1:0] node6095;
	wire [1-1:0] node6096;
	wire [1-1:0] node6100;
	wire [1-1:0] node6101;
	wire [1-1:0] node6102;
	wire [1-1:0] node6107;
	wire [1-1:0] node6108;
	wire [1-1:0] node6109;
	wire [1-1:0] node6110;
	wire [1-1:0] node6117;
	wire [1-1:0] node6118;
	wire [1-1:0] node6119;
	wire [1-1:0] node6120;
	wire [1-1:0] node6121;
	wire [1-1:0] node6122;
	wire [1-1:0] node6124;
	wire [1-1:0] node6127;
	wire [1-1:0] node6128;
	wire [1-1:0] node6131;
	wire [1-1:0] node6134;
	wire [1-1:0] node6135;
	wire [1-1:0] node6136;
	wire [1-1:0] node6141;
	wire [1-1:0] node6142;
	wire [1-1:0] node6143;
	wire [1-1:0] node6148;
	wire [1-1:0] node6149;
	wire [1-1:0] node6150;
	wire [1-1:0] node6151;
	wire [1-1:0] node6152;
	wire [1-1:0] node6159;
	wire [1-1:0] node6160;
	wire [1-1:0] node6161;
	wire [1-1:0] node6162;
	wire [1-1:0] node6163;
	wire [1-1:0] node6164;
	wire [1-1:0] node6172;
	wire [1-1:0] node6173;
	wire [1-1:0] node6174;
	wire [1-1:0] node6175;
	wire [1-1:0] node6176;
	wire [1-1:0] node6177;
	wire [1-1:0] node6178;
	wire [1-1:0] node6180;
	wire [1-1:0] node6182;
	wire [1-1:0] node6185;
	wire [1-1:0] node6187;
	wire [1-1:0] node6188;
	wire [1-1:0] node6192;
	wire [1-1:0] node6193;
	wire [1-1:0] node6194;
	wire [1-1:0] node6196;
	wire [1-1:0] node6199;
	wire [1-1:0] node6200;
	wire [1-1:0] node6204;
	wire [1-1:0] node6205;
	wire [1-1:0] node6206;
	wire [1-1:0] node6211;
	wire [1-1:0] node6212;
	wire [1-1:0] node6213;
	wire [1-1:0] node6214;
	wire [1-1:0] node6216;
	wire [1-1:0] node6219;
	wire [1-1:0] node6220;
	wire [1-1:0] node6224;
	wire [1-1:0] node6225;
	wire [1-1:0] node6226;
	wire [1-1:0] node6231;
	wire [1-1:0] node6232;
	wire [1-1:0] node6233;
	wire [1-1:0] node6234;
	wire [1-1:0] node6240;
	wire [1-1:0] node6241;
	wire [1-1:0] node6242;
	wire [1-1:0] node6243;
	wire [1-1:0] node6244;
	wire [1-1:0] node6246;
	wire [1-1:0] node6249;
	wire [1-1:0] node6250;
	wire [1-1:0] node6254;
	wire [1-1:0] node6255;
	wire [1-1:0] node6256;
	wire [1-1:0] node6261;
	wire [1-1:0] node6262;
	wire [1-1:0] node6263;
	wire [1-1:0] node6264;
	wire [1-1:0] node6270;
	wire [1-1:0] node6271;
	wire [1-1:0] node6272;
	wire [1-1:0] node6273;
	wire [1-1:0] node6279;
	wire [1-1:0] node6280;
	wire [1-1:0] node6281;
	wire [1-1:0] node6282;
	wire [1-1:0] node6283;
	wire [1-1:0] node6284;
	wire [1-1:0] node6286;
	wire [1-1:0] node6289;
	wire [1-1:0] node6290;
	wire [1-1:0] node6294;
	wire [1-1:0] node6295;
	wire [1-1:0] node6296;
	wire [1-1:0] node6301;
	wire [1-1:0] node6302;
	wire [1-1:0] node6303;
	wire [1-1:0] node6304;
	wire [1-1:0] node6310;
	wire [1-1:0] node6311;
	wire [1-1:0] node6312;
	wire [1-1:0] node6313;
	wire [1-1:0] node6314;
	wire [1-1:0] node6321;
	wire [1-1:0] node6322;
	wire [1-1:0] node6323;
	wire [1-1:0] node6324;
	wire [1-1:0] node6325;
	wire [1-1:0] node6326;
	wire [1-1:0] node6334;
	wire [1-1:0] node6335;
	wire [1-1:0] node6336;
	wire [1-1:0] node6337;
	wire [1-1:0] node6338;
	wire [1-1:0] node6339;
	wire [1-1:0] node6341;
	wire [1-1:0] node6343;
	wire [1-1:0] node6346;
	wire [1-1:0] node6347;
	wire [1-1:0] node6348;
	wire [1-1:0] node6353;
	wire [1-1:0] node6354;
	wire [1-1:0] node6355;
	wire [1-1:0] node6356;
	wire [1-1:0] node6362;
	wire [1-1:0] node6363;
	wire [1-1:0] node6364;
	wire [1-1:0] node6365;
	wire [1-1:0] node6366;
	wire [1-1:0] node6373;
	wire [1-1:0] node6374;
	wire [1-1:0] node6375;
	wire [1-1:0] node6376;
	wire [1-1:0] node6377;
	wire [1-1:0] node6384;
	wire [1-1:0] node6385;
	wire [1-1:0] node6386;
	wire [1-1:0] node6387;
	wire [1-1:0] node6388;
	wire [1-1:0] node6389;

	assign outp = (inp[1]) ? node3228 : node1;
		assign node1 = (inp[6]) ? node1473 : node2;
			assign node2 = (inp[0]) ? node602 : node3;
				assign node3 = (inp[12]) ? node227 : node4;
					assign node4 = (inp[14]) ? node70 : node5;
						assign node5 = (inp[4]) ? node19 : node6;
							assign node6 = (inp[13]) ? node8 : 1'b1;
								assign node8 = (inp[11]) ? node10 : 1'b1;
									assign node10 = (inp[10]) ? node12 : 1'b1;
										assign node12 = (inp[5]) ? node14 : 1'b1;
											assign node14 = (inp[8]) ? node16 : 1'b1;
												assign node16 = (inp[2]) ? 1'b0 : 1'b1;
							assign node19 = (inp[13]) ? node33 : node20;
								assign node20 = (inp[7]) ? node22 : 1'b1;
									assign node22 = (inp[9]) ? node24 : 1'b1;
										assign node24 = (inp[2]) ? node26 : 1'b1;
											assign node26 = (inp[5]) ? node28 : 1'b1;
												assign node28 = (inp[11]) ? node30 : 1'b1;
													assign node30 = (inp[10]) ? 1'b0 : 1'b1;
								assign node33 = (inp[3]) ? node45 : node34;
									assign node34 = (inp[11]) ? node36 : 1'b1;
										assign node36 = (inp[5]) ? node38 : 1'b1;
											assign node38 = (inp[2]) ? node40 : 1'b1;
												assign node40 = (inp[8]) ? 1'b0 : node41;
													assign node41 = (inp[9]) ? 1'b0 : 1'b1;
									assign node45 = (inp[9]) ? node55 : node46;
										assign node46 = (inp[11]) ? node48 : 1'b1;
											assign node48 = (inp[8]) ? node50 : 1'b1;
												assign node50 = (inp[5]) ? node52 : 1'b1;
													assign node52 = (inp[10]) ? 1'b0 : 1'b1;
										assign node55 = (inp[7]) ? node63 : node56;
											assign node56 = (inp[2]) ? node58 : 1'b1;
												assign node58 = (inp[10]) ? node60 : 1'b1;
													assign node60 = (inp[11]) ? 1'b0 : 1'b1;
											assign node63 = (inp[2]) ? 1'b0 : node64;
												assign node64 = (inp[11]) ? node66 : 1'b1;
													assign node66 = (inp[5]) ? 1'b0 : 1'b1;
						assign node70 = (inp[9]) ? node124 : node71;
							assign node71 = (inp[11]) ? node83 : node72;
								assign node72 = (inp[2]) ? node74 : 1'b1;
									assign node74 = (inp[4]) ? node76 : 1'b1;
										assign node76 = (inp[10]) ? node78 : 1'b1;
											assign node78 = (inp[5]) ? node80 : 1'b1;
												assign node80 = (inp[13]) ? 1'b0 : 1'b1;
								assign node83 = (inp[4]) ? node95 : node84;
									assign node84 = (inp[10]) ? node86 : 1'b1;
										assign node86 = (inp[5]) ? node88 : 1'b1;
											assign node88 = (inp[13]) ? node90 : 1'b1;
												assign node90 = (inp[3]) ? node92 : 1'b1;
													assign node92 = (inp[8]) ? 1'b0 : 1'b1;
									assign node95 = (inp[8]) ? node105 : node96;
										assign node96 = (inp[7]) ? node98 : 1'b1;
											assign node98 = (inp[13]) ? node100 : 1'b1;
												assign node100 = (inp[10]) ? node102 : 1'b1;
													assign node102 = (inp[3]) ? 1'b0 : 1'b0;
										assign node105 = (inp[10]) ? node113 : node106;
											assign node106 = (inp[13]) ? node108 : 1'b1;
												assign node108 = (inp[5]) ? node110 : 1'b1;
													assign node110 = (inp[2]) ? 1'b0 : 1'b1;
											assign node113 = (inp[3]) ? node119 : node114;
												assign node114 = (inp[7]) ? node116 : 1'b1;
													assign node116 = (inp[2]) ? 1'b0 : 1'b1;
												assign node119 = (inp[7]) ? 1'b0 : node120;
													assign node120 = (inp[2]) ? 1'b0 : 1'b0;
							assign node124 = (inp[10]) ? node166 : node125;
								assign node125 = (inp[7]) ? node137 : node126;
									assign node126 = (inp[5]) ? node128 : 1'b1;
										assign node128 = (inp[8]) ? node130 : 1'b1;
											assign node130 = (inp[11]) ? node132 : 1'b1;
												assign node132 = (inp[4]) ? 1'b0 : node133;
													assign node133 = (inp[3]) ? 1'b1 : 1'b1;
									assign node137 = (inp[3]) ? node147 : node138;
										assign node138 = (inp[5]) ? node140 : 1'b1;
											assign node140 = (inp[13]) ? node142 : 1'b1;
												assign node142 = (inp[4]) ? node144 : 1'b1;
													assign node144 = (inp[8]) ? 1'b0 : 1'b1;
										assign node147 = (inp[2]) ? node155 : node148;
											assign node148 = (inp[4]) ? node150 : 1'b1;
												assign node150 = (inp[11]) ? node152 : 1'b1;
													assign node152 = (inp[13]) ? 1'b0 : 1'b1;
											assign node155 = (inp[13]) ? node161 : node156;
												assign node156 = (inp[5]) ? node158 : 1'b1;
													assign node158 = (inp[11]) ? 1'b0 : 1'b1;
												assign node161 = (inp[4]) ? 1'b0 : node162;
													assign node162 = (inp[8]) ? 1'b0 : 1'b1;
								assign node166 = (inp[8]) ? node194 : node167;
									assign node167 = (inp[7]) ? node177 : node168;
										assign node168 = (inp[11]) ? node170 : 1'b1;
											assign node170 = (inp[3]) ? node172 : 1'b1;
												assign node172 = (inp[4]) ? node174 : 1'b1;
													assign node174 = (inp[5]) ? 1'b0 : 1'b1;
										assign node177 = (inp[3]) ? node187 : node178;
											assign node178 = (inp[13]) ? node180 : 1'b1;
												assign node180 = (inp[11]) ? node184 : node181;
													assign node181 = (inp[2]) ? 1'b1 : 1'b1;
													assign node184 = (inp[5]) ? 1'b0 : 1'b1;
											assign node187 = (inp[5]) ? node189 : 1'b1;
												assign node189 = (inp[4]) ? 1'b0 : node190;
													assign node190 = (inp[13]) ? 1'b0 : 1'b1;
									assign node194 = (inp[2]) ? node208 : node195;
										assign node195 = (inp[7]) ? node197 : 1'b1;
											assign node197 = (inp[5]) ? node203 : node198;
												assign node198 = (inp[11]) ? node200 : 1'b1;
													assign node200 = (inp[3]) ? 1'b0 : 1'b1;
												assign node203 = (inp[13]) ? 1'b0 : node204;
													assign node204 = (inp[4]) ? 1'b0 : 1'b1;
										assign node208 = (inp[13]) ? node220 : node209;
											assign node209 = (inp[4]) ? node215 : node210;
												assign node210 = (inp[5]) ? node212 : 1'b1;
													assign node212 = (inp[3]) ? 1'b0 : 1'b1;
												assign node215 = (inp[7]) ? 1'b0 : node216;
													assign node216 = (inp[5]) ? 1'b0 : 1'b1;
											assign node220 = (inp[3]) ? 1'b0 : node221;
												assign node221 = (inp[7]) ? 1'b0 : node222;
													assign node222 = (inp[5]) ? 1'b0 : 1'b1;
					assign node227 = (inp[14]) ? node377 : node228;
						assign node228 = (inp[13]) ? node282 : node229;
							assign node229 = (inp[4]) ? node243 : node230;
								assign node230 = (inp[5]) ? node232 : 1'b1;
									assign node232 = (inp[8]) ? node234 : 1'b1;
										assign node234 = (inp[10]) ? node236 : 1'b1;
											assign node236 = (inp[7]) ? node238 : 1'b1;
												assign node238 = (inp[2]) ? node240 : 1'b1;
													assign node240 = (inp[9]) ? 1'b0 : 1'b0;
								assign node243 = (inp[8]) ? node257 : node244;
									assign node244 = (inp[9]) ? node246 : 1'b1;
										assign node246 = (inp[7]) ? node248 : 1'b1;
											assign node248 = (inp[10]) ? node250 : 1'b1;
												assign node250 = (inp[3]) ? node254 : node251;
													assign node251 = (inp[2]) ? 1'b1 : 1'b1;
													assign node254 = (inp[2]) ? 1'b0 : 1'b0;
									assign node257 = (inp[3]) ? node267 : node258;
										assign node258 = (inp[5]) ? node260 : 1'b1;
											assign node260 = (inp[9]) ? node262 : 1'b1;
												assign node262 = (inp[10]) ? node264 : 1'b1;
													assign node264 = (inp[7]) ? 1'b0 : 1'b1;
										assign node267 = (inp[7]) ? node275 : node268;
											assign node268 = (inp[2]) ? node270 : 1'b1;
												assign node270 = (inp[11]) ? node272 : 1'b1;
													assign node272 = (inp[10]) ? 1'b0 : 1'b1;
											assign node275 = (inp[11]) ? 1'b0 : node276;
												assign node276 = (inp[5]) ? node278 : 1'b1;
													assign node278 = (inp[10]) ? 1'b0 : 1'b1;
							assign node282 = (inp[2]) ? node320 : node283;
								assign node283 = (inp[9]) ? node293 : node284;
									assign node284 = (inp[4]) ? node286 : 1'b1;
										assign node286 = (inp[3]) ? node288 : 1'b1;
											assign node288 = (inp[10]) ? node290 : 1'b1;
												assign node290 = (inp[8]) ? 1'b0 : 1'b1;
									assign node293 = (inp[8]) ? node303 : node294;
										assign node294 = (inp[4]) ? node296 : 1'b1;
											assign node296 = (inp[7]) ? node298 : 1'b1;
												assign node298 = (inp[10]) ? node300 : 1'b1;
													assign node300 = (inp[5]) ? 1'b0 : 1'b1;
										assign node303 = (inp[11]) ? node309 : node304;
											assign node304 = (inp[5]) ? node306 : 1'b1;
												assign node306 = (inp[4]) ? 1'b0 : 1'b1;
											assign node309 = (inp[4]) ? node315 : node310;
												assign node310 = (inp[3]) ? node312 : 1'b1;
													assign node312 = (inp[7]) ? 1'b0 : 1'b0;
												assign node315 = (inp[10]) ? 1'b0 : node316;
													assign node316 = (inp[3]) ? 1'b0 : 1'b0;
								assign node320 = (inp[11]) ? node348 : node321;
									assign node321 = (inp[3]) ? node331 : node322;
										assign node322 = (inp[10]) ? node324 : 1'b1;
											assign node324 = (inp[8]) ? node326 : 1'b1;
												assign node326 = (inp[9]) ? node328 : 1'b1;
													assign node328 = (inp[7]) ? 1'b0 : 1'b1;
										assign node331 = (inp[4]) ? node339 : node332;
											assign node332 = (inp[9]) ? node334 : 1'b1;
												assign node334 = (inp[10]) ? node336 : 1'b1;
													assign node336 = (inp[7]) ? 1'b0 : 1'b1;
											assign node339 = (inp[8]) ? node343 : node340;
												assign node340 = (inp[9]) ? 1'b0 : 1'b1;
												assign node343 = (inp[10]) ? 1'b0 : node344;
													assign node344 = (inp[7]) ? 1'b0 : 1'b1;
									assign node348 = (inp[7]) ? node364 : node349;
										assign node349 = (inp[4]) ? node357 : node350;
											assign node350 = (inp[8]) ? node352 : 1'b1;
												assign node352 = (inp[10]) ? node354 : 1'b1;
													assign node354 = (inp[5]) ? 1'b0 : 1'b1;
											assign node357 = (inp[10]) ? 1'b0 : node358;
												assign node358 = (inp[9]) ? node360 : 1'b1;
													assign node360 = (inp[5]) ? 1'b0 : 1'b1;
										assign node364 = (inp[8]) ? 1'b0 : node365;
											assign node365 = (inp[9]) ? node371 : node366;
												assign node366 = (inp[10]) ? node368 : 1'b1;
													assign node368 = (inp[5]) ? 1'b0 : 1'b1;
												assign node371 = (inp[5]) ? 1'b0 : node372;
													assign node372 = (inp[4]) ? 1'b0 : 1'b1;
						assign node377 = (inp[7]) ? node479 : node378;
							assign node378 = (inp[9]) ? node414 : node379;
								assign node379 = (inp[10]) ? node389 : node380;
									assign node380 = (inp[5]) ? node382 : 1'b1;
										assign node382 = (inp[8]) ? node384 : 1'b1;
											assign node384 = (inp[2]) ? node386 : 1'b1;
												assign node386 = (inp[4]) ? 1'b0 : 1'b1;
									assign node389 = (inp[13]) ? node399 : node390;
										assign node390 = (inp[4]) ? node392 : 1'b1;
											assign node392 = (inp[8]) ? node394 : 1'b1;
												assign node394 = (inp[3]) ? node396 : 1'b1;
													assign node396 = (inp[11]) ? 1'b0 : 1'b1;
										assign node399 = (inp[8]) ? node407 : node400;
											assign node400 = (inp[4]) ? node402 : 1'b1;
												assign node402 = (inp[5]) ? node404 : 1'b1;
													assign node404 = (inp[3]) ? 1'b0 : 1'b1;
											assign node407 = (inp[2]) ? 1'b0 : node408;
												assign node408 = (inp[4]) ? 1'b0 : node409;
													assign node409 = (inp[11]) ? 1'b0 : 1'b1;
								assign node414 = (inp[2]) ? node440 : node415;
									assign node415 = (inp[8]) ? node425 : node416;
										assign node416 = (inp[5]) ? node418 : 1'b1;
											assign node418 = (inp[10]) ? node420 : 1'b1;
												assign node420 = (inp[13]) ? node422 : 1'b1;
													assign node422 = (inp[3]) ? 1'b0 : 1'b1;
										assign node425 = (inp[13]) ? node433 : node426;
											assign node426 = (inp[4]) ? node428 : 1'b1;
												assign node428 = (inp[3]) ? node430 : 1'b1;
													assign node430 = (inp[5]) ? 1'b0 : 1'b1;
											assign node433 = (inp[11]) ? 1'b0 : node434;
												assign node434 = (inp[10]) ? node436 : 1'b1;
													assign node436 = (inp[3]) ? 1'b0 : 1'b1;
									assign node440 = (inp[5]) ? node460 : node441;
										assign node441 = (inp[13]) ? node449 : node442;
											assign node442 = (inp[4]) ? node444 : 1'b1;
												assign node444 = (inp[8]) ? node446 : 1'b1;
													assign node446 = (inp[11]) ? 1'b0 : 1'b1;
											assign node449 = (inp[11]) ? node455 : node450;
												assign node450 = (inp[4]) ? node452 : 1'b1;
													assign node452 = (inp[10]) ? 1'b0 : 1'b1;
												assign node455 = (inp[8]) ? 1'b0 : node456;
													assign node456 = (inp[10]) ? 1'b0 : 1'b1;
										assign node460 = (inp[3]) ? node472 : node461;
											assign node461 = (inp[10]) ? node467 : node462;
												assign node462 = (inp[4]) ? node464 : 1'b1;
													assign node464 = (inp[13]) ? 1'b0 : 1'b1;
												assign node467 = (inp[4]) ? 1'b0 : node468;
													assign node468 = (inp[8]) ? 1'b0 : 1'b1;
											assign node472 = (inp[10]) ? 1'b0 : node473;
												assign node473 = (inp[11]) ? 1'b0 : node474;
													assign node474 = (inp[4]) ? 1'b0 : 1'b1;
							assign node479 = (inp[11]) ? node547 : node480;
								assign node480 = (inp[8]) ? node508 : node481;
									assign node481 = (inp[4]) ? node491 : node482;
										assign node482 = (inp[2]) ? node484 : 1'b1;
											assign node484 = (inp[3]) ? node486 : 1'b1;
												assign node486 = (inp[10]) ? node488 : 1'b1;
													assign node488 = (inp[9]) ? 1'b0 : 1'b1;
										assign node491 = (inp[5]) ? node501 : node492;
											assign node492 = (inp[9]) ? node494 : 1'b1;
												assign node494 = (inp[10]) ? node498 : node495;
													assign node495 = (inp[2]) ? 1'b1 : 1'b1;
													assign node498 = (inp[3]) ? 1'b0 : 1'b1;
											assign node501 = (inp[2]) ? 1'b0 : node502;
												assign node502 = (inp[3]) ? node504 : 1'b1;
													assign node504 = (inp[10]) ? 1'b0 : 1'b1;
									assign node508 = (inp[3]) ? node528 : node509;
										assign node509 = (inp[13]) ? node517 : node510;
											assign node510 = (inp[5]) ? node512 : 1'b1;
												assign node512 = (inp[2]) ? node514 : 1'b1;
													assign node514 = (inp[10]) ? 1'b0 : 1'b1;
											assign node517 = (inp[9]) ? node523 : node518;
												assign node518 = (inp[10]) ? node520 : 1'b1;
													assign node520 = (inp[4]) ? 1'b0 : 1'b1;
												assign node523 = (inp[5]) ? 1'b0 : node524;
													assign node524 = (inp[10]) ? 1'b0 : 1'b1;
										assign node528 = (inp[2]) ? node540 : node529;
											assign node529 = (inp[10]) ? node535 : node530;
												assign node530 = (inp[5]) ? node532 : 1'b1;
													assign node532 = (inp[13]) ? 1'b0 : 1'b1;
												assign node535 = (inp[4]) ? 1'b0 : node536;
													assign node536 = (inp[5]) ? 1'b0 : 1'b1;
											assign node540 = (inp[5]) ? 1'b0 : node541;
												assign node541 = (inp[4]) ? 1'b0 : node542;
													assign node542 = (inp[9]) ? 1'b0 : 1'b1;
								assign node547 = (inp[10]) ? node581 : node548;
									assign node548 = (inp[4]) ? node568 : node549;
										assign node549 = (inp[2]) ? node557 : node550;
											assign node550 = (inp[5]) ? node552 : 1'b1;
												assign node552 = (inp[3]) ? node554 : 1'b1;
													assign node554 = (inp[8]) ? 1'b0 : 1'b1;
											assign node557 = (inp[8]) ? node563 : node558;
												assign node558 = (inp[5]) ? node560 : 1'b1;
													assign node560 = (inp[13]) ? 1'b0 : 1'b1;
												assign node563 = (inp[9]) ? 1'b0 : node564;
													assign node564 = (inp[13]) ? 1'b0 : 1'b1;
										assign node568 = (inp[8]) ? 1'b0 : node569;
											assign node569 = (inp[3]) ? node575 : node570;
												assign node570 = (inp[9]) ? node572 : 1'b1;
													assign node572 = (inp[13]) ? 1'b0 : 1'b0;
												assign node575 = (inp[5]) ? 1'b0 : node576;
													assign node576 = (inp[9]) ? 1'b0 : 1'b0;
									assign node581 = (inp[9]) ? 1'b0 : node582;
										assign node582 = (inp[3]) ? node594 : node583;
											assign node583 = (inp[8]) ? node589 : node584;
												assign node584 = (inp[4]) ? node586 : 1'b1;
													assign node586 = (inp[13]) ? 1'b0 : 1'b1;
												assign node589 = (inp[2]) ? 1'b0 : node590;
													assign node590 = (inp[5]) ? 1'b0 : 1'b1;
											assign node594 = (inp[4]) ? 1'b0 : node595;
												assign node595 = (inp[5]) ? 1'b0 : node596;
													assign node596 = (inp[2]) ? 1'b0 : 1'b1;
				assign node602 = (inp[8]) ? node988 : node603;
					assign node603 = (inp[7]) ? node739 : node604;
						assign node604 = (inp[11]) ? node650 : node605;
							assign node605 = (inp[3]) ? node607 : 1'b1;
								assign node607 = (inp[10]) ? node619 : node608;
									assign node608 = (inp[2]) ? node610 : 1'b1;
										assign node610 = (inp[13]) ? node612 : 1'b1;
											assign node612 = (inp[12]) ? node614 : 1'b1;
												assign node614 = (inp[9]) ? node616 : 1'b1;
													assign node616 = (inp[14]) ? 1'b0 : 1'b1;
									assign node619 = (inp[12]) ? node629 : node620;
										assign node620 = (inp[5]) ? node622 : 1'b1;
											assign node622 = (inp[9]) ? node624 : 1'b1;
												assign node624 = (inp[13]) ? node626 : 1'b1;
													assign node626 = (inp[4]) ? 1'b0 : 1'b1;
										assign node629 = (inp[14]) ? node637 : node630;
											assign node630 = (inp[5]) ? node632 : 1'b1;
												assign node632 = (inp[4]) ? node634 : 1'b1;
													assign node634 = (inp[13]) ? 1'b0 : 1'b1;
											assign node637 = (inp[9]) ? node645 : node638;
												assign node638 = (inp[5]) ? node642 : node639;
													assign node639 = (inp[13]) ? 1'b1 : 1'b1;
													assign node642 = (inp[13]) ? 1'b0 : 1'b0;
												assign node645 = (inp[5]) ? 1'b0 : node646;
													assign node646 = (inp[2]) ? 1'b0 : 1'b1;
							assign node650 = (inp[4]) ? node686 : node651;
								assign node651 = (inp[2]) ? node661 : node652;
									assign node652 = (inp[14]) ? node654 : 1'b1;
										assign node654 = (inp[3]) ? node656 : 1'b1;
											assign node656 = (inp[13]) ? node658 : 1'b1;
												assign node658 = (inp[9]) ? 1'b0 : 1'b1;
									assign node661 = (inp[13]) ? node671 : node662;
										assign node662 = (inp[12]) ? node664 : 1'b1;
											assign node664 = (inp[10]) ? node666 : 1'b1;
												assign node666 = (inp[14]) ? node668 : 1'b1;
													assign node668 = (inp[9]) ? 1'b0 : 1'b1;
										assign node671 = (inp[3]) ? node679 : node672;
											assign node672 = (inp[10]) ? node674 : 1'b1;
												assign node674 = (inp[9]) ? node676 : 1'b1;
													assign node676 = (inp[5]) ? 1'b0 : 1'b1;
											assign node679 = (inp[14]) ? 1'b0 : node680;
												assign node680 = (inp[5]) ? node682 : 1'b1;
													assign node682 = (inp[10]) ? 1'b0 : 1'b1;
								assign node686 = (inp[13]) ? node710 : node687;
									assign node687 = (inp[12]) ? node689 : 1'b1;
										assign node689 = (inp[9]) ? node699 : node690;
											assign node690 = (inp[3]) ? node692 : 1'b1;
												assign node692 = (inp[5]) ? node696 : node693;
													assign node693 = (inp[10]) ? 1'b1 : 1'b1;
													assign node696 = (inp[10]) ? 1'b0 : 1'b0;
											assign node699 = (inp[14]) ? node705 : node700;
												assign node700 = (inp[2]) ? node702 : 1'b1;
													assign node702 = (inp[10]) ? 1'b0 : 1'b0;
												assign node705 = (inp[10]) ? 1'b0 : node706;
													assign node706 = (inp[5]) ? 1'b0 : 1'b0;
									assign node710 = (inp[14]) ? node726 : node711;
										assign node711 = (inp[10]) ? node719 : node712;
											assign node712 = (inp[9]) ? node714 : 1'b1;
												assign node714 = (inp[2]) ? node716 : 1'b1;
													assign node716 = (inp[3]) ? 1'b0 : 1'b1;
											assign node719 = (inp[5]) ? 1'b0 : node720;
												assign node720 = (inp[2]) ? node722 : 1'b1;
													assign node722 = (inp[3]) ? 1'b0 : 1'b1;
										assign node726 = (inp[2]) ? 1'b0 : node727;
											assign node727 = (inp[9]) ? node733 : node728;
												assign node728 = (inp[12]) ? node730 : 1'b1;
													assign node730 = (inp[3]) ? 1'b0 : 1'b1;
												assign node733 = (inp[10]) ? 1'b0 : node734;
													assign node734 = (inp[5]) ? 1'b1 : 1'b0;
						assign node739 = (inp[4]) ? node847 : node740;
							assign node740 = (inp[10]) ? node782 : node741;
								assign node741 = (inp[13]) ? node753 : node742;
									assign node742 = (inp[3]) ? node744 : 1'b1;
										assign node744 = (inp[2]) ? node746 : 1'b1;
											assign node746 = (inp[14]) ? node748 : 1'b1;
												assign node748 = (inp[5]) ? node750 : 1'b1;
													assign node750 = (inp[9]) ? 1'b0 : 1'b1;
									assign node753 = (inp[5]) ? node763 : node754;
										assign node754 = (inp[11]) ? node756 : 1'b1;
											assign node756 = (inp[2]) ? node758 : 1'b1;
												assign node758 = (inp[14]) ? node760 : 1'b1;
													assign node760 = (inp[9]) ? 1'b0 : 1'b1;
										assign node763 = (inp[11]) ? node771 : node764;
											assign node764 = (inp[3]) ? node766 : 1'b1;
												assign node766 = (inp[12]) ? node768 : 1'b1;
													assign node768 = (inp[9]) ? 1'b0 : 1'b1;
											assign node771 = (inp[14]) ? node777 : node772;
												assign node772 = (inp[3]) ? node774 : 1'b1;
													assign node774 = (inp[12]) ? 1'b0 : 1'b1;
												assign node777 = (inp[2]) ? 1'b0 : node778;
													assign node778 = (inp[9]) ? 1'b0 : 1'b1;
								assign node782 = (inp[11]) ? node808 : node783;
									assign node783 = (inp[9]) ? node793 : node784;
										assign node784 = (inp[3]) ? node786 : 1'b1;
											assign node786 = (inp[12]) ? node788 : 1'b1;
												assign node788 = (inp[13]) ? node790 : 1'b1;
													assign node790 = (inp[14]) ? 1'b0 : 1'b1;
										assign node793 = (inp[13]) ? node801 : node794;
											assign node794 = (inp[2]) ? node796 : 1'b1;
												assign node796 = (inp[3]) ? 1'b0 : node797;
													assign node797 = (inp[5]) ? 1'b1 : 1'b1;
											assign node801 = (inp[5]) ? 1'b0 : node802;
												assign node802 = (inp[3]) ? node804 : 1'b1;
													assign node804 = (inp[14]) ? 1'b0 : 1'b1;
									assign node808 = (inp[2]) ? node828 : node809;
										assign node809 = (inp[13]) ? node817 : node810;
											assign node810 = (inp[12]) ? node812 : 1'b1;
												assign node812 = (inp[5]) ? node814 : 1'b1;
													assign node814 = (inp[3]) ? 1'b0 : 1'b1;
											assign node817 = (inp[5]) ? node823 : node818;
												assign node818 = (inp[9]) ? node820 : 1'b1;
													assign node820 = (inp[3]) ? 1'b0 : 1'b1;
												assign node823 = (inp[9]) ? 1'b0 : node824;
													assign node824 = (inp[14]) ? 1'b0 : 1'b0;
										assign node828 = (inp[14]) ? node840 : node829;
											assign node829 = (inp[12]) ? node835 : node830;
												assign node830 = (inp[13]) ? node832 : 1'b1;
													assign node832 = (inp[5]) ? 1'b0 : 1'b1;
												assign node835 = (inp[5]) ? 1'b0 : node836;
													assign node836 = (inp[9]) ? 1'b0 : 1'b1;
											assign node840 = (inp[9]) ? 1'b0 : node841;
												assign node841 = (inp[3]) ? 1'b0 : node842;
													assign node842 = (inp[5]) ? 1'b0 : 1'b1;
							assign node847 = (inp[11]) ? node917 : node848;
								assign node848 = (inp[2]) ? node880 : node849;
									assign node849 = (inp[9]) ? node859 : node850;
										assign node850 = (inp[13]) ? node852 : 1'b1;
											assign node852 = (inp[12]) ? node854 : 1'b1;
												assign node854 = (inp[14]) ? node856 : 1'b1;
													assign node856 = (inp[10]) ? 1'b0 : 1'b1;
										assign node859 = (inp[14]) ? node867 : node860;
											assign node860 = (inp[10]) ? node862 : 1'b1;
												assign node862 = (inp[13]) ? node864 : 1'b1;
													assign node864 = (inp[3]) ? 1'b0 : 1'b1;
											assign node867 = (inp[13]) ? node873 : node868;
												assign node868 = (inp[3]) ? node870 : 1'b1;
													assign node870 = (inp[12]) ? 1'b0 : 1'b1;
												assign node873 = (inp[10]) ? node877 : node874;
													assign node874 = (inp[12]) ? 1'b0 : 1'b1;
													assign node877 = (inp[5]) ? 1'b0 : 1'b0;
									assign node880 = (inp[5]) ? node900 : node881;
										assign node881 = (inp[13]) ? node889 : node882;
											assign node882 = (inp[10]) ? node884 : 1'b1;
												assign node884 = (inp[9]) ? node886 : 1'b1;
													assign node886 = (inp[12]) ? 1'b0 : 1'b1;
											assign node889 = (inp[12]) ? node895 : node890;
												assign node890 = (inp[9]) ? node892 : 1'b1;
													assign node892 = (inp[10]) ? 1'b0 : 1'b1;
												assign node895 = (inp[3]) ? 1'b0 : node896;
													assign node896 = (inp[10]) ? 1'b0 : 1'b1;
										assign node900 = (inp[12]) ? node910 : node901;
											assign node901 = (inp[9]) ? node905 : node902;
												assign node902 = (inp[3]) ? 1'b0 : 1'b1;
												assign node905 = (inp[13]) ? 1'b0 : node906;
													assign node906 = (inp[10]) ? 1'b0 : 1'b1;
											assign node910 = (inp[14]) ? 1'b0 : node911;
												assign node911 = (inp[13]) ? 1'b0 : node912;
													assign node912 = (inp[10]) ? 1'b0 : 1'b1;
								assign node917 = (inp[10]) ? node959 : node918;
									assign node918 = (inp[12]) ? node940 : node919;
										assign node919 = (inp[13]) ? node927 : node920;
											assign node920 = (inp[3]) ? node922 : 1'b1;
												assign node922 = (inp[2]) ? node924 : 1'b1;
													assign node924 = (inp[14]) ? 1'b0 : 1'b1;
											assign node927 = (inp[14]) ? node935 : node928;
												assign node928 = (inp[9]) ? node932 : node929;
													assign node929 = (inp[3]) ? 1'b1 : 1'b1;
													assign node932 = (inp[2]) ? 1'b0 : 1'b0;
												assign node935 = (inp[3]) ? 1'b0 : node936;
													assign node936 = (inp[5]) ? 1'b0 : 1'b1;
										assign node940 = (inp[9]) ? node952 : node941;
											assign node941 = (inp[3]) ? node947 : node942;
												assign node942 = (inp[5]) ? node944 : 1'b1;
													assign node944 = (inp[13]) ? 1'b0 : 1'b1;
												assign node947 = (inp[2]) ? 1'b0 : node948;
													assign node948 = (inp[14]) ? 1'b0 : 1'b1;
											assign node952 = (inp[2]) ? 1'b0 : node953;
												assign node953 = (inp[14]) ? 1'b0 : node954;
													assign node954 = (inp[3]) ? 1'b0 : 1'b1;
									assign node959 = (inp[14]) ? node979 : node960;
										assign node960 = (inp[12]) ? node972 : node961;
											assign node961 = (inp[3]) ? node967 : node962;
												assign node962 = (inp[9]) ? node964 : 1'b1;
													assign node964 = (inp[13]) ? 1'b0 : 1'b1;
												assign node967 = (inp[13]) ? 1'b0 : node968;
													assign node968 = (inp[2]) ? 1'b0 : 1'b1;
											assign node972 = (inp[2]) ? 1'b0 : node973;
												assign node973 = (inp[3]) ? 1'b0 : node974;
													assign node974 = (inp[5]) ? 1'b0 : 1'b1;
										assign node979 = (inp[3]) ? 1'b0 : node980;
											assign node980 = (inp[9]) ? 1'b0 : node981;
												assign node981 = (inp[5]) ? 1'b0 : node982;
													assign node982 = (inp[2]) ? 1'b0 : 1'b1;
					assign node988 = (inp[5]) ? node1224 : node989;
						assign node989 = (inp[11]) ? node1097 : node990;
							assign node990 = (inp[10]) ? node1032 : node991;
								assign node991 = (inp[13]) ? node1003 : node992;
									assign node992 = (inp[4]) ? node994 : 1'b1;
										assign node994 = (inp[2]) ? node996 : 1'b1;
											assign node996 = (inp[7]) ? node998 : 1'b1;
												assign node998 = (inp[9]) ? node1000 : 1'b1;
													assign node1000 = (inp[12]) ? 1'b0 : 1'b1;
									assign node1003 = (inp[2]) ? node1013 : node1004;
										assign node1004 = (inp[9]) ? node1006 : 1'b1;
											assign node1006 = (inp[3]) ? node1008 : 1'b1;
												assign node1008 = (inp[7]) ? node1010 : 1'b1;
													assign node1010 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1013 = (inp[3]) ? node1021 : node1014;
											assign node1014 = (inp[7]) ? node1016 : 1'b1;
												assign node1016 = (inp[12]) ? node1018 : 1'b1;
													assign node1018 = (inp[9]) ? 1'b0 : 1'b1;
											assign node1021 = (inp[14]) ? node1027 : node1022;
												assign node1022 = (inp[7]) ? node1024 : 1'b1;
													assign node1024 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1027 = (inp[7]) ? 1'b0 : node1028;
													assign node1028 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1032 = (inp[9]) ? node1064 : node1033;
									assign node1033 = (inp[3]) ? node1043 : node1034;
										assign node1034 = (inp[13]) ? node1036 : 1'b1;
											assign node1036 = (inp[7]) ? node1038 : 1'b1;
												assign node1038 = (inp[14]) ? node1040 : 1'b1;
													assign node1040 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1043 = (inp[4]) ? node1051 : node1044;
											assign node1044 = (inp[2]) ? node1046 : 1'b1;
												assign node1046 = (inp[14]) ? node1048 : 1'b1;
													assign node1048 = (inp[13]) ? 1'b0 : 1'b0;
											assign node1051 = (inp[2]) ? node1059 : node1052;
												assign node1052 = (inp[13]) ? node1056 : node1053;
													assign node1053 = (inp[14]) ? 1'b1 : 1'b1;
													assign node1056 = (inp[7]) ? 1'b0 : 1'b0;
												assign node1059 = (inp[7]) ? 1'b0 : node1060;
													assign node1060 = (inp[14]) ? 1'b0 : 1'b0;
									assign node1064 = (inp[12]) ? node1078 : node1065;
										assign node1065 = (inp[7]) ? node1067 : 1'b1;
											assign node1067 = (inp[2]) ? node1073 : node1068;
												assign node1068 = (inp[13]) ? node1070 : 1'b1;
													assign node1070 = (inp[4]) ? 1'b0 : 1'b1;
												assign node1073 = (inp[13]) ? 1'b0 : node1074;
													assign node1074 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1078 = (inp[13]) ? node1090 : node1079;
											assign node1079 = (inp[4]) ? node1085 : node1080;
												assign node1080 = (inp[3]) ? node1082 : 1'b1;
													assign node1082 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1085 = (inp[3]) ? 1'b0 : node1086;
													assign node1086 = (inp[2]) ? 1'b0 : 1'b1;
											assign node1090 = (inp[2]) ? 1'b0 : node1091;
												assign node1091 = (inp[3]) ? 1'b0 : node1092;
													assign node1092 = (inp[7]) ? 1'b0 : 1'b1;
							assign node1097 = (inp[14]) ? node1161 : node1098;
								assign node1098 = (inp[9]) ? node1122 : node1099;
									assign node1099 = (inp[7]) ? node1109 : node1100;
										assign node1100 = (inp[3]) ? node1102 : 1'b1;
											assign node1102 = (inp[12]) ? node1104 : 1'b1;
												assign node1104 = (inp[4]) ? node1106 : 1'b1;
													assign node1106 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1109 = (inp[10]) ? node1115 : node1110;
											assign node1110 = (inp[3]) ? node1112 : 1'b1;
												assign node1112 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1115 = (inp[13]) ? 1'b0 : node1116;
												assign node1116 = (inp[2]) ? node1118 : 1'b1;
													assign node1118 = (inp[4]) ? 1'b0 : 1'b1;
									assign node1122 = (inp[4]) ? node1142 : node1123;
										assign node1123 = (inp[10]) ? node1131 : node1124;
											assign node1124 = (inp[13]) ? node1126 : 1'b1;
												assign node1126 = (inp[7]) ? node1128 : 1'b1;
													assign node1128 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1131 = (inp[2]) ? node1137 : node1132;
												assign node1132 = (inp[3]) ? node1134 : 1'b1;
													assign node1134 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1137 = (inp[12]) ? 1'b0 : node1138;
													assign node1138 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1142 = (inp[2]) ? node1154 : node1143;
											assign node1143 = (inp[7]) ? node1149 : node1144;
												assign node1144 = (inp[13]) ? node1146 : 1'b1;
													assign node1146 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1149 = (inp[3]) ? 1'b0 : node1150;
													assign node1150 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1154 = (inp[12]) ? 1'b0 : node1155;
												assign node1155 = (inp[7]) ? 1'b0 : node1156;
													assign node1156 = (inp[3]) ? 1'b0 : 1'b0;
								assign node1161 = (inp[3]) ? node1195 : node1162;
									assign node1162 = (inp[10]) ? node1176 : node1163;
										assign node1163 = (inp[13]) ? node1165 : 1'b1;
											assign node1165 = (inp[2]) ? node1171 : node1166;
												assign node1166 = (inp[4]) ? node1168 : 1'b1;
													assign node1168 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1171 = (inp[9]) ? 1'b0 : node1172;
													assign node1172 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1176 = (inp[12]) ? node1188 : node1177;
											assign node1177 = (inp[4]) ? node1183 : node1178;
												assign node1178 = (inp[2]) ? node1180 : 1'b1;
													assign node1180 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1183 = (inp[9]) ? 1'b0 : node1184;
													assign node1184 = (inp[13]) ? 1'b0 : 1'b0;
											assign node1188 = (inp[7]) ? 1'b0 : node1189;
												assign node1189 = (inp[9]) ? 1'b0 : node1190;
													assign node1190 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1195 = (inp[9]) ? node1215 : node1196;
										assign node1196 = (inp[2]) ? node1208 : node1197;
											assign node1197 = (inp[4]) ? node1203 : node1198;
												assign node1198 = (inp[13]) ? node1200 : 1'b1;
													assign node1200 = (inp[12]) ? 1'b0 : 1'b1;
												assign node1203 = (inp[7]) ? 1'b0 : node1204;
													assign node1204 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1208 = (inp[7]) ? 1'b0 : node1209;
												assign node1209 = (inp[12]) ? 1'b0 : node1210;
													assign node1210 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1215 = (inp[12]) ? 1'b0 : node1216;
											assign node1216 = (inp[10]) ? 1'b0 : node1217;
												assign node1217 = (inp[2]) ? 1'b0 : node1218;
													assign node1218 = (inp[4]) ? 1'b0 : 1'b1;
						assign node1224 = (inp[12]) ? node1364 : node1225;
							assign node1225 = (inp[10]) ? node1295 : node1226;
								assign node1226 = (inp[14]) ? node1256 : node1227;
									assign node1227 = (inp[3]) ? node1237 : node1228;
										assign node1228 = (inp[7]) ? node1230 : 1'b1;
											assign node1230 = (inp[13]) ? node1232 : 1'b1;
												assign node1232 = (inp[2]) ? node1234 : 1'b1;
													assign node1234 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1237 = (inp[11]) ? node1245 : node1238;
											assign node1238 = (inp[13]) ? node1240 : 1'b1;
												assign node1240 = (inp[2]) ? node1242 : 1'b1;
													assign node1242 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1245 = (inp[9]) ? node1251 : node1246;
												assign node1246 = (inp[7]) ? node1248 : 1'b1;
													assign node1248 = (inp[4]) ? 1'b0 : 1'b1;
												assign node1251 = (inp[2]) ? 1'b0 : node1252;
													assign node1252 = (inp[7]) ? 1'b0 : 1'b0;
									assign node1256 = (inp[3]) ? node1276 : node1257;
										assign node1257 = (inp[7]) ? node1265 : node1258;
											assign node1258 = (inp[2]) ? node1260 : 1'b1;
												assign node1260 = (inp[9]) ? node1262 : 1'b1;
													assign node1262 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1265 = (inp[9]) ? node1271 : node1266;
												assign node1266 = (inp[4]) ? node1268 : 1'b1;
													assign node1268 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1271 = (inp[11]) ? 1'b0 : node1272;
													assign node1272 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1276 = (inp[13]) ? node1288 : node1277;
											assign node1277 = (inp[11]) ? node1283 : node1278;
												assign node1278 = (inp[4]) ? node1280 : 1'b1;
													assign node1280 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1283 = (inp[4]) ? 1'b0 : node1284;
													assign node1284 = (inp[9]) ? 1'b0 : 1'b1;
											assign node1288 = (inp[9]) ? 1'b0 : node1289;
												assign node1289 = (inp[7]) ? 1'b0 : node1290;
													assign node1290 = (inp[2]) ? 1'b0 : 1'b1;
								assign node1295 = (inp[2]) ? node1335 : node1296;
									assign node1296 = (inp[14]) ? node1316 : node1297;
										assign node1297 = (inp[9]) ? node1305 : node1298;
											assign node1298 = (inp[13]) ? node1300 : 1'b1;
												assign node1300 = (inp[11]) ? node1302 : 1'b1;
													assign node1302 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1305 = (inp[3]) ? node1311 : node1306;
												assign node1306 = (inp[13]) ? node1308 : 1'b1;
													assign node1308 = (inp[4]) ? 1'b0 : 1'b1;
												assign node1311 = (inp[11]) ? 1'b0 : node1312;
													assign node1312 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1316 = (inp[4]) ? node1328 : node1317;
											assign node1317 = (inp[3]) ? node1323 : node1318;
												assign node1318 = (inp[9]) ? node1320 : 1'b1;
													assign node1320 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1323 = (inp[11]) ? 1'b0 : node1324;
													assign node1324 = (inp[13]) ? 1'b1 : 1'b0;
											assign node1328 = (inp[13]) ? 1'b0 : node1329;
												assign node1329 = (inp[11]) ? 1'b0 : node1330;
													assign node1330 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1335 = (inp[11]) ? node1355 : node1336;
										assign node1336 = (inp[7]) ? node1348 : node1337;
											assign node1337 = (inp[9]) ? node1343 : node1338;
												assign node1338 = (inp[14]) ? node1340 : 1'b1;
													assign node1340 = (inp[4]) ? 1'b0 : 1'b1;
												assign node1343 = (inp[13]) ? 1'b0 : node1344;
													assign node1344 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1348 = (inp[9]) ? 1'b0 : node1349;
												assign node1349 = (inp[14]) ? 1'b0 : node1350;
													assign node1350 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1355 = (inp[3]) ? 1'b0 : node1356;
											assign node1356 = (inp[13]) ? 1'b0 : node1357;
												assign node1357 = (inp[14]) ? 1'b0 : node1358;
													assign node1358 = (inp[4]) ? 1'b0 : 1'b1;
							assign node1364 = (inp[11]) ? node1432 : node1365;
								assign node1365 = (inp[13]) ? node1405 : node1366;
									assign node1366 = (inp[10]) ? node1386 : node1367;
										assign node1367 = (inp[9]) ? node1375 : node1368;
											assign node1368 = (inp[3]) ? node1370 : 1'b1;
												assign node1370 = (inp[7]) ? node1372 : 1'b1;
													assign node1372 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1375 = (inp[2]) ? node1381 : node1376;
												assign node1376 = (inp[7]) ? node1378 : 1'b1;
													assign node1378 = (inp[14]) ? 1'b0 : 1'b1;
												assign node1381 = (inp[4]) ? 1'b0 : node1382;
													assign node1382 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1386 = (inp[14]) ? node1398 : node1387;
											assign node1387 = (inp[3]) ? node1393 : node1388;
												assign node1388 = (inp[9]) ? node1390 : 1'b1;
													assign node1390 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1393 = (inp[2]) ? 1'b0 : node1394;
													assign node1394 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1398 = (inp[7]) ? 1'b0 : node1399;
												assign node1399 = (inp[3]) ? 1'b0 : node1400;
													assign node1400 = (inp[4]) ? 1'b0 : 1'b1;
									assign node1405 = (inp[9]) ? node1423 : node1406;
										assign node1406 = (inp[10]) ? node1418 : node1407;
											assign node1407 = (inp[4]) ? node1413 : node1408;
												assign node1408 = (inp[7]) ? node1410 : 1'b1;
													assign node1410 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1413 = (inp[3]) ? 1'b0 : node1414;
													assign node1414 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1418 = (inp[3]) ? 1'b0 : node1419;
												assign node1419 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1423 = (inp[14]) ? 1'b0 : node1424;
											assign node1424 = (inp[4]) ? 1'b0 : node1425;
												assign node1425 = (inp[2]) ? 1'b0 : node1426;
													assign node1426 = (inp[3]) ? 1'b0 : 1'b1;
								assign node1432 = (inp[3]) ? node1462 : node1433;
									assign node1433 = (inp[14]) ? node1453 : node1434;
										assign node1434 = (inp[2]) ? node1446 : node1435;
											assign node1435 = (inp[13]) ? node1441 : node1436;
												assign node1436 = (inp[9]) ? node1438 : 1'b1;
													assign node1438 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1441 = (inp[10]) ? 1'b0 : node1442;
													assign node1442 = (inp[9]) ? 1'b0 : 1'b1;
											assign node1446 = (inp[9]) ? 1'b0 : node1447;
												assign node1447 = (inp[10]) ? 1'b0 : node1448;
													assign node1448 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1453 = (inp[4]) ? 1'b0 : node1454;
											assign node1454 = (inp[7]) ? 1'b0 : node1455;
												assign node1455 = (inp[2]) ? 1'b0 : node1456;
													assign node1456 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1462 = (inp[7]) ? 1'b0 : node1463;
										assign node1463 = (inp[14]) ? 1'b0 : node1464;
											assign node1464 = (inp[10]) ? 1'b0 : node1465;
												assign node1465 = (inp[13]) ? 1'b0 : node1466;
													assign node1466 = (inp[9]) ? 1'b0 : 1'b1;
			assign node1473 = (inp[13]) ? node2357 : node1474;
				assign node1474 = (inp[9]) ? node1874 : node1475;
					assign node1475 = (inp[4]) ? node1639 : node1476;
						assign node1476 = (inp[0]) ? node1534 : node1477;
							assign node1477 = (inp[8]) ? node1491 : node1478;
								assign node1478 = (inp[3]) ? node1480 : 1'b1;
									assign node1480 = (inp[5]) ? node1482 : 1'b1;
										assign node1482 = (inp[10]) ? node1484 : 1'b1;
											assign node1484 = (inp[7]) ? node1486 : 1'b1;
												assign node1486 = (inp[2]) ? node1488 : 1'b1;
													assign node1488 = (inp[14]) ? 1'b0 : 1'b1;
								assign node1491 = (inp[2]) ? node1503 : node1492;
									assign node1492 = (inp[11]) ? node1494 : 1'b1;
										assign node1494 = (inp[10]) ? node1496 : 1'b1;
											assign node1496 = (inp[12]) ? node1498 : 1'b1;
												assign node1498 = (inp[3]) ? node1500 : 1'b1;
													assign node1500 = (inp[14]) ? 1'b0 : 1'b1;
									assign node1503 = (inp[12]) ? node1513 : node1504;
										assign node1504 = (inp[11]) ? node1506 : 1'b1;
											assign node1506 = (inp[5]) ? node1508 : 1'b1;
												assign node1508 = (inp[10]) ? node1510 : 1'b1;
													assign node1510 = (inp[3]) ? 1'b1 : 1'b0;
										assign node1513 = (inp[11]) ? node1521 : node1514;
											assign node1514 = (inp[10]) ? node1516 : 1'b1;
												assign node1516 = (inp[14]) ? node1518 : 1'b1;
													assign node1518 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1521 = (inp[5]) ? node1529 : node1522;
												assign node1522 = (inp[10]) ? node1526 : node1523;
													assign node1523 = (inp[3]) ? 1'b1 : 1'b1;
													assign node1526 = (inp[14]) ? 1'b0 : 1'b1;
												assign node1529 = (inp[10]) ? 1'b0 : node1530;
													assign node1530 = (inp[3]) ? 1'b0 : 1'b1;
							assign node1534 = (inp[7]) ? node1570 : node1535;
								assign node1535 = (inp[3]) ? node1547 : node1536;
									assign node1536 = (inp[11]) ? node1538 : 1'b1;
										assign node1538 = (inp[14]) ? node1540 : 1'b1;
											assign node1540 = (inp[10]) ? node1542 : 1'b1;
												assign node1542 = (inp[5]) ? node1544 : 1'b1;
													assign node1544 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1547 = (inp[12]) ? node1557 : node1548;
										assign node1548 = (inp[5]) ? node1550 : 1'b1;
											assign node1550 = (inp[14]) ? node1552 : 1'b1;
												assign node1552 = (inp[11]) ? node1554 : 1'b1;
													assign node1554 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1557 = (inp[11]) ? node1565 : node1558;
											assign node1558 = (inp[8]) ? node1560 : 1'b1;
												assign node1560 = (inp[5]) ? node1562 : 1'b1;
													assign node1562 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1565 = (inp[14]) ? 1'b0 : node1566;
												assign node1566 = (inp[5]) ? 1'b0 : 1'b1;
								assign node1570 = (inp[8]) ? node1600 : node1571;
									assign node1571 = (inp[12]) ? node1581 : node1572;
										assign node1572 = (inp[10]) ? node1574 : 1'b1;
											assign node1574 = (inp[11]) ? node1576 : 1'b1;
												assign node1576 = (inp[5]) ? node1578 : 1'b1;
													assign node1578 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1581 = (inp[2]) ? node1589 : node1582;
											assign node1582 = (inp[14]) ? node1584 : 1'b1;
												assign node1584 = (inp[5]) ? node1586 : 1'b1;
													assign node1586 = (inp[3]) ? 1'b0 : 1'b0;
											assign node1589 = (inp[3]) ? node1595 : node1590;
												assign node1590 = (inp[14]) ? node1592 : 1'b1;
													assign node1592 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1595 = (inp[14]) ? 1'b0 : node1596;
													assign node1596 = (inp[10]) ? 1'b0 : 1'b0;
									assign node1600 = (inp[11]) ? node1620 : node1601;
										assign node1601 = (inp[5]) ? node1609 : node1602;
											assign node1602 = (inp[3]) ? node1604 : 1'b1;
												assign node1604 = (inp[10]) ? node1606 : 1'b1;
													assign node1606 = (inp[2]) ? 1'b0 : 1'b1;
											assign node1609 = (inp[10]) ? node1615 : node1610;
												assign node1610 = (inp[2]) ? node1612 : 1'b1;
													assign node1612 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1615 = (inp[2]) ? 1'b0 : node1616;
													assign node1616 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1620 = (inp[5]) ? node1632 : node1621;
											assign node1621 = (inp[10]) ? node1627 : node1622;
												assign node1622 = (inp[12]) ? node1624 : 1'b1;
													assign node1624 = (inp[14]) ? 1'b0 : 1'b1;
												assign node1627 = (inp[3]) ? 1'b0 : node1628;
													assign node1628 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1632 = (inp[2]) ? 1'b0 : node1633;
												assign node1633 = (inp[14]) ? 1'b0 : node1634;
													assign node1634 = (inp[3]) ? 1'b0 : 1'b1;
						assign node1639 = (inp[14]) ? node1747 : node1640;
							assign node1640 = (inp[12]) ? node1678 : node1641;
								assign node1641 = (inp[2]) ? node1653 : node1642;
									assign node1642 = (inp[3]) ? node1644 : 1'b1;
										assign node1644 = (inp[7]) ? node1646 : 1'b1;
											assign node1646 = (inp[5]) ? node1648 : 1'b1;
												assign node1648 = (inp[0]) ? node1650 : 1'b1;
													assign node1650 = (inp[8]) ? 1'b0 : 1'b1;
									assign node1653 = (inp[3]) ? node1663 : node1654;
										assign node1654 = (inp[10]) ? node1656 : 1'b1;
											assign node1656 = (inp[8]) ? node1658 : 1'b1;
												assign node1658 = (inp[0]) ? node1660 : 1'b1;
													assign node1660 = (inp[11]) ? 1'b0 : 1'b0;
										assign node1663 = (inp[0]) ? node1671 : node1664;
											assign node1664 = (inp[5]) ? node1666 : 1'b1;
												assign node1666 = (inp[7]) ? node1668 : 1'b1;
													assign node1668 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1671 = (inp[10]) ? 1'b0 : node1672;
												assign node1672 = (inp[11]) ? node1674 : 1'b1;
													assign node1674 = (inp[5]) ? 1'b0 : 1'b1;
								assign node1678 = (inp[8]) ? node1708 : node1679;
									assign node1679 = (inp[7]) ? node1689 : node1680;
										assign node1680 = (inp[2]) ? node1682 : 1'b1;
											assign node1682 = (inp[5]) ? node1684 : 1'b1;
												assign node1684 = (inp[3]) ? node1686 : 1'b1;
													assign node1686 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1689 = (inp[2]) ? node1697 : node1690;
											assign node1690 = (inp[0]) ? node1692 : 1'b1;
												assign node1692 = (inp[10]) ? node1694 : 1'b1;
													assign node1694 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1697 = (inp[5]) ? node1703 : node1698;
												assign node1698 = (inp[3]) ? node1700 : 1'b1;
													assign node1700 = (inp[0]) ? 1'b0 : 1'b1;
												assign node1703 = (inp[10]) ? 1'b0 : node1704;
													assign node1704 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1708 = (inp[7]) ? node1728 : node1709;
										assign node1709 = (inp[10]) ? node1717 : node1710;
											assign node1710 = (inp[3]) ? node1712 : 1'b1;
												assign node1712 = (inp[0]) ? node1714 : 1'b1;
													assign node1714 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1717 = (inp[11]) ? node1723 : node1718;
												assign node1718 = (inp[0]) ? node1720 : 1'b1;
													assign node1720 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1723 = (inp[2]) ? 1'b0 : node1724;
													assign node1724 = (inp[5]) ? 1'b0 : 1'b1;
										assign node1728 = (inp[2]) ? node1740 : node1729;
											assign node1729 = (inp[5]) ? node1735 : node1730;
												assign node1730 = (inp[3]) ? node1732 : 1'b1;
													assign node1732 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1735 = (inp[3]) ? 1'b0 : node1736;
													assign node1736 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1740 = (inp[0]) ? 1'b0 : node1741;
												assign node1741 = (inp[3]) ? 1'b0 : node1742;
													assign node1742 = (inp[11]) ? 1'b0 : 1'b1;
							assign node1747 = (inp[10]) ? node1807 : node1748;
								assign node1748 = (inp[5]) ? node1770 : node1749;
									assign node1749 = (inp[0]) ? node1751 : 1'b1;
										assign node1751 = (inp[8]) ? node1759 : node1752;
											assign node1752 = (inp[3]) ? node1754 : 1'b1;
												assign node1754 = (inp[7]) ? node1756 : 1'b1;
													assign node1756 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1759 = (inp[12]) ? node1765 : node1760;
												assign node1760 = (inp[2]) ? node1762 : 1'b1;
													assign node1762 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1765 = (inp[3]) ? 1'b0 : node1766;
													assign node1766 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1770 = (inp[8]) ? node1790 : node1771;
										assign node1771 = (inp[12]) ? node1779 : node1772;
											assign node1772 = (inp[11]) ? node1774 : 1'b1;
												assign node1774 = (inp[3]) ? node1776 : 1'b1;
													assign node1776 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1779 = (inp[0]) ? node1785 : node1780;
												assign node1780 = (inp[7]) ? node1782 : 1'b1;
													assign node1782 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1785 = (inp[11]) ? 1'b0 : node1786;
													assign node1786 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1790 = (inp[11]) ? node1802 : node1791;
											assign node1791 = (inp[12]) ? node1797 : node1792;
												assign node1792 = (inp[0]) ? node1794 : 1'b1;
													assign node1794 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1797 = (inp[3]) ? 1'b0 : node1798;
													assign node1798 = (inp[2]) ? 1'b0 : 1'b1;
											assign node1802 = (inp[3]) ? 1'b0 : node1803;
												assign node1803 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1807 = (inp[5]) ? node1847 : node1808;
									assign node1808 = (inp[3]) ? node1828 : node1809;
										assign node1809 = (inp[2]) ? node1817 : node1810;
											assign node1810 = (inp[8]) ? node1812 : 1'b1;
												assign node1812 = (inp[7]) ? node1814 : 1'b1;
													assign node1814 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1817 = (inp[11]) ? node1823 : node1818;
												assign node1818 = (inp[12]) ? node1820 : 1'b1;
													assign node1820 = (inp[0]) ? 1'b0 : 1'b1;
												assign node1823 = (inp[7]) ? 1'b0 : node1824;
													assign node1824 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1828 = (inp[11]) ? node1840 : node1829;
											assign node1829 = (inp[0]) ? node1835 : node1830;
												assign node1830 = (inp[8]) ? node1832 : 1'b1;
													assign node1832 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1835 = (inp[7]) ? 1'b0 : node1836;
													assign node1836 = (inp[2]) ? 1'b0 : 1'b1;
											assign node1840 = (inp[2]) ? 1'b0 : node1841;
												assign node1841 = (inp[0]) ? 1'b0 : node1842;
													assign node1842 = (inp[8]) ? 1'b0 : 1'b1;
									assign node1847 = (inp[2]) ? node1867 : node1848;
										assign node1848 = (inp[8]) ? node1860 : node1849;
											assign node1849 = (inp[7]) ? node1855 : node1850;
												assign node1850 = (inp[3]) ? node1852 : 1'b1;
													assign node1852 = (inp[12]) ? 1'b0 : 1'b1;
												assign node1855 = (inp[3]) ? 1'b0 : node1856;
													assign node1856 = (inp[11]) ? 1'b0 : 1'b0;
											assign node1860 = (inp[11]) ? 1'b0 : node1861;
												assign node1861 = (inp[0]) ? 1'b0 : node1862;
													assign node1862 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1867 = (inp[11]) ? 1'b0 : node1868;
											assign node1868 = (inp[8]) ? 1'b0 : node1869;
												assign node1869 = (inp[12]) ? 1'b0 : 1'b1;
					assign node1874 = (inp[12]) ? node2112 : node1875;
						assign node1875 = (inp[8]) ? node1981 : node1876;
							assign node1876 = (inp[3]) ? node1916 : node1877;
								assign node1877 = (inp[4]) ? node1889 : node1878;
									assign node1878 = (inp[10]) ? node1880 : 1'b1;
										assign node1880 = (inp[11]) ? node1882 : 1'b1;
											assign node1882 = (inp[5]) ? node1884 : 1'b1;
												assign node1884 = (inp[14]) ? node1886 : 1'b1;
													assign node1886 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1889 = (inp[0]) ? node1897 : node1890;
										assign node1890 = (inp[7]) ? node1892 : 1'b1;
											assign node1892 = (inp[2]) ? node1894 : 1'b1;
												assign node1894 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1897 = (inp[11]) ? node1905 : node1898;
											assign node1898 = (inp[2]) ? node1900 : 1'b1;
												assign node1900 = (inp[10]) ? node1902 : 1'b1;
													assign node1902 = (inp[5]) ? 1'b0 : 1'b1;
											assign node1905 = (inp[10]) ? node1911 : node1906;
												assign node1906 = (inp[5]) ? node1908 : 1'b1;
													assign node1908 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1911 = (inp[5]) ? 1'b0 : node1912;
													assign node1912 = (inp[14]) ? 1'b0 : 1'b1;
								assign node1916 = (inp[14]) ? node1948 : node1917;
									assign node1917 = (inp[10]) ? node1927 : node1918;
										assign node1918 = (inp[11]) ? node1920 : 1'b1;
											assign node1920 = (inp[5]) ? node1922 : 1'b1;
												assign node1922 = (inp[0]) ? node1924 : 1'b1;
													assign node1924 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1927 = (inp[7]) ? node1935 : node1928;
											assign node1928 = (inp[2]) ? node1930 : 1'b1;
												assign node1930 = (inp[5]) ? node1932 : 1'b1;
													assign node1932 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1935 = (inp[0]) ? node1943 : node1936;
												assign node1936 = (inp[4]) ? node1940 : node1937;
													assign node1937 = (inp[2]) ? 1'b1 : 1'b1;
													assign node1940 = (inp[5]) ? 1'b0 : 1'b1;
												assign node1943 = (inp[5]) ? 1'b0 : node1944;
													assign node1944 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1948 = (inp[5]) ? node1968 : node1949;
										assign node1949 = (inp[4]) ? node1957 : node1950;
											assign node1950 = (inp[10]) ? node1952 : 1'b1;
												assign node1952 = (inp[11]) ? node1954 : 1'b1;
													assign node1954 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1957 = (inp[0]) ? node1963 : node1958;
												assign node1958 = (inp[7]) ? node1960 : 1'b1;
													assign node1960 = (inp[10]) ? 1'b0 : 1'b1;
												assign node1963 = (inp[11]) ? 1'b0 : node1964;
													assign node1964 = (inp[10]) ? 1'b0 : 1'b0;
										assign node1968 = (inp[2]) ? 1'b0 : node1969;
											assign node1969 = (inp[11]) ? node1975 : node1970;
												assign node1970 = (inp[0]) ? node1972 : 1'b1;
													assign node1972 = (inp[4]) ? 1'b0 : 1'b1;
												assign node1975 = (inp[7]) ? 1'b0 : node1976;
													assign node1976 = (inp[0]) ? 1'b0 : 1'b1;
							assign node1981 = (inp[4]) ? node2043 : node1982;
								assign node1982 = (inp[0]) ? node2010 : node1983;
									assign node1983 = (inp[2]) ? node1993 : node1984;
										assign node1984 = (inp[11]) ? node1986 : 1'b1;
											assign node1986 = (inp[3]) ? node1988 : 1'b1;
												assign node1988 = (inp[5]) ? node1990 : 1'b1;
													assign node1990 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1993 = (inp[14]) ? node1999 : node1994;
											assign node1994 = (inp[11]) ? node1996 : 1'b1;
												assign node1996 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1999 = (inp[3]) ? node2005 : node2000;
												assign node2000 = (inp[10]) ? node2002 : 1'b1;
													assign node2002 = (inp[5]) ? 1'b0 : 1'b1;
												assign node2005 = (inp[11]) ? 1'b0 : node2006;
													assign node2006 = (inp[10]) ? 1'b0 : 1'b1;
									assign node2010 = (inp[3]) ? node2030 : node2011;
										assign node2011 = (inp[10]) ? node2019 : node2012;
											assign node2012 = (inp[14]) ? node2014 : 1'b1;
												assign node2014 = (inp[11]) ? node2016 : 1'b1;
													assign node2016 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2019 = (inp[14]) ? node2025 : node2020;
												assign node2020 = (inp[11]) ? node2022 : 1'b1;
													assign node2022 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2025 = (inp[7]) ? 1'b0 : node2026;
													assign node2026 = (inp[5]) ? 1'b0 : 1'b1;
										assign node2030 = (inp[10]) ? 1'b0 : node2031;
											assign node2031 = (inp[14]) ? node2037 : node2032;
												assign node2032 = (inp[11]) ? node2034 : 1'b1;
													assign node2034 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2037 = (inp[7]) ? 1'b0 : node2038;
													assign node2038 = (inp[5]) ? 1'b0 : 1'b1;
								assign node2043 = (inp[5]) ? node2083 : node2044;
									assign node2044 = (inp[0]) ? node2062 : node2045;
										assign node2045 = (inp[14]) ? node2053 : node2046;
											assign node2046 = (inp[10]) ? node2048 : 1'b1;
												assign node2048 = (inp[2]) ? 1'b1 : node2049;
													assign node2049 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2053 = (inp[3]) ? node2057 : node2054;
												assign node2054 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2057 = (inp[2]) ? 1'b0 : node2058;
													assign node2058 = (inp[7]) ? 1'b0 : 1'b1;
										assign node2062 = (inp[11]) ? node2076 : node2063;
											assign node2063 = (inp[10]) ? node2069 : node2064;
												assign node2064 = (inp[2]) ? node2066 : 1'b1;
													assign node2066 = (inp[3]) ? 1'b0 : 1'b1;
												assign node2069 = (inp[2]) ? node2073 : node2070;
													assign node2070 = (inp[3]) ? 1'b0 : 1'b1;
													assign node2073 = (inp[7]) ? 1'b0 : 1'b0;
											assign node2076 = (inp[10]) ? 1'b0 : node2077;
												assign node2077 = (inp[7]) ? 1'b0 : node2078;
													assign node2078 = (inp[2]) ? 1'b0 : 1'b1;
									assign node2083 = (inp[0]) ? node2103 : node2084;
										assign node2084 = (inp[11]) ? node2096 : node2085;
											assign node2085 = (inp[3]) ? node2091 : node2086;
												assign node2086 = (inp[7]) ? node2088 : 1'b1;
													assign node2088 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2091 = (inp[7]) ? 1'b0 : node2092;
													assign node2092 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2096 = (inp[10]) ? 1'b0 : node2097;
												assign node2097 = (inp[7]) ? 1'b0 : node2098;
													assign node2098 = (inp[2]) ? 1'b0 : 1'b0;
										assign node2103 = (inp[14]) ? 1'b0 : node2104;
											assign node2104 = (inp[11]) ? 1'b0 : node2105;
												assign node2105 = (inp[7]) ? 1'b0 : node2106;
													assign node2106 = (inp[3]) ? 1'b0 : 1'b1;
						assign node2112 = (inp[5]) ? node2248 : node2113;
							assign node2113 = (inp[4]) ? node2183 : node2114;
								assign node2114 = (inp[8]) ? node2144 : node2115;
									assign node2115 = (inp[11]) ? node2125 : node2116;
										assign node2116 = (inp[2]) ? node2118 : 1'b1;
											assign node2118 = (inp[3]) ? node2120 : 1'b1;
												assign node2120 = (inp[14]) ? node2122 : 1'b1;
													assign node2122 = (inp[0]) ? 1'b0 : 1'b1;
										assign node2125 = (inp[3]) ? node2133 : node2126;
											assign node2126 = (inp[7]) ? node2128 : 1'b1;
												assign node2128 = (inp[10]) ? node2130 : 1'b1;
													assign node2130 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2133 = (inp[14]) ? node2139 : node2134;
												assign node2134 = (inp[10]) ? node2136 : 1'b1;
													assign node2136 = (inp[7]) ? 1'b0 : 1'b0;
												assign node2139 = (inp[2]) ? 1'b0 : node2140;
													assign node2140 = (inp[0]) ? 1'b0 : 1'b1;
									assign node2144 = (inp[2]) ? node2164 : node2145;
										assign node2145 = (inp[3]) ? node2153 : node2146;
											assign node2146 = (inp[14]) ? node2148 : 1'b1;
												assign node2148 = (inp[10]) ? node2150 : 1'b1;
													assign node2150 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2153 = (inp[10]) ? node2159 : node2154;
												assign node2154 = (inp[11]) ? node2156 : 1'b1;
													assign node2156 = (inp[14]) ? 1'b0 : 1'b1;
												assign node2159 = (inp[7]) ? 1'b0 : node2160;
													assign node2160 = (inp[0]) ? 1'b0 : 1'b1;
										assign node2164 = (inp[7]) ? node2176 : node2165;
											assign node2165 = (inp[11]) ? node2171 : node2166;
												assign node2166 = (inp[3]) ? node2168 : 1'b1;
													assign node2168 = (inp[14]) ? 1'b0 : 1'b1;
												assign node2171 = (inp[10]) ? 1'b0 : node2172;
													assign node2172 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2176 = (inp[10]) ? 1'b0 : node2177;
												assign node2177 = (inp[0]) ? 1'b0 : node2178;
													assign node2178 = (inp[14]) ? 1'b0 : 1'b1;
								assign node2183 = (inp[2]) ? node2225 : node2184;
									assign node2184 = (inp[11]) ? node2204 : node2185;
										assign node2185 = (inp[3]) ? node2193 : node2186;
											assign node2186 = (inp[7]) ? node2188 : 1'b1;
												assign node2188 = (inp[14]) ? node2190 : 1'b1;
													assign node2190 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2193 = (inp[0]) ? node2199 : node2194;
												assign node2194 = (inp[14]) ? node2196 : 1'b1;
													assign node2196 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2199 = (inp[7]) ? 1'b0 : node2200;
													assign node2200 = (inp[10]) ? 1'b0 : 1'b0;
										assign node2204 = (inp[14]) ? node2218 : node2205;
											assign node2205 = (inp[8]) ? node2213 : node2206;
												assign node2206 = (inp[7]) ? node2210 : node2207;
													assign node2207 = (inp[10]) ? 1'b1 : 1'b1;
													assign node2210 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2213 = (inp[0]) ? 1'b0 : node2214;
													assign node2214 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2218 = (inp[3]) ? 1'b0 : node2219;
												assign node2219 = (inp[8]) ? 1'b0 : node2220;
													assign node2220 = (inp[7]) ? 1'b0 : 1'b1;
									assign node2225 = (inp[0]) ? node2241 : node2226;
										assign node2226 = (inp[11]) ? node2234 : node2227;
											assign node2227 = (inp[14]) ? node2229 : 1'b1;
												assign node2229 = (inp[3]) ? 1'b0 : node2230;
													assign node2230 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2234 = (inp[10]) ? 1'b0 : node2235;
												assign node2235 = (inp[3]) ? 1'b0 : node2236;
													assign node2236 = (inp[8]) ? 1'b0 : 1'b1;
										assign node2241 = (inp[3]) ? 1'b0 : node2242;
											assign node2242 = (inp[14]) ? 1'b0 : node2243;
												assign node2243 = (inp[8]) ? 1'b0 : 1'b1;
							assign node2248 = (inp[7]) ? node2316 : node2249;
								assign node2249 = (inp[2]) ? node2289 : node2250;
									assign node2250 = (inp[10]) ? node2270 : node2251;
										assign node2251 = (inp[14]) ? node2259 : node2252;
											assign node2252 = (inp[0]) ? node2254 : 1'b1;
												assign node2254 = (inp[11]) ? node2256 : 1'b1;
													assign node2256 = (inp[4]) ? 1'b0 : 1'b1;
											assign node2259 = (inp[3]) ? node2265 : node2260;
												assign node2260 = (inp[11]) ? node2262 : 1'b1;
													assign node2262 = (inp[4]) ? 1'b0 : 1'b1;
												assign node2265 = (inp[4]) ? 1'b0 : node2266;
													assign node2266 = (inp[8]) ? 1'b0 : 1'b1;
										assign node2270 = (inp[11]) ? node2282 : node2271;
											assign node2271 = (inp[8]) ? node2277 : node2272;
												assign node2272 = (inp[4]) ? node2274 : 1'b1;
													assign node2274 = (inp[0]) ? 1'b0 : 1'b1;
												assign node2277 = (inp[14]) ? 1'b0 : node2278;
													assign node2278 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2282 = (inp[4]) ? 1'b0 : node2283;
												assign node2283 = (inp[0]) ? 1'b0 : node2284;
													assign node2284 = (inp[14]) ? 1'b0 : 1'b1;
									assign node2289 = (inp[8]) ? node2309 : node2290;
										assign node2290 = (inp[11]) ? node2302 : node2291;
											assign node2291 = (inp[0]) ? node2297 : node2292;
												assign node2292 = (inp[4]) ? node2294 : 1'b1;
													assign node2294 = (inp[3]) ? 1'b0 : 1'b1;
												assign node2297 = (inp[14]) ? 1'b0 : node2298;
													assign node2298 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2302 = (inp[10]) ? 1'b0 : node2303;
												assign node2303 = (inp[3]) ? 1'b0 : node2304;
													assign node2304 = (inp[0]) ? 1'b0 : 1'b1;
										assign node2309 = (inp[10]) ? 1'b0 : node2310;
											assign node2310 = (inp[11]) ? 1'b0 : node2311;
												assign node2311 = (inp[0]) ? 1'b0 : 1'b1;
								assign node2316 = (inp[14]) ? node2346 : node2317;
									assign node2317 = (inp[8]) ? node2337 : node2318;
										assign node2318 = (inp[11]) ? node2330 : node2319;
											assign node2319 = (inp[10]) ? node2325 : node2320;
												assign node2320 = (inp[2]) ? node2322 : 1'b1;
													assign node2322 = (inp[4]) ? 1'b0 : 1'b1;
												assign node2325 = (inp[3]) ? 1'b0 : node2326;
													assign node2326 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2330 = (inp[4]) ? 1'b0 : node2331;
												assign node2331 = (inp[10]) ? 1'b0 : node2332;
													assign node2332 = (inp[0]) ? 1'b0 : 1'b1;
										assign node2337 = (inp[11]) ? 1'b0 : node2338;
											assign node2338 = (inp[0]) ? 1'b0 : node2339;
												assign node2339 = (inp[3]) ? 1'b0 : node2340;
													assign node2340 = (inp[10]) ? 1'b0 : 1'b1;
									assign node2346 = (inp[0]) ? 1'b0 : node2347;
										assign node2347 = (inp[10]) ? 1'b0 : node2348;
											assign node2348 = (inp[2]) ? 1'b0 : node2349;
												assign node2349 = (inp[3]) ? 1'b0 : node2350;
													assign node2350 = (inp[4]) ? 1'b0 : 1'b1;
				assign node2357 = (inp[7]) ? node2815 : node2358;
					assign node2358 = (inp[8]) ? node2596 : node2359;
						assign node2359 = (inp[14]) ? node2467 : node2360;
							assign node2360 = (inp[11]) ? node2402 : node2361;
								assign node2361 = (inp[4]) ? node2373 : node2362;
									assign node2362 = (inp[10]) ? node2364 : 1'b1;
										assign node2364 = (inp[5]) ? node2366 : 1'b1;
											assign node2366 = (inp[3]) ? node2368 : 1'b1;
												assign node2368 = (inp[2]) ? node2370 : 1'b1;
													assign node2370 = (inp[0]) ? 1'b0 : 1'b1;
									assign node2373 = (inp[12]) ? node2383 : node2374;
										assign node2374 = (inp[5]) ? node2376 : 1'b1;
											assign node2376 = (inp[0]) ? node2378 : 1'b1;
												assign node2378 = (inp[10]) ? node2380 : 1'b1;
													assign node2380 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2383 = (inp[10]) ? node2391 : node2384;
											assign node2384 = (inp[9]) ? node2386 : 1'b1;
												assign node2386 = (inp[3]) ? node2388 : 1'b1;
													assign node2388 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2391 = (inp[2]) ? node2397 : node2392;
												assign node2392 = (inp[0]) ? node2394 : 1'b1;
													assign node2394 = (inp[3]) ? 1'b0 : 1'b1;
												assign node2397 = (inp[9]) ? 1'b0 : node2398;
													assign node2398 = (inp[5]) ? 1'b0 : 1'b1;
								assign node2402 = (inp[2]) ? node2432 : node2403;
									assign node2403 = (inp[0]) ? node2413 : node2404;
										assign node2404 = (inp[4]) ? node2406 : 1'b1;
											assign node2406 = (inp[10]) ? node2408 : 1'b1;
												assign node2408 = (inp[5]) ? node2410 : 1'b1;
													assign node2410 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2413 = (inp[5]) ? node2421 : node2414;
											assign node2414 = (inp[9]) ? node2416 : 1'b1;
												assign node2416 = (inp[4]) ? node2418 : 1'b1;
													assign node2418 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2421 = (inp[12]) ? node2427 : node2422;
												assign node2422 = (inp[9]) ? node2424 : 1'b1;
													assign node2424 = (inp[3]) ? 1'b0 : 1'b1;
												assign node2427 = (inp[10]) ? 1'b0 : node2428;
													assign node2428 = (inp[3]) ? 1'b0 : 1'b1;
									assign node2432 = (inp[5]) ? node2450 : node2433;
										assign node2433 = (inp[9]) ? node2439 : node2434;
											assign node2434 = (inp[3]) ? node2436 : 1'b1;
												assign node2436 = (inp[4]) ? 1'b0 : 1'b1;
											assign node2439 = (inp[3]) ? node2445 : node2440;
												assign node2440 = (inp[10]) ? node2442 : 1'b1;
													assign node2442 = (inp[4]) ? 1'b0 : 1'b1;
												assign node2445 = (inp[0]) ? 1'b0 : node2446;
													assign node2446 = (inp[12]) ? 1'b0 : 1'b1;
										assign node2450 = (inp[0]) ? node2460 : node2451;
											assign node2451 = (inp[12]) ? node2455 : node2452;
												assign node2452 = (inp[4]) ? 1'b0 : 1'b1;
												assign node2455 = (inp[3]) ? 1'b0 : node2456;
													assign node2456 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2460 = (inp[4]) ? 1'b0 : node2461;
												assign node2461 = (inp[3]) ? 1'b0 : node2462;
													assign node2462 = (inp[9]) ? 1'b0 : 1'b1;
							assign node2467 = (inp[12]) ? node2529 : node2468;
								assign node2468 = (inp[11]) ? node2490 : node2469;
									assign node2469 = (inp[9]) ? node2471 : 1'b1;
										assign node2471 = (inp[2]) ? node2479 : node2472;
											assign node2472 = (inp[10]) ? node2474 : 1'b1;
												assign node2474 = (inp[0]) ? node2476 : 1'b1;
													assign node2476 = (inp[5]) ? 1'b0 : 1'b1;
											assign node2479 = (inp[3]) ? node2485 : node2480;
												assign node2480 = (inp[0]) ? node2482 : 1'b1;
													assign node2482 = (inp[4]) ? 1'b0 : 1'b1;
												assign node2485 = (inp[4]) ? 1'b0 : node2486;
													assign node2486 = (inp[0]) ? 1'b0 : 1'b1;
									assign node2490 = (inp[10]) ? node2510 : node2491;
										assign node2491 = (inp[2]) ? node2499 : node2492;
											assign node2492 = (inp[9]) ? node2494 : 1'b1;
												assign node2494 = (inp[5]) ? node2496 : 1'b1;
													assign node2496 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2499 = (inp[0]) ? node2505 : node2500;
												assign node2500 = (inp[3]) ? node2502 : 1'b1;
													assign node2502 = (inp[9]) ? 1'b1 : 1'b0;
												assign node2505 = (inp[4]) ? 1'b0 : node2506;
													assign node2506 = (inp[5]) ? 1'b0 : 1'b1;
										assign node2510 = (inp[9]) ? node2522 : node2511;
											assign node2511 = (inp[4]) ? node2517 : node2512;
												assign node2512 = (inp[2]) ? node2514 : 1'b1;
													assign node2514 = (inp[0]) ? 1'b0 : 1'b1;
												assign node2517 = (inp[0]) ? 1'b0 : node2518;
													assign node2518 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2522 = (inp[0]) ? 1'b0 : node2523;
												assign node2523 = (inp[2]) ? 1'b0 : node2524;
													assign node2524 = (inp[3]) ? 1'b0 : 1'b1;
								assign node2529 = (inp[10]) ? node2569 : node2530;
									assign node2530 = (inp[3]) ? node2550 : node2531;
										assign node2531 = (inp[4]) ? node2539 : node2532;
											assign node2532 = (inp[0]) ? node2534 : 1'b1;
												assign node2534 = (inp[2]) ? node2536 : 1'b1;
													assign node2536 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2539 = (inp[5]) ? node2545 : node2540;
												assign node2540 = (inp[11]) ? node2542 : 1'b1;
													assign node2542 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2545 = (inp[9]) ? 1'b0 : node2546;
													assign node2546 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2550 = (inp[9]) ? node2562 : node2551;
											assign node2551 = (inp[0]) ? node2557 : node2552;
												assign node2552 = (inp[5]) ? node2554 : 1'b1;
													assign node2554 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2557 = (inp[5]) ? 1'b0 : node2558;
													assign node2558 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2562 = (inp[11]) ? 1'b0 : node2563;
												assign node2563 = (inp[5]) ? 1'b0 : node2564;
													assign node2564 = (inp[0]) ? 1'b0 : 1'b1;
									assign node2569 = (inp[5]) ? node2589 : node2570;
										assign node2570 = (inp[2]) ? node2582 : node2571;
											assign node2571 = (inp[0]) ? node2577 : node2572;
												assign node2572 = (inp[11]) ? node2574 : 1'b1;
													assign node2574 = (inp[4]) ? 1'b0 : 1'b1;
												assign node2577 = (inp[3]) ? 1'b0 : node2578;
													assign node2578 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2582 = (inp[9]) ? 1'b0 : node2583;
												assign node2583 = (inp[11]) ? 1'b0 : node2584;
													assign node2584 = (inp[4]) ? 1'b0 : 1'b1;
										assign node2589 = (inp[0]) ? 1'b0 : node2590;
											assign node2590 = (inp[2]) ? 1'b0 : node2591;
												assign node2591 = (inp[9]) ? 1'b0 : 1'b1;
						assign node2596 = (inp[12]) ? node2730 : node2597;
							assign node2597 = (inp[9]) ? node2667 : node2598;
								assign node2598 = (inp[14]) ? node2628 : node2599;
									assign node2599 = (inp[3]) ? node2609 : node2600;
										assign node2600 = (inp[4]) ? node2602 : 1'b1;
											assign node2602 = (inp[11]) ? node2604 : 1'b1;
												assign node2604 = (inp[0]) ? node2606 : 1'b1;
													assign node2606 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2609 = (inp[10]) ? node2617 : node2610;
											assign node2610 = (inp[11]) ? node2612 : 1'b1;
												assign node2612 = (inp[0]) ? node2614 : 1'b1;
													assign node2614 = (inp[4]) ? 1'b0 : 1'b1;
											assign node2617 = (inp[5]) ? node2623 : node2618;
												assign node2618 = (inp[0]) ? node2620 : 1'b1;
													assign node2620 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2623 = (inp[11]) ? 1'b0 : node2624;
													assign node2624 = (inp[0]) ? 1'b0 : 1'b1;
									assign node2628 = (inp[3]) ? node2648 : node2629;
										assign node2629 = (inp[10]) ? node2637 : node2630;
											assign node2630 = (inp[5]) ? node2632 : 1'b1;
												assign node2632 = (inp[0]) ? node2634 : 1'b1;
													assign node2634 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2637 = (inp[5]) ? node2643 : node2638;
												assign node2638 = (inp[11]) ? node2640 : 1'b1;
													assign node2640 = (inp[4]) ? 1'b0 : 1'b1;
												assign node2643 = (inp[4]) ? 1'b0 : node2644;
													assign node2644 = (inp[2]) ? 1'b0 : 1'b0;
										assign node2648 = (inp[4]) ? node2660 : node2649;
											assign node2649 = (inp[2]) ? node2655 : node2650;
												assign node2650 = (inp[10]) ? node2652 : 1'b1;
													assign node2652 = (inp[0]) ? 1'b0 : 1'b1;
												assign node2655 = (inp[11]) ? 1'b0 : node2656;
													assign node2656 = (inp[5]) ? 1'b0 : 1'b1;
											assign node2660 = (inp[11]) ? 1'b0 : node2661;
												assign node2661 = (inp[0]) ? 1'b0 : node2662;
													assign node2662 = (inp[5]) ? 1'b0 : 1'b1;
								assign node2667 = (inp[10]) ? node2701 : node2668;
									assign node2668 = (inp[11]) ? node2688 : node2669;
										assign node2669 = (inp[3]) ? node2677 : node2670;
											assign node2670 = (inp[0]) ? node2672 : 1'b1;
												assign node2672 = (inp[4]) ? node2674 : 1'b1;
													assign node2674 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2677 = (inp[4]) ? node2683 : node2678;
												assign node2678 = (inp[0]) ? node2680 : 1'b1;
													assign node2680 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2683 = (inp[5]) ? 1'b0 : node2684;
													assign node2684 = (inp[0]) ? 1'b0 : 1'b1;
										assign node2688 = (inp[5]) ? 1'b0 : node2689;
											assign node2689 = (inp[0]) ? node2695 : node2690;
												assign node2690 = (inp[14]) ? node2692 : 1'b1;
													assign node2692 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2695 = (inp[2]) ? 1'b0 : node2696;
													assign node2696 = (inp[3]) ? 1'b0 : 1'b0;
									assign node2701 = (inp[0]) ? node2721 : node2702;
										assign node2702 = (inp[11]) ? node2714 : node2703;
											assign node2703 = (inp[2]) ? node2709 : node2704;
												assign node2704 = (inp[4]) ? node2706 : 1'b1;
													assign node2706 = (inp[3]) ? 1'b0 : 1'b1;
												assign node2709 = (inp[14]) ? 1'b0 : node2710;
													assign node2710 = (inp[5]) ? 1'b0 : 1'b1;
											assign node2714 = (inp[5]) ? 1'b0 : node2715;
												assign node2715 = (inp[3]) ? 1'b0 : node2716;
													assign node2716 = (inp[2]) ? 1'b0 : 1'b1;
										assign node2721 = (inp[3]) ? 1'b0 : node2722;
											assign node2722 = (inp[2]) ? 1'b0 : node2723;
												assign node2723 = (inp[14]) ? 1'b0 : node2724;
													assign node2724 = (inp[4]) ? 1'b0 : 1'b1;
							assign node2730 = (inp[5]) ? node2784 : node2731;
								assign node2731 = (inp[11]) ? node2765 : node2732;
									assign node2732 = (inp[14]) ? node2748 : node2733;
										assign node2733 = (inp[0]) ? node2741 : node2734;
											assign node2734 = (inp[9]) ? node2736 : 1'b1;
												assign node2736 = (inp[2]) ? node2738 : 1'b1;
													assign node2738 = (inp[4]) ? 1'b0 : 1'b1;
											assign node2741 = (inp[3]) ? 1'b0 : node2742;
												assign node2742 = (inp[9]) ? node2744 : 1'b1;
													assign node2744 = (inp[2]) ? 1'b0 : 1'b1;
										assign node2748 = (inp[4]) ? node2758 : node2749;
											assign node2749 = (inp[0]) ? node2751 : 1'b1;
												assign node2751 = (inp[10]) ? node2755 : node2752;
													assign node2752 = (inp[9]) ? 1'b0 : 1'b1;
													assign node2755 = (inp[3]) ? 1'b0 : 1'b0;
											assign node2758 = (inp[3]) ? 1'b0 : node2759;
												assign node2759 = (inp[9]) ? 1'b0 : node2760;
													assign node2760 = (inp[0]) ? 1'b0 : 1'b1;
									assign node2765 = (inp[4]) ? 1'b0 : node2766;
										assign node2766 = (inp[10]) ? node2778 : node2767;
											assign node2767 = (inp[3]) ? node2773 : node2768;
												assign node2768 = (inp[9]) ? node2770 : 1'b1;
													assign node2770 = (inp[0]) ? 1'b0 : 1'b1;
												assign node2773 = (inp[9]) ? 1'b0 : node2774;
													assign node2774 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2778 = (inp[0]) ? 1'b0 : node2779;
												assign node2779 = (inp[14]) ? 1'b1 : 1'b0;
								assign node2784 = (inp[0]) ? 1'b0 : node2785;
									assign node2785 = (inp[3]) ? node2805 : node2786;
										assign node2786 = (inp[9]) ? node2798 : node2787;
											assign node2787 = (inp[4]) ? node2793 : node2788;
												assign node2788 = (inp[11]) ? node2790 : 1'b1;
													assign node2790 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2793 = (inp[10]) ? 1'b0 : node2794;
													assign node2794 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2798 = (inp[14]) ? 1'b0 : node2799;
												assign node2799 = (inp[4]) ? 1'b0 : node2800;
													assign node2800 = (inp[2]) ? 1'b0 : 1'b1;
										assign node2805 = (inp[2]) ? 1'b0 : node2806;
											assign node2806 = (inp[4]) ? 1'b0 : node2807;
												assign node2807 = (inp[14]) ? 1'b0 : node2808;
													assign node2808 = (inp[9]) ? 1'b0 : 1'b1;
					assign node2815 = (inp[5]) ? node3063 : node2816;
						assign node2816 = (inp[3]) ? node2956 : node2817;
							assign node2817 = (inp[9]) ? node2887 : node2818;
								assign node2818 = (inp[2]) ? node2848 : node2819;
									assign node2819 = (inp[12]) ? node2829 : node2820;
										assign node2820 = (inp[8]) ? node2822 : 1'b1;
											assign node2822 = (inp[0]) ? node2824 : 1'b1;
												assign node2824 = (inp[10]) ? node2826 : 1'b1;
													assign node2826 = (inp[4]) ? 1'b0 : 1'b0;
										assign node2829 = (inp[4]) ? node2837 : node2830;
											assign node2830 = (inp[8]) ? node2832 : 1'b1;
												assign node2832 = (inp[0]) ? node2834 : 1'b1;
													assign node2834 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2837 = (inp[14]) ? node2843 : node2838;
												assign node2838 = (inp[10]) ? node2840 : 1'b1;
													assign node2840 = (inp[8]) ? 1'b0 : 1'b1;
												assign node2843 = (inp[11]) ? 1'b0 : node2844;
													assign node2844 = (inp[8]) ? 1'b0 : 1'b1;
									assign node2848 = (inp[4]) ? node2868 : node2849;
										assign node2849 = (inp[11]) ? node2857 : node2850;
											assign node2850 = (inp[10]) ? node2852 : 1'b1;
												assign node2852 = (inp[14]) ? node2854 : 1'b1;
													assign node2854 = (inp[0]) ? 1'b0 : 1'b1;
											assign node2857 = (inp[0]) ? node2863 : node2858;
												assign node2858 = (inp[8]) ? node2860 : 1'b1;
													assign node2860 = (inp[14]) ? 1'b0 : 1'b1;
												assign node2863 = (inp[12]) ? 1'b0 : node2864;
													assign node2864 = (inp[14]) ? 1'b0 : 1'b1;
										assign node2868 = (inp[0]) ? node2880 : node2869;
											assign node2869 = (inp[10]) ? node2875 : node2870;
												assign node2870 = (inp[14]) ? node2872 : 1'b1;
													assign node2872 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2875 = (inp[12]) ? 1'b0 : node2876;
													assign node2876 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2880 = (inp[8]) ? 1'b0 : node2881;
												assign node2881 = (inp[11]) ? 1'b0 : node2882;
													assign node2882 = (inp[12]) ? 1'b0 : 1'b1;
								assign node2887 = (inp[14]) ? node2927 : node2888;
									assign node2888 = (inp[4]) ? node2908 : node2889;
										assign node2889 = (inp[0]) ? node2897 : node2890;
											assign node2890 = (inp[10]) ? node2892 : 1'b1;
												assign node2892 = (inp[12]) ? node2894 : 1'b1;
													assign node2894 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2897 = (inp[8]) ? node2903 : node2898;
												assign node2898 = (inp[12]) ? node2900 : 1'b1;
													assign node2900 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2903 = (inp[2]) ? 1'b0 : node2904;
													assign node2904 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2908 = (inp[8]) ? node2920 : node2909;
											assign node2909 = (inp[0]) ? node2915 : node2910;
												assign node2910 = (inp[2]) ? node2912 : 1'b1;
													assign node2912 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2915 = (inp[11]) ? 1'b0 : node2916;
													assign node2916 = (inp[12]) ? 1'b0 : 1'b1;
											assign node2920 = (inp[11]) ? 1'b0 : node2921;
												assign node2921 = (inp[2]) ? 1'b0 : node2922;
													assign node2922 = (inp[12]) ? 1'b0 : 1'b1;
									assign node2927 = (inp[4]) ? node2947 : node2928;
										assign node2928 = (inp[8]) ? node2940 : node2929;
											assign node2929 = (inp[12]) ? node2935 : node2930;
												assign node2930 = (inp[11]) ? node2932 : 1'b1;
													assign node2932 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2935 = (inp[2]) ? 1'b0 : node2936;
													assign node2936 = (inp[0]) ? 1'b0 : 1'b1;
											assign node2940 = (inp[11]) ? 1'b0 : node2941;
												assign node2941 = (inp[2]) ? 1'b0 : node2942;
													assign node2942 = (inp[12]) ? 1'b0 : 1'b1;
										assign node2947 = (inp[11]) ? 1'b0 : node2948;
											assign node2948 = (inp[8]) ? 1'b0 : node2949;
												assign node2949 = (inp[12]) ? 1'b0 : node2950;
													assign node2950 = (inp[0]) ? 1'b0 : 1'b1;
							assign node2956 = (inp[11]) ? node3022 : node2957;
								assign node2957 = (inp[4]) ? node2993 : node2958;
									assign node2958 = (inp[9]) ? node2976 : node2959;
										assign node2959 = (inp[8]) ? node2967 : node2960;
											assign node2960 = (inp[2]) ? node2962 : 1'b1;
												assign node2962 = (inp[14]) ? node2964 : 1'b1;
													assign node2964 = (inp[0]) ? 1'b0 : 1'b1;
											assign node2967 = (inp[12]) ? node2971 : node2968;
												assign node2968 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2971 = (inp[10]) ? 1'b0 : node2972;
													assign node2972 = (inp[2]) ? 1'b0 : 1'b1;
										assign node2976 = (inp[0]) ? node2988 : node2977;
											assign node2977 = (inp[12]) ? node2983 : node2978;
												assign node2978 = (inp[14]) ? node2980 : 1'b1;
													assign node2980 = (inp[8]) ? 1'b0 : 1'b1;
												assign node2983 = (inp[8]) ? 1'b0 : node2984;
													assign node2984 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2988 = (inp[10]) ? 1'b0 : node2989;
												assign node2989 = (inp[2]) ? 1'b0 : 1'b1;
									assign node2993 = (inp[12]) ? node3013 : node2994;
										assign node2994 = (inp[9]) ? node3006 : node2995;
											assign node2995 = (inp[10]) ? node3001 : node2996;
												assign node2996 = (inp[8]) ? node2998 : 1'b1;
													assign node2998 = (inp[14]) ? 1'b0 : 1'b1;
												assign node3001 = (inp[2]) ? 1'b0 : node3002;
													assign node3002 = (inp[14]) ? 1'b0 : 1'b1;
											assign node3006 = (inp[0]) ? 1'b0 : node3007;
												assign node3007 = (inp[10]) ? 1'b0 : node3008;
													assign node3008 = (inp[8]) ? 1'b0 : 1'b1;
										assign node3013 = (inp[8]) ? 1'b0 : node3014;
											assign node3014 = (inp[14]) ? 1'b0 : node3015;
												assign node3015 = (inp[10]) ? 1'b0 : node3016;
													assign node3016 = (inp[9]) ? 1'b0 : 1'b1;
								assign node3022 = (inp[0]) ? node3052 : node3023;
									assign node3023 = (inp[8]) ? node3043 : node3024;
										assign node3024 = (inp[14]) ? node3036 : node3025;
											assign node3025 = (inp[10]) ? node3031 : node3026;
												assign node3026 = (inp[9]) ? node3028 : 1'b1;
													assign node3028 = (inp[4]) ? 1'b0 : 1'b1;
												assign node3031 = (inp[9]) ? 1'b0 : node3032;
													assign node3032 = (inp[12]) ? 1'b0 : 1'b1;
											assign node3036 = (inp[2]) ? 1'b0 : node3037;
												assign node3037 = (inp[4]) ? node3039 : 1'b1;
													assign node3039 = (inp[12]) ? 1'b0 : 1'b0;
										assign node3043 = (inp[10]) ? 1'b0 : node3044;
											assign node3044 = (inp[12]) ? 1'b0 : node3045;
												assign node3045 = (inp[14]) ? 1'b0 : node3046;
													assign node3046 = (inp[9]) ? 1'b0 : 1'b1;
									assign node3052 = (inp[8]) ? 1'b0 : node3053;
										assign node3053 = (inp[2]) ? 1'b0 : node3054;
											assign node3054 = (inp[9]) ? 1'b0 : node3055;
												assign node3055 = (inp[4]) ? 1'b0 : node3056;
													assign node3056 = (inp[10]) ? 1'b0 : 1'b0;
						assign node3063 = (inp[4]) ? node3173 : node3064;
							assign node3064 = (inp[14]) ? node3132 : node3065;
								assign node3065 = (inp[0]) ? node3103 : node3066;
									assign node3066 = (inp[10]) ? node3084 : node3067;
										assign node3067 = (inp[8]) ? node3073 : node3068;
											assign node3068 = (inp[9]) ? node3070 : 1'b1;
												assign node3070 = (inp[12]) ? 1'b0 : 1'b1;
											assign node3073 = (inp[3]) ? node3079 : node3074;
												assign node3074 = (inp[11]) ? node3076 : 1'b1;
													assign node3076 = (inp[9]) ? 1'b0 : 1'b1;
												assign node3079 = (inp[2]) ? 1'b0 : node3080;
													assign node3080 = (inp[9]) ? 1'b0 : 1'b1;
										assign node3084 = (inp[8]) ? node3098 : node3085;
											assign node3085 = (inp[2]) ? node3091 : node3086;
												assign node3086 = (inp[12]) ? node3088 : 1'b1;
													assign node3088 = (inp[3]) ? 1'b0 : 1'b1;
												assign node3091 = (inp[11]) ? node3095 : node3092;
													assign node3092 = (inp[12]) ? 1'b0 : 1'b1;
													assign node3095 = (inp[3]) ? 1'b0 : 1'b0;
											assign node3098 = (inp[11]) ? 1'b0 : node3099;
												assign node3099 = (inp[3]) ? 1'b0 : 1'b1;
									assign node3103 = (inp[11]) ? node3123 : node3104;
										assign node3104 = (inp[10]) ? node3116 : node3105;
											assign node3105 = (inp[3]) ? node3111 : node3106;
												assign node3106 = (inp[12]) ? node3108 : 1'b1;
													assign node3108 = (inp[2]) ? 1'b0 : 1'b1;
												assign node3111 = (inp[2]) ? 1'b0 : node3112;
													assign node3112 = (inp[9]) ? 1'b0 : 1'b1;
											assign node3116 = (inp[12]) ? 1'b0 : node3117;
												assign node3117 = (inp[9]) ? 1'b0 : node3118;
													assign node3118 = (inp[8]) ? 1'b0 : 1'b1;
										assign node3123 = (inp[2]) ? 1'b0 : node3124;
											assign node3124 = (inp[12]) ? 1'b0 : node3125;
												assign node3125 = (inp[8]) ? 1'b0 : node3126;
													assign node3126 = (inp[9]) ? 1'b0 : 1'b1;
								assign node3132 = (inp[9]) ? node3162 : node3133;
									assign node3133 = (inp[12]) ? node3153 : node3134;
										assign node3134 = (inp[3]) ? node3146 : node3135;
											assign node3135 = (inp[11]) ? node3141 : node3136;
												assign node3136 = (inp[2]) ? node3138 : 1'b1;
													assign node3138 = (inp[0]) ? 1'b0 : 1'b1;
												assign node3141 = (inp[8]) ? 1'b0 : node3142;
													assign node3142 = (inp[2]) ? 1'b0 : 1'b1;
											assign node3146 = (inp[11]) ? 1'b0 : node3147;
												assign node3147 = (inp[8]) ? 1'b0 : node3148;
													assign node3148 = (inp[10]) ? 1'b0 : 1'b1;
										assign node3153 = (inp[2]) ? 1'b0 : node3154;
											assign node3154 = (inp[0]) ? 1'b0 : node3155;
												assign node3155 = (inp[10]) ? node3157 : 1'b1;
													assign node3157 = (inp[3]) ? 1'b0 : 1'b0;
									assign node3162 = (inp[11]) ? 1'b0 : node3163;
										assign node3163 = (inp[3]) ? 1'b0 : node3164;
											assign node3164 = (inp[8]) ? 1'b0 : node3165;
												assign node3165 = (inp[10]) ? node3167 : 1'b1;
													assign node3167 = (inp[2]) ? 1'b0 : 1'b0;
							assign node3173 = (inp[14]) ? node3215 : node3174;
								assign node3174 = (inp[0]) ? node3204 : node3175;
									assign node3175 = (inp[10]) ? node3195 : node3176;
										assign node3176 = (inp[2]) ? node3188 : node3177;
											assign node3177 = (inp[11]) ? node3183 : node3178;
												assign node3178 = (inp[8]) ? node3180 : 1'b1;
													assign node3180 = (inp[3]) ? 1'b0 : 1'b1;
												assign node3183 = (inp[12]) ? 1'b0 : node3184;
													assign node3184 = (inp[3]) ? 1'b0 : 1'b1;
											assign node3188 = (inp[12]) ? 1'b0 : node3189;
												assign node3189 = (inp[3]) ? 1'b0 : node3190;
													assign node3190 = (inp[11]) ? 1'b0 : 1'b1;
										assign node3195 = (inp[2]) ? 1'b0 : node3196;
											assign node3196 = (inp[9]) ? 1'b0 : node3197;
												assign node3197 = (inp[11]) ? 1'b0 : node3198;
													assign node3198 = (inp[8]) ? 1'b0 : 1'b1;
									assign node3204 = (inp[12]) ? 1'b0 : node3205;
										assign node3205 = (inp[9]) ? 1'b0 : node3206;
											assign node3206 = (inp[2]) ? 1'b0 : node3207;
												assign node3207 = (inp[3]) ? 1'b0 : node3208;
													assign node3208 = (inp[8]) ? 1'b0 : 1'b1;
								assign node3215 = (inp[0]) ? node3217 : 1'b0;
									assign node3217 = (inp[10]) ? 1'b0 : node3218;
										assign node3218 = (inp[12]) ? 1'b0 : node3219;
											assign node3219 = (inp[3]) ? 1'b0 : node3220;
												assign node3220 = (inp[8]) ? 1'b0 : node3221;
													assign node3221 = (inp[9]) ? 1'b0 : 1'b0;
		assign node3228 = (inp[3]) ? node4934 : node3229;
			assign node3229 = (inp[11]) ? node4081 : node3230;
				assign node3230 = (inp[4]) ? node3606 : node3231;
					assign node3231 = (inp[10]) ? node3391 : node3232;
						assign node3232 = (inp[12]) ? node3288 : node3233;
							assign node3233 = (inp[8]) ? node3247 : node3234;
								assign node3234 = (inp[7]) ? node3236 : 1'b1;
									assign node3236 = (inp[0]) ? node3238 : 1'b1;
										assign node3238 = (inp[2]) ? node3240 : 1'b1;
											assign node3240 = (inp[6]) ? node3242 : 1'b1;
												assign node3242 = (inp[13]) ? node3244 : 1'b1;
													assign node3244 = (inp[5]) ? 1'b0 : 1'b1;
								assign node3247 = (inp[13]) ? node3259 : node3248;
									assign node3248 = (inp[5]) ? node3250 : 1'b1;
										assign node3250 = (inp[0]) ? node3252 : 1'b1;
											assign node3252 = (inp[6]) ? node3254 : 1'b1;
												assign node3254 = (inp[9]) ? node3256 : 1'b1;
													assign node3256 = (inp[14]) ? 1'b0 : 1'b1;
									assign node3259 = (inp[9]) ? node3269 : node3260;
										assign node3260 = (inp[6]) ? node3262 : 1'b1;
											assign node3262 = (inp[0]) ? node3264 : 1'b1;
												assign node3264 = (inp[7]) ? node3266 : 1'b1;
													assign node3266 = (inp[2]) ? 1'b0 : 1'b1;
										assign node3269 = (inp[2]) ? node3277 : node3270;
											assign node3270 = (inp[0]) ? node3272 : 1'b1;
												assign node3272 = (inp[7]) ? node3274 : 1'b1;
													assign node3274 = (inp[14]) ? 1'b0 : 1'b1;
											assign node3277 = (inp[7]) ? node3283 : node3278;
												assign node3278 = (inp[14]) ? node3280 : 1'b1;
													assign node3280 = (inp[6]) ? 1'b0 : 1'b0;
												assign node3283 = (inp[6]) ? 1'b0 : node3284;
													assign node3284 = (inp[14]) ? 1'b0 : 1'b1;
							assign node3288 = (inp[14]) ? node3330 : node3289;
								assign node3289 = (inp[5]) ? node3301 : node3290;
									assign node3290 = (inp[0]) ? node3292 : 1'b1;
										assign node3292 = (inp[8]) ? node3294 : 1'b1;
											assign node3294 = (inp[13]) ? node3296 : 1'b1;
												assign node3296 = (inp[9]) ? node3298 : 1'b1;
													assign node3298 = (inp[6]) ? 1'b0 : 1'b1;
									assign node3301 = (inp[6]) ? node3311 : node3302;
										assign node3302 = (inp[9]) ? node3304 : 1'b1;
											assign node3304 = (inp[8]) ? node3306 : 1'b1;
												assign node3306 = (inp[13]) ? node3308 : 1'b1;
													assign node3308 = (inp[2]) ? 1'b0 : 1'b1;
										assign node3311 = (inp[0]) ? node3319 : node3312;
											assign node3312 = (inp[9]) ? node3314 : 1'b1;
												assign node3314 = (inp[13]) ? node3316 : 1'b1;
													assign node3316 = (inp[2]) ? 1'b0 : 1'b1;
											assign node3319 = (inp[13]) ? node3325 : node3320;
												assign node3320 = (inp[7]) ? node3322 : 1'b1;
													assign node3322 = (inp[2]) ? 1'b0 : 1'b0;
												assign node3325 = (inp[8]) ? 1'b0 : node3326;
													assign node3326 = (inp[2]) ? 1'b0 : 1'b1;
								assign node3330 = (inp[8]) ? node3356 : node3331;
									assign node3331 = (inp[13]) ? node3341 : node3332;
										assign node3332 = (inp[7]) ? node3334 : 1'b1;
											assign node3334 = (inp[9]) ? node3336 : 1'b1;
												assign node3336 = (inp[2]) ? node3338 : 1'b1;
													assign node3338 = (inp[6]) ? 1'b0 : 1'b1;
										assign node3341 = (inp[5]) ? node3349 : node3342;
											assign node3342 = (inp[6]) ? node3344 : 1'b1;
												assign node3344 = (inp[2]) ? node3346 : 1'b1;
													assign node3346 = (inp[9]) ? 1'b1 : 1'b0;
											assign node3349 = (inp[0]) ? 1'b0 : node3350;
												assign node3350 = (inp[2]) ? node3352 : 1'b1;
													assign node3352 = (inp[7]) ? 1'b0 : 1'b1;
									assign node3356 = (inp[0]) ? node3376 : node3357;
										assign node3357 = (inp[2]) ? node3365 : node3358;
											assign node3358 = (inp[13]) ? 1'b1 : node3359;
												assign node3359 = (inp[9]) ? node3361 : 1'b1;
													assign node3361 = (inp[7]) ? 1'b0 : 1'b1;
											assign node3365 = (inp[5]) ? node3371 : node3366;
												assign node3366 = (inp[6]) ? node3368 : 1'b1;
													assign node3368 = (inp[9]) ? 1'b0 : 1'b1;
												assign node3371 = (inp[13]) ? 1'b0 : node3372;
													assign node3372 = (inp[6]) ? 1'b0 : 1'b1;
										assign node3376 = (inp[6]) ? node3384 : node3377;
											assign node3377 = (inp[2]) ? node3379 : 1'b1;
												assign node3379 = (inp[9]) ? 1'b0 : node3380;
													assign node3380 = (inp[5]) ? 1'b0 : 1'b1;
											assign node3384 = (inp[9]) ? 1'b0 : node3385;
												assign node3385 = (inp[5]) ? 1'b0 : node3386;
													assign node3386 = (inp[13]) ? 1'b0 : 1'b1;
						assign node3391 = (inp[12]) ? node3493 : node3392;
							assign node3392 = (inp[14]) ? node3430 : node3393;
								assign node3393 = (inp[8]) ? node3405 : node3394;
									assign node3394 = (inp[9]) ? node3396 : 1'b1;
										assign node3396 = (inp[6]) ? node3398 : 1'b1;
											assign node3398 = (inp[5]) ? node3400 : 1'b1;
												assign node3400 = (inp[2]) ? node3402 : 1'b1;
													assign node3402 = (inp[0]) ? 1'b0 : 1'b1;
									assign node3405 = (inp[5]) ? node3415 : node3406;
										assign node3406 = (inp[0]) ? node3408 : 1'b1;
											assign node3408 = (inp[7]) ? node3410 : 1'b1;
												assign node3410 = (inp[6]) ? node3412 : 1'b1;
													assign node3412 = (inp[13]) ? 1'b0 : 1'b1;
										assign node3415 = (inp[9]) ? node3423 : node3416;
											assign node3416 = (inp[6]) ? node3418 : 1'b1;
												assign node3418 = (inp[13]) ? node3420 : 1'b1;
													assign node3420 = (inp[0]) ? 1'b0 : 1'b0;
											assign node3423 = (inp[7]) ? 1'b0 : node3424;
												assign node3424 = (inp[0]) ? node3426 : 1'b1;
													assign node3426 = (inp[6]) ? 1'b0 : 1'b1;
								assign node3430 = (inp[5]) ? node3458 : node3431;
									assign node3431 = (inp[13]) ? node3439 : node3432;
										assign node3432 = (inp[9]) ? node3434 : 1'b1;
											assign node3434 = (inp[6]) ? node3436 : 1'b1;
												assign node3436 = (inp[2]) ? 1'b0 : 1'b1;
										assign node3439 = (inp[0]) ? node3447 : node3440;
											assign node3440 = (inp[6]) ? node3442 : 1'b1;
												assign node3442 = (inp[8]) ? node3444 : 1'b1;
													assign node3444 = (inp[9]) ? 1'b0 : 1'b0;
											assign node3447 = (inp[7]) ? node3453 : node3448;
												assign node3448 = (inp[6]) ? node3450 : 1'b1;
													assign node3450 = (inp[8]) ? 1'b0 : 1'b1;
												assign node3453 = (inp[6]) ? 1'b0 : node3454;
													assign node3454 = (inp[9]) ? 1'b0 : 1'b0;
									assign node3458 = (inp[2]) ? node3476 : node3459;
										assign node3459 = (inp[8]) ? node3465 : node3460;
											assign node3460 = (inp[13]) ? node3462 : 1'b1;
												assign node3462 = (inp[6]) ? 1'b0 : 1'b1;
											assign node3465 = (inp[0]) ? node3471 : node3466;
												assign node3466 = (inp[7]) ? node3468 : 1'b1;
													assign node3468 = (inp[6]) ? 1'b0 : 1'b1;
												assign node3471 = (inp[9]) ? 1'b0 : node3472;
													assign node3472 = (inp[7]) ? 1'b0 : 1'b1;
										assign node3476 = (inp[0]) ? node3488 : node3477;
											assign node3477 = (inp[7]) ? node3483 : node3478;
												assign node3478 = (inp[13]) ? node3480 : 1'b1;
													assign node3480 = (inp[8]) ? 1'b0 : 1'b1;
												assign node3483 = (inp[8]) ? 1'b0 : node3484;
													assign node3484 = (inp[9]) ? 1'b0 : 1'b1;
											assign node3488 = (inp[9]) ? 1'b0 : node3489;
												assign node3489 = (inp[6]) ? 1'b0 : 1'b1;
							assign node3493 = (inp[2]) ? node3555 : node3494;
								assign node3494 = (inp[8]) ? node3516 : node3495;
									assign node3495 = (inp[7]) ? node3497 : 1'b1;
										assign node3497 = (inp[6]) ? node3505 : node3498;
											assign node3498 = (inp[5]) ? node3500 : 1'b1;
												assign node3500 = (inp[13]) ? node3502 : 1'b1;
													assign node3502 = (inp[0]) ? 1'b0 : 1'b1;
											assign node3505 = (inp[13]) ? node3511 : node3506;
												assign node3506 = (inp[9]) ? node3508 : 1'b1;
													assign node3508 = (inp[5]) ? 1'b0 : 1'b1;
												assign node3511 = (inp[0]) ? 1'b0 : node3512;
													assign node3512 = (inp[9]) ? 1'b0 : 1'b1;
									assign node3516 = (inp[9]) ? node3538 : node3517;
										assign node3517 = (inp[6]) ? node3527 : node3518;
											assign node3518 = (inp[5]) ? node3520 : 1'b1;
												assign node3520 = (inp[7]) ? node3524 : node3521;
													assign node3521 = (inp[0]) ? 1'b1 : 1'b1;
													assign node3524 = (inp[13]) ? 1'b0 : 1'b0;
											assign node3527 = (inp[5]) ? node3533 : node3528;
												assign node3528 = (inp[7]) ? node3530 : 1'b1;
													assign node3530 = (inp[14]) ? 1'b0 : 1'b0;
												assign node3533 = (inp[14]) ? 1'b0 : node3534;
													assign node3534 = (inp[7]) ? 1'b0 : 1'b1;
										assign node3538 = (inp[7]) ? node3548 : node3539;
											assign node3539 = (inp[0]) ? node3543 : node3540;
												assign node3540 = (inp[13]) ? 1'b0 : 1'b1;
												assign node3543 = (inp[5]) ? 1'b0 : node3544;
													assign node3544 = (inp[14]) ? 1'b0 : 1'b1;
											assign node3548 = (inp[14]) ? 1'b0 : node3549;
												assign node3549 = (inp[0]) ? 1'b0 : node3550;
													assign node3550 = (inp[13]) ? 1'b0 : 1'b1;
								assign node3555 = (inp[14]) ? node3585 : node3556;
									assign node3556 = (inp[13]) ? node3566 : node3557;
										assign node3557 = (inp[6]) ? node3559 : 1'b1;
											assign node3559 = (inp[0]) ? node3561 : 1'b1;
												assign node3561 = (inp[9]) ? 1'b0 : node3562;
													assign node3562 = (inp[8]) ? 1'b0 : 1'b1;
										assign node3566 = (inp[7]) ? node3578 : node3567;
											assign node3567 = (inp[9]) ? node3573 : node3568;
												assign node3568 = (inp[5]) ? node3570 : 1'b1;
													assign node3570 = (inp[8]) ? 1'b0 : 1'b1;
												assign node3573 = (inp[6]) ? 1'b0 : node3574;
													assign node3574 = (inp[0]) ? 1'b0 : 1'b1;
											assign node3578 = (inp[8]) ? 1'b0 : node3579;
												assign node3579 = (inp[6]) ? 1'b0 : node3580;
													assign node3580 = (inp[0]) ? 1'b0 : 1'b1;
									assign node3585 = (inp[6]) ? 1'b0 : node3586;
										assign node3586 = (inp[8]) ? node3598 : node3587;
											assign node3587 = (inp[5]) ? node3593 : node3588;
												assign node3588 = (inp[13]) ? node3590 : 1'b1;
													assign node3590 = (inp[9]) ? 1'b0 : 1'b1;
												assign node3593 = (inp[7]) ? 1'b0 : node3594;
													assign node3594 = (inp[13]) ? 1'b0 : 1'b1;
											assign node3598 = (inp[9]) ? 1'b0 : node3599;
												assign node3599 = (inp[0]) ? 1'b0 : node3600;
													assign node3600 = (inp[7]) ? 1'b0 : 1'b1;
					assign node3606 = (inp[9]) ? node3844 : node3607;
						assign node3607 = (inp[13]) ? node3717 : node3608;
							assign node3608 = (inp[2]) ? node3652 : node3609;
								assign node3609 = (inp[12]) ? node3621 : node3610;
									assign node3610 = (inp[8]) ? node3612 : 1'b1;
										assign node3612 = (inp[5]) ? node3614 : 1'b1;
											assign node3614 = (inp[0]) ? node3616 : 1'b1;
												assign node3616 = (inp[7]) ? node3618 : 1'b1;
													assign node3618 = (inp[10]) ? 1'b0 : 1'b1;
									assign node3621 = (inp[7]) ? node3631 : node3622;
										assign node3622 = (inp[14]) ? node3624 : 1'b1;
											assign node3624 = (inp[8]) ? node3626 : 1'b1;
												assign node3626 = (inp[10]) ? node3628 : 1'b1;
													assign node3628 = (inp[0]) ? 1'b0 : 1'b1;
										assign node3631 = (inp[6]) ? node3641 : node3632;
											assign node3632 = (inp[0]) ? node3634 : 1'b1;
												assign node3634 = (inp[8]) ? node3638 : node3635;
													assign node3635 = (inp[14]) ? 1'b1 : 1'b1;
													assign node3638 = (inp[10]) ? 1'b0 : 1'b1;
											assign node3641 = (inp[5]) ? node3647 : node3642;
												assign node3642 = (inp[14]) ? node3644 : 1'b1;
													assign node3644 = (inp[8]) ? 1'b0 : 1'b1;
												assign node3647 = (inp[0]) ? 1'b0 : node3648;
													assign node3648 = (inp[14]) ? 1'b0 : 1'b1;
								assign node3652 = (inp[6]) ? node3678 : node3653;
									assign node3653 = (inp[14]) ? node3663 : node3654;
										assign node3654 = (inp[12]) ? node3656 : 1'b1;
											assign node3656 = (inp[0]) ? node3658 : 1'b1;
												assign node3658 = (inp[8]) ? node3660 : 1'b1;
													assign node3660 = (inp[7]) ? 1'b0 : 1'b1;
										assign node3663 = (inp[7]) ? node3671 : node3664;
											assign node3664 = (inp[8]) ? node3666 : 1'b1;
												assign node3666 = (inp[0]) ? node3668 : 1'b1;
													assign node3668 = (inp[5]) ? 1'b0 : 1'b1;
											assign node3671 = (inp[0]) ? 1'b0 : node3672;
												assign node3672 = (inp[12]) ? node3674 : 1'b1;
													assign node3674 = (inp[8]) ? 1'b0 : 1'b1;
									assign node3678 = (inp[10]) ? node3696 : node3679;
										assign node3679 = (inp[8]) ? node3685 : node3680;
											assign node3680 = (inp[0]) ? node3682 : 1'b1;
												assign node3682 = (inp[5]) ? 1'b0 : 1'b1;
											assign node3685 = (inp[5]) ? node3691 : node3686;
												assign node3686 = (inp[0]) ? node3688 : 1'b1;
													assign node3688 = (inp[7]) ? 1'b0 : 1'b1;
												assign node3691 = (inp[14]) ? 1'b0 : node3692;
													assign node3692 = (inp[0]) ? 1'b0 : 1'b1;
										assign node3696 = (inp[14]) ? node3710 : node3697;
											assign node3697 = (inp[8]) ? node3703 : node3698;
												assign node3698 = (inp[12]) ? node3700 : 1'b1;
													assign node3700 = (inp[0]) ? 1'b0 : 1'b1;
												assign node3703 = (inp[7]) ? node3707 : node3704;
													assign node3704 = (inp[5]) ? 1'b0 : 1'b1;
													assign node3707 = (inp[5]) ? 1'b0 : 1'b0;
											assign node3710 = (inp[8]) ? 1'b0 : node3711;
												assign node3711 = (inp[12]) ? 1'b0 : node3712;
													assign node3712 = (inp[7]) ? 1'b0 : 1'b1;
							assign node3717 = (inp[0]) ? node3775 : node3718;
								assign node3718 = (inp[10]) ? node3748 : node3719;
									assign node3719 = (inp[6]) ? node3729 : node3720;
										assign node3720 = (inp[14]) ? node3722 : 1'b1;
											assign node3722 = (inp[5]) ? node3724 : 1'b1;
												assign node3724 = (inp[12]) ? node3726 : 1'b1;
													assign node3726 = (inp[8]) ? 1'b1 : 1'b0;
										assign node3729 = (inp[2]) ? node3737 : node3730;
											assign node3730 = (inp[7]) ? node3732 : 1'b1;
												assign node3732 = (inp[14]) ? node3734 : 1'b1;
													assign node3734 = (inp[12]) ? 1'b0 : 1'b1;
											assign node3737 = (inp[5]) ? node3743 : node3738;
												assign node3738 = (inp[8]) ? node3740 : 1'b1;
													assign node3740 = (inp[12]) ? 1'b0 : 1'b1;
												assign node3743 = (inp[14]) ? 1'b0 : node3744;
													assign node3744 = (inp[7]) ? 1'b0 : 1'b1;
									assign node3748 = (inp[14]) ? node3766 : node3749;
										assign node3749 = (inp[2]) ? node3757 : node3750;
											assign node3750 = (inp[7]) ? node3752 : 1'b1;
												assign node3752 = (inp[6]) ? node3754 : 1'b1;
													assign node3754 = (inp[5]) ? 1'b0 : 1'b1;
											assign node3757 = (inp[7]) ? node3761 : node3758;
												assign node3758 = (inp[12]) ? 1'b0 : 1'b1;
												assign node3761 = (inp[5]) ? 1'b0 : node3762;
													assign node3762 = (inp[8]) ? 1'b0 : 1'b0;
										assign node3766 = (inp[12]) ? 1'b0 : node3767;
											assign node3767 = (inp[5]) ? 1'b0 : node3768;
												assign node3768 = (inp[8]) ? node3770 : 1'b1;
													assign node3770 = (inp[7]) ? 1'b0 : 1'b1;
								assign node3775 = (inp[8]) ? node3815 : node3776;
									assign node3776 = (inp[6]) ? node3796 : node3777;
										assign node3777 = (inp[10]) ? node3785 : node3778;
											assign node3778 = (inp[5]) ? node3780 : 1'b1;
												assign node3780 = (inp[14]) ? node3782 : 1'b1;
													assign node3782 = (inp[2]) ? 1'b0 : 1'b1;
											assign node3785 = (inp[5]) ? node3791 : node3786;
												assign node3786 = (inp[7]) ? node3788 : 1'b1;
													assign node3788 = (inp[2]) ? 1'b0 : 1'b1;
												assign node3791 = (inp[14]) ? 1'b0 : node3792;
													assign node3792 = (inp[12]) ? 1'b0 : 1'b1;
										assign node3796 = (inp[12]) ? node3808 : node3797;
											assign node3797 = (inp[10]) ? node3803 : node3798;
												assign node3798 = (inp[5]) ? node3800 : 1'b1;
													assign node3800 = (inp[7]) ? 1'b0 : 1'b1;
												assign node3803 = (inp[5]) ? 1'b0 : node3804;
													assign node3804 = (inp[14]) ? 1'b0 : 1'b1;
											assign node3808 = (inp[14]) ? 1'b0 : node3809;
												assign node3809 = (inp[5]) ? node3811 : 1'b1;
													assign node3811 = (inp[10]) ? 1'b0 : 1'b0;
									assign node3815 = (inp[12]) ? node3835 : node3816;
										assign node3816 = (inp[5]) ? node3828 : node3817;
											assign node3817 = (inp[7]) ? node3823 : node3818;
												assign node3818 = (inp[14]) ? node3820 : 1'b1;
													assign node3820 = (inp[2]) ? 1'b0 : 1'b1;
												assign node3823 = (inp[2]) ? 1'b0 : node3824;
													assign node3824 = (inp[10]) ? 1'b0 : 1'b1;
											assign node3828 = (inp[10]) ? 1'b0 : node3829;
												assign node3829 = (inp[14]) ? 1'b0 : node3830;
													assign node3830 = (inp[2]) ? 1'b0 : 1'b1;
										assign node3835 = (inp[7]) ? 1'b0 : node3836;
											assign node3836 = (inp[6]) ? 1'b0 : node3837;
												assign node3837 = (inp[5]) ? 1'b0 : node3838;
													assign node3838 = (inp[14]) ? 1'b0 : 1'b1;
						assign node3844 = (inp[2]) ? node3976 : node3845;
							assign node3845 = (inp[12]) ? node3911 : node3846;
								assign node3846 = (inp[13]) ? node3876 : node3847;
									assign node3847 = (inp[7]) ? node3857 : node3848;
										assign node3848 = (inp[5]) ? node3850 : 1'b1;
											assign node3850 = (inp[14]) ? node3852 : 1'b1;
												assign node3852 = (inp[10]) ? node3854 : 1'b1;
													assign node3854 = (inp[6]) ? 1'b0 : 1'b1;
										assign node3857 = (inp[8]) ? node3865 : node3858;
											assign node3858 = (inp[14]) ? node3860 : 1'b1;
												assign node3860 = (inp[6]) ? node3862 : 1'b1;
													assign node3862 = (inp[5]) ? 1'b0 : 1'b1;
											assign node3865 = (inp[14]) ? node3871 : node3866;
												assign node3866 = (inp[0]) ? node3868 : 1'b1;
													assign node3868 = (inp[5]) ? 1'b0 : 1'b1;
												assign node3871 = (inp[5]) ? 1'b0 : node3872;
													assign node3872 = (inp[10]) ? 1'b0 : 1'b1;
									assign node3876 = (inp[0]) ? node3892 : node3877;
										assign node3877 = (inp[5]) ? node3885 : node3878;
											assign node3878 = (inp[7]) ? node3880 : 1'b1;
												assign node3880 = (inp[10]) ? node3882 : 1'b1;
													assign node3882 = (inp[6]) ? 1'b0 : 1'b1;
											assign node3885 = (inp[10]) ? 1'b0 : node3886;
												assign node3886 = (inp[14]) ? node3888 : 1'b1;
													assign node3888 = (inp[6]) ? 1'b0 : 1'b1;
										assign node3892 = (inp[6]) ? node3904 : node3893;
											assign node3893 = (inp[7]) ? node3899 : node3894;
												assign node3894 = (inp[10]) ? node3896 : 1'b1;
													assign node3896 = (inp[14]) ? 1'b0 : 1'b1;
												assign node3899 = (inp[8]) ? 1'b0 : node3900;
													assign node3900 = (inp[14]) ? 1'b0 : 1'b1;
											assign node3904 = (inp[5]) ? 1'b0 : node3905;
												assign node3905 = (inp[8]) ? 1'b0 : node3906;
													assign node3906 = (inp[7]) ? 1'b0 : 1'b1;
								assign node3911 = (inp[5]) ? node3947 : node3912;
									assign node3912 = (inp[8]) ? node3928 : node3913;
										assign node3913 = (inp[7]) ? node3921 : node3914;
											assign node3914 = (inp[10]) ? node3916 : 1'b1;
												assign node3916 = (inp[14]) ? node3918 : 1'b1;
													assign node3918 = (inp[6]) ? 1'b0 : 1'b1;
											assign node3921 = (inp[13]) ? 1'b0 : node3922;
												assign node3922 = (inp[6]) ? node3924 : 1'b1;
													assign node3924 = (inp[0]) ? 1'b0 : 1'b1;
										assign node3928 = (inp[13]) ? node3940 : node3929;
											assign node3929 = (inp[14]) ? node3935 : node3930;
												assign node3930 = (inp[7]) ? node3932 : 1'b1;
													assign node3932 = (inp[0]) ? 1'b0 : 1'b1;
												assign node3935 = (inp[0]) ? 1'b0 : node3936;
													assign node3936 = (inp[7]) ? 1'b0 : 1'b1;
											assign node3940 = (inp[0]) ? 1'b0 : node3941;
												assign node3941 = (inp[6]) ? 1'b0 : node3942;
													assign node3942 = (inp[10]) ? 1'b0 : 1'b1;
									assign node3947 = (inp[6]) ? node3967 : node3948;
										assign node3948 = (inp[10]) ? node3960 : node3949;
											assign node3949 = (inp[13]) ? node3955 : node3950;
												assign node3950 = (inp[0]) ? node3952 : 1'b1;
													assign node3952 = (inp[8]) ? 1'b0 : 1'b1;
												assign node3955 = (inp[14]) ? node3957 : 1'b1;
													assign node3957 = (inp[8]) ? 1'b0 : 1'b0;
											assign node3960 = (inp[0]) ? 1'b0 : node3961;
												assign node3961 = (inp[14]) ? 1'b0 : node3962;
													assign node3962 = (inp[7]) ? 1'b0 : 1'b1;
										assign node3967 = (inp[10]) ? 1'b0 : node3968;
											assign node3968 = (inp[14]) ? 1'b0 : node3969;
												assign node3969 = (inp[0]) ? 1'b0 : node3970;
													assign node3970 = (inp[7]) ? 1'b0 : 1'b1;
							assign node3976 = (inp[0]) ? node4042 : node3977;
								assign node3977 = (inp[8]) ? node4013 : node3978;
									assign node3978 = (inp[10]) ? node3994 : node3979;
										assign node3979 = (inp[13]) ? node3987 : node3980;
											assign node3980 = (inp[12]) ? node3982 : 1'b1;
												assign node3982 = (inp[14]) ? node3984 : 1'b1;
													assign node3984 = (inp[5]) ? 1'b0 : 1'b1;
											assign node3987 = (inp[7]) ? 1'b0 : node3988;
												assign node3988 = (inp[14]) ? node3990 : 1'b1;
													assign node3990 = (inp[5]) ? 1'b0 : 1'b1;
										assign node3994 = (inp[6]) ? node4006 : node3995;
											assign node3995 = (inp[5]) ? node4001 : node3996;
												assign node3996 = (inp[7]) ? node3998 : 1'b1;
													assign node3998 = (inp[12]) ? 1'b0 : 1'b1;
												assign node4001 = (inp[14]) ? 1'b0 : node4002;
													assign node4002 = (inp[12]) ? 1'b0 : 1'b1;
											assign node4006 = (inp[12]) ? 1'b0 : node4007;
												assign node4007 = (inp[5]) ? node4009 : 1'b1;
													assign node4009 = (inp[13]) ? 1'b0 : 1'b0;
									assign node4013 = (inp[7]) ? node4033 : node4014;
										assign node4014 = (inp[14]) ? node4026 : node4015;
											assign node4015 = (inp[13]) ? node4021 : node4016;
												assign node4016 = (inp[5]) ? node4018 : 1'b1;
													assign node4018 = (inp[10]) ? 1'b0 : 1'b1;
												assign node4021 = (inp[6]) ? node4023 : 1'b1;
													assign node4023 = (inp[10]) ? 1'b0 : 1'b0;
											assign node4026 = (inp[6]) ? 1'b0 : node4027;
												assign node4027 = (inp[10]) ? node4029 : 1'b1;
													assign node4029 = (inp[12]) ? 1'b0 : 1'b0;
										assign node4033 = (inp[14]) ? 1'b0 : node4034;
											assign node4034 = (inp[6]) ? 1'b0 : node4035;
												assign node4035 = (inp[13]) ? 1'b0 : node4036;
													assign node4036 = (inp[5]) ? 1'b0 : 1'b1;
								assign node4042 = (inp[13]) ? node4070 : node4043;
									assign node4043 = (inp[12]) ? node4063 : node4044;
										assign node4044 = (inp[8]) ? node4056 : node4045;
											assign node4045 = (inp[5]) ? node4051 : node4046;
												assign node4046 = (inp[10]) ? node4048 : 1'b1;
													assign node4048 = (inp[14]) ? 1'b0 : 1'b1;
												assign node4051 = (inp[6]) ? 1'b0 : node4052;
													assign node4052 = (inp[7]) ? 1'b0 : 1'b1;
											assign node4056 = (inp[14]) ? 1'b0 : node4057;
												assign node4057 = (inp[6]) ? 1'b0 : node4058;
													assign node4058 = (inp[7]) ? 1'b0 : 1'b1;
										assign node4063 = (inp[7]) ? 1'b0 : node4064;
											assign node4064 = (inp[14]) ? 1'b0 : node4065;
												assign node4065 = (inp[10]) ? 1'b0 : 1'b1;
									assign node4070 = (inp[10]) ? 1'b0 : node4071;
										assign node4071 = (inp[14]) ? 1'b0 : node4072;
											assign node4072 = (inp[5]) ? 1'b0 : node4073;
												assign node4073 = (inp[12]) ? 1'b0 : node4074;
													assign node4074 = (inp[6]) ? 1'b0 : 1'b0;
				assign node4081 = (inp[13]) ? node4539 : node4082;
					assign node4082 = (inp[0]) ? node4296 : node4083;
						assign node4083 = (inp[9]) ? node4181 : node4084;
							assign node4084 = (inp[5]) ? node4118 : node4085;
								assign node4085 = (inp[12]) ? node4097 : node4086;
									assign node4086 = (inp[4]) ? node4088 : 1'b1;
										assign node4088 = (inp[14]) ? node4090 : 1'b1;
											assign node4090 = (inp[10]) ? node4092 : 1'b1;
												assign node4092 = (inp[2]) ? node4094 : 1'b1;
													assign node4094 = (inp[6]) ? 1'b0 : 1'b0;
									assign node4097 = (inp[6]) ? node4105 : node4098;
										assign node4098 = (inp[7]) ? node4100 : 1'b1;
											assign node4100 = (inp[4]) ? node4102 : 1'b1;
												assign node4102 = (inp[14]) ? 1'b0 : 1'b1;
										assign node4105 = (inp[2]) ? node4113 : node4106;
											assign node4106 = (inp[8]) ? node4108 : 1'b1;
												assign node4108 = (inp[4]) ? node4110 : 1'b1;
													assign node4110 = (inp[7]) ? 1'b0 : 1'b0;
											assign node4113 = (inp[8]) ? 1'b0 : node4114;
												assign node4114 = (inp[4]) ? 1'b0 : 1'b1;
								assign node4118 = (inp[4]) ? node4148 : node4119;
									assign node4119 = (inp[7]) ? node4129 : node4120;
										assign node4120 = (inp[14]) ? node4122 : 1'b1;
											assign node4122 = (inp[12]) ? node4124 : 1'b1;
												assign node4124 = (inp[6]) ? node4126 : 1'b1;
													assign node4126 = (inp[8]) ? 1'b0 : 1'b1;
										assign node4129 = (inp[2]) ? node4137 : node4130;
											assign node4130 = (inp[12]) ? node4132 : 1'b1;
												assign node4132 = (inp[10]) ? node4134 : 1'b1;
													assign node4134 = (inp[14]) ? 1'b0 : 1'b1;
											assign node4137 = (inp[6]) ? node4143 : node4138;
												assign node4138 = (inp[10]) ? node4140 : 1'b1;
													assign node4140 = (inp[8]) ? 1'b0 : 1'b1;
												assign node4143 = (inp[8]) ? 1'b0 : node4144;
													assign node4144 = (inp[10]) ? 1'b0 : 1'b1;
									assign node4148 = (inp[14]) ? node4162 : node4149;
										assign node4149 = (inp[8]) ? node4151 : 1'b1;
											assign node4151 = (inp[12]) ? node4157 : node4152;
												assign node4152 = (inp[7]) ? node4154 : 1'b1;
													assign node4154 = (inp[10]) ? 1'b0 : 1'b1;
												assign node4157 = (inp[10]) ? 1'b0 : node4158;
													assign node4158 = (inp[7]) ? 1'b0 : 1'b1;
										assign node4162 = (inp[2]) ? node4174 : node4163;
											assign node4163 = (inp[6]) ? node4169 : node4164;
												assign node4164 = (inp[12]) ? node4166 : 1'b1;
													assign node4166 = (inp[7]) ? 1'b0 : 1'b1;
												assign node4169 = (inp[10]) ? 1'b0 : node4170;
													assign node4170 = (inp[7]) ? 1'b0 : 1'b1;
											assign node4174 = (inp[12]) ? 1'b0 : node4175;
												assign node4175 = (inp[10]) ? 1'b0 : node4176;
													assign node4176 = (inp[8]) ? 1'b0 : 1'b1;
							assign node4181 = (inp[7]) ? node4239 : node4182;
								assign node4182 = (inp[2]) ? node4208 : node4183;
									assign node4183 = (inp[12]) ? node4193 : node4184;
										assign node4184 = (inp[10]) ? node4186 : 1'b1;
											assign node4186 = (inp[5]) ? node4188 : 1'b1;
												assign node4188 = (inp[6]) ? node4190 : 1'b1;
													assign node4190 = (inp[8]) ? 1'b0 : 1'b1;
										assign node4193 = (inp[4]) ? node4201 : node4194;
											assign node4194 = (inp[10]) ? node4196 : 1'b1;
												assign node4196 = (inp[8]) ? node4198 : 1'b1;
													assign node4198 = (inp[6]) ? 1'b0 : 1'b1;
											assign node4201 = (inp[6]) ? 1'b0 : node4202;
												assign node4202 = (inp[14]) ? node4204 : 1'b1;
													assign node4204 = (inp[5]) ? 1'b0 : 1'b0;
									assign node4208 = (inp[8]) ? node4226 : node4209;
										assign node4209 = (inp[5]) ? node4215 : node4210;
											assign node4210 = (inp[6]) ? node4212 : 1'b1;
												assign node4212 = (inp[14]) ? 1'b1 : 1'b0;
											assign node4215 = (inp[4]) ? node4221 : node4216;
												assign node4216 = (inp[10]) ? node4218 : 1'b1;
													assign node4218 = (inp[12]) ? 1'b0 : 1'b1;
												assign node4221 = (inp[6]) ? 1'b0 : node4222;
													assign node4222 = (inp[12]) ? 1'b0 : 1'b1;
										assign node4226 = (inp[5]) ? 1'b0 : node4227;
											assign node4227 = (inp[4]) ? node4233 : node4228;
												assign node4228 = (inp[12]) ? node4230 : 1'b1;
													assign node4230 = (inp[14]) ? 1'b0 : 1'b1;
												assign node4233 = (inp[14]) ? 1'b0 : node4234;
													assign node4234 = (inp[6]) ? 1'b0 : 1'b1;
								assign node4239 = (inp[6]) ? node4267 : node4240;
									assign node4240 = (inp[12]) ? node4254 : node4241;
										assign node4241 = (inp[4]) ? node4243 : 1'b1;
											assign node4243 = (inp[10]) ? node4249 : node4244;
												assign node4244 = (inp[5]) ? node4246 : 1'b1;
													assign node4246 = (inp[8]) ? 1'b0 : 1'b1;
												assign node4249 = (inp[14]) ? 1'b0 : node4250;
													assign node4250 = (inp[8]) ? 1'b0 : 1'b1;
										assign node4254 = (inp[4]) ? 1'b0 : node4255;
											assign node4255 = (inp[2]) ? node4261 : node4256;
												assign node4256 = (inp[10]) ? node4258 : 1'b1;
													assign node4258 = (inp[5]) ? 1'b0 : 1'b1;
												assign node4261 = (inp[5]) ? 1'b0 : node4262;
													assign node4262 = (inp[8]) ? 1'b0 : 1'b1;
									assign node4267 = (inp[14]) ? node4287 : node4268;
										assign node4268 = (inp[8]) ? node4280 : node4269;
											assign node4269 = (inp[12]) ? node4275 : node4270;
												assign node4270 = (inp[4]) ? node4272 : 1'b1;
													assign node4272 = (inp[2]) ? 1'b0 : 1'b1;
												assign node4275 = (inp[2]) ? 1'b0 : node4276;
													assign node4276 = (inp[10]) ? 1'b0 : 1'b1;
											assign node4280 = (inp[10]) ? 1'b0 : node4281;
												assign node4281 = (inp[5]) ? 1'b0 : node4282;
													assign node4282 = (inp[4]) ? 1'b0 : 1'b1;
										assign node4287 = (inp[5]) ? 1'b0 : node4288;
											assign node4288 = (inp[12]) ? 1'b0 : node4289;
												assign node4289 = (inp[8]) ? 1'b0 : node4290;
													assign node4290 = (inp[10]) ? 1'b0 : 1'b1;
						assign node4296 = (inp[2]) ? node4428 : node4297;
							assign node4297 = (inp[14]) ? node4357 : node4298;
								assign node4298 = (inp[6]) ? node4324 : node4299;
									assign node4299 = (inp[4]) ? node4307 : node4300;
										assign node4300 = (inp[5]) ? node4302 : 1'b1;
											assign node4302 = (inp[10]) ? node4304 : 1'b1;
												assign node4304 = (inp[9]) ? 1'b0 : 1'b1;
										assign node4307 = (inp[12]) ? node4315 : node4308;
											assign node4308 = (inp[7]) ? node4310 : 1'b1;
												assign node4310 = (inp[5]) ? node4312 : 1'b1;
													assign node4312 = (inp[8]) ? 1'b0 : 1'b1;
											assign node4315 = (inp[10]) ? node4319 : node4316;
												assign node4316 = (inp[8]) ? 1'b0 : 1'b1;
												assign node4319 = (inp[9]) ? 1'b0 : node4320;
													assign node4320 = (inp[7]) ? 1'b0 : 1'b1;
									assign node4324 = (inp[5]) ? node4344 : node4325;
										assign node4325 = (inp[9]) ? node4333 : node4326;
											assign node4326 = (inp[4]) ? node4328 : 1'b1;
												assign node4328 = (inp[7]) ? node4330 : 1'b1;
													assign node4330 = (inp[8]) ? 1'b0 : 1'b1;
											assign node4333 = (inp[10]) ? node4339 : node4334;
												assign node4334 = (inp[4]) ? node4336 : 1'b1;
													assign node4336 = (inp[12]) ? 1'b0 : 1'b1;
												assign node4339 = (inp[12]) ? 1'b0 : node4340;
													assign node4340 = (inp[4]) ? 1'b1 : 1'b0;
										assign node4344 = (inp[12]) ? 1'b0 : node4345;
											assign node4345 = (inp[7]) ? node4351 : node4346;
												assign node4346 = (inp[10]) ? node4348 : 1'b1;
													assign node4348 = (inp[8]) ? 1'b0 : 1'b1;
												assign node4351 = (inp[8]) ? 1'b0 : node4352;
													assign node4352 = (inp[10]) ? 1'b0 : 1'b1;
								assign node4357 = (inp[12]) ? node4397 : node4358;
									assign node4358 = (inp[10]) ? node4378 : node4359;
										assign node4359 = (inp[8]) ? node4367 : node4360;
											assign node4360 = (inp[4]) ? node4362 : 1'b1;
												assign node4362 = (inp[9]) ? node4364 : 1'b1;
													assign node4364 = (inp[7]) ? 1'b0 : 1'b1;
											assign node4367 = (inp[7]) ? node4373 : node4368;
												assign node4368 = (inp[9]) ? node4370 : 1'b1;
													assign node4370 = (inp[4]) ? 1'b0 : 1'b1;
												assign node4373 = (inp[5]) ? 1'b0 : node4374;
													assign node4374 = (inp[9]) ? 1'b0 : 1'b1;
										assign node4378 = (inp[8]) ? node4390 : node4379;
											assign node4379 = (inp[7]) ? node4385 : node4380;
												assign node4380 = (inp[9]) ? node4382 : 1'b1;
													assign node4382 = (inp[4]) ? 1'b0 : 1'b1;
												assign node4385 = (inp[5]) ? 1'b0 : node4386;
													assign node4386 = (inp[6]) ? 1'b0 : 1'b1;
											assign node4390 = (inp[9]) ? 1'b0 : node4391;
												assign node4391 = (inp[4]) ? 1'b0 : node4392;
													assign node4392 = (inp[5]) ? 1'b0 : 1'b1;
									assign node4397 = (inp[6]) ? node4419 : node4398;
										assign node4398 = (inp[10]) ? node4412 : node4399;
											assign node4399 = (inp[5]) ? node4405 : node4400;
												assign node4400 = (inp[8]) ? node4402 : 1'b1;
													assign node4402 = (inp[4]) ? 1'b0 : 1'b1;
												assign node4405 = (inp[8]) ? node4409 : node4406;
													assign node4406 = (inp[7]) ? 1'b0 : 1'b1;
													assign node4409 = (inp[9]) ? 1'b0 : 1'b0;
											assign node4412 = (inp[4]) ? 1'b0 : node4413;
												assign node4413 = (inp[7]) ? 1'b0 : node4414;
													assign node4414 = (inp[5]) ? 1'b0 : 1'b1;
										assign node4419 = (inp[4]) ? 1'b0 : node4420;
											assign node4420 = (inp[10]) ? 1'b0 : node4421;
												assign node4421 = (inp[8]) ? 1'b0 : node4422;
													assign node4422 = (inp[9]) ? 1'b0 : 1'b1;
							assign node4428 = (inp[14]) ? node4498 : node4429;
								assign node4429 = (inp[10]) ? node4469 : node4430;
									assign node4430 = (inp[6]) ? node4450 : node4431;
										assign node4431 = (inp[4]) ? node4439 : node4432;
											assign node4432 = (inp[5]) ? node4434 : 1'b1;
												assign node4434 = (inp[9]) ? node4436 : 1'b1;
													assign node4436 = (inp[8]) ? 1'b0 : 1'b1;
											assign node4439 = (inp[9]) ? node4445 : node4440;
												assign node4440 = (inp[5]) ? node4442 : 1'b1;
													assign node4442 = (inp[8]) ? 1'b0 : 1'b1;
												assign node4445 = (inp[12]) ? 1'b0 : node4446;
													assign node4446 = (inp[8]) ? 1'b0 : 1'b1;
										assign node4450 = (inp[5]) ? node4462 : node4451;
											assign node4451 = (inp[7]) ? node4457 : node4452;
												assign node4452 = (inp[9]) ? node4454 : 1'b1;
													assign node4454 = (inp[8]) ? 1'b0 : 1'b1;
												assign node4457 = (inp[4]) ? 1'b0 : node4458;
													assign node4458 = (inp[12]) ? 1'b0 : 1'b1;
											assign node4462 = (inp[9]) ? 1'b0 : node4463;
												assign node4463 = (inp[8]) ? 1'b0 : node4464;
													assign node4464 = (inp[12]) ? 1'b0 : 1'b1;
									assign node4469 = (inp[8]) ? node4489 : node4470;
										assign node4470 = (inp[9]) ? node4482 : node4471;
											assign node4471 = (inp[4]) ? node4477 : node4472;
												assign node4472 = (inp[6]) ? node4474 : 1'b1;
													assign node4474 = (inp[12]) ? 1'b0 : 1'b1;
												assign node4477 = (inp[5]) ? 1'b0 : node4478;
													assign node4478 = (inp[7]) ? 1'b0 : 1'b1;
											assign node4482 = (inp[5]) ? 1'b0 : node4483;
												assign node4483 = (inp[12]) ? 1'b0 : node4484;
													assign node4484 = (inp[4]) ? 1'b0 : 1'b1;
										assign node4489 = (inp[7]) ? 1'b0 : node4490;
											assign node4490 = (inp[6]) ? 1'b0 : node4491;
												assign node4491 = (inp[12]) ? 1'b0 : node4492;
													assign node4492 = (inp[9]) ? 1'b0 : 1'b0;
								assign node4498 = (inp[9]) ? node4528 : node4499;
									assign node4499 = (inp[8]) ? node4519 : node4500;
										assign node4500 = (inp[5]) ? node4512 : node4501;
											assign node4501 = (inp[7]) ? node4507 : node4502;
												assign node4502 = (inp[6]) ? node4504 : 1'b1;
													assign node4504 = (inp[4]) ? 1'b0 : 1'b1;
												assign node4507 = (inp[10]) ? 1'b0 : node4508;
													assign node4508 = (inp[4]) ? 1'b0 : 1'b1;
											assign node4512 = (inp[10]) ? 1'b0 : node4513;
												assign node4513 = (inp[4]) ? 1'b0 : node4514;
													assign node4514 = (inp[6]) ? 1'b0 : 1'b1;
										assign node4519 = (inp[12]) ? 1'b0 : node4520;
											assign node4520 = (inp[6]) ? 1'b0 : node4521;
												assign node4521 = (inp[7]) ? 1'b0 : node4522;
													assign node4522 = (inp[4]) ? 1'b0 : 1'b1;
									assign node4528 = (inp[6]) ? 1'b0 : node4529;
										assign node4529 = (inp[12]) ? 1'b0 : node4530;
											assign node4530 = (inp[5]) ? 1'b0 : node4531;
												assign node4531 = (inp[4]) ? 1'b0 : node4532;
													assign node4532 = (inp[7]) ? 1'b0 : 1'b1;
					assign node4539 = (inp[14]) ? node4785 : node4540;
						assign node4540 = (inp[5]) ? node4678 : node4541;
							assign node4541 = (inp[7]) ? node4611 : node4542;
								assign node4542 = (inp[9]) ? node4572 : node4543;
									assign node4543 = (inp[4]) ? node4553 : node4544;
										assign node4544 = (inp[8]) ? node4546 : 1'b1;
											assign node4546 = (inp[12]) ? node4548 : 1'b1;
												assign node4548 = (inp[6]) ? node4550 : 1'b1;
													assign node4550 = (inp[2]) ? 1'b0 : 1'b1;
										assign node4553 = (inp[0]) ? node4561 : node4554;
											assign node4554 = (inp[10]) ? node4556 : 1'b1;
												assign node4556 = (inp[2]) ? node4558 : 1'b1;
													assign node4558 = (inp[12]) ? 1'b0 : 1'b1;
											assign node4561 = (inp[12]) ? node4567 : node4562;
												assign node4562 = (inp[10]) ? node4564 : 1'b1;
													assign node4564 = (inp[6]) ? 1'b0 : 1'b1;
												assign node4567 = (inp[6]) ? 1'b0 : node4568;
													assign node4568 = (inp[10]) ? 1'b0 : 1'b1;
									assign node4572 = (inp[8]) ? node4592 : node4573;
										assign node4573 = (inp[6]) ? node4581 : node4574;
											assign node4574 = (inp[4]) ? node4576 : 1'b1;
												assign node4576 = (inp[2]) ? node4578 : 1'b1;
													assign node4578 = (inp[10]) ? 1'b0 : 1'b1;
											assign node4581 = (inp[12]) ? node4587 : node4582;
												assign node4582 = (inp[0]) ? node4584 : 1'b1;
													assign node4584 = (inp[2]) ? 1'b0 : 1'b1;
												assign node4587 = (inp[0]) ? 1'b0 : node4588;
													assign node4588 = (inp[2]) ? 1'b0 : 1'b1;
										assign node4592 = (inp[12]) ? node4604 : node4593;
											assign node4593 = (inp[0]) ? node4601 : node4594;
												assign node4594 = (inp[10]) ? node4598 : node4595;
													assign node4595 = (inp[2]) ? 1'b1 : 1'b1;
													assign node4598 = (inp[2]) ? 1'b0 : 1'b1;
												assign node4601 = (inp[6]) ? 1'b0 : 1'b1;
											assign node4604 = (inp[2]) ? 1'b0 : node4605;
												assign node4605 = (inp[0]) ? 1'b0 : node4606;
													assign node4606 = (inp[10]) ? 1'b0 : 1'b1;
								assign node4611 = (inp[2]) ? node4649 : node4612;
									assign node4612 = (inp[9]) ? node4632 : node4613;
										assign node4613 = (inp[12]) ? node4621 : node4614;
											assign node4614 = (inp[10]) ? node4616 : 1'b1;
												assign node4616 = (inp[8]) ? node4618 : 1'b1;
													assign node4618 = (inp[4]) ? 1'b0 : 1'b1;
											assign node4621 = (inp[4]) ? node4627 : node4622;
												assign node4622 = (inp[0]) ? node4624 : 1'b1;
													assign node4624 = (inp[8]) ? 1'b0 : 1'b1;
												assign node4627 = (inp[8]) ? 1'b0 : node4628;
													assign node4628 = (inp[10]) ? 1'b0 : 1'b1;
										assign node4632 = (inp[10]) ? node4642 : node4633;
											assign node4633 = (inp[0]) ? node4639 : node4634;
												assign node4634 = (inp[4]) ? node4636 : 1'b1;
													assign node4636 = (inp[8]) ? 1'b0 : 1'b1;
												assign node4639 = (inp[6]) ? 1'b0 : 1'b1;
											assign node4642 = (inp[12]) ? 1'b0 : node4643;
												assign node4643 = (inp[8]) ? 1'b0 : node4644;
													assign node4644 = (inp[6]) ? 1'b0 : 1'b1;
									assign node4649 = (inp[10]) ? node4669 : node4650;
										assign node4650 = (inp[6]) ? node4662 : node4651;
											assign node4651 = (inp[4]) ? node4657 : node4652;
												assign node4652 = (inp[9]) ? node4654 : 1'b1;
													assign node4654 = (inp[8]) ? 1'b0 : 1'b1;
												assign node4657 = (inp[0]) ? 1'b0 : node4658;
													assign node4658 = (inp[8]) ? 1'b0 : 1'b1;
											assign node4662 = (inp[8]) ? 1'b0 : node4663;
												assign node4663 = (inp[12]) ? 1'b0 : node4664;
													assign node4664 = (inp[0]) ? 1'b0 : 1'b1;
										assign node4669 = (inp[4]) ? 1'b0 : node4670;
											assign node4670 = (inp[0]) ? 1'b0 : node4671;
												assign node4671 = (inp[9]) ? 1'b0 : node4672;
													assign node4672 = (inp[8]) ? 1'b0 : 1'b1;
							assign node4678 = (inp[10]) ? node4746 : node4679;
								assign node4679 = (inp[9]) ? node4717 : node4680;
									assign node4680 = (inp[8]) ? node4700 : node4681;
										assign node4681 = (inp[12]) ? node4689 : node4682;
											assign node4682 = (inp[6]) ? node4684 : 1'b1;
												assign node4684 = (inp[7]) ? node4686 : 1'b1;
													assign node4686 = (inp[2]) ? 1'b0 : 1'b1;
											assign node4689 = (inp[7]) ? node4695 : node4690;
												assign node4690 = (inp[0]) ? node4692 : 1'b1;
													assign node4692 = (inp[6]) ? 1'b0 : 1'b1;
												assign node4695 = (inp[6]) ? 1'b0 : node4696;
													assign node4696 = (inp[2]) ? 1'b0 : 1'b1;
										assign node4700 = (inp[7]) ? node4710 : node4701;
											assign node4701 = (inp[0]) ? node4705 : node4702;
												assign node4702 = (inp[6]) ? 1'b0 : 1'b1;
												assign node4705 = (inp[4]) ? 1'b0 : node4706;
													assign node4706 = (inp[2]) ? 1'b0 : 1'b1;
											assign node4710 = (inp[2]) ? 1'b0 : node4711;
												assign node4711 = (inp[4]) ? 1'b0 : node4712;
													assign node4712 = (inp[12]) ? 1'b0 : 1'b1;
									assign node4717 = (inp[2]) ? node4737 : node4718;
										assign node4718 = (inp[0]) ? node4730 : node4719;
											assign node4719 = (inp[4]) ? node4725 : node4720;
												assign node4720 = (inp[8]) ? node4722 : 1'b1;
													assign node4722 = (inp[7]) ? 1'b0 : 1'b1;
												assign node4725 = (inp[7]) ? 1'b0 : node4726;
													assign node4726 = (inp[6]) ? 1'b0 : 1'b1;
											assign node4730 = (inp[7]) ? 1'b0 : node4731;
												assign node4731 = (inp[6]) ? 1'b0 : node4732;
													assign node4732 = (inp[8]) ? 1'b0 : 1'b1;
										assign node4737 = (inp[6]) ? 1'b0 : node4738;
											assign node4738 = (inp[8]) ? 1'b0 : node4739;
												assign node4739 = (inp[7]) ? 1'b0 : node4740;
													assign node4740 = (inp[4]) ? 1'b0 : 1'b1;
								assign node4746 = (inp[12]) ? node4774 : node4747;
									assign node4747 = (inp[9]) ? node4765 : node4748;
										assign node4748 = (inp[0]) ? node4760 : node4749;
											assign node4749 = (inp[8]) ? node4755 : node4750;
												assign node4750 = (inp[6]) ? node4752 : 1'b1;
													assign node4752 = (inp[4]) ? 1'b1 : 1'b0;
												assign node4755 = (inp[4]) ? 1'b0 : node4756;
													assign node4756 = (inp[7]) ? 1'b0 : 1'b1;
											assign node4760 = (inp[2]) ? 1'b0 : node4761;
												assign node4761 = (inp[8]) ? 1'b0 : 1'b1;
										assign node4765 = (inp[6]) ? 1'b0 : node4766;
											assign node4766 = (inp[8]) ? 1'b0 : node4767;
												assign node4767 = (inp[7]) ? 1'b0 : node4768;
													assign node4768 = (inp[0]) ? 1'b0 : 1'b1;
									assign node4774 = (inp[4]) ? 1'b0 : node4775;
										assign node4775 = (inp[0]) ? 1'b0 : node4776;
											assign node4776 = (inp[8]) ? 1'b0 : node4777;
												assign node4777 = (inp[2]) ? 1'b0 : node4778;
													assign node4778 = (inp[7]) ? 1'b0 : 1'b1;
						assign node4785 = (inp[10]) ? node4883 : node4786;
							assign node4786 = (inp[7]) ? node4856 : node4787;
								assign node4787 = (inp[6]) ? node4827 : node4788;
									assign node4788 = (inp[0]) ? node4808 : node4789;
										assign node4789 = (inp[8]) ? node4797 : node4790;
											assign node4790 = (inp[2]) ? node4792 : 1'b1;
												assign node4792 = (inp[4]) ? node4794 : 1'b1;
													assign node4794 = (inp[12]) ? 1'b0 : 1'b1;
											assign node4797 = (inp[4]) ? node4803 : node4798;
												assign node4798 = (inp[9]) ? node4800 : 1'b1;
													assign node4800 = (inp[2]) ? 1'b0 : 1'b1;
												assign node4803 = (inp[5]) ? 1'b0 : node4804;
													assign node4804 = (inp[2]) ? 1'b0 : 1'b1;
										assign node4808 = (inp[2]) ? node4820 : node4809;
											assign node4809 = (inp[5]) ? node4815 : node4810;
												assign node4810 = (inp[9]) ? node4812 : 1'b1;
													assign node4812 = (inp[12]) ? 1'b1 : 1'b0;
												assign node4815 = (inp[4]) ? 1'b0 : node4816;
													assign node4816 = (inp[12]) ? 1'b0 : 1'b1;
											assign node4820 = (inp[4]) ? 1'b0 : node4821;
												assign node4821 = (inp[9]) ? 1'b0 : node4822;
													assign node4822 = (inp[5]) ? 1'b1 : 1'b0;
									assign node4827 = (inp[5]) ? node4847 : node4828;
										assign node4828 = (inp[12]) ? node4840 : node4829;
											assign node4829 = (inp[9]) ? node4835 : node4830;
												assign node4830 = (inp[2]) ? node4832 : 1'b1;
													assign node4832 = (inp[4]) ? 1'b0 : 1'b1;
												assign node4835 = (inp[4]) ? 1'b0 : node4836;
													assign node4836 = (inp[0]) ? 1'b0 : 1'b1;
											assign node4840 = (inp[4]) ? 1'b0 : node4841;
												assign node4841 = (inp[8]) ? 1'b0 : node4842;
													assign node4842 = (inp[2]) ? 1'b0 : 1'b1;
										assign node4847 = (inp[8]) ? 1'b0 : node4848;
											assign node4848 = (inp[4]) ? 1'b0 : node4849;
												assign node4849 = (inp[0]) ? 1'b0 : node4850;
													assign node4850 = (inp[12]) ? 1'b0 : 1'b1;
								assign node4856 = (inp[12]) ? 1'b0 : node4857;
									assign node4857 = (inp[5]) ? node4873 : node4858;
										assign node4858 = (inp[9]) ? node4866 : node4859;
											assign node4859 = (inp[6]) ? node4861 : 1'b1;
												assign node4861 = (inp[2]) ? 1'b0 : node4862;
													assign node4862 = (inp[4]) ? 1'b0 : 1'b1;
											assign node4866 = (inp[0]) ? 1'b0 : node4867;
												assign node4867 = (inp[8]) ? node4869 : 1'b1;
													assign node4869 = (inp[4]) ? 1'b0 : 1'b0;
										assign node4873 = (inp[6]) ? 1'b0 : node4874;
											assign node4874 = (inp[0]) ? 1'b0 : node4875;
												assign node4875 = (inp[2]) ? 1'b0 : node4876;
													assign node4876 = (inp[4]) ? 1'b0 : 1'b1;
							assign node4883 = (inp[0]) ? node4921 : node4884;
								assign node4884 = (inp[4]) ? node4912 : node4885;
									assign node4885 = (inp[6]) ? node4905 : node4886;
										assign node4886 = (inp[8]) ? node4898 : node4887;
											assign node4887 = (inp[9]) ? node4893 : node4888;
												assign node4888 = (inp[5]) ? node4890 : 1'b1;
													assign node4890 = (inp[7]) ? 1'b0 : 1'b1;
												assign node4893 = (inp[7]) ? 1'b0 : node4894;
													assign node4894 = (inp[12]) ? 1'b0 : 1'b1;
											assign node4898 = (inp[7]) ? 1'b0 : node4899;
												assign node4899 = (inp[2]) ? 1'b0 : node4900;
													assign node4900 = (inp[9]) ? 1'b0 : 1'b1;
										assign node4905 = (inp[7]) ? 1'b0 : node4906;
											assign node4906 = (inp[5]) ? 1'b0 : node4907;
												assign node4907 = (inp[2]) ? 1'b0 : 1'b1;
									assign node4912 = (inp[12]) ? 1'b0 : node4913;
										assign node4913 = (inp[8]) ? 1'b0 : node4914;
											assign node4914 = (inp[5]) ? 1'b0 : node4915;
												assign node4915 = (inp[7]) ? 1'b0 : 1'b1;
								assign node4921 = (inp[8]) ? 1'b0 : node4922;
									assign node4922 = (inp[9]) ? 1'b0 : node4923;
										assign node4923 = (inp[5]) ? 1'b0 : node4924;
											assign node4924 = (inp[2]) ? 1'b0 : node4925;
												assign node4925 = (inp[4]) ? 1'b0 : node4926;
													assign node4926 = (inp[6]) ? 1'b0 : 1'b1;
			assign node4934 = (inp[8]) ? node5796 : node4935;
				assign node4935 = (inp[6]) ? node5409 : node4936;
					assign node4936 = (inp[2]) ? node5180 : node4937;
						assign node4937 = (inp[5]) ? node5049 : node4938;
							assign node4938 = (inp[13]) ? node4980 : node4939;
								assign node4939 = (inp[4]) ? node4951 : node4940;
									assign node4940 = (inp[12]) ? node4942 : 1'b1;
										assign node4942 = (inp[14]) ? node4944 : 1'b1;
											assign node4944 = (inp[11]) ? node4946 : 1'b1;
												assign node4946 = (inp[9]) ? node4948 : 1'b1;
													assign node4948 = (inp[7]) ? 1'b0 : 1'b1;
									assign node4951 = (inp[10]) ? node4961 : node4952;
										assign node4952 = (inp[0]) ? node4954 : 1'b1;
											assign node4954 = (inp[9]) ? node4956 : 1'b1;
												assign node4956 = (inp[14]) ? node4958 : 1'b1;
													assign node4958 = (inp[11]) ? 1'b0 : 1'b1;
										assign node4961 = (inp[11]) ? node4969 : node4962;
											assign node4962 = (inp[9]) ? node4964 : 1'b1;
												assign node4964 = (inp[0]) ? node4966 : 1'b1;
													assign node4966 = (inp[7]) ? 1'b0 : 1'b1;
											assign node4969 = (inp[0]) ? node4975 : node4970;
												assign node4970 = (inp[14]) ? node4972 : 1'b1;
													assign node4972 = (inp[9]) ? 1'b0 : 1'b1;
												assign node4975 = (inp[12]) ? 1'b0 : node4976;
													assign node4976 = (inp[14]) ? 1'b0 : 1'b1;
								assign node4980 = (inp[10]) ? node5010 : node4981;
									assign node4981 = (inp[9]) ? node4991 : node4982;
										assign node4982 = (inp[12]) ? node4984 : 1'b1;
											assign node4984 = (inp[11]) ? node4986 : 1'b1;
												assign node4986 = (inp[4]) ? node4988 : 1'b1;
													assign node4988 = (inp[14]) ? 1'b0 : 1'b1;
										assign node4991 = (inp[0]) ? node4999 : node4992;
											assign node4992 = (inp[4]) ? node4994 : 1'b1;
												assign node4994 = (inp[11]) ? node4996 : 1'b1;
													assign node4996 = (inp[14]) ? 1'b1 : 1'b0;
											assign node4999 = (inp[12]) ? node5005 : node5000;
												assign node5000 = (inp[7]) ? 1'b0 : node5001;
													assign node5001 = (inp[11]) ? 1'b1 : 1'b1;
												assign node5005 = (inp[14]) ? 1'b0 : node5006;
													assign node5006 = (inp[7]) ? 1'b1 : 1'b0;
									assign node5010 = (inp[11]) ? node5030 : node5011;
										assign node5011 = (inp[4]) ? node5019 : node5012;
											assign node5012 = (inp[0]) ? node5014 : 1'b1;
												assign node5014 = (inp[7]) ? node5016 : 1'b1;
													assign node5016 = (inp[9]) ? 1'b0 : 1'b1;
											assign node5019 = (inp[9]) ? node5025 : node5020;
												assign node5020 = (inp[14]) ? node5022 : 1'b1;
													assign node5022 = (inp[0]) ? 1'b0 : 1'b1;
												assign node5025 = (inp[14]) ? 1'b0 : node5026;
													assign node5026 = (inp[0]) ? 1'b0 : 1'b1;
										assign node5030 = (inp[14]) ? node5042 : node5031;
											assign node5031 = (inp[9]) ? node5037 : node5032;
												assign node5032 = (inp[4]) ? node5034 : 1'b1;
													assign node5034 = (inp[7]) ? 1'b0 : 1'b1;
												assign node5037 = (inp[12]) ? 1'b0 : node5038;
													assign node5038 = (inp[0]) ? 1'b0 : 1'b1;
											assign node5042 = (inp[7]) ? 1'b0 : node5043;
												assign node5043 = (inp[0]) ? 1'b0 : node5044;
													assign node5044 = (inp[9]) ? 1'b0 : 1'b1;
							assign node5049 = (inp[4]) ? node5115 : node5050;
								assign node5050 = (inp[11]) ? node5080 : node5051;
									assign node5051 = (inp[14]) ? node5061 : node5052;
										assign node5052 = (inp[10]) ? node5054 : 1'b1;
											assign node5054 = (inp[0]) ? node5056 : 1'b1;
												assign node5056 = (inp[12]) ? node5058 : 1'b1;
													assign node5058 = (inp[13]) ? 1'b0 : 1'b1;
										assign node5061 = (inp[12]) ? node5069 : node5062;
											assign node5062 = (inp[0]) ? node5064 : 1'b1;
												assign node5064 = (inp[13]) ? node5066 : 1'b1;
													assign node5066 = (inp[7]) ? 1'b0 : 1'b1;
											assign node5069 = (inp[10]) ? node5075 : node5070;
												assign node5070 = (inp[9]) ? node5072 : 1'b1;
													assign node5072 = (inp[7]) ? 1'b0 : 1'b1;
												assign node5075 = (inp[0]) ? 1'b0 : node5076;
													assign node5076 = (inp[9]) ? 1'b0 : 1'b1;
									assign node5080 = (inp[7]) ? node5096 : node5081;
										assign node5081 = (inp[13]) ? node5089 : node5082;
											assign node5082 = (inp[10]) ? node5084 : 1'b1;
												assign node5084 = (inp[14]) ? node5086 : 1'b1;
													assign node5086 = (inp[9]) ? 1'b0 : 1'b1;
											assign node5089 = (inp[9]) ? 1'b0 : node5090;
												assign node5090 = (inp[10]) ? node5092 : 1'b1;
													assign node5092 = (inp[0]) ? 1'b0 : 1'b1;
										assign node5096 = (inp[12]) ? node5108 : node5097;
											assign node5097 = (inp[13]) ? node5103 : node5098;
												assign node5098 = (inp[9]) ? node5100 : 1'b1;
													assign node5100 = (inp[10]) ? 1'b0 : 1'b1;
												assign node5103 = (inp[0]) ? 1'b0 : node5104;
													assign node5104 = (inp[10]) ? 1'b0 : 1'b1;
											assign node5108 = (inp[13]) ? 1'b0 : node5109;
												assign node5109 = (inp[10]) ? 1'b0 : node5110;
													assign node5110 = (inp[9]) ? 1'b0 : 1'b1;
								assign node5115 = (inp[10]) ? node5151 : node5116;
									assign node5116 = (inp[11]) ? node5134 : node5117;
										assign node5117 = (inp[12]) ? node5125 : node5118;
											assign node5118 = (inp[0]) ? node5120 : 1'b1;
												assign node5120 = (inp[14]) ? node5122 : 1'b1;
													assign node5122 = (inp[9]) ? 1'b0 : 1'b1;
											assign node5125 = (inp[14]) ? 1'b0 : node5126;
												assign node5126 = (inp[7]) ? node5130 : node5127;
													assign node5127 = (inp[13]) ? 1'b1 : 1'b1;
													assign node5130 = (inp[9]) ? 1'b0 : 1'b1;
										assign node5134 = (inp[0]) ? node5144 : node5135;
											assign node5135 = (inp[14]) ? node5141 : node5136;
												assign node5136 = (inp[12]) ? node5138 : 1'b1;
													assign node5138 = (inp[7]) ? 1'b0 : 1'b1;
												assign node5141 = (inp[9]) ? 1'b0 : 1'b1;
											assign node5144 = (inp[13]) ? 1'b0 : node5145;
												assign node5145 = (inp[7]) ? 1'b0 : node5146;
													assign node5146 = (inp[12]) ? 1'b0 : 1'b1;
									assign node5151 = (inp[13]) ? node5171 : node5152;
										assign node5152 = (inp[12]) ? node5164 : node5153;
											assign node5153 = (inp[14]) ? node5159 : node5154;
												assign node5154 = (inp[0]) ? node5156 : 1'b1;
													assign node5156 = (inp[7]) ? 1'b0 : 1'b1;
												assign node5159 = (inp[11]) ? 1'b0 : node5160;
													assign node5160 = (inp[0]) ? 1'b0 : 1'b1;
											assign node5164 = (inp[9]) ? 1'b0 : node5165;
												assign node5165 = (inp[14]) ? 1'b0 : node5166;
													assign node5166 = (inp[0]) ? 1'b0 : 1'b1;
										assign node5171 = (inp[9]) ? 1'b0 : node5172;
											assign node5172 = (inp[0]) ? 1'b0 : node5173;
												assign node5173 = (inp[7]) ? 1'b0 : node5174;
													assign node5174 = (inp[11]) ? 1'b0 : 1'b1;
						assign node5180 = (inp[11]) ? node5302 : node5181;
							assign node5181 = (inp[10]) ? node5239 : node5182;
								assign node5182 = (inp[0]) ? node5200 : node5183;
									assign node5183 = (inp[9]) ? node5185 : 1'b1;
										assign node5185 = (inp[4]) ? node5193 : node5186;
											assign node5186 = (inp[14]) ? node5188 : 1'b1;
												assign node5188 = (inp[13]) ? node5190 : 1'b1;
													assign node5190 = (inp[7]) ? 1'b0 : 1'b1;
											assign node5193 = (inp[13]) ? 1'b0 : node5194;
												assign node5194 = (inp[5]) ? node5196 : 1'b1;
													assign node5196 = (inp[14]) ? 1'b0 : 1'b1;
									assign node5200 = (inp[12]) ? node5220 : node5201;
										assign node5201 = (inp[7]) ? node5209 : node5202;
											assign node5202 = (inp[9]) ? node5204 : 1'b1;
												assign node5204 = (inp[4]) ? node5206 : 1'b1;
													assign node5206 = (inp[13]) ? 1'b0 : 1'b1;
											assign node5209 = (inp[14]) ? node5215 : node5210;
												assign node5210 = (inp[5]) ? node5212 : 1'b1;
													assign node5212 = (inp[4]) ? 1'b0 : 1'b1;
												assign node5215 = (inp[13]) ? 1'b0 : node5216;
													assign node5216 = (inp[5]) ? 1'b0 : 1'b1;
										assign node5220 = (inp[13]) ? node5232 : node5221;
											assign node5221 = (inp[4]) ? node5227 : node5222;
												assign node5222 = (inp[7]) ? node5224 : 1'b1;
													assign node5224 = (inp[9]) ? 1'b0 : 1'b1;
												assign node5227 = (inp[9]) ? 1'b0 : node5228;
													assign node5228 = (inp[14]) ? 1'b0 : 1'b1;
											assign node5232 = (inp[9]) ? 1'b0 : node5233;
												assign node5233 = (inp[4]) ? 1'b0 : node5234;
													assign node5234 = (inp[14]) ? 1'b0 : 1'b1;
								assign node5239 = (inp[14]) ? node5273 : node5240;
									assign node5240 = (inp[12]) ? node5254 : node5241;
										assign node5241 = (inp[4]) ? node5243 : 1'b1;
											assign node5243 = (inp[13]) ? node5249 : node5244;
												assign node5244 = (inp[0]) ? node5246 : 1'b1;
													assign node5246 = (inp[9]) ? 1'b0 : 1'b1;
												assign node5249 = (inp[9]) ? 1'b0 : node5250;
													assign node5250 = (inp[5]) ? 1'b0 : 1'b1;
										assign node5254 = (inp[7]) ? node5266 : node5255;
											assign node5255 = (inp[0]) ? node5261 : node5256;
												assign node5256 = (inp[5]) ? node5258 : 1'b1;
													assign node5258 = (inp[4]) ? 1'b0 : 1'b1;
												assign node5261 = (inp[9]) ? 1'b0 : node5262;
													assign node5262 = (inp[4]) ? 1'b0 : 1'b1;
											assign node5266 = (inp[5]) ? 1'b0 : node5267;
												assign node5267 = (inp[4]) ? 1'b0 : node5268;
													assign node5268 = (inp[0]) ? 1'b0 : 1'b0;
									assign node5273 = (inp[9]) ? node5293 : node5274;
										assign node5274 = (inp[7]) ? node5286 : node5275;
											assign node5275 = (inp[0]) ? node5281 : node5276;
												assign node5276 = (inp[5]) ? node5278 : 1'b1;
													assign node5278 = (inp[12]) ? 1'b0 : 1'b1;
												assign node5281 = (inp[13]) ? 1'b0 : node5282;
													assign node5282 = (inp[12]) ? 1'b0 : 1'b1;
											assign node5286 = (inp[13]) ? 1'b0 : node5287;
												assign node5287 = (inp[4]) ? 1'b0 : node5288;
													assign node5288 = (inp[0]) ? 1'b0 : 1'b1;
										assign node5293 = (inp[0]) ? 1'b0 : node5294;
											assign node5294 = (inp[5]) ? 1'b0 : node5295;
												assign node5295 = (inp[13]) ? 1'b0 : node5296;
													assign node5296 = (inp[7]) ? 1'b0 : 1'b1;
							assign node5302 = (inp[4]) ? node5372 : node5303;
								assign node5303 = (inp[0]) ? node5343 : node5304;
									assign node5304 = (inp[7]) ? node5324 : node5305;
										assign node5305 = (inp[12]) ? node5313 : node5306;
											assign node5306 = (inp[13]) ? node5308 : 1'b1;
												assign node5308 = (inp[14]) ? node5310 : 1'b1;
													assign node5310 = (inp[5]) ? 1'b1 : 1'b0;
											assign node5313 = (inp[5]) ? node5319 : node5314;
												assign node5314 = (inp[14]) ? node5316 : 1'b1;
													assign node5316 = (inp[13]) ? 1'b0 : 1'b1;
												assign node5319 = (inp[10]) ? 1'b0 : node5320;
													assign node5320 = (inp[14]) ? 1'b0 : 1'b1;
										assign node5324 = (inp[14]) ? node5336 : node5325;
											assign node5325 = (inp[13]) ? node5331 : node5326;
												assign node5326 = (inp[12]) ? node5328 : 1'b1;
													assign node5328 = (inp[9]) ? 1'b0 : 1'b1;
												assign node5331 = (inp[12]) ? 1'b0 : node5332;
													assign node5332 = (inp[9]) ? 1'b0 : 1'b1;
											assign node5336 = (inp[10]) ? 1'b0 : node5337;
												assign node5337 = (inp[9]) ? 1'b0 : node5338;
													assign node5338 = (inp[5]) ? 1'b0 : 1'b1;
									assign node5343 = (inp[5]) ? node5363 : node5344;
										assign node5344 = (inp[12]) ? node5356 : node5345;
											assign node5345 = (inp[9]) ? node5351 : node5346;
												assign node5346 = (inp[14]) ? node5348 : 1'b1;
													assign node5348 = (inp[13]) ? 1'b0 : 1'b1;
												assign node5351 = (inp[13]) ? 1'b0 : node5352;
													assign node5352 = (inp[7]) ? 1'b0 : 1'b1;
											assign node5356 = (inp[14]) ? 1'b0 : node5357;
												assign node5357 = (inp[10]) ? 1'b0 : node5358;
													assign node5358 = (inp[7]) ? 1'b0 : 1'b1;
										assign node5363 = (inp[7]) ? 1'b0 : node5364;
											assign node5364 = (inp[14]) ? 1'b0 : node5365;
												assign node5365 = (inp[13]) ? 1'b0 : node5366;
													assign node5366 = (inp[10]) ? 1'b0 : 1'b1;
								assign node5372 = (inp[9]) ? node5398 : node5373;
									assign node5373 = (inp[14]) ? node5389 : node5374;
										assign node5374 = (inp[5]) ? node5382 : node5375;
											assign node5375 = (inp[13]) ? node5377 : 1'b1;
												assign node5377 = (inp[0]) ? 1'b0 : node5378;
													assign node5378 = (inp[7]) ? 1'b0 : 1'b1;
											assign node5382 = (inp[10]) ? 1'b0 : node5383;
												assign node5383 = (inp[13]) ? 1'b0 : node5384;
													assign node5384 = (inp[0]) ? 1'b0 : 1'b1;
										assign node5389 = (inp[10]) ? 1'b0 : node5390;
											assign node5390 = (inp[12]) ? 1'b0 : node5391;
												assign node5391 = (inp[5]) ? 1'b0 : node5392;
													assign node5392 = (inp[0]) ? 1'b0 : 1'b1;
									assign node5398 = (inp[5]) ? 1'b0 : node5399;
										assign node5399 = (inp[12]) ? 1'b0 : node5400;
											assign node5400 = (inp[10]) ? 1'b0 : node5401;
												assign node5401 = (inp[7]) ? 1'b0 : node5402;
													assign node5402 = (inp[13]) ? 1'b0 : 1'b1;
					assign node5409 = (inp[4]) ? node5641 : node5410;
						assign node5410 = (inp[5]) ? node5550 : node5411;
							assign node5411 = (inp[2]) ? node5481 : node5412;
								assign node5412 = (inp[10]) ? node5442 : node5413;
									assign node5413 = (inp[11]) ? node5423 : node5414;
										assign node5414 = (inp[9]) ? node5416 : 1'b1;
											assign node5416 = (inp[13]) ? node5418 : 1'b1;
												assign node5418 = (inp[14]) ? node5420 : 1'b1;
													assign node5420 = (inp[7]) ? 1'b0 : 1'b1;
										assign node5423 = (inp[7]) ? node5431 : node5424;
											assign node5424 = (inp[14]) ? node5426 : 1'b1;
												assign node5426 = (inp[0]) ? node5428 : 1'b1;
													assign node5428 = (inp[13]) ? 1'b0 : 1'b1;
											assign node5431 = (inp[0]) ? node5437 : node5432;
												assign node5432 = (inp[12]) ? node5434 : 1'b1;
													assign node5434 = (inp[14]) ? 1'b0 : 1'b1;
												assign node5437 = (inp[9]) ? 1'b0 : node5438;
													assign node5438 = (inp[12]) ? 1'b0 : 1'b1;
									assign node5442 = (inp[11]) ? node5462 : node5443;
										assign node5443 = (inp[0]) ? node5451 : node5444;
											assign node5444 = (inp[13]) ? node5446 : 1'b1;
												assign node5446 = (inp[12]) ? node5448 : 1'b1;
													assign node5448 = (inp[7]) ? 1'b0 : 1'b1;
											assign node5451 = (inp[9]) ? node5457 : node5452;
												assign node5452 = (inp[7]) ? node5454 : 1'b1;
													assign node5454 = (inp[12]) ? 1'b0 : 1'b1;
												assign node5457 = (inp[12]) ? 1'b0 : node5458;
													assign node5458 = (inp[13]) ? 1'b0 : 1'b1;
										assign node5462 = (inp[7]) ? node5474 : node5463;
											assign node5463 = (inp[12]) ? node5469 : node5464;
												assign node5464 = (inp[13]) ? node5466 : 1'b1;
													assign node5466 = (inp[0]) ? 1'b0 : 1'b1;
												assign node5469 = (inp[14]) ? 1'b0 : node5470;
													assign node5470 = (inp[13]) ? 1'b0 : 1'b1;
											assign node5474 = (inp[14]) ? 1'b0 : node5475;
												assign node5475 = (inp[13]) ? 1'b0 : node5476;
													assign node5476 = (inp[12]) ? 1'b0 : 1'b0;
								assign node5481 = (inp[9]) ? node5521 : node5482;
									assign node5482 = (inp[0]) ? node5502 : node5483;
										assign node5483 = (inp[13]) ? node5491 : node5484;
											assign node5484 = (inp[12]) ? node5486 : 1'b1;
												assign node5486 = (inp[7]) ? node5488 : 1'b1;
													assign node5488 = (inp[11]) ? 1'b0 : 1'b1;
											assign node5491 = (inp[7]) ? node5497 : node5492;
												assign node5492 = (inp[11]) ? node5494 : 1'b1;
													assign node5494 = (inp[10]) ? 1'b0 : 1'b1;
												assign node5497 = (inp[14]) ? 1'b0 : node5498;
													assign node5498 = (inp[11]) ? 1'b0 : 1'b1;
										assign node5502 = (inp[7]) ? node5514 : node5503;
											assign node5503 = (inp[13]) ? node5509 : node5504;
												assign node5504 = (inp[11]) ? node5506 : 1'b1;
													assign node5506 = (inp[10]) ? 1'b0 : 1'b1;
												assign node5509 = (inp[10]) ? 1'b0 : node5510;
													assign node5510 = (inp[12]) ? 1'b0 : 1'b1;
											assign node5514 = (inp[14]) ? 1'b0 : node5515;
												assign node5515 = (inp[12]) ? 1'b0 : node5516;
													assign node5516 = (inp[13]) ? 1'b0 : 1'b1;
									assign node5521 = (inp[7]) ? node5541 : node5522;
										assign node5522 = (inp[0]) ? node5534 : node5523;
											assign node5523 = (inp[11]) ? node5529 : node5524;
												assign node5524 = (inp[13]) ? node5526 : 1'b1;
													assign node5526 = (inp[12]) ? 1'b0 : 1'b1;
												assign node5529 = (inp[14]) ? 1'b0 : node5530;
													assign node5530 = (inp[12]) ? 1'b0 : 1'b1;
											assign node5534 = (inp[14]) ? 1'b0 : node5535;
												assign node5535 = (inp[11]) ? 1'b0 : node5536;
													assign node5536 = (inp[10]) ? 1'b0 : 1'b1;
										assign node5541 = (inp[10]) ? 1'b0 : node5542;
											assign node5542 = (inp[12]) ? 1'b0 : node5543;
												assign node5543 = (inp[11]) ? 1'b0 : node5544;
													assign node5544 = (inp[14]) ? 1'b0 : 1'b1;
							assign node5550 = (inp[13]) ? node5612 : node5551;
								assign node5551 = (inp[9]) ? node5587 : node5552;
									assign node5552 = (inp[2]) ? node5568 : node5553;
										assign node5553 = (inp[0]) ? node5561 : node5554;
											assign node5554 = (inp[7]) ? node5556 : 1'b1;
												assign node5556 = (inp[11]) ? node5558 : 1'b1;
													assign node5558 = (inp[14]) ? 1'b0 : 1'b1;
											assign node5561 = (inp[10]) ? node5563 : 1'b1;
												assign node5563 = (inp[14]) ? 1'b0 : node5564;
													assign node5564 = (inp[12]) ? 1'b0 : 1'b1;
										assign node5568 = (inp[14]) ? node5580 : node5569;
											assign node5569 = (inp[11]) ? node5575 : node5570;
												assign node5570 = (inp[10]) ? node5572 : 1'b1;
													assign node5572 = (inp[0]) ? 1'b0 : 1'b1;
												assign node5575 = (inp[7]) ? 1'b0 : node5576;
													assign node5576 = (inp[10]) ? 1'b0 : 1'b0;
											assign node5580 = (inp[12]) ? 1'b0 : node5581;
												assign node5581 = (inp[7]) ? 1'b0 : node5582;
													assign node5582 = (inp[10]) ? 1'b0 : 1'b1;
									assign node5587 = (inp[11]) ? node5603 : node5588;
										assign node5588 = (inp[12]) ? node5596 : node5589;
											assign node5589 = (inp[7]) ? node5591 : 1'b1;
												assign node5591 = (inp[0]) ? 1'b0 : node5592;
													assign node5592 = (inp[10]) ? 1'b0 : 1'b1;
											assign node5596 = (inp[10]) ? 1'b0 : node5597;
												assign node5597 = (inp[2]) ? 1'b0 : node5598;
													assign node5598 = (inp[14]) ? 1'b0 : 1'b1;
										assign node5603 = (inp[12]) ? 1'b0 : node5604;
											assign node5604 = (inp[14]) ? 1'b0 : node5605;
												assign node5605 = (inp[0]) ? 1'b0 : node5606;
													assign node5606 = (inp[2]) ? 1'b0 : 1'b0;
								assign node5612 = (inp[14]) ? 1'b0 : node5613;
									assign node5613 = (inp[7]) ? node5633 : node5614;
										assign node5614 = (inp[0]) ? node5626 : node5615;
											assign node5615 = (inp[10]) ? node5621 : node5616;
												assign node5616 = (inp[9]) ? node5618 : 1'b1;
													assign node5618 = (inp[2]) ? 1'b0 : 1'b1;
												assign node5621 = (inp[9]) ? 1'b0 : node5622;
													assign node5622 = (inp[12]) ? 1'b0 : 1'b1;
											assign node5626 = (inp[10]) ? 1'b0 : node5627;
												assign node5627 = (inp[9]) ? 1'b0 : node5628;
													assign node5628 = (inp[2]) ? 1'b0 : 1'b1;
										assign node5633 = (inp[10]) ? 1'b0 : node5634;
											assign node5634 = (inp[9]) ? 1'b0 : node5635;
												assign node5635 = (inp[11]) ? 1'b0 : 1'b1;
						assign node5641 = (inp[14]) ? node5743 : node5642;
							assign node5642 = (inp[0]) ? node5702 : node5643;
								assign node5643 = (inp[9]) ? node5677 : node5644;
									assign node5644 = (inp[5]) ? node5664 : node5645;
										assign node5645 = (inp[7]) ? node5653 : node5646;
											assign node5646 = (inp[2]) ? node5648 : 1'b1;
												assign node5648 = (inp[12]) ? node5650 : 1'b1;
													assign node5650 = (inp[11]) ? 1'b1 : 1'b0;
											assign node5653 = (inp[12]) ? node5659 : node5654;
												assign node5654 = (inp[11]) ? node5656 : 1'b1;
													assign node5656 = (inp[13]) ? 1'b0 : 1'b1;
												assign node5659 = (inp[11]) ? 1'b0 : node5660;
													assign node5660 = (inp[13]) ? 1'b0 : 1'b1;
										assign node5664 = (inp[2]) ? 1'b0 : node5665;
											assign node5665 = (inp[11]) ? node5671 : node5666;
												assign node5666 = (inp[10]) ? node5668 : 1'b1;
													assign node5668 = (inp[13]) ? 1'b0 : 1'b1;
												assign node5671 = (inp[10]) ? 1'b0 : node5672;
													assign node5672 = (inp[13]) ? 1'b0 : 1'b1;
									assign node5677 = (inp[13]) ? node5693 : node5678;
										assign node5678 = (inp[11]) ? node5686 : node5679;
											assign node5679 = (inp[10]) ? node5681 : 1'b1;
												assign node5681 = (inp[2]) ? 1'b0 : node5682;
													assign node5682 = (inp[7]) ? 1'b0 : 1'b1;
											assign node5686 = (inp[7]) ? 1'b0 : node5687;
												assign node5687 = (inp[10]) ? 1'b0 : node5688;
													assign node5688 = (inp[2]) ? 1'b0 : 1'b0;
										assign node5693 = (inp[2]) ? 1'b0 : node5694;
											assign node5694 = (inp[7]) ? 1'b0 : node5695;
												assign node5695 = (inp[10]) ? 1'b0 : node5696;
													assign node5696 = (inp[12]) ? 1'b0 : 1'b1;
								assign node5702 = (inp[7]) ? node5732 : node5703;
									assign node5703 = (inp[12]) ? node5723 : node5704;
										assign node5704 = (inp[13]) ? node5716 : node5705;
											assign node5705 = (inp[10]) ? node5711 : node5706;
												assign node5706 = (inp[2]) ? node5708 : 1'b1;
													assign node5708 = (inp[9]) ? 1'b0 : 1'b1;
												assign node5711 = (inp[11]) ? 1'b0 : node5712;
													assign node5712 = (inp[9]) ? 1'b0 : 1'b1;
											assign node5716 = (inp[9]) ? 1'b0 : node5717;
												assign node5717 = (inp[5]) ? 1'b0 : node5718;
													assign node5718 = (inp[11]) ? 1'b0 : 1'b1;
										assign node5723 = (inp[9]) ? 1'b0 : node5724;
											assign node5724 = (inp[2]) ? 1'b0 : node5725;
												assign node5725 = (inp[5]) ? 1'b0 : node5726;
													assign node5726 = (inp[10]) ? 1'b0 : 1'b1;
									assign node5732 = (inp[2]) ? 1'b0 : node5733;
										assign node5733 = (inp[12]) ? 1'b0 : node5734;
											assign node5734 = (inp[10]) ? 1'b0 : node5735;
												assign node5735 = (inp[5]) ? 1'b0 : node5736;
													assign node5736 = (inp[11]) ? 1'b0 : 1'b0;
							assign node5743 = (inp[2]) ? node5785 : node5744;
								assign node5744 = (inp[12]) ? node5774 : node5745;
									assign node5745 = (inp[11]) ? node5765 : node5746;
										assign node5746 = (inp[7]) ? node5758 : node5747;
											assign node5747 = (inp[10]) ? node5753 : node5748;
												assign node5748 = (inp[13]) ? node5750 : 1'b1;
													assign node5750 = (inp[5]) ? 1'b0 : 1'b1;
												assign node5753 = (inp[5]) ? 1'b0 : node5754;
													assign node5754 = (inp[9]) ? 1'b0 : 1'b1;
											assign node5758 = (inp[5]) ? 1'b0 : node5759;
												assign node5759 = (inp[0]) ? 1'b0 : node5760;
													assign node5760 = (inp[9]) ? 1'b0 : 1'b1;
										assign node5765 = (inp[9]) ? 1'b0 : node5766;
											assign node5766 = (inp[0]) ? 1'b0 : node5767;
												assign node5767 = (inp[13]) ? 1'b0 : node5768;
													assign node5768 = (inp[10]) ? 1'b0 : 1'b1;
									assign node5774 = (inp[13]) ? 1'b0 : node5775;
										assign node5775 = (inp[5]) ? 1'b0 : node5776;
											assign node5776 = (inp[9]) ? 1'b0 : node5777;
												assign node5777 = (inp[7]) ? 1'b0 : node5778;
													assign node5778 = (inp[0]) ? 1'b0 : 1'b1;
								assign node5785 = (inp[5]) ? 1'b0 : node5786;
									assign node5786 = (inp[13]) ? 1'b0 : node5787;
										assign node5787 = (inp[0]) ? 1'b0 : node5788;
											assign node5788 = (inp[7]) ? 1'b0 : node5789;
												assign node5789 = (inp[11]) ? 1'b0 : 1'b1;
				assign node5796 = (inp[11]) ? node6172 : node5797;
					assign node5797 = (inp[6]) ? node6021 : node5798;
						assign node5798 = (inp[4]) ? node5920 : node5799;
							assign node5799 = (inp[12]) ? node5859 : node5800;
								assign node5800 = (inp[5]) ? node5830 : node5801;
									assign node5801 = (inp[14]) ? node5811 : node5802;
										assign node5802 = (inp[9]) ? node5804 : 1'b1;
											assign node5804 = (inp[10]) ? node5806 : 1'b1;
												assign node5806 = (inp[0]) ? node5808 : 1'b1;
													assign node5808 = (inp[2]) ? 1'b0 : 1'b1;
										assign node5811 = (inp[2]) ? node5819 : node5812;
											assign node5812 = (inp[7]) ? node5814 : 1'b1;
												assign node5814 = (inp[0]) ? node5816 : 1'b1;
													assign node5816 = (inp[10]) ? 1'b0 : 1'b1;
											assign node5819 = (inp[9]) ? node5825 : node5820;
												assign node5820 = (inp[13]) ? node5822 : 1'b1;
													assign node5822 = (inp[0]) ? 1'b0 : 1'b0;
												assign node5825 = (inp[7]) ? 1'b0 : node5826;
													assign node5826 = (inp[0]) ? 1'b0 : 1'b1;
									assign node5830 = (inp[13]) ? node5844 : node5831;
										assign node5831 = (inp[2]) ? node5833 : 1'b1;
											assign node5833 = (inp[10]) ? node5839 : node5834;
												assign node5834 = (inp[14]) ? node5836 : 1'b1;
													assign node5836 = (inp[0]) ? 1'b0 : 1'b1;
												assign node5839 = (inp[7]) ? 1'b0 : node5840;
													assign node5840 = (inp[0]) ? 1'b0 : 1'b1;
										assign node5844 = (inp[14]) ? node5852 : node5845;
											assign node5845 = (inp[10]) ? node5847 : 1'b1;
												assign node5847 = (inp[7]) ? 1'b0 : node5848;
													assign node5848 = (inp[2]) ? 1'b0 : 1'b1;
											assign node5852 = (inp[0]) ? 1'b0 : node5853;
												assign node5853 = (inp[7]) ? 1'b0 : node5854;
													assign node5854 = (inp[2]) ? 1'b0 : 1'b1;
								assign node5859 = (inp[2]) ? node5893 : node5860;
									assign node5860 = (inp[9]) ? node5874 : node5861;
										assign node5861 = (inp[14]) ? node5863 : 1'b1;
											assign node5863 = (inp[10]) ? node5869 : node5864;
												assign node5864 = (inp[0]) ? node5866 : 1'b1;
													assign node5866 = (inp[13]) ? 1'b0 : 1'b1;
												assign node5869 = (inp[7]) ? 1'b0 : node5870;
													assign node5870 = (inp[0]) ? 1'b0 : 1'b1;
										assign node5874 = (inp[5]) ? node5886 : node5875;
											assign node5875 = (inp[13]) ? node5881 : node5876;
												assign node5876 = (inp[14]) ? node5878 : 1'b1;
													assign node5878 = (inp[10]) ? 1'b0 : 1'b1;
												assign node5881 = (inp[10]) ? 1'b0 : node5882;
													assign node5882 = (inp[7]) ? 1'b0 : 1'b1;
											assign node5886 = (inp[10]) ? 1'b0 : node5887;
												assign node5887 = (inp[0]) ? node5889 : 1'b1;
													assign node5889 = (inp[13]) ? 1'b0 : 1'b0;
									assign node5893 = (inp[5]) ? node5911 : node5894;
										assign node5894 = (inp[0]) ? node5902 : node5895;
											assign node5895 = (inp[9]) ? node5897 : 1'b1;
												assign node5897 = (inp[10]) ? 1'b0 : node5898;
													assign node5898 = (inp[7]) ? 1'b0 : 1'b1;
											assign node5902 = (inp[10]) ? 1'b0 : node5903;
												assign node5903 = (inp[13]) ? node5907 : node5904;
													assign node5904 = (inp[7]) ? 1'b0 : 1'b1;
													assign node5907 = (inp[7]) ? 1'b0 : 1'b0;
										assign node5911 = (inp[13]) ? 1'b0 : node5912;
											assign node5912 = (inp[9]) ? 1'b0 : node5913;
												assign node5913 = (inp[7]) ? 1'b0 : node5914;
													assign node5914 = (inp[10]) ? 1'b0 : 1'b1;
							assign node5920 = (inp[10]) ? node5984 : node5921;
								assign node5921 = (inp[7]) ? node5959 : node5922;
									assign node5922 = (inp[5]) ? node5942 : node5923;
										assign node5923 = (inp[13]) ? node5931 : node5924;
											assign node5924 = (inp[9]) ? node5926 : 1'b1;
												assign node5926 = (inp[0]) ? node5928 : 1'b1;
													assign node5928 = (inp[12]) ? 1'b0 : 1'b1;
											assign node5931 = (inp[12]) ? node5937 : node5932;
												assign node5932 = (inp[9]) ? node5934 : 1'b1;
													assign node5934 = (inp[0]) ? 1'b0 : 1'b1;
												assign node5937 = (inp[0]) ? 1'b0 : node5938;
													assign node5938 = (inp[14]) ? 1'b0 : 1'b1;
										assign node5942 = (inp[0]) ? node5954 : node5943;
											assign node5943 = (inp[9]) ? node5949 : node5944;
												assign node5944 = (inp[13]) ? node5946 : 1'b1;
													assign node5946 = (inp[14]) ? 1'b0 : 1'b1;
												assign node5949 = (inp[13]) ? 1'b0 : node5950;
													assign node5950 = (inp[2]) ? 1'b0 : 1'b1;
											assign node5954 = (inp[14]) ? 1'b0 : node5955;
												assign node5955 = (inp[12]) ? 1'b0 : 1'b1;
									assign node5959 = (inp[0]) ? node5975 : node5960;
										assign node5960 = (inp[9]) ? node5968 : node5961;
											assign node5961 = (inp[2]) ? node5963 : 1'b1;
												assign node5963 = (inp[13]) ? 1'b0 : node5964;
													assign node5964 = (inp[12]) ? 1'b0 : 1'b1;
											assign node5968 = (inp[12]) ? 1'b0 : node5969;
												assign node5969 = (inp[2]) ? 1'b0 : node5970;
													assign node5970 = (inp[14]) ? 1'b0 : 1'b1;
										assign node5975 = (inp[12]) ? 1'b0 : node5976;
											assign node5976 = (inp[14]) ? 1'b0 : node5977;
												assign node5977 = (inp[5]) ? 1'b0 : node5978;
													assign node5978 = (inp[2]) ? 1'b0 : 1'b1;
								assign node5984 = (inp[2]) ? node6010 : node5985;
									assign node5985 = (inp[9]) ? node6001 : node5986;
										assign node5986 = (inp[0]) ? node5994 : node5987;
											assign node5987 = (inp[12]) ? node5989 : 1'b1;
												assign node5989 = (inp[14]) ? 1'b0 : node5990;
													assign node5990 = (inp[13]) ? 1'b0 : 1'b1;
											assign node5994 = (inp[14]) ? 1'b0 : node5995;
												assign node5995 = (inp[5]) ? 1'b0 : node5996;
													assign node5996 = (inp[7]) ? 1'b0 : 1'b1;
										assign node6001 = (inp[12]) ? 1'b0 : node6002;
											assign node6002 = (inp[13]) ? 1'b0 : node6003;
												assign node6003 = (inp[7]) ? 1'b0 : node6004;
													assign node6004 = (inp[5]) ? 1'b0 : 1'b1;
									assign node6010 = (inp[0]) ? 1'b0 : node6011;
										assign node6011 = (inp[9]) ? 1'b0 : node6012;
											assign node6012 = (inp[12]) ? 1'b0 : node6013;
												assign node6013 = (inp[13]) ? 1'b0 : node6014;
													assign node6014 = (inp[7]) ? 1'b0 : 1'b1;
						assign node6021 = (inp[12]) ? node6117 : node6022;
							assign node6022 = (inp[5]) ? node6086 : node6023;
								assign node6023 = (inp[7]) ? node6059 : node6024;
									assign node6024 = (inp[2]) ? node6040 : node6025;
										assign node6025 = (inp[14]) ? node6033 : node6026;
											assign node6026 = (inp[9]) ? node6028 : 1'b1;
												assign node6028 = (inp[0]) ? node6030 : 1'b1;
													assign node6030 = (inp[13]) ? 1'b0 : 1'b1;
											assign node6033 = (inp[0]) ? 1'b0 : node6034;
												assign node6034 = (inp[10]) ? node6036 : 1'b1;
													assign node6036 = (inp[13]) ? 1'b0 : 1'b1;
										assign node6040 = (inp[10]) ? node6052 : node6041;
											assign node6041 = (inp[0]) ? node6047 : node6042;
												assign node6042 = (inp[13]) ? node6044 : 1'b1;
													assign node6044 = (inp[4]) ? 1'b0 : 1'b1;
												assign node6047 = (inp[9]) ? 1'b0 : node6048;
													assign node6048 = (inp[13]) ? 1'b0 : 1'b1;
											assign node6052 = (inp[14]) ? 1'b0 : node6053;
												assign node6053 = (inp[0]) ? 1'b0 : node6054;
													assign node6054 = (inp[13]) ? 1'b0 : 1'b1;
									assign node6059 = (inp[0]) ? node6079 : node6060;
										assign node6060 = (inp[10]) ? node6072 : node6061;
											assign node6061 = (inp[2]) ? node6067 : node6062;
												assign node6062 = (inp[9]) ? node6064 : 1'b1;
													assign node6064 = (inp[14]) ? 1'b0 : 1'b1;
												assign node6067 = (inp[13]) ? 1'b0 : node6068;
													assign node6068 = (inp[14]) ? 1'b0 : 1'b1;
											assign node6072 = (inp[9]) ? 1'b0 : node6073;
												assign node6073 = (inp[2]) ? 1'b0 : node6074;
													assign node6074 = (inp[14]) ? 1'b0 : 1'b1;
										assign node6079 = (inp[2]) ? 1'b0 : node6080;
											assign node6080 = (inp[10]) ? 1'b0 : node6081;
												assign node6081 = (inp[13]) ? 1'b0 : 1'b1;
								assign node6086 = (inp[10]) ? 1'b0 : node6087;
									assign node6087 = (inp[13]) ? node6107 : node6088;
										assign node6088 = (inp[7]) ? node6100 : node6089;
											assign node6089 = (inp[0]) ? node6095 : node6090;
												assign node6090 = (inp[14]) ? node6092 : 1'b1;
													assign node6092 = (inp[2]) ? 1'b0 : 1'b1;
												assign node6095 = (inp[9]) ? 1'b0 : node6096;
													assign node6096 = (inp[14]) ? 1'b0 : 1'b1;
											assign node6100 = (inp[2]) ? 1'b0 : node6101;
												assign node6101 = (inp[9]) ? 1'b0 : node6102;
													assign node6102 = (inp[0]) ? 1'b0 : 1'b1;
										assign node6107 = (inp[7]) ? 1'b0 : node6108;
											assign node6108 = (inp[0]) ? 1'b0 : node6109;
												assign node6109 = (inp[14]) ? 1'b0 : node6110;
													assign node6110 = (inp[2]) ? 1'b0 : 1'b1;
							assign node6117 = (inp[9]) ? node6159 : node6118;
								assign node6118 = (inp[13]) ? node6148 : node6119;
									assign node6119 = (inp[4]) ? node6141 : node6120;
										assign node6120 = (inp[5]) ? node6134 : node6121;
											assign node6121 = (inp[7]) ? node6127 : node6122;
												assign node6122 = (inp[14]) ? node6124 : 1'b1;
													assign node6124 = (inp[0]) ? 1'b0 : 1'b1;
												assign node6127 = (inp[0]) ? node6131 : node6128;
													assign node6128 = (inp[14]) ? 1'b0 : 1'b1;
													assign node6131 = (inp[10]) ? 1'b0 : 1'b0;
											assign node6134 = (inp[14]) ? 1'b0 : node6135;
												assign node6135 = (inp[0]) ? 1'b0 : node6136;
													assign node6136 = (inp[10]) ? 1'b0 : 1'b1;
										assign node6141 = (inp[0]) ? 1'b0 : node6142;
											assign node6142 = (inp[7]) ? 1'b0 : node6143;
												assign node6143 = (inp[2]) ? 1'b0 : 1'b1;
									assign node6148 = (inp[10]) ? 1'b0 : node6149;
										assign node6149 = (inp[5]) ? 1'b0 : node6150;
											assign node6150 = (inp[4]) ? 1'b0 : node6151;
												assign node6151 = (inp[2]) ? 1'b0 : node6152;
													assign node6152 = (inp[0]) ? 1'b0 : 1'b1;
								assign node6159 = (inp[2]) ? 1'b0 : node6160;
									assign node6160 = (inp[5]) ? 1'b0 : node6161;
										assign node6161 = (inp[7]) ? 1'b0 : node6162;
											assign node6162 = (inp[0]) ? 1'b0 : node6163;
												assign node6163 = (inp[14]) ? 1'b0 : node6164;
													assign node6164 = (inp[10]) ? 1'b0 : 1'b1;
					assign node6172 = (inp[0]) ? node6334 : node6173;
						assign node6173 = (inp[9]) ? node6279 : node6174;
							assign node6174 = (inp[4]) ? node6240 : node6175;
								assign node6175 = (inp[14]) ? node6211 : node6176;
									assign node6176 = (inp[12]) ? node6192 : node6177;
										assign node6177 = (inp[7]) ? node6185 : node6178;
											assign node6178 = (inp[13]) ? node6180 : 1'b1;
												assign node6180 = (inp[5]) ? node6182 : 1'b1;
													assign node6182 = (inp[2]) ? 1'b0 : 1'b1;
											assign node6185 = (inp[6]) ? node6187 : 1'b1;
												assign node6187 = (inp[5]) ? 1'b0 : node6188;
													assign node6188 = (inp[2]) ? 1'b0 : 1'b1;
										assign node6192 = (inp[2]) ? node6204 : node6193;
											assign node6193 = (inp[13]) ? node6199 : node6194;
												assign node6194 = (inp[10]) ? node6196 : 1'b1;
													assign node6196 = (inp[7]) ? 1'b0 : 1'b1;
												assign node6199 = (inp[6]) ? 1'b0 : node6200;
													assign node6200 = (inp[7]) ? 1'b0 : 1'b1;
											assign node6204 = (inp[10]) ? 1'b0 : node6205;
												assign node6205 = (inp[6]) ? 1'b0 : node6206;
													assign node6206 = (inp[13]) ? 1'b0 : 1'b1;
									assign node6211 = (inp[10]) ? node6231 : node6212;
										assign node6212 = (inp[13]) ? node6224 : node6213;
											assign node6213 = (inp[12]) ? node6219 : node6214;
												assign node6214 = (inp[5]) ? node6216 : 1'b1;
													assign node6216 = (inp[7]) ? 1'b0 : 1'b1;
												assign node6219 = (inp[6]) ? 1'b0 : node6220;
													assign node6220 = (inp[5]) ? 1'b0 : 1'b1;
											assign node6224 = (inp[7]) ? 1'b0 : node6225;
												assign node6225 = (inp[6]) ? 1'b0 : node6226;
													assign node6226 = (inp[5]) ? 1'b0 : 1'b1;
										assign node6231 = (inp[2]) ? 1'b0 : node6232;
											assign node6232 = (inp[5]) ? 1'b0 : node6233;
												assign node6233 = (inp[7]) ? 1'b0 : node6234;
													assign node6234 = (inp[6]) ? 1'b0 : 1'b1;
								assign node6240 = (inp[2]) ? node6270 : node6241;
									assign node6241 = (inp[12]) ? node6261 : node6242;
										assign node6242 = (inp[13]) ? node6254 : node6243;
											assign node6243 = (inp[5]) ? node6249 : node6244;
												assign node6244 = (inp[7]) ? node6246 : 1'b1;
													assign node6246 = (inp[6]) ? 1'b0 : 1'b1;
												assign node6249 = (inp[14]) ? 1'b0 : node6250;
													assign node6250 = (inp[7]) ? 1'b0 : 1'b1;
											assign node6254 = (inp[6]) ? 1'b0 : node6255;
												assign node6255 = (inp[10]) ? 1'b0 : node6256;
													assign node6256 = (inp[7]) ? 1'b0 : 1'b0;
										assign node6261 = (inp[10]) ? 1'b0 : node6262;
											assign node6262 = (inp[14]) ? 1'b0 : node6263;
												assign node6263 = (inp[6]) ? 1'b0 : node6264;
													assign node6264 = (inp[13]) ? 1'b0 : 1'b1;
									assign node6270 = (inp[10]) ? 1'b0 : node6271;
										assign node6271 = (inp[5]) ? 1'b0 : node6272;
											assign node6272 = (inp[7]) ? 1'b0 : node6273;
												assign node6273 = (inp[13]) ? 1'b0 : 1'b1;
							assign node6279 = (inp[7]) ? node6321 : node6280;
								assign node6280 = (inp[10]) ? node6310 : node6281;
									assign node6281 = (inp[12]) ? node6301 : node6282;
										assign node6282 = (inp[5]) ? node6294 : node6283;
											assign node6283 = (inp[6]) ? node6289 : node6284;
												assign node6284 = (inp[13]) ? node6286 : 1'b1;
													assign node6286 = (inp[2]) ? 1'b0 : 1'b1;
												assign node6289 = (inp[14]) ? 1'b0 : node6290;
													assign node6290 = (inp[13]) ? 1'b0 : 1'b1;
											assign node6294 = (inp[2]) ? 1'b0 : node6295;
												assign node6295 = (inp[4]) ? 1'b0 : node6296;
													assign node6296 = (inp[14]) ? 1'b0 : 1'b1;
										assign node6301 = (inp[14]) ? 1'b0 : node6302;
											assign node6302 = (inp[5]) ? 1'b0 : node6303;
												assign node6303 = (inp[4]) ? 1'b0 : node6304;
													assign node6304 = (inp[2]) ? 1'b0 : 1'b1;
									assign node6310 = (inp[6]) ? 1'b0 : node6311;
										assign node6311 = (inp[13]) ? 1'b0 : node6312;
											assign node6312 = (inp[2]) ? 1'b0 : node6313;
												assign node6313 = (inp[5]) ? 1'b0 : node6314;
													assign node6314 = (inp[12]) ? 1'b0 : 1'b1;
								assign node6321 = (inp[12]) ? 1'b0 : node6322;
									assign node6322 = (inp[6]) ? 1'b0 : node6323;
										assign node6323 = (inp[4]) ? 1'b0 : node6324;
											assign node6324 = (inp[2]) ? 1'b0 : node6325;
												assign node6325 = (inp[14]) ? 1'b0 : node6326;
													assign node6326 = (inp[10]) ? 1'b0 : 1'b1;
						assign node6334 = (inp[12]) ? node6384 : node6335;
							assign node6335 = (inp[7]) ? node6373 : node6336;
								assign node6336 = (inp[9]) ? node6362 : node6337;
									assign node6337 = (inp[5]) ? node6353 : node6338;
										assign node6338 = (inp[6]) ? node6346 : node6339;
											assign node6339 = (inp[4]) ? node6341 : 1'b1;
												assign node6341 = (inp[14]) ? node6343 : 1'b1;
													assign node6343 = (inp[10]) ? 1'b0 : 1'b0;
											assign node6346 = (inp[14]) ? 1'b0 : node6347;
												assign node6347 = (inp[2]) ? 1'b0 : node6348;
													assign node6348 = (inp[4]) ? 1'b0 : 1'b1;
										assign node6353 = (inp[4]) ? 1'b0 : node6354;
											assign node6354 = (inp[14]) ? 1'b0 : node6355;
												assign node6355 = (inp[13]) ? 1'b0 : node6356;
													assign node6356 = (inp[10]) ? 1'b0 : 1'b1;
									assign node6362 = (inp[10]) ? 1'b0 : node6363;
										assign node6363 = (inp[2]) ? 1'b0 : node6364;
											assign node6364 = (inp[14]) ? 1'b0 : node6365;
												assign node6365 = (inp[6]) ? 1'b0 : node6366;
													assign node6366 = (inp[13]) ? 1'b0 : 1'b1;
								assign node6373 = (inp[10]) ? 1'b0 : node6374;
									assign node6374 = (inp[2]) ? 1'b0 : node6375;
										assign node6375 = (inp[4]) ? 1'b0 : node6376;
											assign node6376 = (inp[14]) ? 1'b0 : node6377;
												assign node6377 = (inp[13]) ? 1'b0 : 1'b1;
							assign node6384 = (inp[6]) ? 1'b0 : node6385;
								assign node6385 = (inp[2]) ? 1'b0 : node6386;
									assign node6386 = (inp[9]) ? 1'b0 : node6387;
										assign node6387 = (inp[13]) ? 1'b0 : node6388;
											assign node6388 = (inp[4]) ? 1'b0 : node6389;
												assign node6389 = (inp[10]) ? 1'b0 : 1'b1;

endmodule