module dtc_split05_bm57 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node121;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node217;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node229;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node253;

	assign outp = (inp[8]) ? node126 : node1;
		assign node1 = (inp[5]) ? node67 : node2;
			assign node2 = (inp[6]) ? node28 : node3;
				assign node3 = (inp[4]) ? node15 : node4;
					assign node4 = (inp[9]) ? node12 : node5;
						assign node5 = (inp[11]) ? node9 : node6;
							assign node6 = (inp[0]) ? 3'b010 : 3'b000;
							assign node9 = (inp[0]) ? 3'b001 : 3'b011;
						assign node12 = (inp[10]) ? 3'b001 : 3'b011;
					assign node15 = (inp[11]) ? node23 : node16;
						assign node16 = (inp[10]) ? 3'b111 : node17;
							assign node17 = (inp[0]) ? node19 : 3'b101;
								assign node19 = (inp[2]) ? 3'b100 : 3'b101;
						assign node23 = (inp[10]) ? node25 : 3'b110;
							assign node25 = (inp[0]) ? 3'b100 : 3'b101;
				assign node28 = (inp[10]) ? node42 : node29;
					assign node29 = (inp[2]) ? node31 : 3'b101;
						assign node31 = (inp[9]) ? node37 : node32;
							assign node32 = (inp[7]) ? node34 : 3'b111;
								assign node34 = (inp[0]) ? 3'b111 : 3'b101;
							assign node37 = (inp[0]) ? node39 : 3'b111;
								assign node39 = (inp[1]) ? 3'b100 : 3'b110;
					assign node42 = (inp[11]) ? node56 : node43;
						assign node43 = (inp[7]) ? node49 : node44;
							assign node44 = (inp[2]) ? 3'b110 : node45;
								assign node45 = (inp[4]) ? 3'b111 : 3'b110;
							assign node49 = (inp[9]) ? node53 : node50;
								assign node50 = (inp[3]) ? 3'b110 : 3'b111;
								assign node53 = (inp[3]) ? 3'b111 : 3'b101;
						assign node56 = (inp[3]) ? node64 : node57;
							assign node57 = (inp[4]) ? 3'b101 : node58;
								assign node58 = (inp[2]) ? node60 : 3'b110;
									assign node60 = (inp[1]) ? 3'b110 : 3'b111;
							assign node64 = (inp[7]) ? 3'b100 : 3'b101;
			assign node67 = (inp[4]) ? node89 : node68;
				assign node68 = (inp[6]) ? node82 : node69;
					assign node69 = (inp[11]) ? node79 : node70;
						assign node70 = (inp[9]) ? node72 : 3'b101;
							assign node72 = (inp[7]) ? node76 : node73;
								assign node73 = (inp[10]) ? 3'b101 : 3'b111;
								assign node76 = (inp[10]) ? 3'b111 : 3'b101;
						assign node79 = (inp[3]) ? 3'b110 : 3'b100;
					assign node82 = (inp[0]) ? node86 : node83;
						assign node83 = (inp[1]) ? 3'b011 : 3'b010;
						assign node86 = (inp[10]) ? 3'b000 : 3'b010;
				assign node89 = (inp[11]) ? node105 : node90;
					assign node90 = (inp[9]) ? node96 : node91;
						assign node91 = (inp[3]) ? 3'b011 : node92;
							assign node92 = (inp[10]) ? 3'b011 : 3'b000;
						assign node96 = (inp[3]) ? node102 : node97;
							assign node97 = (inp[2]) ? 3'b001 : node98;
								assign node98 = (inp[7]) ? 3'b001 : 3'b011;
							assign node102 = (inp[0]) ? 3'b000 : 3'b001;
					assign node105 = (inp[10]) ? node111 : node106;
						assign node106 = (inp[7]) ? node108 : 3'b000;
							assign node108 = (inp[0]) ? 3'b010 : 3'b011;
						assign node111 = (inp[7]) ? node119 : node112;
							assign node112 = (inp[3]) ? node116 : node113;
								assign node113 = (inp[6]) ? 3'b000 : 3'b010;
								assign node116 = (inp[9]) ? 3'b001 : 3'b011;
							assign node119 = (inp[3]) ? node121 : 3'b001;
								assign node121 = (inp[9]) ? node123 : 3'b000;
									assign node123 = (inp[1]) ? 3'b001 : 3'b000;
		assign node126 = (inp[6]) ? node188 : node127;
			assign node127 = (inp[4]) ? node159 : node128;
				assign node128 = (inp[2]) ? node154 : node129;
					assign node129 = (inp[1]) ? node141 : node130;
						assign node130 = (inp[11]) ? node136 : node131;
							assign node131 = (inp[5]) ? 3'b101 : node132;
								assign node132 = (inp[9]) ? 3'b111 : 3'b101;
							assign node136 = (inp[0]) ? node138 : 3'b100;
								assign node138 = (inp[3]) ? 3'b111 : 3'b110;
						assign node141 = (inp[0]) ? node149 : node142;
							assign node142 = (inp[5]) ? 3'b101 : node143;
								assign node143 = (inp[11]) ? 3'b100 : node144;
									assign node144 = (inp[7]) ? 3'b110 : 3'b100;
							assign node149 = (inp[7]) ? 3'b101 : node150;
								assign node150 = (inp[10]) ? 3'b100 : 3'b101;
					assign node154 = (inp[9]) ? node156 : 3'b100;
						assign node156 = (inp[5]) ? 3'b111 : 3'b110;
				assign node159 = (inp[7]) ? node179 : node160;
					assign node160 = (inp[2]) ? node166 : node161;
						assign node161 = (inp[5]) ? 3'b011 : node162;
							assign node162 = (inp[11]) ? 3'b011 : 3'b001;
						assign node166 = (inp[0]) ? node172 : node167;
							assign node167 = (inp[5]) ? node169 : 3'b000;
								assign node169 = (inp[9]) ? 3'b011 : 3'b010;
							assign node172 = (inp[9]) ? node176 : node173;
								assign node173 = (inp[3]) ? 3'b001 : 3'b011;
								assign node176 = (inp[5]) ? 3'b010 : 3'b011;
					assign node179 = (inp[11]) ? node183 : node180;
						assign node180 = (inp[5]) ? 3'b001 : 3'b011;
						assign node183 = (inp[1]) ? 3'b000 : node184;
							assign node184 = (inp[10]) ? 3'b000 : 3'b001;
			assign node188 = (inp[5]) ? node224 : node189;
				assign node189 = (inp[11]) ? node205 : node190;
					assign node190 = (inp[4]) ? node196 : node191;
						assign node191 = (inp[0]) ? 3'b001 : node192;
							assign node192 = (inp[10]) ? 3'b000 : 3'b001;
						assign node196 = (inp[3]) ? node198 : 3'b011;
							assign node198 = (inp[0]) ? node200 : 3'b010;
								assign node200 = (inp[2]) ? 3'b011 : node201;
									assign node201 = (inp[10]) ? 3'b011 : 3'b010;
					assign node205 = (inp[3]) ? node217 : node206;
						assign node206 = (inp[4]) ? node212 : node207;
							assign node207 = (inp[2]) ? node209 : 3'b010;
								assign node209 = (inp[1]) ? 3'b010 : 3'b011;
							assign node212 = (inp[2]) ? 3'b000 : node213;
								assign node213 = (inp[7]) ? 3'b001 : 3'b000;
						assign node217 = (inp[1]) ? node219 : 3'b000;
							assign node219 = (inp[0]) ? 3'b001 : node220;
								assign node220 = (inp[7]) ? 3'b000 : 3'b001;
				assign node224 = (inp[3]) ? node242 : node225;
					assign node225 = (inp[4]) ? node233 : node226;
						assign node226 = (inp[7]) ? 3'b010 : node227;
							assign node227 = (inp[1]) ? node229 : 3'b011;
								assign node229 = (inp[11]) ? 3'b011 : 3'b010;
						assign node233 = (inp[1]) ? node235 : 3'b000;
							assign node235 = (inp[0]) ? 3'b000 : node236;
								assign node236 = (inp[10]) ? 3'b001 : node237;
									assign node237 = (inp[7]) ? 3'b001 : 3'b000;
					assign node242 = (inp[9]) ? node252 : node243;
						assign node243 = (inp[7]) ? node249 : node244;
							assign node244 = (inp[4]) ? node246 : 3'b000;
								assign node246 = (inp[0]) ? 3'b000 : 3'b001;
							assign node249 = (inp[1]) ? 3'b001 : 3'b000;
						assign node252 = (inp[0]) ? 3'b000 : node253;
							assign node253 = (inp[10]) ? 3'b000 : 3'b001;

endmodule