module dtc_split5_bm87 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node114;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node169;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node219;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node242;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node281;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node291;
	wire [3-1:0] node293;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node321;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node357;
	wire [3-1:0] node360;
	wire [3-1:0] node362;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node373;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node397;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node409;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node424;
	wire [3-1:0] node426;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node436;
	wire [3-1:0] node438;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node447;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node453;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node462;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node504;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node509;
	wire [3-1:0] node512;
	wire [3-1:0] node514;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node540;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node547;
	wire [3-1:0] node549;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node558;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node565;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node581;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node594;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node603;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node618;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node626;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node634;
	wire [3-1:0] node636;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node654;
	wire [3-1:0] node657;
	wire [3-1:0] node659;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node684;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node694;
	wire [3-1:0] node695;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node700;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node720;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node731;
	wire [3-1:0] node734;
	wire [3-1:0] node735;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node762;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node770;
	wire [3-1:0] node774;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node783;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node789;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node803;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node812;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node819;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node826;
	wire [3-1:0] node829;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node839;
	wire [3-1:0] node842;
	wire [3-1:0] node844;
	wire [3-1:0] node847;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node857;
	wire [3-1:0] node858;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node869;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node882;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node887;
	wire [3-1:0] node890;
	wire [3-1:0] node893;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node899;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node907;
	wire [3-1:0] node908;

	assign outp = (inp[6]) ? node186 : node1;
		assign node1 = (inp[7]) ? node33 : node2;
			assign node2 = (inp[9]) ? 3'b000 : node3;
				assign node3 = (inp[1]) ? 3'b000 : node4;
					assign node4 = (inp[8]) ? node6 : 3'b000;
						assign node6 = (inp[10]) ? 3'b000 : node7;
							assign node7 = (inp[0]) ? node9 : 3'b000;
								assign node9 = (inp[3]) ? node21 : node10;
									assign node10 = (inp[4]) ? node16 : node11;
										assign node11 = (inp[2]) ? node13 : 3'b100;
											assign node13 = (inp[11]) ? 3'b100 : 3'b000;
										assign node16 = (inp[2]) ? 3'b000 : node17;
											assign node17 = (inp[11]) ? 3'b000 : 3'b100;
									assign node21 = (inp[5]) ? 3'b000 : node22;
										assign node22 = (inp[2]) ? node26 : node23;
											assign node23 = (inp[11]) ? 3'b000 : 3'b100;
											assign node26 = (inp[11]) ? 3'b100 : 3'b000;
			assign node33 = (inp[9]) ? node151 : node34;
				assign node34 = (inp[0]) ? node90 : node35;
					assign node35 = (inp[10]) ? node73 : node36;
						assign node36 = (inp[1]) ? node40 : node37;
							assign node37 = (inp[11]) ? 3'b001 : 3'b101;
							assign node40 = (inp[8]) ? node58 : node41;
								assign node41 = (inp[3]) ? node51 : node42;
									assign node42 = (inp[2]) ? node44 : 3'b110;
										assign node44 = (inp[11]) ? node48 : node45;
											assign node45 = (inp[4]) ? 3'b010 : 3'b110;
											assign node48 = (inp[4]) ? 3'b110 : 3'b010;
									assign node51 = (inp[2]) ? node55 : node52;
										assign node52 = (inp[11]) ? 3'b010 : 3'b110;
										assign node55 = (inp[11]) ? 3'b110 : 3'b010;
								assign node58 = (inp[11]) ? node68 : node59;
									assign node59 = (inp[2]) ? node61 : 3'b001;
										assign node61 = (inp[5]) ? 3'b110 : node62;
											assign node62 = (inp[4]) ? 3'b001 : node63;
												assign node63 = (inp[3]) ? 3'b110 : 3'b001;
									assign node68 = (inp[3]) ? 3'b110 : node69;
										assign node69 = (inp[5]) ? 3'b110 : 3'b001;
						assign node73 = (inp[1]) ? node75 : 3'b110;
							assign node75 = (inp[8]) ? node79 : node76;
								assign node76 = (inp[11]) ? 3'b000 : 3'b100;
								assign node79 = (inp[11]) ? node85 : node80;
									assign node80 = (inp[2]) ? node82 : 3'b010;
										assign node82 = (inp[3]) ? 3'b100 : 3'b110;
									assign node85 = (inp[4]) ? 3'b100 : node86;
										assign node86 = (inp[5]) ? 3'b000 : 3'b110;
					assign node90 = (inp[10]) ? node142 : node91;
						assign node91 = (inp[1]) ? node117 : node92;
							assign node92 = (inp[3]) ? node108 : node93;
								assign node93 = (inp[11]) ? node101 : node94;
									assign node94 = (inp[8]) ? node96 : 3'b010;
										assign node96 = (inp[2]) ? node98 : 3'b110;
											assign node98 = (inp[4]) ? 3'b010 : 3'b110;
									assign node101 = (inp[2]) ? node105 : node102;
										assign node102 = (inp[8]) ? 3'b010 : 3'b100;
										assign node105 = (inp[8]) ? 3'b100 : 3'b010;
								assign node108 = (inp[8]) ? node114 : node109;
									assign node109 = (inp[11]) ? node111 : 3'b100;
										assign node111 = (inp[2]) ? 3'b010 : 3'b100;
									assign node114 = (inp[2]) ? 3'b100 : 3'b010;
							assign node117 = (inp[8]) ? node125 : node118;
								assign node118 = (inp[3]) ? 3'b000 : node119;
									assign node119 = (inp[2]) ? 3'b000 : node120;
										assign node120 = (inp[11]) ? 3'b000 : 3'b100;
								assign node125 = (inp[4]) ? node135 : node126;
									assign node126 = (inp[5]) ? 3'b100 : node127;
										assign node127 = (inp[3]) ? 3'b010 : node128;
											assign node128 = (inp[11]) ? 3'b100 : node129;
												assign node129 = (inp[2]) ? 3'b100 : 3'b010;
									assign node135 = (inp[3]) ? node139 : node136;
										assign node136 = (inp[11]) ? 3'b100 : 3'b010;
										assign node139 = (inp[11]) ? 3'b000 : 3'b100;
						assign node142 = (inp[11]) ? 3'b000 : node143;
							assign node143 = (inp[8]) ? node145 : 3'b000;
								assign node145 = (inp[2]) ? 3'b000 : node146;
									assign node146 = (inp[1]) ? 3'b000 : 3'b100;
				assign node151 = (inp[10]) ? 3'b000 : node152;
					assign node152 = (inp[0]) ? 3'b000 : node153;
						assign node153 = (inp[1]) ? node161 : node154;
							assign node154 = (inp[2]) ? node158 : node155;
								assign node155 = (inp[11]) ? 3'b110 : 3'b010;
								assign node158 = (inp[11]) ? 3'b000 : 3'b100;
							assign node161 = (inp[8]) ? node163 : 3'b000;
								assign node163 = (inp[3]) ? node173 : node164;
									assign node164 = (inp[4]) ? 3'b000 : node165;
										assign node165 = (inp[2]) ? node169 : node166;
											assign node166 = (inp[11]) ? 3'b000 : 3'b100;
											assign node169 = (inp[11]) ? 3'b100 : 3'b000;
									assign node173 = (inp[11]) ? node179 : node174;
										assign node174 = (inp[4]) ? node176 : 3'b000;
											assign node176 = (inp[2]) ? 3'b100 : 3'b000;
										assign node179 = (inp[2]) ? node181 : 3'b100;
											assign node181 = (inp[4]) ? 3'b000 : 3'b100;
		assign node186 = (inp[9]) ? node646 : node187;
			assign node187 = (inp[0]) ? node401 : node188;
				assign node188 = (inp[7]) ? node330 : node189;
					assign node189 = (inp[10]) ? node255 : node190;
						assign node190 = (inp[11]) ? node222 : node191;
							assign node191 = (inp[1]) ? node205 : node192;
								assign node192 = (inp[4]) ? node198 : node193;
									assign node193 = (inp[8]) ? node195 : 3'b011;
										assign node195 = (inp[3]) ? 3'b111 : 3'b011;
									assign node198 = (inp[8]) ? node202 : node199;
										assign node199 = (inp[3]) ? 3'b011 : 3'b111;
										assign node202 = (inp[2]) ? 3'b111 : 3'b011;
								assign node205 = (inp[8]) ? node213 : node206;
									assign node206 = (inp[2]) ? node208 : 3'b101;
										assign node208 = (inp[4]) ? node210 : 3'b001;
											assign node210 = (inp[3]) ? 3'b001 : 3'b101;
									assign node213 = (inp[4]) ? node217 : node214;
										assign node214 = (inp[3]) ? 3'b011 : 3'b101;
										assign node217 = (inp[3]) ? node219 : 3'b011;
											assign node219 = (inp[2]) ? 3'b101 : 3'b011;
							assign node222 = (inp[8]) ? node238 : node223;
								assign node223 = (inp[1]) ? node229 : node224;
									assign node224 = (inp[3]) ? 3'b101 : node225;
										assign node225 = (inp[2]) ? 3'b101 : 3'b001;
									assign node229 = (inp[4]) ? node231 : 3'b001;
										assign node231 = (inp[5]) ? node233 : 3'b110;
											assign node233 = (inp[2]) ? node235 : 3'b001;
												assign node235 = (inp[3]) ? 3'b110 : 3'b001;
								assign node238 = (inp[1]) ? node246 : node239;
									assign node239 = (inp[2]) ? 3'b011 : node240;
										assign node240 = (inp[3]) ? node242 : 3'b111;
											assign node242 = (inp[5]) ? 3'b011 : 3'b111;
									assign node246 = (inp[2]) ? node250 : node247;
										assign node247 = (inp[4]) ? 3'b101 : 3'b011;
										assign node250 = (inp[4]) ? node252 : 3'b101;
											assign node252 = (inp[3]) ? 3'b001 : 3'b101;
						assign node255 = (inp[8]) ? node297 : node256;
							assign node256 = (inp[1]) ? node274 : node257;
								assign node257 = (inp[5]) ? node269 : node258;
									assign node258 = (inp[3]) ? 3'b101 : node259;
										assign node259 = (inp[4]) ? node261 : 3'b001;
											assign node261 = (inp[11]) ? node265 : node262;
												assign node262 = (inp[2]) ? 3'b001 : 3'b101;
												assign node265 = (inp[2]) ? 3'b101 : 3'b001;
									assign node269 = (inp[11]) ? node271 : 3'b001;
										assign node271 = (inp[4]) ? 3'b110 : 3'b010;
								assign node274 = (inp[11]) ? node284 : node275;
									assign node275 = (inp[3]) ? node279 : node276;
										assign node276 = (inp[4]) ? 3'b110 : 3'b001;
										assign node279 = (inp[2]) ? node281 : 3'b110;
											assign node281 = (inp[4]) ? 3'b010 : 3'b110;
									assign node284 = (inp[5]) ? 3'b010 : node285;
										assign node285 = (inp[2]) ? node291 : node286;
											assign node286 = (inp[3]) ? 3'b010 : node287;
												assign node287 = (inp[4]) ? 3'b010 : 3'b110;
											assign node291 = (inp[4]) ? node293 : 3'b010;
												assign node293 = (inp[3]) ? 3'b100 : 3'b010;
							assign node297 = (inp[4]) ? node309 : node298;
								assign node298 = (inp[1]) ? node306 : node299;
									assign node299 = (inp[11]) ? node303 : node300;
										assign node300 = (inp[2]) ? 3'b101 : 3'b011;
										assign node303 = (inp[2]) ? 3'b001 : 3'b101;
									assign node306 = (inp[11]) ? 3'b110 : 3'b001;
								assign node309 = (inp[1]) ? node321 : node310;
									assign node310 = (inp[11]) ? node316 : node311;
										assign node311 = (inp[2]) ? 3'b101 : node312;
											assign node312 = (inp[5]) ? 3'b101 : 3'b011;
										assign node316 = (inp[3]) ? 3'b001 : node317;
											assign node317 = (inp[2]) ? 3'b011 : 3'b101;
									assign node321 = (inp[3]) ? node323 : 3'b001;
										assign node323 = (inp[2]) ? node327 : node324;
											assign node324 = (inp[11]) ? 3'b101 : 3'b001;
											assign node327 = (inp[5]) ? 3'b010 : 3'b001;
					assign node330 = (inp[10]) ? node346 : node331;
						assign node331 = (inp[1]) ? node333 : 3'b111;
							assign node333 = (inp[8]) ? 3'b111 : node334;
								assign node334 = (inp[11]) ? node340 : node335;
									assign node335 = (inp[3]) ? 3'b111 : node336;
										assign node336 = (inp[2]) ? 3'b111 : 3'b011;
									assign node340 = (inp[2]) ? 3'b011 : node341;
										assign node341 = (inp[3]) ? 3'b011 : 3'b111;
						assign node346 = (inp[1]) ? node376 : node347;
							assign node347 = (inp[11]) ? node353 : node348;
								assign node348 = (inp[8]) ? 3'b111 : node349;
									assign node349 = (inp[2]) ? 3'b011 : 3'b111;
								assign node353 = (inp[5]) ? node365 : node354;
									assign node354 = (inp[4]) ? node360 : node355;
										assign node355 = (inp[8]) ? node357 : 3'b011;
											assign node357 = (inp[2]) ? 3'b011 : 3'b111;
										assign node360 = (inp[2]) ? node362 : 3'b011;
											assign node362 = (inp[8]) ? 3'b011 : 3'b111;
									assign node365 = (inp[8]) ? node373 : node366;
										assign node366 = (inp[4]) ? 3'b101 : node367;
											assign node367 = (inp[2]) ? 3'b001 : node368;
												assign node368 = (inp[3]) ? 3'b001 : 3'b011;
										assign node373 = (inp[2]) ? 3'b011 : 3'b111;
							assign node376 = (inp[11]) ? node388 : node377;
								assign node377 = (inp[8]) ? node383 : node378;
									assign node378 = (inp[2]) ? 3'b101 : node379;
										assign node379 = (inp[4]) ? 3'b011 : 3'b101;
									assign node383 = (inp[2]) ? 3'b011 : node384;
										assign node384 = (inp[3]) ? 3'b011 : 3'b111;
								assign node388 = (inp[8]) ? node394 : node389;
									assign node389 = (inp[3]) ? 3'b001 : node390;
										assign node390 = (inp[2]) ? 3'b001 : 3'b101;
									assign node394 = (inp[2]) ? 3'b101 : node395;
										assign node395 = (inp[3]) ? node397 : 3'b001;
											assign node397 = (inp[5]) ? 3'b101 : 3'b001;
				assign node401 = (inp[7]) ? node517 : node402;
					assign node402 = (inp[10]) ? node456 : node403;
						assign node403 = (inp[1]) ? node429 : node404;
							assign node404 = (inp[8]) ? node416 : node405;
								assign node405 = (inp[11]) ? node409 : node406;
									assign node406 = (inp[4]) ? 3'b110 : 3'b001;
									assign node409 = (inp[2]) ? node411 : 3'b110;
										assign node411 = (inp[3]) ? 3'b010 : node412;
											assign node412 = (inp[4]) ? 3'b010 : 3'b110;
								assign node416 = (inp[11]) ? node424 : node417;
									assign node417 = (inp[2]) ? node419 : 3'b101;
										assign node419 = (inp[3]) ? 3'b001 : node420;
											assign node420 = (inp[4]) ? 3'b001 : 3'b101;
									assign node424 = (inp[2]) ? node426 : 3'b001;
										assign node426 = (inp[3]) ? 3'b110 : 3'b101;
							assign node429 = (inp[8]) ? node443 : node430;
								assign node430 = (inp[2]) ? node436 : node431;
									assign node431 = (inp[11]) ? 3'b010 : node432;
										assign node432 = (inp[4]) ? 3'b010 : 3'b110;
									assign node436 = (inp[11]) ? node438 : 3'b010;
										assign node438 = (inp[4]) ? node440 : 3'b100;
											assign node440 = (inp[5]) ? 3'b100 : 3'b010;
								assign node443 = (inp[11]) ? node447 : node444;
									assign node444 = (inp[2]) ? 3'b110 : 3'b001;
									assign node447 = (inp[4]) ? node449 : 3'b110;
										assign node449 = (inp[3]) ? node453 : node450;
											assign node450 = (inp[2]) ? 3'b010 : 3'b110;
											assign node453 = (inp[2]) ? 3'b001 : 3'b010;
						assign node456 = (inp[1]) ? node484 : node457;
							assign node457 = (inp[11]) ? node469 : node458;
								assign node458 = (inp[8]) ? node462 : node459;
									assign node459 = (inp[2]) ? 3'b100 : 3'b010;
									assign node462 = (inp[2]) ? node464 : 3'b110;
										assign node464 = (inp[4]) ? 3'b010 : node465;
											assign node465 = (inp[5]) ? 3'b010 : 3'b110;
								assign node469 = (inp[8]) ? node477 : node470;
									assign node470 = (inp[2]) ? 3'b000 : node471;
										assign node471 = (inp[4]) ? 3'b100 : node472;
											assign node472 = (inp[3]) ? 3'b100 : 3'b000;
									assign node477 = (inp[2]) ? 3'b100 : node478;
										assign node478 = (inp[3]) ? 3'b010 : node479;
											assign node479 = (inp[4]) ? 3'b010 : 3'b110;
							assign node484 = (inp[4]) ? node494 : node485;
								assign node485 = (inp[8]) ? node487 : 3'b100;
									assign node487 = (inp[11]) ? node491 : node488;
										assign node488 = (inp[2]) ? 3'b100 : 3'b010;
										assign node491 = (inp[2]) ? 3'b000 : 3'b100;
								assign node494 = (inp[8]) ? node504 : node495;
									assign node495 = (inp[11]) ? 3'b000 : node496;
										assign node496 = (inp[5]) ? node498 : 3'b000;
											assign node498 = (inp[3]) ? 3'b000 : node499;
												assign node499 = (inp[2]) ? 3'b000 : 3'b100;
									assign node504 = (inp[5]) ? node506 : 3'b100;
										assign node506 = (inp[3]) ? node512 : node507;
											assign node507 = (inp[2]) ? node509 : 3'b010;
												assign node509 = (inp[11]) ? 3'b000 : 3'b100;
											assign node512 = (inp[2]) ? node514 : 3'b100;
												assign node514 = (inp[11]) ? 3'b000 : 3'b100;
					assign node517 = (inp[10]) ? node585 : node518;
						assign node518 = (inp[1]) ? node552 : node519;
							assign node519 = (inp[8]) ? node543 : node520;
								assign node520 = (inp[2]) ? node534 : node521;
									assign node521 = (inp[11]) ? node527 : node522;
										assign node522 = (inp[4]) ? 3'b011 : node523;
											assign node523 = (inp[5]) ? 3'b001 : 3'b101;
										assign node527 = (inp[3]) ? 3'b101 : node528;
											assign node528 = (inp[4]) ? 3'b101 : node529;
												assign node529 = (inp[5]) ? 3'b111 : 3'b011;
									assign node534 = (inp[11]) ? node540 : node535;
										assign node535 = (inp[4]) ? 3'b101 : node536;
											assign node536 = (inp[5]) ? 3'b111 : 3'b101;
										assign node540 = (inp[4]) ? 3'b001 : 3'b101;
								assign node543 = (inp[2]) ? node547 : node544;
									assign node544 = (inp[11]) ? 3'b011 : 3'b111;
									assign node547 = (inp[11]) ? node549 : 3'b011;
										assign node549 = (inp[3]) ? 3'b011 : 3'b101;
							assign node552 = (inp[3]) ? node568 : node553;
								assign node553 = (inp[11]) ? node561 : node554;
									assign node554 = (inp[8]) ? node558 : node555;
										assign node555 = (inp[2]) ? 3'b001 : 3'b101;
										assign node558 = (inp[2]) ? 3'b101 : 3'b011;
									assign node561 = (inp[8]) ? node565 : node562;
										assign node562 = (inp[2]) ? 3'b111 : 3'b001;
										assign node565 = (inp[2]) ? 3'b001 : 3'b101;
								assign node568 = (inp[11]) ? node574 : node569;
									assign node569 = (inp[8]) ? 3'b101 : node570;
										assign node570 = (inp[2]) ? 3'b001 : 3'b101;
									assign node574 = (inp[2]) ? node578 : node575;
										assign node575 = (inp[8]) ? 3'b101 : 3'b001;
										assign node578 = (inp[8]) ? 3'b001 : node579;
											assign node579 = (inp[4]) ? node581 : 3'b111;
												assign node581 = (inp[5]) ? 3'b110 : 3'b111;
						assign node585 = (inp[1]) ? node621 : node586;
							assign node586 = (inp[2]) ? node606 : node587;
								assign node587 = (inp[4]) ? node597 : node588;
									assign node588 = (inp[8]) ? node594 : node589;
										assign node589 = (inp[5]) ? 3'b101 : node590;
											assign node590 = (inp[11]) ? 3'b101 : 3'b001;
										assign node594 = (inp[11]) ? 3'b001 : 3'b101;
									assign node597 = (inp[5]) ? node603 : node598;
										assign node598 = (inp[8]) ? 3'b101 : node599;
											assign node599 = (inp[11]) ? 3'b101 : 3'b001;
										assign node603 = (inp[3]) ? 3'b110 : 3'b101;
								assign node606 = (inp[4]) ? node614 : node607;
									assign node607 = (inp[8]) ? node611 : node608;
										assign node608 = (inp[11]) ? 3'b101 : 3'b001;
										assign node611 = (inp[11]) ? 3'b010 : 3'b101;
									assign node614 = (inp[11]) ? node618 : node615;
										assign node615 = (inp[8]) ? 3'b001 : 3'b110;
										assign node618 = (inp[8]) ? 3'b110 : 3'b010;
							assign node621 = (inp[8]) ? node629 : node622;
								assign node622 = (inp[2]) ? node626 : node623;
									assign node623 = (inp[11]) ? 3'b010 : 3'b110;
									assign node626 = (inp[11]) ? 3'b100 : 3'b010;
								assign node629 = (inp[11]) ? node639 : node630;
									assign node630 = (inp[2]) ? node634 : node631;
										assign node631 = (inp[3]) ? 3'b001 : 3'b000;
										assign node634 = (inp[3]) ? node636 : 3'b111;
											assign node636 = (inp[5]) ? 3'b111 : 3'b110;
									assign node639 = (inp[2]) ? 3'b010 : node640;
										assign node640 = (inp[3]) ? 3'b110 : node641;
											assign node641 = (inp[4]) ? 3'b110 : 3'b111;
			assign node646 = (inp[0]) ? node832 : node647;
				assign node647 = (inp[7]) ? node725 : node648;
					assign node648 = (inp[10]) ? node694 : node649;
						assign node649 = (inp[11]) ? node673 : node650;
							assign node650 = (inp[1]) ? node662 : node651;
								assign node651 = (inp[2]) ? node657 : node652;
									assign node652 = (inp[3]) ? node654 : 3'b110;
										assign node654 = (inp[4]) ? 3'b010 : 3'b110;
									assign node657 = (inp[8]) ? node659 : 3'b010;
										assign node659 = (inp[4]) ? 3'b010 : 3'b110;
								assign node662 = (inp[8]) ? node668 : node663;
									assign node663 = (inp[3]) ? 3'b100 : node664;
										assign node664 = (inp[5]) ? 3'b100 : 3'b010;
									assign node668 = (inp[3]) ? 3'b010 : node669;
										assign node669 = (inp[2]) ? 3'b010 : 3'b110;
							assign node673 = (inp[8]) ? node687 : node674;
								assign node674 = (inp[4]) ? node684 : node675;
									assign node675 = (inp[3]) ? 3'b000 : node676;
										assign node676 = (inp[5]) ? 3'b000 : node677;
											assign node677 = (inp[2]) ? 3'b000 : node678;
												assign node678 = (inp[1]) ? 3'b100 : 3'b000;
									assign node684 = (inp[1]) ? 3'b000 : 3'b100;
								assign node687 = (inp[1]) ? 3'b100 : node688;
									assign node688 = (inp[2]) ? 3'b010 : node689;
										assign node689 = (inp[4]) ? 3'b110 : 3'b101;
						assign node694 = (inp[1]) ? 3'b000 : node695;
							assign node695 = (inp[11]) ? node703 : node696;
								assign node696 = (inp[8]) ? node700 : node697;
									assign node697 = (inp[2]) ? 3'b000 : 3'b100;
									assign node700 = (inp[2]) ? 3'b100 : 3'b010;
								assign node703 = (inp[3]) ? node715 : node704;
									assign node704 = (inp[5]) ? node710 : node705;
										assign node705 = (inp[8]) ? 3'b000 : node706;
											assign node706 = (inp[2]) ? 3'b100 : 3'b000;
										assign node710 = (inp[2]) ? 3'b000 : node711;
											assign node711 = (inp[8]) ? 3'b100 : 3'b000;
									assign node715 = (inp[5]) ? 3'b000 : node716;
										assign node716 = (inp[2]) ? node720 : node717;
											assign node717 = (inp[8]) ? 3'b100 : 3'b000;
											assign node720 = (inp[8]) ? 3'b000 : 3'b100;
					assign node725 = (inp[10]) ? node777 : node726;
						assign node726 = (inp[1]) ? node754 : node727;
							assign node727 = (inp[8]) ? node743 : node728;
								assign node728 = (inp[5]) ? node734 : node729;
									assign node729 = (inp[2]) ? node731 : 3'b101;
										assign node731 = (inp[11]) ? 3'b110 : 3'b101;
									assign node734 = (inp[2]) ? node738 : node735;
										assign node735 = (inp[3]) ? 3'b001 : 3'b101;
										assign node738 = (inp[11]) ? 3'b110 : node739;
											assign node739 = (inp[4]) ? 3'b001 : 3'b101;
								assign node743 = (inp[2]) ? node747 : node744;
									assign node744 = (inp[11]) ? 3'b101 : 3'b011;
									assign node747 = (inp[11]) ? 3'b001 : node748;
										assign node748 = (inp[4]) ? 3'b101 : node749;
											assign node749 = (inp[3]) ? 3'b101 : 3'b011;
							assign node754 = (inp[8]) ? node766 : node755;
								assign node755 = (inp[11]) ? node757 : 3'b110;
									assign node757 = (inp[5]) ? 3'b110 : node758;
										assign node758 = (inp[3]) ? node762 : node759;
											assign node759 = (inp[2]) ? 3'b010 : 3'b110;
											assign node762 = (inp[4]) ? 3'b010 : 3'b001;
								assign node766 = (inp[11]) ? node774 : node767;
									assign node767 = (inp[2]) ? 3'b001 : node768;
										assign node768 = (inp[3]) ? node770 : 3'b101;
											assign node770 = (inp[5]) ? 3'b101 : 3'b001;
									assign node774 = (inp[2]) ? 3'b110 : 3'b010;
						assign node777 = (inp[1]) ? node793 : node778;
							assign node778 = (inp[2]) ? node786 : node779;
								assign node779 = (inp[11]) ? node783 : node780;
									assign node780 = (inp[8]) ? 3'b001 : 3'b110;
									assign node783 = (inp[8]) ? 3'b110 : 3'b010;
								assign node786 = (inp[11]) ? 3'b010 : node787;
									assign node787 = (inp[8]) ? node789 : 3'b010;
										assign node789 = (inp[4]) ? 3'b110 : 3'b111;
							assign node793 = (inp[8]) ? node807 : node794;
								assign node794 = (inp[11]) ? node800 : node795;
									assign node795 = (inp[2]) ? 3'b100 : node796;
										assign node796 = (inp[4]) ? 3'b010 : 3'b000;
									assign node800 = (inp[2]) ? 3'b000 : node801;
										assign node801 = (inp[4]) ? node803 : 3'b100;
											assign node803 = (inp[3]) ? 3'b000 : 3'b100;
								assign node807 = (inp[4]) ? node823 : node808;
									assign node808 = (inp[3]) ? 3'b100 : node809;
										assign node809 = (inp[5]) ? node815 : node810;
											assign node810 = (inp[11]) ? node812 : 3'b010;
												assign node812 = (inp[2]) ? 3'b100 : 3'b010;
											assign node815 = (inp[11]) ? node819 : node816;
												assign node816 = (inp[2]) ? 3'b010 : 3'b100;
												assign node819 = (inp[2]) ? 3'b100 : 3'b010;
									assign node823 = (inp[2]) ? node829 : node824;
										assign node824 = (inp[5]) ? node826 : 3'b010;
											assign node826 = (inp[11]) ? 3'b010 : 3'b110;
										assign node829 = (inp[5]) ? 3'b010 : 3'b100;
				assign node832 = (inp[7]) ? node852 : node833;
					assign node833 = (inp[8]) ? node835 : 3'b000;
						assign node835 = (inp[1]) ? 3'b000 : node836;
							assign node836 = (inp[10]) ? 3'b000 : node837;
								assign node837 = (inp[11]) ? node847 : node838;
									assign node838 = (inp[4]) ? node842 : node839;
										assign node839 = (inp[3]) ? 3'b100 : 3'b010;
										assign node842 = (inp[2]) ? node844 : 3'b100;
											assign node844 = (inp[3]) ? 3'b000 : 3'b100;
									assign node847 = (inp[4]) ? 3'b000 : 3'b010;
					assign node852 = (inp[10]) ? node896 : node853;
						assign node853 = (inp[1]) ? node877 : node854;
							assign node854 = (inp[8]) ? node866 : node855;
								assign node855 = (inp[4]) ? node857 : 3'b010;
									assign node857 = (inp[2]) ? node861 : node858;
										assign node858 = (inp[5]) ? 3'b100 : 3'b010;
										assign node861 = (inp[11]) ? 3'b000 : node862;
											assign node862 = (inp[3]) ? 3'b000 : 3'b100;
								assign node866 = (inp[2]) ? node872 : node867;
									assign node867 = (inp[4]) ? node869 : 3'b110;
										assign node869 = (inp[11]) ? 3'b010 : 3'b110;
									assign node872 = (inp[11]) ? 3'b100 : node873;
										assign node873 = (inp[4]) ? 3'b010 : 3'b110;
							assign node877 = (inp[8]) ? node885 : node878;
								assign node878 = (inp[2]) ? node882 : node879;
									assign node879 = (inp[11]) ? 3'b000 : 3'b100;
									assign node882 = (inp[11]) ? 3'b100 : 3'b000;
								assign node885 = (inp[11]) ? node893 : node886;
									assign node886 = (inp[2]) ? node890 : node887;
										assign node887 = (inp[4]) ? 3'b010 : 3'b000;
										assign node890 = (inp[4]) ? 3'b100 : 3'b110;
									assign node893 = (inp[2]) ? 3'b000 : 3'b100;
						assign node896 = (inp[1]) ? 3'b000 : node897;
							assign node897 = (inp[8]) ? node899 : 3'b000;
								assign node899 = (inp[11]) ? node907 : node900;
									assign node900 = (inp[2]) ? 3'b100 : node901;
										assign node901 = (inp[3]) ? 3'b100 : node902;
											assign node902 = (inp[4]) ? 3'b010 : 3'b000;
									assign node907 = (inp[2]) ? 3'b000 : node908;
										assign node908 = (inp[4]) ? 3'b000 : 3'b100;

endmodule