module dtc_split125_bm78 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node35;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node192;

	assign outp = (inp[3]) ? node130 : node1;
		assign node1 = (inp[4]) ? node73 : node2;
			assign node2 = (inp[0]) ? node50 : node3;
				assign node3 = (inp[6]) ? node31 : node4;
					assign node4 = (inp[1]) ? node18 : node5;
						assign node5 = (inp[9]) ? node11 : node6;
							assign node6 = (inp[11]) ? 3'b100 : node7;
								assign node7 = (inp[8]) ? 3'b100 : 3'b000;
							assign node11 = (inp[5]) ? node15 : node12;
								assign node12 = (inp[8]) ? 3'b010 : 3'b110;
								assign node15 = (inp[2]) ? 3'b010 : 3'b000;
						assign node18 = (inp[9]) ? node24 : node19;
							assign node19 = (inp[2]) ? node21 : 3'b010;
								assign node21 = (inp[10]) ? 3'b110 : 3'b010;
							assign node24 = (inp[2]) ? node28 : node25;
								assign node25 = (inp[7]) ? 3'b100 : 3'b010;
								assign node28 = (inp[5]) ? 3'b101 : 3'b011;
					assign node31 = (inp[9]) ? node39 : node32;
						assign node32 = (inp[1]) ? 3'b011 : node33;
							assign node33 = (inp[2]) ? node35 : 3'b010;
								assign node35 = (inp[11]) ? 3'b011 : 3'b010;
						assign node39 = (inp[5]) ? node45 : node40;
							assign node40 = (inp[2]) ? 3'b111 : node41;
								assign node41 = (inp[10]) ? 3'b111 : 3'b011;
							assign node45 = (inp[1]) ? 3'b011 : node46;
								assign node46 = (inp[2]) ? 3'b001 : 3'b001;
				assign node50 = (inp[6]) ? 3'b111 : node51;
					assign node51 = (inp[7]) ? node67 : node52;
						assign node52 = (inp[8]) ? node60 : node53;
							assign node53 = (inp[1]) ? node57 : node54;
								assign node54 = (inp[2]) ? 3'b111 : 3'b110;
								assign node57 = (inp[5]) ? 3'b101 : 3'b111;
							assign node60 = (inp[5]) ? node64 : node61;
								assign node61 = (inp[1]) ? 3'b111 : 3'b011;
								assign node64 = (inp[9]) ? 3'b001 : 3'b010;
						assign node67 = (inp[8]) ? 3'b111 : node68;
							assign node68 = (inp[9]) ? 3'b111 : 3'b101;
			assign node73 = (inp[0]) ? node97 : node74;
				assign node74 = (inp[9]) ? node76 : 3'b000;
					assign node76 = (inp[6]) ? node90 : node77;
						assign node77 = (inp[7]) ? node83 : node78;
							assign node78 = (inp[1]) ? node80 : 3'b000;
								assign node80 = (inp[5]) ? 3'b000 : 3'b100;
							assign node83 = (inp[5]) ? node87 : node84;
								assign node84 = (inp[1]) ? 3'b010 : 3'b100;
								assign node87 = (inp[1]) ? 3'b100 : 3'b000;
						assign node90 = (inp[1]) ? node92 : 3'b000;
							assign node92 = (inp[11]) ? 3'b001 : node93;
								assign node93 = (inp[7]) ? 3'b001 : 3'b000;
				assign node97 = (inp[9]) ? node109 : node98;
					assign node98 = (inp[6]) ? 3'b000 : node99;
						assign node99 = (inp[7]) ? 3'b110 : node100;
							assign node100 = (inp[5]) ? node104 : node101;
								assign node101 = (inp[8]) ? 3'b001 : 3'b100;
								assign node104 = (inp[1]) ? 3'b010 : 3'b000;
					assign node109 = (inp[6]) ? node125 : node110;
						assign node110 = (inp[1]) ? node118 : node111;
							assign node111 = (inp[7]) ? node115 : node112;
								assign node112 = (inp[10]) ? 3'b000 : 3'b110;
								assign node115 = (inp[11]) ? 3'b010 : 3'b101;
							assign node118 = (inp[5]) ? node122 : node119;
								assign node119 = (inp[7]) ? 3'b111 : 3'b101;
								assign node122 = (inp[11]) ? 3'b011 : 3'b001;
						assign node125 = (inp[1]) ? 3'b111 : node126;
							assign node126 = (inp[7]) ? 3'b111 : 3'b011;
		assign node130 = (inp[0]) ? node142 : node131;
			assign node131 = (inp[2]) ? 3'b000 : node132;
				assign node132 = (inp[9]) ? node134 : 3'b000;
					assign node134 = (inp[8]) ? node136 : 3'b000;
						assign node136 = (inp[11]) ? node138 : 3'b000;
							assign node138 = (inp[6]) ? 3'b000 : 3'b100;
			assign node142 = (inp[4]) ? node176 : node143;
				assign node143 = (inp[7]) ? node165 : node144;
					assign node144 = (inp[9]) ? node152 : node145;
						assign node145 = (inp[1]) ? node147 : 3'b000;
							assign node147 = (inp[11]) ? 3'b000 : node148;
								assign node148 = (inp[8]) ? 3'b100 : 3'b000;
						assign node152 = (inp[6]) ? node160 : node153;
							assign node153 = (inp[11]) ? node157 : node154;
								assign node154 = (inp[10]) ? 3'b000 : 3'b000;
								assign node157 = (inp[2]) ? 3'b100 : 3'b000;
							assign node160 = (inp[1]) ? 3'b001 : node161;
								assign node161 = (inp[10]) ? 3'b011 : 3'b010;
					assign node165 = (inp[6]) ? node173 : node166;
						assign node166 = (inp[9]) ? node168 : 3'b100;
							assign node168 = (inp[1]) ? 3'b010 : node169;
								assign node169 = (inp[5]) ? 3'b000 : 3'b100;
						assign node173 = (inp[9]) ? 3'b101 : 3'b000;
				assign node176 = (inp[9]) ? node178 : 3'b000;
					assign node178 = (inp[11]) ? node186 : node179;
						assign node179 = (inp[2]) ? node181 : 3'b000;
							assign node181 = (inp[7]) ? node183 : 3'b000;
								assign node183 = (inp[5]) ? 3'b010 : 3'b000;
						assign node186 = (inp[1]) ? node188 : 3'b000;
							assign node188 = (inp[6]) ? node192 : node189;
								assign node189 = (inp[2]) ? 3'b100 : 3'b000;
								assign node192 = (inp[7]) ? 3'b010 : 3'b000;

endmodule