module dtc_split05_bm41 (
	input  wire [5-1:0] inp,
	output wire [3-1:0] outp
);



endmodule