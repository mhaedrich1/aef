module dtc_split125_bm45 (
	input  wire [16-1:0] inp,
	output wire [46-1:0] outp
);

	wire [46-1:0] node1;
	wire [46-1:0] node2;
	wire [46-1:0] node4;
	wire [46-1:0] node6;
	wire [46-1:0] node8;
	wire [46-1:0] node9;
	wire [46-1:0] node11;
	wire [46-1:0] node13;
	wire [46-1:0] node15;
	wire [46-1:0] node17;
	wire [46-1:0] node19;
	wire [46-1:0] node23;
	wire [46-1:0] node25;
	wire [46-1:0] node26;
	wire [46-1:0] node27;
	wire [46-1:0] node28;
	wire [46-1:0] node29;
	wire [46-1:0] node32;
	wire [46-1:0] node35;
	wire [46-1:0] node36;
	wire [46-1:0] node39;
	wire [46-1:0] node42;
	wire [46-1:0] node43;
	wire [46-1:0] node45;
	wire [46-1:0] node47;
	wire [46-1:0] node49;
	wire [46-1:0] node51;
	wire [46-1:0] node52;
	wire [46-1:0] node55;
	wire [46-1:0] node58;
	wire [46-1:0] node59;
	wire [46-1:0] node62;
	wire [46-1:0] node64;
	wire [46-1:0] node66;
	wire [46-1:0] node67;
	wire [46-1:0] node68;
	wire [46-1:0] node73;
	wire [46-1:0] node74;
	wire [46-1:0] node76;
	wire [46-1:0] node78;
	wire [46-1:0] node80;
	wire [46-1:0] node81;
	wire [46-1:0] node83;
	wire [46-1:0] node87;
	wire [46-1:0] node89;
	wire [46-1:0] node90;
	wire [46-1:0] node93;
	wire [46-1:0] node95;
	wire [46-1:0] node96;
	wire [46-1:0] node97;
	wire [46-1:0] node99;
	wire [46-1:0] node101;
	wire [46-1:0] node104;
	wire [46-1:0] node108;
	wire [46-1:0] node109;
	wire [46-1:0] node110;
	wire [46-1:0] node113;
	wire [46-1:0] node114;
	wire [46-1:0] node115;
	wire [46-1:0] node116;
	wire [46-1:0] node117;
	wire [46-1:0] node120;
	wire [46-1:0] node123;
	wire [46-1:0] node124;
	wire [46-1:0] node127;
	wire [46-1:0] node130;
	wire [46-1:0] node131;
	wire [46-1:0] node132;
	wire [46-1:0] node135;
	wire [46-1:0] node138;
	wire [46-1:0] node139;
	wire [46-1:0] node142;
	wire [46-1:0] node145;
	wire [46-1:0] node146;
	wire [46-1:0] node147;
	wire [46-1:0] node148;
	wire [46-1:0] node151;
	wire [46-1:0] node154;
	wire [46-1:0] node155;
	wire [46-1:0] node158;
	wire [46-1:0] node161;
	wire [46-1:0] node162;
	wire [46-1:0] node163;
	wire [46-1:0] node166;
	wire [46-1:0] node169;
	wire [46-1:0] node170;
	wire [46-1:0] node173;
	wire [46-1:0] node176;
	wire [46-1:0] node177;
	wire [46-1:0] node180;
	wire [46-1:0] node182;
	wire [46-1:0] node183;
	wire [46-1:0] node184;
	wire [46-1:0] node185;
	wire [46-1:0] node186;
	wire [46-1:0] node187;
	wire [46-1:0] node188;
	wire [46-1:0] node189;
	wire [46-1:0] node190;
	wire [46-1:0] node194;
	wire [46-1:0] node195;
	wire [46-1:0] node198;
	wire [46-1:0] node199;
	wire [46-1:0] node203;
	wire [46-1:0] node204;
	wire [46-1:0] node205;
	wire [46-1:0] node208;
	wire [46-1:0] node211;
	wire [46-1:0] node214;
	wire [46-1:0] node215;
	wire [46-1:0] node217;
	wire [46-1:0] node220;
	wire [46-1:0] node221;
	wire [46-1:0] node223;
	wire [46-1:0] node226;
	wire [46-1:0] node229;
	wire [46-1:0] node230;
	wire [46-1:0] node231;
	wire [46-1:0] node232;
	wire [46-1:0] node233;
	wire [46-1:0] node237;
	wire [46-1:0] node239;
	wire [46-1:0] node242;
	wire [46-1:0] node243;
	wire [46-1:0] node244;
	wire [46-1:0] node247;
	wire [46-1:0] node250;
	wire [46-1:0] node252;
	wire [46-1:0] node255;
	wire [46-1:0] node256;
	wire [46-1:0] node257;
	wire [46-1:0] node258;
	wire [46-1:0] node259;
	wire [46-1:0] node264;
	wire [46-1:0] node265;
	wire [46-1:0] node269;
	wire [46-1:0] node270;
	wire [46-1:0] node271;
	wire [46-1:0] node276;
	wire [46-1:0] node277;
	wire [46-1:0] node279;
	wire [46-1:0] node280;
	wire [46-1:0] node281;
	wire [46-1:0] node282;
	wire [46-1:0] node286;
	wire [46-1:0] node291;
	wire [46-1:0] node292;
	wire [46-1:0] node293;
	wire [46-1:0] node295;
	wire [46-1:0] node296;
	wire [46-1:0] node298;
	wire [46-1:0] node300;
	wire [46-1:0] node302;
	wire [46-1:0] node303;
	wire [46-1:0] node307;
	wire [46-1:0] node308;
	wire [46-1:0] node310;
	wire [46-1:0] node314;
	wire [46-1:0] node315;
	wire [46-1:0] node316;
	wire [46-1:0] node317;
	wire [46-1:0] node320;
	wire [46-1:0] node321;
	wire [46-1:0] node324;
	wire [46-1:0] node327;
	wire [46-1:0] node328;
	wire [46-1:0] node329;
	wire [46-1:0] node333;
	wire [46-1:0] node335;
	wire [46-1:0] node338;
	wire [46-1:0] node339;
	wire [46-1:0] node341;
	wire [46-1:0] node342;
	wire [46-1:0] node345;
	wire [46-1:0] node348;
	wire [46-1:0] node349;
	wire [46-1:0] node351;
	wire [46-1:0] node352;
	wire [46-1:0] node356;
	wire [46-1:0] node357;
	wire [46-1:0] node358;
	wire [46-1:0] node362;
	wire [46-1:0] node365;
	wire [46-1:0] node366;
	wire [46-1:0] node367;
	wire [46-1:0] node368;
	wire [46-1:0] node369;
	wire [46-1:0] node371;
	wire [46-1:0] node374;
	wire [46-1:0] node377;
	wire [46-1:0] node378;
	wire [46-1:0] node379;
	wire [46-1:0] node381;
	wire [46-1:0] node384;
	wire [46-1:0] node387;
	wire [46-1:0] node388;
	wire [46-1:0] node392;
	wire [46-1:0] node393;
	wire [46-1:0] node394;
	wire [46-1:0] node395;
	wire [46-1:0] node397;
	wire [46-1:0] node401;
	wire [46-1:0] node402;
	wire [46-1:0] node403;
	wire [46-1:0] node404;
	wire [46-1:0] node407;
	wire [46-1:0] node410;
	wire [46-1:0] node414;
	wire [46-1:0] node415;
	wire [46-1:0] node416;
	wire [46-1:0] node419;
	wire [46-1:0] node422;
	wire [46-1:0] node425;
	wire [46-1:0] node426;
	wire [46-1:0] node427;
	wire [46-1:0] node428;
	wire [46-1:0] node432;
	wire [46-1:0] node433;
	wire [46-1:0] node435;
	wire [46-1:0] node436;
	wire [46-1:0] node440;
	wire [46-1:0] node442;
	wire [46-1:0] node445;
	wire [46-1:0] node446;
	wire [46-1:0] node447;
	wire [46-1:0] node448;
	wire [46-1:0] node452;
	wire [46-1:0] node453;
	wire [46-1:0] node456;
	wire [46-1:0] node459;
	wire [46-1:0] node460;
	wire [46-1:0] node461;
	wire [46-1:0] node463;
	wire [46-1:0] node467;
	wire [46-1:0] node469;
	wire [46-1:0] node470;
	wire [46-1:0] node472;
	wire [46-1:0] node476;
	wire [46-1:0] node477;
	wire [46-1:0] node478;
	wire [46-1:0] node479;
	wire [46-1:0] node481;
	wire [46-1:0] node483;
	wire [46-1:0] node485;
	wire [46-1:0] node488;
	wire [46-1:0] node489;
	wire [46-1:0] node491;
	wire [46-1:0] node492;
	wire [46-1:0] node495;
	wire [46-1:0] node498;
	wire [46-1:0] node499;
	wire [46-1:0] node501;
	wire [46-1:0] node503;
	wire [46-1:0] node504;
	wire [46-1:0] node506;
	wire [46-1:0] node507;
	wire [46-1:0] node511;
	wire [46-1:0] node512;
	wire [46-1:0] node516;
	wire [46-1:0] node517;
	wire [46-1:0] node518;
	wire [46-1:0] node519;
	wire [46-1:0] node523;
	wire [46-1:0] node526;
	wire [46-1:0] node527;
	wire [46-1:0] node528;
	wire [46-1:0] node530;
	wire [46-1:0] node533;
	wire [46-1:0] node537;
	wire [46-1:0] node538;
	wire [46-1:0] node539;
	wire [46-1:0] node540;
	wire [46-1:0] node541;
	wire [46-1:0] node542;
	wire [46-1:0] node546;
	wire [46-1:0] node547;
	wire [46-1:0] node549;
	wire [46-1:0] node552;
	wire [46-1:0] node555;
	wire [46-1:0] node557;
	wire [46-1:0] node558;
	wire [46-1:0] node559;
	wire [46-1:0] node560;
	wire [46-1:0] node564;
	wire [46-1:0] node567;
	wire [46-1:0] node570;
	wire [46-1:0] node571;
	wire [46-1:0] node572;
	wire [46-1:0] node575;
	wire [46-1:0] node576;
	wire [46-1:0] node579;
	wire [46-1:0] node581;
	wire [46-1:0] node584;
	wire [46-1:0] node585;
	wire [46-1:0] node586;
	wire [46-1:0] node587;
	wire [46-1:0] node592;
	wire [46-1:0] node593;
	wire [46-1:0] node595;
	wire [46-1:0] node598;
	wire [46-1:0] node601;
	wire [46-1:0] node602;
	wire [46-1:0] node603;
	wire [46-1:0] node604;
	wire [46-1:0] node605;
	wire [46-1:0] node609;
	wire [46-1:0] node610;
	wire [46-1:0] node613;
	wire [46-1:0] node615;
	wire [46-1:0] node618;
	wire [46-1:0] node619;
	wire [46-1:0] node622;
	wire [46-1:0] node624;
	wire [46-1:0] node627;
	wire [46-1:0] node628;
	wire [46-1:0] node629;
	wire [46-1:0] node630;
	wire [46-1:0] node634;
	wire [46-1:0] node635;
	wire [46-1:0] node636;
	wire [46-1:0] node637;
	wire [46-1:0] node642;
	wire [46-1:0] node645;
	wire [46-1:0] node646;
	wire [46-1:0] node647;
	wire [46-1:0] node650;
	wire [46-1:0] node653;
	wire [46-1:0] node655;
	wire [46-1:0] node658;
	wire [46-1:0] node659;
	wire [46-1:0] node660;
	wire [46-1:0] node661;
	wire [46-1:0] node663;
	wire [46-1:0] node664;
	wire [46-1:0] node667;
	wire [46-1:0] node670;
	wire [46-1:0] node671;
	wire [46-1:0] node672;
	wire [46-1:0] node675;
	wire [46-1:0] node679;
	wire [46-1:0] node680;
	wire [46-1:0] node682;
	wire [46-1:0] node683;
	wire [46-1:0] node686;
	wire [46-1:0] node689;
	wire [46-1:0] node690;
	wire [46-1:0] node691;
	wire [46-1:0] node694;
	wire [46-1:0] node698;
	wire [46-1:0] node699;
	wire [46-1:0] node700;
	wire [46-1:0] node702;
	wire [46-1:0] node703;
	wire [46-1:0] node706;
	wire [46-1:0] node709;
	wire [46-1:0] node710;
	wire [46-1:0] node711;

	assign outp = (inp[1]) ? node108 : node1;
		assign node1 = (inp[15]) ? node23 : node2;
			assign node2 = (inp[11]) ? node4 : 46'b0000000000000000000000000000000000000000000000;
				assign node4 = (inp[12]) ? node6 : 46'b0000000000000000000000000000000000000000000000;
					assign node6 = (inp[4]) ? node8 : 46'b0000000000000000000000000000000000000000000000;
						assign node8 = (inp[13]) ? 46'b0000000000000000000000000000000000000000000000 : node9;
							assign node9 = (inp[5]) ? node11 : 46'b0000000000000000000000000000000000000000000000;
								assign node11 = (inp[8]) ? node13 : 46'b0000000000000000000000000000000000000000000000;
									assign node13 = (inp[6]) ? node15 : 46'b0000000000000000000000000000000000000000000000;
										assign node15 = (inp[7]) ? node17 : 46'b0000000000000000000000000000000000000000000000;
											assign node17 = (inp[9]) ? node19 : 46'b0000000000000000000000000000000000000000000000;
												assign node19 = (inp[3]) ? 46'b0000000000000000100000000000000000000000000000 : 46'b0000000000000000000000000000000000000000000000;
			assign node23 = (inp[3]) ? node25 : 46'b0000000000000000000000000000001000000000000000;
				assign node25 = (inp[2]) ? node73 : node26;
					assign node26 = (inp[13]) ? node42 : node27;
						assign node27 = (inp[11]) ? node35 : node28;
							assign node28 = (inp[0]) ? node32 : node29;
								assign node29 = (inp[9]) ? 46'b0000000100001000000000000000000000000000000000 : 46'b0000001000001000000000000000000000000000000000;
								assign node32 = (inp[9]) ? 46'b0010001000000000000000000000000000000000010000 : 46'b0000000000001000000000000010000000000000000000;
							assign node35 = (inp[0]) ? node39 : node36;
								assign node36 = (inp[9]) ? 46'b0000010100000000000000000000000000000000000000 : 46'b0000011000000000000000000000000000000000000000;
								assign node39 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000010000000000000000000010000000000000000000;
						assign node42 = (inp[11]) ? node58 : node43;
							assign node43 = (inp[5]) ? node45 : 46'b0000000000000000000000000000000000000000000000;
								assign node45 = (inp[14]) ? node47 : 46'b0000000000000000000000000000000000000000000000;
									assign node47 = (inp[10]) ? node49 : 46'b0000000000000000000000000000000000000000000000;
										assign node49 = (inp[6]) ? node51 : 46'b0000000000000000000000000000000000000000000000;
											assign node51 = (inp[12]) ? node55 : node52;
												assign node52 = (inp[4]) ? 46'b0000000000011000010000000000000000000000010000 : 46'b0000000000000000000000000000000000000000000000;
												assign node55 = (inp[8]) ? 46'b0000010000000000010000010000000000000000010100 : 46'b0000010000010000010000000000000000000000010100;
							assign node58 = (inp[9]) ? node62 : node59;
								assign node59 = (inp[0]) ? 46'b0000001000000000011000000100000000000000010000 : 46'b0000001000000000010000000100000000000000010010;
								assign node62 = (inp[6]) ? node64 : 46'b0000000000000000000000000000000000000000000000;
									assign node64 = (inp[4]) ? node66 : 46'b0000000000000000000000000000000000000000000000;
										assign node66 = (inp[10]) ? 46'b0000000000000000000000000000000000000000000000 : node67;
											assign node67 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node68;
												assign node68 = (inp[8]) ? 46'b0000010000000000011000000100000100000000010000 : 46'b0000000000000000000000000000000000000000000000;
					assign node73 = (inp[11]) ? node87 : node74;
						assign node74 = (inp[6]) ? node76 : 46'b0000000000000000000000000000000000000000000000;
							assign node76 = (inp[10]) ? node78 : 46'b0000000000000000000000000000000000000000000000;
								assign node78 = (inp[5]) ? node80 : 46'b0000000000000000000000000000000000000000000000;
									assign node80 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node81;
										assign node81 = (inp[9]) ? node83 : 46'b0000000000000000000000000000000000000000000000;
											assign node83 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0010000000010000000000000000000000000010000000;
						assign node87 = (inp[13]) ? node89 : 46'b0000000000000000000000000000000000000000000000;
							assign node89 = (inp[9]) ? node93 : node90;
								assign node90 = (inp[0]) ? 46'b0000001000000000010010000000010000000010000000 : 46'b0000001000000000010010100000000000000010000000;
								assign node93 = (inp[14]) ? node95 : 46'b0000000000000000000000000000000000000000000000;
									assign node95 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : node96;
										assign node96 = (inp[10]) ? node104 : node97;
											assign node97 = (inp[7]) ? node99 : 46'b0000000000000000000000000000000000000000000000;
												assign node99 = (inp[4]) ? node101 : 46'b0000000000000000000000000000000000000000000000;
													assign node101 = (inp[0]) ? 46'b0000000000001000010010000000010100000010000000 : 46'b0000000000000000000000000000000000000000000000;
											assign node104 = (inp[8]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0010000000010000000010100000000000000010000000;
		assign node108 = (inp[15]) ? node176 : node109;
			assign node109 = (inp[13]) ? node113 : node110;
				assign node110 = (inp[3]) ? 46'b0000100000000000000000000000001000000000000000 : 46'b0000100000000000000000000000000000000000000000;
				assign node113 = (inp[2]) ? node145 : node114;
					assign node114 = (inp[9]) ? node130 : node115;
						assign node115 = (inp[0]) ? node123 : node116;
							assign node116 = (inp[11]) ? node120 : node117;
								assign node117 = (inp[3]) ? 46'b0000100000001000010000010100001000000000010010 : 46'b0000100000001000010000010100000000000000010010;
								assign node120 = (inp[3]) ? 46'b0000100000001000011000010100001000000000010000 : 46'b0000100000001000011000010100000000000000010000;
							assign node123 = (inp[11]) ? node127 : node124;
								assign node124 = (inp[3]) ? 46'b0000100000001000010000000100001100000000010010 : 46'b0000100000001000010000000100000100000000010010;
								assign node127 = (inp[3]) ? 46'b0000100000001000011000000100001100000000010000 : 46'b0000100000001000011000000100000100000000010000;
						assign node130 = (inp[0]) ? node138 : node131;
							assign node131 = (inp[11]) ? node135 : node132;
								assign node132 = (inp[3]) ? 46'b0000110000000000010000010100001000000000010010 : 46'b0000110000000000010000010100000000000000010010;
								assign node135 = (inp[3]) ? 46'b0000110000000000011000010100001000000000010000 : 46'b0000110000000000011000010100000000000000010000;
							assign node138 = (inp[11]) ? node142 : node139;
								assign node139 = (inp[3]) ? 46'b0000110000000000010000000100001100000000010010 : 46'b0000110000000000010000000100000100000000010010;
								assign node142 = (inp[3]) ? 46'b0000110000000000011000000100001100000000010000 : 46'b0000110000000000011000000100000100000000010000;
					assign node145 = (inp[11]) ? node161 : node146;
						assign node146 = (inp[0]) ? node154 : node147;
							assign node147 = (inp[9]) ? node151 : node148;
								assign node148 = (inp[3]) ? 46'b0000100000001000010010110000001000000010000000 : 46'b0000100000001000010010110000000000000010000000;
								assign node151 = (inp[3]) ? 46'b0000110000000000010010110000001000000010000000 : 46'b0000110000000000010010110000000000000010000000;
							assign node154 = (inp[9]) ? node158 : node155;
								assign node155 = (inp[3]) ? 46'b0000100000001000010010100000001100000010000000 : 46'b0000100000001000010010100000000100000010000000;
								assign node158 = (inp[3]) ? 46'b0000110000000000010010100000001100000010000000 : 46'b0000110000000000010010100000000100000010000000;
						assign node161 = (inp[9]) ? node169 : node162;
							assign node162 = (inp[0]) ? node166 : node163;
								assign node163 = (inp[3]) ? 46'b0000100000001000010010010000011000000010000000 : 46'b0000100000001000010010010000010000000010000000;
								assign node166 = (inp[3]) ? 46'b0000100000001000010010000000011100000010000000 : 46'b0000100000001000010010000000010100000010000000;
							assign node169 = (inp[0]) ? node173 : node170;
								assign node170 = (inp[3]) ? 46'b0000110000000000010010010000011000000010000000 : 46'b0000110000000000010010010000010000000010000000;
								assign node173 = (inp[3]) ? 46'b0000110000000000010010000000011100000010000000 : 46'b0000110000000000010010000000010100000010000000;
			assign node176 = (inp[3]) ? node180 : node177;
				assign node177 = (inp[13]) ? 46'b0000000000000000000000000000001000000000000000 : 46'b0000000000000000000000000000001000000000001000;
				assign node180 = (inp[13]) ? node182 : 46'b0000000000000000000000000000000000000000001000;
					assign node182 = (inp[2]) ? node476 : node183;
						assign node183 = (inp[11]) ? node291 : node184;
							assign node184 = (inp[9]) ? node276 : node185;
								assign node185 = (inp[12]) ? node229 : node186;
									assign node186 = (inp[7]) ? node214 : node187;
										assign node187 = (inp[4]) ? node203 : node188;
											assign node188 = (inp[10]) ? node194 : node189;
												assign node189 = (inp[6]) ? 46'b0011000000000100000000010000100010010000010000 : node190;
													assign node190 = (inp[14]) ? 46'b0011000000000110000000010000100010110000010000 : 46'b0011000000000100000000010001100010110000010010;
												assign node194 = (inp[6]) ? node198 : node195;
													assign node195 = (inp[14]) ? 46'b0011000000000000001000010001100010110000010010 : 46'b0011000000000100000000010001100010110001010010;
													assign node198 = (inp[14]) ? 46'b0011000000000010000000010001100010010000010010 : node199;
														assign node199 = (inp[8]) ? 46'b0011000000000000000000010001100010010001010010 : 46'b0011000000000100000000010001100010010000010010;
											assign node203 = (inp[14]) ? node211 : node204;
												assign node204 = (inp[0]) ? node208 : node205;
													assign node205 = (inp[6]) ? 46'b0010000000000010000000010001100010010001010010 : 46'b0011000000000010000000010001100010110001010010;
													assign node208 = (inp[5]) ? 46'b0010000000000010000000010001100010110000010010 : 46'b0011000000000010000000010001100010010000010010;
												assign node211 = (inp[0]) ? 46'b0011000000000010001000010001100010010000010000 : 46'b0011000000000010001000010001100010010001010000;
										assign node214 = (inp[0]) ? node220 : node215;
											assign node215 = (inp[6]) ? node217 : 46'b0011000000000010000000010001000010110001010010;
												assign node217 = (inp[4]) ? 46'b0010000000000100001000010001000010010001010000 : 46'b0010000000000000001000010001000010010001010010;
											assign node220 = (inp[10]) ? node226 : node221;
												assign node221 = (inp[14]) ? node223 : 46'b0010000000000100000000010000000010010000010000;
													assign node223 = (inp[6]) ? 46'b0010000000000110000000010000000010010000010000 : 46'b0010000000000110000000010000000010110000010000;
												assign node226 = (inp[14]) ? 46'b0011000000000010000000010000000010110000010000 : 46'b0011000000000100000000010001000010110000010010;
									assign node229 = (inp[0]) ? node255 : node230;
										assign node230 = (inp[6]) ? node242 : node231;
											assign node231 = (inp[14]) ? node237 : node232;
												assign node232 = (inp[4]) ? 46'b0010000000000100001000010001100000110001010000 : node233;
													assign node233 = (inp[10]) ? 46'b0011000000000100000000010001000000110001010010 : 46'b0010000000000100000000010000000000110001010000;
												assign node237 = (inp[4]) ? node239 : 46'b0011000000000110000000010000100000110001010000;
													assign node239 = (inp[10]) ? 46'b0011000000000010001000010001100000110001010000 : 46'b0011000000000010001000010001000000110001010000;
											assign node242 = (inp[10]) ? node250 : node243;
												assign node243 = (inp[8]) ? node247 : node244;
													assign node244 = (inp[7]) ? 46'b0011000000000100001000010001000000010001010000 : 46'b0010000000000100001000010001100000010001010000;
													assign node247 = (inp[14]) ? 46'b0010000000000110000000010000100000010001010000 : 46'b0010000000000100000000010001100000010001010010;
												assign node250 = (inp[14]) ? node252 : 46'b0010000000000010000000010001000000010001010010;
													assign node252 = (inp[4]) ? 46'b0010000000000010001000010001000000010001010000 : 46'b0010000000000000001000010001000000010001010010;
										assign node255 = (inp[8]) ? node269 : node256;
											assign node256 = (inp[7]) ? node264 : node257;
												assign node257 = (inp[10]) ? 46'b0011000000000010001000010001100000010000010000 : node258;
													assign node258 = (inp[6]) ? 46'b0011000000000100001000010001100000010000010000 : node259;
														assign node259 = (inp[14]) ? 46'b0011000000000000001000010001100000110000010000 : 46'b0011000000000100001000010001100000110000010000;
												assign node264 = (inp[6]) ? 46'b0010000000000000001000010001000000010000010000 : node265;
													assign node265 = (inp[5]) ? 46'b0010000000000100001000010001000000110000010000 : 46'b0011000000000100001000010001000000110000010000;
											assign node269 = (inp[14]) ? 46'b0010000000000110000000010000000000110000010000 : node270;
												assign node270 = (inp[4]) ? 46'b0010000000000000001000010001100000110000010010 : node271;
													assign node271 = (inp[5]) ? 46'b0010000000000100000000010001100000110000010010 : 46'b0011000000000100000000010001100000110000010010;
								assign node276 = (inp[0]) ? 46'b0000000000000000000000000000000000000000000000 : node277;
									assign node277 = (inp[5]) ? node279 : 46'b0000000000000000000000000000000000000000000000;
										assign node279 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node280;
											assign node280 = (inp[8]) ? node286 : node281;
												assign node281 = (inp[4]) ? 46'b0000000000000000000000000000000000000000000000 : node282;
													assign node282 = (inp[10]) ? 46'b0000000000000000001000001001100000000000000010 : 46'b0000000000000000000000000000000000000000000000;
												assign node286 = (inp[6]) ? 46'b0000000000000000000000001001100010000000000010 : 46'b0000000000000000000000001001100000100000000010;
							assign node291 = (inp[0]) ? node365 : node292;
								assign node292 = (inp[9]) ? node314 : node293;
									assign node293 = (inp[7]) ? node295 : 46'b0000000000000000000000000000000000000000000000;
										assign node295 = (inp[12]) ? node307 : node296;
											assign node296 = (inp[6]) ? node298 : 46'b0000000000000000000000000000000000000000000000;
												assign node298 = (inp[4]) ? node300 : 46'b0000000000000000000000000000000000000000000000;
													assign node300 = (inp[14]) ? node302 : 46'b0000000000000010000001000001000010000000000010;
														assign node302 = (inp[8]) ? 46'b0000000000000010001001000001000010000000000000 : node303;
															assign node303 = (inp[10]) ? 46'b0000000000000010001001000001000010000000000000 : 46'b0000000000000000001001000001000010000000000000;
											assign node307 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : node308;
												assign node308 = (inp[8]) ? node310 : 46'b0000000000000100001001000001000000100000000000;
													assign node310 = (inp[10]) ? 46'b0000000000000010000001000001000000100000000010 : 46'b0000000000000010001001000001000000100000000000;
									assign node314 = (inp[10]) ? node338 : node315;
										assign node315 = (inp[7]) ? node327 : node316;
											assign node316 = (inp[6]) ? node320 : node317;
												assign node317 = (inp[14]) ? 46'b1001000000000100001000000001100000100000000000 : 46'b1001000000000100000000000000100010100000000000;
												assign node320 = (inp[14]) ? node324 : node321;
													assign node321 = (inp[4]) ? 46'b1001000000000000001000000001100010000000000010 : 46'b1001000000000100000000000001100010000000000010;
													assign node324 = (inp[4]) ? 46'b1000000000000000001000000001100010000000000000 : 46'b1001000000000100001000000001100010000000000000;
											assign node327 = (inp[12]) ? node333 : node328;
												assign node328 = (inp[5]) ? 46'b1000000000000100001000000001000010100000000000 : node329;
													assign node329 = (inp[8]) ? 46'b1001000000000010001000000001000010100000000000 : 46'b1001000000000000001000000001000010100000000000;
												assign node333 = (inp[4]) ? node335 : 46'b1001000000000100000000000001000000100000000010;
													assign node335 = (inp[14]) ? 46'b1001000000000010001000000001000000000000000000 : 46'b1001000000000100001000000001000000000000000000;
										assign node338 = (inp[4]) ? node348 : node339;
											assign node339 = (inp[8]) ? node341 : 46'b1000000000000000001000000001000010100000000010;
												assign node341 = (inp[12]) ? node345 : node342;
													assign node342 = (inp[7]) ? 46'b1001000000000010000000000001000010000000000010 : 46'b1001000000000010000000000001100010100000000010;
													assign node345 = (inp[14]) ? 46'b1000000000000010000000000001000000100000000010 : 46'b1001000000000000000000000001000000100000000010;
											assign node348 = (inp[5]) ? node356 : node349;
												assign node349 = (inp[7]) ? node351 : 46'b1001000000000010000000000000100010100000000000;
													assign node351 = (inp[12]) ? 46'b1001000000000010000000000000000000100000000000 : node352;
														assign node352 = (inp[6]) ? 46'b1001000000000010000000000000000010000000000000 : 46'b1001000000000010000000000000000010100000000000;
												assign node356 = (inp[12]) ? node362 : node357;
													assign node357 = (inp[6]) ? 46'b1000000000000110000000000000100010000000000000 : node358;
														assign node358 = (inp[8]) ? 46'b1000000000000010000000000000100010100000000000 : 46'b1000000000000010001000000001100010100000000000;
													assign node362 = (inp[8]) ? 46'b1000000000000010000000000001100000100000000010 : 46'b1000000000000010001000000001100000000000000000;
								assign node365 = (inp[9]) ? node425 : node366;
									assign node366 = (inp[5]) ? node392 : node367;
										assign node367 = (inp[12]) ? node377 : node368;
											assign node368 = (inp[6]) ? node374 : node369;
												assign node369 = (inp[14]) ? node371 : 46'b0101000000000000001000000001000010100000000010;
													assign node371 = (inp[7]) ? 46'b0101000000000010001000000001000010100000000000 : 46'b0101000000000010001000000001100010100000000000;
												assign node374 = (inp[8]) ? 46'b0101000000000010001000000001100010000000000000 : 46'b0101000000000100001000000001100010000000000000;
											assign node377 = (inp[7]) ? node387 : node378;
												assign node378 = (inp[4]) ? node384 : node379;
													assign node379 = (inp[8]) ? node381 : 46'b0101000000000100000000000001100000100000000010;
														assign node381 = (inp[6]) ? 46'b0101000000000010000000000001100000000000000010 : 46'b0101000000000010000000000001100000100000000010;
													assign node384 = (inp[6]) ? 46'b0101000000000000001000000001100000000000000000 : 46'b0101000000000010001000000001100000100000000000;
												assign node387 = (inp[8]) ? 46'b0101000000000110000000000000000000100000000000 : node388;
													assign node388 = (inp[4]) ? 46'b0101000000000100001000000001000000100000000000 : 46'b0101000000000100000000000001000000000000000010;
										assign node392 = (inp[6]) ? node414 : node393;
											assign node393 = (inp[12]) ? node401 : node394;
												assign node394 = (inp[14]) ? 46'b0100000000000110000000000000000010100000000000 : node395;
													assign node395 = (inp[4]) ? node397 : 46'b0100000000000100000000000001000010100000000010;
														assign node397 = (inp[7]) ? 46'b0100000000000000001000000001000010100000000010 : 46'b0100000000000000001000000001100010100000000010;
												assign node401 = (inp[8]) ? 46'b0100000000000010000000000001100000100000000010 : node402;
													assign node402 = (inp[14]) ? node410 : node403;
														assign node403 = (inp[4]) ? node407 : node404;
															assign node404 = (inp[10]) ? 46'b0100000000000100000000000001100000100000000010 : 46'b0100000000000100000000000000100000100000000000;
															assign node407 = (inp[7]) ? 46'b0100000000000110000000000000000000100000000000 : 46'b0100000000000110000000000000100000100000000000;
														assign node410 = (inp[7]) ? 46'b0100000000000000001000000001000000100000000000 : 46'b0100000000000010001000000001100000100000000000;
											assign node414 = (inp[4]) ? node422 : node415;
												assign node415 = (inp[14]) ? node419 : node416;
													assign node416 = (inp[10]) ? 46'b0100000000000000000000000001000000000000000010 : 46'b0100000000000100000000000001100000000000000010;
													assign node419 = (inp[12]) ? 46'b0100000000000010000000000001000000000000000010 : 46'b0100000000000010000000000001100010000000000010;
												assign node422 = (inp[8]) ? 46'b0100000000000010000000000000000010000000000000 : 46'b0100000000000110000000000000100010000000000000;
									assign node425 = (inp[10]) ? node445 : node426;
										assign node426 = (inp[12]) ? node432 : node427;
											assign node427 = (inp[5]) ? 46'b0000000000000000001000000001000010101000000000 : node428;
												assign node428 = (inp[4]) ? 46'b0001000000000000001000000001100010101000000000 : 46'b0001000000000100001000000001100010101000000000;
											assign node432 = (inp[7]) ? node440 : node433;
												assign node433 = (inp[4]) ? node435 : 46'b0000000000000100000000000000100000101000000000;
													assign node435 = (inp[6]) ? 46'b0000000000000100001000000001100000001000000000 : node436;
														assign node436 = (inp[14]) ? 46'b0000000000000000001000000001100000101000000000 : 46'b0000000000000000001000000001100000101000000010;
												assign node440 = (inp[5]) ? node442 : 46'b0001000000000100001000000001000000101000000000;
													assign node442 = (inp[6]) ? 46'b0000000000000100001000000001000000001000000000 : 46'b0000000000000100001000000001000000101000000000;
										assign node445 = (inp[4]) ? node459 : node446;
											assign node446 = (inp[7]) ? node452 : node447;
												assign node447 = (inp[5]) ? 46'b0000000000000100000000000001100010101000000010 : node448;
													assign node448 = (inp[6]) ? 46'b0001000000000010000000000001100010001000000010 : 46'b0001000000000000000000000001100010101000000010;
												assign node452 = (inp[12]) ? node456 : node453;
													assign node453 = (inp[5]) ? 46'b0000000000000100000000000001000010001000000010 : 46'b0001000000000100000000000001000010001000000010;
													assign node456 = (inp[5]) ? 46'b0000000000000000000000000001000000001000000010 : 46'b0001000000000010000000000001000000001000000010;
											assign node459 = (inp[12]) ? node467 : node460;
												assign node460 = (inp[5]) ? 46'b0000000000000110000000000000100010001000000000 : node461;
													assign node461 = (inp[7]) ? node463 : 46'b0001000000000010000000000000100010101000000000;
														assign node463 = (inp[6]) ? 46'b0001000000000010000000000000000010001000000000 : 46'b0001000000000110000000000000000010101000000000;
												assign node467 = (inp[6]) ? node469 : 46'b0001000000000010000000000001000000101000000010;
													assign node469 = (inp[5]) ? 46'b0000000000000010001000000001100000001000000000 : node470;
														assign node470 = (inp[14]) ? node472 : 46'b0001000000000110000000000000100000001000000000;
															assign node472 = (inp[8]) ? 46'b0001000000000010000000000000000000001000000000 : 46'b0001000000000010001000000001000000001000000000;
						assign node476 = (inp[11]) ? node658 : node477;
							assign node477 = (inp[9]) ? node537 : node478;
								assign node478 = (inp[7]) ? node488 : node479;
									assign node479 = (inp[0]) ? node481 : 46'b0000000000000000000000000000000000000000000000;
										assign node481 = (inp[14]) ? node483 : 46'b0000000000000000000000000000000000000000000000;
											assign node483 = (inp[5]) ? node485 : 46'b0000000000000000000000000000000000000000000000;
												assign node485 = (inp[10]) ? 46'b0000000000000011000000000000100000000000100000 : 46'b0000000000000001001000000001100000000000100000;
									assign node488 = (inp[0]) ? node498 : node489;
										assign node489 = (inp[5]) ? node491 : 46'b0000000000000000000000000000000000000000000000;
											assign node491 = (inp[8]) ? node495 : node492;
												assign node492 = (inp[4]) ? 46'b0000000000100110000001000000000010000000000000 : 46'b0000000000100100000001000001000010000000000010;
												assign node495 = (inp[14]) ? 46'b0000000000100010000001000001000000000000000010 : 46'b0000000000100000001001000001000000100000000010;
										assign node498 = (inp[6]) ? node516 : node499;
											assign node499 = (inp[12]) ? node501 : 46'b0000000000000000000000000000000000000000000000;
												assign node501 = (inp[5]) ? node503 : 46'b0000000000000000000000000000000000000000000000;
													assign node503 = (inp[14]) ? node511 : node504;
														assign node504 = (inp[8]) ? node506 : 46'b0000000000000111000000000000000000100000100000;
															assign node506 = (inp[4]) ? 46'b0000000000000001001000000001000000100000100010 : node507;
																assign node507 = (inp[10]) ? 46'b0000000000000001000000000001000000100000100010 : 46'b0000000000000101000000000001000000100000100010;
														assign node511 = (inp[8]) ? 46'b0000000000000111000000000000000000100000100000 : node512;
															assign node512 = (inp[4]) ? 46'b0000000000000011001000000001000000100000100000 : 46'b0000000000000101001000000001000000100000100000;
											assign node516 = (inp[10]) ? node526 : node517;
												assign node517 = (inp[5]) ? node523 : node518;
													assign node518 = (inp[14]) ? 46'b0001000000000111000000000000000000000000100000 : node519;
														assign node519 = (inp[8]) ? 46'b0001000000000101000000000001000000000000100010 : 46'b0001000000000101000000000000000000000000100000;
													assign node523 = (inp[12]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0000000000000111000000000000000010000000100000;
												assign node526 = (inp[14]) ? 46'b0000000000000000000000000000000000000000000000 : node527;
													assign node527 = (inp[12]) ? node533 : node528;
														assign node528 = (inp[5]) ? node530 : 46'b0000000000000000000000000000000000000000000000;
															assign node530 = (inp[4]) ? 46'b0000000000000011000000000001000010000000100010 : 46'b0000000000000001000000000001000010000000100010;
														assign node533 = (inp[5]) ? 46'b0000000000000000000000000000000000000000000000 : 46'b0001000000000101000000000001000000000000100010;
								assign node537 = (inp[7]) ? node601 : node538;
									assign node538 = (inp[0]) ? node570 : node539;
										assign node539 = (inp[4]) ? node555 : node540;
											assign node540 = (inp[14]) ? node546 : node541;
												assign node541 = (inp[6]) ? 46'b0000000000100100000000000000100010000000100000 : node542;
													assign node542 = (inp[10]) ? 46'b0001000000100000000000000001100010100000100010 : 46'b0000000000100100000000000001100000100000100010;
												assign node546 = (inp[6]) ? node552 : node547;
													assign node547 = (inp[5]) ? node549 : 46'b0001000000100110000000000000100010100000100000;
														assign node549 = (inp[12]) ? 46'b0000000000100110000000000000100000100000100000 : 46'b0000000000100110000000000000100010100000100000;
													assign node552 = (inp[12]) ? 46'b0000000000100110000000000000100000000000100000 : 46'b0000000000100110000000000000100010000000100000;
											assign node555 = (inp[5]) ? node557 : 46'b0001000000100110000000000000100000000000100000;
												assign node557 = (inp[6]) ? node567 : node558;
													assign node558 = (inp[8]) ? node564 : node559;
														assign node559 = (inp[14]) ? 46'b0000000000100000001000000001100010100000100000 : node560;
															assign node560 = (inp[12]) ? 46'b0000000000100100001000000001100000100000100000 : 46'b0000000000100100001000000001100010100000100000;
														assign node564 = (inp[10]) ? 46'b0000000000100010000000000001100010100000100010 : 46'b0000000000100000001000000001100010100000100010;
													assign node567 = (inp[12]) ? 46'b0000000000100000001000000001100000000000100010 : 46'b0000000000100010001000000001100010000000100000;
										assign node570 = (inp[5]) ? node584 : node571;
											assign node571 = (inp[12]) ? node575 : node572;
												assign node572 = (inp[4]) ? 46'b0001000000000010000000000000100010000000100000 : 46'b0001000000000100000000000000100010100000100000;
												assign node575 = (inp[14]) ? node579 : node576;
													assign node576 = (inp[4]) ? 46'b0001000000000100001000000001100000100000100000 : 46'b0001000000000100000000000000100000000000100000;
													assign node579 = (inp[4]) ? node581 : 46'b0001000000000100001000000001100000000000100000;
														assign node581 = (inp[8]) ? 46'b0001000000000010001000000001100000000000100000 : 46'b0001000000000000001000000001100000000000100000;
											assign node584 = (inp[10]) ? node592 : node585;
												assign node585 = (inp[4]) ? 46'b0000000000000100001000000001100010100000100000 : node586;
													assign node586 = (inp[14]) ? 46'b0000000000000110000000000000100010000000100000 : node587;
														assign node587 = (inp[8]) ? 46'b0000000000000100000000000001100010000000100010 : 46'b0000000000000100000000000000100010000000100000;
												assign node592 = (inp[12]) ? node598 : node593;
													assign node593 = (inp[6]) ? node595 : 46'b0000000000000010000000000001100010100000100010;
														assign node595 = (inp[8]) ? 46'b0000000000000000000000000001100010000000100010 : 46'b0000000000000100000000000001100010000000100010;
													assign node598 = (inp[14]) ? 46'b0000000000000010000000000001100000000000100010 : 46'b0000000000000010000000000001100000100000100010;
									assign node601 = (inp[12]) ? node627 : node602;
										assign node602 = (inp[8]) ? node618 : node603;
											assign node603 = (inp[0]) ? node609 : node604;
												assign node604 = (inp[4]) ? 46'b0001000000100100001000000001000010000000100000 : node605;
													assign node605 = (inp[5]) ? 46'b0000000000100100000000000001000010000000100010 : 46'b0001000000100100000000000001000010000000100010;
												assign node609 = (inp[14]) ? node613 : node610;
													assign node610 = (inp[10]) ? 46'b0000000000000110000000000000000010000000100000 : 46'b0000000000000100000000000000000010100000100000;
													assign node613 = (inp[4]) ? node615 : 46'b0000000000000000001000000001000010000000100010;
														assign node615 = (inp[6]) ? 46'b0000000000000000001000000001000010000000100000 : 46'b0000000000000000001000000001000010100000100000;
											assign node618 = (inp[10]) ? node622 : node619;
												assign node619 = (inp[6]) ? 46'b0001000000000010001000000001000010000000100000 : 46'b0001000000000010001000000001000010100000100000;
												assign node622 = (inp[0]) ? node624 : 46'b0001000000100010000000000000000010100000100000;
													assign node624 = (inp[14]) ? 46'b0001000000000010000000000000000010000000100000 : 46'b0001000000000010000000000001000010000000100010;
										assign node627 = (inp[8]) ? node645 : node628;
											assign node628 = (inp[14]) ? node634 : node629;
												assign node629 = (inp[0]) ? 46'b0001000000000100000000000001000000000000100010 : node630;
													assign node630 = (inp[4]) ? 46'b0001000000100110000000000000000000000000100000 : 46'b0000000000100100000000000000000000000000100000;
												assign node634 = (inp[10]) ? node642 : node635;
													assign node635 = (inp[6]) ? 46'b0001000000000100001000000001000000000000100000 : node636;
														assign node636 = (inp[5]) ? 46'b0000000000100100001000000001000000100000100000 : node637;
															assign node637 = (inp[4]) ? 46'b0001000000100000001000000001000000100000100000 : 46'b0001000000100100001000000001000000100000100000;
													assign node642 = (inp[6]) ? 46'b0001000000100000001000000001000000000000100010 : 46'b0001000000100000001000000001000000100000100010;
											assign node645 = (inp[6]) ? node653 : node646;
												assign node646 = (inp[10]) ? node650 : node647;
													assign node647 = (inp[0]) ? 46'b0000000000000000001000000001000000100000100010 : 46'b0000000000100010001000000001000000100000100000;
													assign node650 = (inp[5]) ? 46'b0000000000000010000000000001000000100000100010 : 46'b0001000000000010000000000001000000100000100010;
												assign node653 = (inp[10]) ? node655 : 46'b0000000000100100000000000001000000000000100010;
													assign node655 = (inp[5]) ? 46'b0000000000100010000000000001000000000000100010 : 46'b0001000000100010000000000001000000000000100010;
							assign node658 = (inp[0]) ? node698 : node659;
								assign node659 = (inp[9]) ? node679 : node660;
									assign node660 = (inp[12]) ? node670 : node661;
										assign node661 = (inp[6]) ? node663 : 46'b0000000000000000000000000000000000000000000000;
											assign node663 = (inp[5]) ? node667 : node664;
												assign node664 = (inp[7]) ? 46'b0001000000100010000000000000000010000000100000 : 46'b0001000000100010000000000000100010000000100000;
												assign node667 = (inp[7]) ? 46'b0000000000100010000000000000000010000000100000 : 46'b0000000000100010000000000000100010000000100000;
										assign node670 = (inp[6]) ? 46'b0000000000000000000000000000000000000000000000 : node671;
											assign node671 = (inp[5]) ? node675 : node672;
												assign node672 = (inp[7]) ? 46'b0001000000100000001000000001000000100000100000 : 46'b0001000000100000001000000001100000100000100000;
												assign node675 = (inp[7]) ? 46'b0000000000100000001000000001000000100000100000 : 46'b0000000000100000001000000001100000100000100000;
									assign node679 = (inp[5]) ? node689 : node680;
										assign node680 = (inp[7]) ? node682 : 46'b0000000000000000000000000000000000000000000000;
											assign node682 = (inp[12]) ? node686 : node683;
												assign node683 = (inp[6]) ? 46'b0001000010000100000000000000000010000001000000 : 46'b0001000010000100000000000000000010100001000000;
												assign node686 = (inp[10]) ? 46'b0001000010000100000000000000000000000001000000 : 46'b0001000010000100000000000000000000100001000000;
										assign node689 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node690;
											assign node690 = (inp[6]) ? node694 : node691;
												assign node691 = (inp[12]) ? 46'b0000000010000000000000000001100000100001000010 : 46'b0000000010000000000000000001100010100001000010;
												assign node694 = (inp[14]) ? 46'b0000000010000000000000000001100000000001000010 : 46'b0000000010000000000000000001100010000001000010;
								assign node698 = (inp[9]) ? 46'b0000000000000000000000000000000000000000000000 : node699;
									assign node699 = (inp[5]) ? node709 : node700;
										assign node700 = (inp[7]) ? node702 : 46'b0000000000000000000000000000000000000000000000;
											assign node702 = (inp[12]) ? node706 : node703;
												assign node703 = (inp[6]) ? 46'b0001000010000100000000000000000010000000000000 : 46'b0001000010000100000000000000000010100000000000;
												assign node706 = (inp[6]) ? 46'b0001000010000100000000000000000000000000000000 : 46'b0001000010000100000000000000000000100000000000;
										assign node709 = (inp[7]) ? 46'b0000000000000000000000000000000000000000000000 : node710;
											assign node710 = (inp[6]) ? 46'b0000000010000000000000000001100000000000000010 : node711;
												assign node711 = (inp[12]) ? 46'b0000000010000000000000000001100000100000000010 : 46'b0000000010000000000000000001100010100000000010;

endmodule