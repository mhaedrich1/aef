module dtc_split33_bm63 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node14;
	wire [4-1:0] node17;
	wire [4-1:0] node18;
	wire [4-1:0] node20;
	wire [4-1:0] node23;
	wire [4-1:0] node26;
	wire [4-1:0] node27;
	wire [4-1:0] node28;
	wire [4-1:0] node32;
	wire [4-1:0] node34;
	wire [4-1:0] node35;
	wire [4-1:0] node39;
	wire [4-1:0] node40;
	wire [4-1:0] node41;
	wire [4-1:0] node42;
	wire [4-1:0] node43;
	wire [4-1:0] node48;
	wire [4-1:0] node49;
	wire [4-1:0] node51;
	wire [4-1:0] node54;
	wire [4-1:0] node55;
	wire [4-1:0] node59;
	wire [4-1:0] node60;
	wire [4-1:0] node62;
	wire [4-1:0] node63;
	wire [4-1:0] node67;
	wire [4-1:0] node70;
	wire [4-1:0] node71;
	wire [4-1:0] node72;
	wire [4-1:0] node75;
	wire [4-1:0] node77;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node82;
	wire [4-1:0] node83;
	wire [4-1:0] node85;
	wire [4-1:0] node88;
	wire [4-1:0] node89;
	wire [4-1:0] node93;
	wire [4-1:0] node94;
	wire [4-1:0] node96;
	wire [4-1:0] node100;
	wire [4-1:0] node101;
	wire [4-1:0] node102;
	wire [4-1:0] node104;
	wire [4-1:0] node108;
	wire [4-1:0] node109;
	wire [4-1:0] node110;
	wire [4-1:0] node114;
	wire [4-1:0] node117;
	wire [4-1:0] node118;
	wire [4-1:0] node119;
	wire [4-1:0] node120;
	wire [4-1:0] node121;
	wire [4-1:0] node122;
	wire [4-1:0] node125;
	wire [4-1:0] node128;
	wire [4-1:0] node129;
	wire [4-1:0] node132;
	wire [4-1:0] node135;
	wire [4-1:0] node136;
	wire [4-1:0] node137;
	wire [4-1:0] node138;
	wire [4-1:0] node142;
	wire [4-1:0] node143;
	wire [4-1:0] node148;
	wire [4-1:0] node149;
	wire [4-1:0] node150;
	wire [4-1:0] node153;
	wire [4-1:0] node155;
	wire [4-1:0] node158;
	wire [4-1:0] node159;
	wire [4-1:0] node160;
	wire [4-1:0] node161;
	wire [4-1:0] node164;
	wire [4-1:0] node167;
	wire [4-1:0] node170;
	wire [4-1:0] node173;
	wire [4-1:0] node174;
	wire [4-1:0] node175;
	wire [4-1:0] node176;
	wire [4-1:0] node178;
	wire [4-1:0] node181;
	wire [4-1:0] node182;
	wire [4-1:0] node183;
	wire [4-1:0] node186;
	wire [4-1:0] node190;
	wire [4-1:0] node191;
	wire [4-1:0] node192;
	wire [4-1:0] node193;
	wire [4-1:0] node197;
	wire [4-1:0] node200;
	wire [4-1:0] node201;
	wire [4-1:0] node202;
	wire [4-1:0] node207;
	wire [4-1:0] node208;
	wire [4-1:0] node209;
	wire [4-1:0] node210;
	wire [4-1:0] node214;
	wire [4-1:0] node215;
	wire [4-1:0] node216;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node224;
	wire [4-1:0] node226;
	wire [4-1:0] node229;
	wire [4-1:0] node232;
	wire [4-1:0] node233;
	wire [4-1:0] node234;
	wire [4-1:0] node235;
	wire [4-1:0] node236;
	wire [4-1:0] node237;
	wire [4-1:0] node239;
	wire [4-1:0] node242;
	wire [4-1:0] node244;
	wire [4-1:0] node247;
	wire [4-1:0] node249;
	wire [4-1:0] node252;
	wire [4-1:0] node253;
	wire [4-1:0] node254;
	wire [4-1:0] node255;
	wire [4-1:0] node256;
	wire [4-1:0] node259;
	wire [4-1:0] node262;
	wire [4-1:0] node265;
	wire [4-1:0] node266;
	wire [4-1:0] node267;
	wire [4-1:0] node270;
	wire [4-1:0] node273;
	wire [4-1:0] node275;
	wire [4-1:0] node278;
	wire [4-1:0] node279;
	wire [4-1:0] node282;
	wire [4-1:0] node283;
	wire [4-1:0] node284;
	wire [4-1:0] node289;
	wire [4-1:0] node290;
	wire [4-1:0] node291;
	wire [4-1:0] node292;
	wire [4-1:0] node293;
	wire [4-1:0] node294;
	wire [4-1:0] node298;
	wire [4-1:0] node301;
	wire [4-1:0] node302;
	wire [4-1:0] node303;
	wire [4-1:0] node306;
	wire [4-1:0] node310;
	wire [4-1:0] node311;
	wire [4-1:0] node312;
	wire [4-1:0] node313;
	wire [4-1:0] node316;
	wire [4-1:0] node320;
	wire [4-1:0] node322;
	wire [4-1:0] node323;
	wire [4-1:0] node327;
	wire [4-1:0] node328;
	wire [4-1:0] node329;
	wire [4-1:0] node331;
	wire [4-1:0] node333;
	wire [4-1:0] node336;
	wire [4-1:0] node337;
	wire [4-1:0] node338;
	wire [4-1:0] node343;
	wire [4-1:0] node344;
	wire [4-1:0] node346;
	wire [4-1:0] node349;
	wire [4-1:0] node352;
	wire [4-1:0] node353;
	wire [4-1:0] node354;
	wire [4-1:0] node355;
	wire [4-1:0] node356;
	wire [4-1:0] node357;
	wire [4-1:0] node358;
	wire [4-1:0] node362;
	wire [4-1:0] node365;
	wire [4-1:0] node366;
	wire [4-1:0] node368;
	wire [4-1:0] node371;
	wire [4-1:0] node372;
	wire [4-1:0] node375;
	wire [4-1:0] node378;
	wire [4-1:0] node379;
	wire [4-1:0] node381;
	wire [4-1:0] node384;
	wire [4-1:0] node386;
	wire [4-1:0] node389;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node392;
	wire [4-1:0] node395;
	wire [4-1:0] node398;
	wire [4-1:0] node399;
	wire [4-1:0] node403;
	wire [4-1:0] node404;
	wire [4-1:0] node407;
	wire [4-1:0] node408;
	wire [4-1:0] node409;
	wire [4-1:0] node414;
	wire [4-1:0] node415;
	wire [4-1:0] node416;
	wire [4-1:0] node417;
	wire [4-1:0] node418;
	wire [4-1:0] node422;
	wire [4-1:0] node423;
	wire [4-1:0] node427;
	wire [4-1:0] node428;
	wire [4-1:0] node429;
	wire [4-1:0] node431;
	wire [4-1:0] node436;
	wire [4-1:0] node437;
	wire [4-1:0] node438;
	wire [4-1:0] node439;
	wire [4-1:0] node443;
	wire [4-1:0] node444;
	wire [4-1:0] node446;
	wire [4-1:0] node449;
	wire [4-1:0] node452;
	wire [4-1:0] node453;
	wire [4-1:0] node454;
	wire [4-1:0] node456;
	wire [4-1:0] node459;
	wire [4-1:0] node461;
	wire [4-1:0] node464;
	wire [4-1:0] node465;
	wire [4-1:0] node469;
	wire [4-1:0] node470;
	wire [4-1:0] node471;
	wire [4-1:0] node472;
	wire [4-1:0] node473;
	wire [4-1:0] node474;
	wire [4-1:0] node475;
	wire [4-1:0] node478;
	wire [4-1:0] node479;
	wire [4-1:0] node482;
	wire [4-1:0] node485;
	wire [4-1:0] node486;
	wire [4-1:0] node487;
	wire [4-1:0] node488;
	wire [4-1:0] node491;
	wire [4-1:0] node495;
	wire [4-1:0] node497;
	wire [4-1:0] node498;
	wire [4-1:0] node502;
	wire [4-1:0] node503;
	wire [4-1:0] node504;
	wire [4-1:0] node505;
	wire [4-1:0] node507;
	wire [4-1:0] node510;
	wire [4-1:0] node512;
	wire [4-1:0] node516;
	wire [4-1:0] node517;
	wire [4-1:0] node518;
	wire [4-1:0] node520;
	wire [4-1:0] node523;
	wire [4-1:0] node526;
	wire [4-1:0] node527;
	wire [4-1:0] node529;
	wire [4-1:0] node533;
	wire [4-1:0] node534;
	wire [4-1:0] node535;
	wire [4-1:0] node536;
	wire [4-1:0] node537;
	wire [4-1:0] node540;
	wire [4-1:0] node542;
	wire [4-1:0] node545;
	wire [4-1:0] node546;
	wire [4-1:0] node550;
	wire [4-1:0] node551;
	wire [4-1:0] node552;
	wire [4-1:0] node554;
	wire [4-1:0] node557;
	wire [4-1:0] node560;
	wire [4-1:0] node561;
	wire [4-1:0] node563;
	wire [4-1:0] node566;
	wire [4-1:0] node569;
	wire [4-1:0] node570;
	wire [4-1:0] node571;
	wire [4-1:0] node572;
	wire [4-1:0] node573;
	wire [4-1:0] node577;
	wire [4-1:0] node579;
	wire [4-1:0] node582;
	wire [4-1:0] node583;
	wire [4-1:0] node585;
	wire [4-1:0] node588;
	wire [4-1:0] node591;
	wire [4-1:0] node592;
	wire [4-1:0] node593;
	wire [4-1:0] node597;
	wire [4-1:0] node600;
	wire [4-1:0] node601;
	wire [4-1:0] node602;
	wire [4-1:0] node603;
	wire [4-1:0] node604;
	wire [4-1:0] node605;
	wire [4-1:0] node609;
	wire [4-1:0] node610;
	wire [4-1:0] node613;
	wire [4-1:0] node616;
	wire [4-1:0] node617;
	wire [4-1:0] node618;
	wire [4-1:0] node621;
	wire [4-1:0] node624;
	wire [4-1:0] node625;
	wire [4-1:0] node627;
	wire [4-1:0] node630;
	wire [4-1:0] node633;
	wire [4-1:0] node634;
	wire [4-1:0] node635;
	wire [4-1:0] node636;
	wire [4-1:0] node638;
	wire [4-1:0] node642;
	wire [4-1:0] node645;
	wire [4-1:0] node648;
	wire [4-1:0] node649;
	wire [4-1:0] node650;
	wire [4-1:0] node651;
	wire [4-1:0] node652;
	wire [4-1:0] node653;
	wire [4-1:0] node656;
	wire [4-1:0] node660;
	wire [4-1:0] node661;
	wire [4-1:0] node663;
	wire [4-1:0] node667;
	wire [4-1:0] node668;
	wire [4-1:0] node669;
	wire [4-1:0] node672;
	wire [4-1:0] node675;
	wire [4-1:0] node676;
	wire [4-1:0] node677;
	wire [4-1:0] node681;
	wire [4-1:0] node683;
	wire [4-1:0] node686;
	wire [4-1:0] node687;
	wire [4-1:0] node688;
	wire [4-1:0] node689;
	wire [4-1:0] node690;
	wire [4-1:0] node693;
	wire [4-1:0] node697;
	wire [4-1:0] node700;
	wire [4-1:0] node701;
	wire [4-1:0] node702;
	wire [4-1:0] node705;
	wire [4-1:0] node706;
	wire [4-1:0] node709;
	wire [4-1:0] node712;
	wire [4-1:0] node714;
	wire [4-1:0] node717;
	wire [4-1:0] node718;
	wire [4-1:0] node719;
	wire [4-1:0] node720;
	wire [4-1:0] node721;
	wire [4-1:0] node722;
	wire [4-1:0] node723;
	wire [4-1:0] node725;
	wire [4-1:0] node728;
	wire [4-1:0] node731;
	wire [4-1:0] node734;
	wire [4-1:0] node735;
	wire [4-1:0] node737;
	wire [4-1:0] node740;
	wire [4-1:0] node742;
	wire [4-1:0] node743;
	wire [4-1:0] node747;
	wire [4-1:0] node748;
	wire [4-1:0] node749;
	wire [4-1:0] node750;
	wire [4-1:0] node751;
	wire [4-1:0] node754;
	wire [4-1:0] node758;
	wire [4-1:0] node759;
	wire [4-1:0] node761;
	wire [4-1:0] node764;
	wire [4-1:0] node765;
	wire [4-1:0] node769;
	wire [4-1:0] node770;
	wire [4-1:0] node771;
	wire [4-1:0] node772;
	wire [4-1:0] node775;
	wire [4-1:0] node778;
	wire [4-1:0] node781;
	wire [4-1:0] node782;
	wire [4-1:0] node784;
	wire [4-1:0] node787;
	wire [4-1:0] node788;
	wire [4-1:0] node792;
	wire [4-1:0] node793;
	wire [4-1:0] node794;
	wire [4-1:0] node795;
	wire [4-1:0] node796;
	wire [4-1:0] node797;
	wire [4-1:0] node801;
	wire [4-1:0] node804;
	wire [4-1:0] node806;
	wire [4-1:0] node807;
	wire [4-1:0] node810;
	wire [4-1:0] node813;
	wire [4-1:0] node814;
	wire [4-1:0] node815;
	wire [4-1:0] node819;
	wire [4-1:0] node821;
	wire [4-1:0] node823;
	wire [4-1:0] node826;
	wire [4-1:0] node827;
	wire [4-1:0] node828;
	wire [4-1:0] node830;
	wire [4-1:0] node832;
	wire [4-1:0] node835;
	wire [4-1:0] node836;
	wire [4-1:0] node839;
	wire [4-1:0] node840;
	wire [4-1:0] node844;
	wire [4-1:0] node845;
	wire [4-1:0] node846;
	wire [4-1:0] node849;
	wire [4-1:0] node851;
	wire [4-1:0] node854;
	wire [4-1:0] node855;
	wire [4-1:0] node859;
	wire [4-1:0] node860;
	wire [4-1:0] node861;
	wire [4-1:0] node862;
	wire [4-1:0] node864;
	wire [4-1:0] node865;
	wire [4-1:0] node867;
	wire [4-1:0] node870;
	wire [4-1:0] node872;
	wire [4-1:0] node875;
	wire [4-1:0] node876;
	wire [4-1:0] node878;
	wire [4-1:0] node881;
	wire [4-1:0] node882;
	wire [4-1:0] node883;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node891;
	wire [4-1:0] node892;
	wire [4-1:0] node893;
	wire [4-1:0] node896;
	wire [4-1:0] node899;
	wire [4-1:0] node900;
	wire [4-1:0] node903;
	wire [4-1:0] node906;
	wire [4-1:0] node907;
	wire [4-1:0] node908;
	wire [4-1:0] node911;
	wire [4-1:0] node915;
	wire [4-1:0] node916;
	wire [4-1:0] node917;
	wire [4-1:0] node918;
	wire [4-1:0] node919;
	wire [4-1:0] node921;
	wire [4-1:0] node925;
	wire [4-1:0] node926;
	wire [4-1:0] node928;
	wire [4-1:0] node931;
	wire [4-1:0] node934;
	wire [4-1:0] node935;
	wire [4-1:0] node936;
	wire [4-1:0] node938;
	wire [4-1:0] node941;
	wire [4-1:0] node944;
	wire [4-1:0] node947;
	wire [4-1:0] node948;
	wire [4-1:0] node949;
	wire [4-1:0] node950;
	wire [4-1:0] node951;
	wire [4-1:0] node954;
	wire [4-1:0] node957;
	wire [4-1:0] node958;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node965;
	wire [4-1:0] node968;
	wire [4-1:0] node971;
	wire [4-1:0] node972;
	wire [4-1:0] node973;
	wire [4-1:0] node975;
	wire [4-1:0] node979;
	wire [4-1:0] node980;
	wire [4-1:0] node982;
	wire [4-1:0] node985;
	wire [4-1:0] node988;
	wire [4-1:0] node989;
	wire [4-1:0] node990;
	wire [4-1:0] node991;
	wire [4-1:0] node992;
	wire [4-1:0] node993;
	wire [4-1:0] node994;
	wire [4-1:0] node995;
	wire [4-1:0] node996;
	wire [4-1:0] node1000;
	wire [4-1:0] node1001;
	wire [4-1:0] node1003;
	wire [4-1:0] node1007;
	wire [4-1:0] node1008;
	wire [4-1:0] node1009;
	wire [4-1:0] node1010;
	wire [4-1:0] node1014;
	wire [4-1:0] node1015;
	wire [4-1:0] node1018;
	wire [4-1:0] node1021;
	wire [4-1:0] node1022;
	wire [4-1:0] node1024;
	wire [4-1:0] node1027;
	wire [4-1:0] node1028;
	wire [4-1:0] node1032;
	wire [4-1:0] node1033;
	wire [4-1:0] node1034;
	wire [4-1:0] node1035;
	wire [4-1:0] node1037;
	wire [4-1:0] node1041;
	wire [4-1:0] node1043;
	wire [4-1:0] node1045;
	wire [4-1:0] node1048;
	wire [4-1:0] node1050;
	wire [4-1:0] node1053;
	wire [4-1:0] node1054;
	wire [4-1:0] node1055;
	wire [4-1:0] node1056;
	wire [4-1:0] node1058;
	wire [4-1:0] node1061;
	wire [4-1:0] node1062;
	wire [4-1:0] node1063;
	wire [4-1:0] node1068;
	wire [4-1:0] node1069;
	wire [4-1:0] node1070;
	wire [4-1:0] node1071;
	wire [4-1:0] node1074;
	wire [4-1:0] node1077;
	wire [4-1:0] node1080;
	wire [4-1:0] node1081;
	wire [4-1:0] node1082;
	wire [4-1:0] node1085;
	wire [4-1:0] node1088;
	wire [4-1:0] node1089;
	wire [4-1:0] node1093;
	wire [4-1:0] node1094;
	wire [4-1:0] node1095;
	wire [4-1:0] node1097;
	wire [4-1:0] node1100;
	wire [4-1:0] node1102;
	wire [4-1:0] node1105;
	wire [4-1:0] node1107;
	wire [4-1:0] node1108;
	wire [4-1:0] node1111;
	wire [4-1:0] node1113;
	wire [4-1:0] node1116;
	wire [4-1:0] node1117;
	wire [4-1:0] node1118;
	wire [4-1:0] node1119;
	wire [4-1:0] node1120;
	wire [4-1:0] node1122;
	wire [4-1:0] node1123;
	wire [4-1:0] node1126;
	wire [4-1:0] node1129;
	wire [4-1:0] node1130;
	wire [4-1:0] node1132;
	wire [4-1:0] node1136;
	wire [4-1:0] node1137;
	wire [4-1:0] node1140;
	wire [4-1:0] node1141;
	wire [4-1:0] node1145;
	wire [4-1:0] node1146;
	wire [4-1:0] node1148;
	wire [4-1:0] node1149;
	wire [4-1:0] node1153;
	wire [4-1:0] node1154;
	wire [4-1:0] node1155;
	wire [4-1:0] node1159;
	wire [4-1:0] node1161;
	wire [4-1:0] node1164;
	wire [4-1:0] node1165;
	wire [4-1:0] node1166;
	wire [4-1:0] node1167;
	wire [4-1:0] node1168;
	wire [4-1:0] node1170;
	wire [4-1:0] node1174;
	wire [4-1:0] node1176;
	wire [4-1:0] node1177;
	wire [4-1:0] node1180;
	wire [4-1:0] node1183;
	wire [4-1:0] node1184;
	wire [4-1:0] node1185;
	wire [4-1:0] node1188;
	wire [4-1:0] node1191;
	wire [4-1:0] node1192;
	wire [4-1:0] node1196;
	wire [4-1:0] node1197;
	wire [4-1:0] node1198;
	wire [4-1:0] node1200;
	wire [4-1:0] node1201;
	wire [4-1:0] node1204;
	wire [4-1:0] node1207;
	wire [4-1:0] node1209;
	wire [4-1:0] node1212;
	wire [4-1:0] node1213;
	wire [4-1:0] node1215;
	wire [4-1:0] node1218;
	wire [4-1:0] node1219;
	wire [4-1:0] node1220;
	wire [4-1:0] node1223;
	wire [4-1:0] node1227;
	wire [4-1:0] node1228;
	wire [4-1:0] node1229;
	wire [4-1:0] node1230;
	wire [4-1:0] node1231;
	wire [4-1:0] node1232;
	wire [4-1:0] node1234;
	wire [4-1:0] node1238;
	wire [4-1:0] node1239;
	wire [4-1:0] node1240;
	wire [4-1:0] node1244;
	wire [4-1:0] node1245;
	wire [4-1:0] node1246;
	wire [4-1:0] node1249;
	wire [4-1:0] node1253;
	wire [4-1:0] node1254;
	wire [4-1:0] node1255;
	wire [4-1:0] node1256;
	wire [4-1:0] node1257;
	wire [4-1:0] node1262;
	wire [4-1:0] node1263;
	wire [4-1:0] node1266;
	wire [4-1:0] node1269;
	wire [4-1:0] node1271;
	wire [4-1:0] node1272;
	wire [4-1:0] node1274;
	wire [4-1:0] node1278;
	wire [4-1:0] node1279;
	wire [4-1:0] node1280;
	wire [4-1:0] node1281;
	wire [4-1:0] node1283;
	wire [4-1:0] node1286;
	wire [4-1:0] node1287;
	wire [4-1:0] node1288;
	wire [4-1:0] node1291;
	wire [4-1:0] node1295;
	wire [4-1:0] node1296;
	wire [4-1:0] node1299;
	wire [4-1:0] node1300;
	wire [4-1:0] node1302;
	wire [4-1:0] node1306;
	wire [4-1:0] node1307;
	wire [4-1:0] node1309;
	wire [4-1:0] node1310;
	wire [4-1:0] node1312;
	wire [4-1:0] node1315;
	wire [4-1:0] node1317;
	wire [4-1:0] node1320;
	wire [4-1:0] node1321;
	wire [4-1:0] node1322;
	wire [4-1:0] node1325;
	wire [4-1:0] node1328;
	wire [4-1:0] node1329;
	wire [4-1:0] node1330;
	wire [4-1:0] node1333;
	wire [4-1:0] node1337;
	wire [4-1:0] node1338;
	wire [4-1:0] node1339;
	wire [4-1:0] node1340;
	wire [4-1:0] node1342;
	wire [4-1:0] node1343;
	wire [4-1:0] node1347;
	wire [4-1:0] node1348;
	wire [4-1:0] node1351;
	wire [4-1:0] node1353;
	wire [4-1:0] node1354;
	wire [4-1:0] node1357;
	wire [4-1:0] node1360;
	wire [4-1:0] node1361;
	wire [4-1:0] node1362;
	wire [4-1:0] node1363;
	wire [4-1:0] node1364;
	wire [4-1:0] node1369;
	wire [4-1:0] node1371;
	wire [4-1:0] node1374;
	wire [4-1:0] node1375;
	wire [4-1:0] node1376;
	wire [4-1:0] node1379;
	wire [4-1:0] node1381;
	wire [4-1:0] node1384;
	wire [4-1:0] node1385;
	wire [4-1:0] node1389;
	wire [4-1:0] node1390;
	wire [4-1:0] node1391;
	wire [4-1:0] node1392;
	wire [4-1:0] node1393;
	wire [4-1:0] node1397;
	wire [4-1:0] node1399;
	wire [4-1:0] node1401;
	wire [4-1:0] node1404;
	wire [4-1:0] node1405;
	wire [4-1:0] node1408;
	wire [4-1:0] node1410;
	wire [4-1:0] node1411;
	wire [4-1:0] node1415;
	wire [4-1:0] node1416;
	wire [4-1:0] node1417;
	wire [4-1:0] node1420;
	wire [4-1:0] node1421;
	wire [4-1:0] node1425;
	wire [4-1:0] node1426;
	wire [4-1:0] node1428;
	wire [4-1:0] node1429;
	wire [4-1:0] node1433;
	wire [4-1:0] node1435;
	wire [4-1:0] node1436;
	wire [4-1:0] node1440;
	wire [4-1:0] node1441;
	wire [4-1:0] node1442;
	wire [4-1:0] node1443;
	wire [4-1:0] node1444;
	wire [4-1:0] node1445;
	wire [4-1:0] node1446;
	wire [4-1:0] node1448;
	wire [4-1:0] node1450;
	wire [4-1:0] node1453;
	wire [4-1:0] node1454;
	wire [4-1:0] node1455;
	wire [4-1:0] node1458;
	wire [4-1:0] node1462;
	wire [4-1:0] node1463;
	wire [4-1:0] node1464;
	wire [4-1:0] node1465;
	wire [4-1:0] node1470;
	wire [4-1:0] node1472;
	wire [4-1:0] node1475;
	wire [4-1:0] node1476;
	wire [4-1:0] node1477;
	wire [4-1:0] node1478;
	wire [4-1:0] node1480;
	wire [4-1:0] node1485;
	wire [4-1:0] node1486;
	wire [4-1:0] node1488;
	wire [4-1:0] node1491;
	wire [4-1:0] node1494;
	wire [4-1:0] node1495;
	wire [4-1:0] node1496;
	wire [4-1:0] node1497;
	wire [4-1:0] node1498;
	wire [4-1:0] node1499;
	wire [4-1:0] node1502;
	wire [4-1:0] node1506;
	wire [4-1:0] node1508;
	wire [4-1:0] node1511;
	wire [4-1:0] node1512;
	wire [4-1:0] node1513;
	wire [4-1:0] node1516;
	wire [4-1:0] node1519;
	wire [4-1:0] node1520;
	wire [4-1:0] node1524;
	wire [4-1:0] node1525;
	wire [4-1:0] node1526;
	wire [4-1:0] node1528;
	wire [4-1:0] node1529;
	wire [4-1:0] node1533;
	wire [4-1:0] node1534;
	wire [4-1:0] node1536;
	wire [4-1:0] node1539;
	wire [4-1:0] node1542;
	wire [4-1:0] node1543;
	wire [4-1:0] node1545;
	wire [4-1:0] node1546;
	wire [4-1:0] node1549;
	wire [4-1:0] node1552;
	wire [4-1:0] node1553;
	wire [4-1:0] node1554;
	wire [4-1:0] node1557;
	wire [4-1:0] node1560;
	wire [4-1:0] node1561;
	wire [4-1:0] node1564;
	wire [4-1:0] node1567;
	wire [4-1:0] node1568;
	wire [4-1:0] node1569;
	wire [4-1:0] node1570;
	wire [4-1:0] node1571;
	wire [4-1:0] node1572;
	wire [4-1:0] node1573;
	wire [4-1:0] node1578;
	wire [4-1:0] node1581;
	wire [4-1:0] node1582;
	wire [4-1:0] node1583;
	wire [4-1:0] node1586;
	wire [4-1:0] node1589;
	wire [4-1:0] node1590;
	wire [4-1:0] node1591;
	wire [4-1:0] node1594;
	wire [4-1:0] node1598;
	wire [4-1:0] node1599;
	wire [4-1:0] node1600;
	wire [4-1:0] node1601;
	wire [4-1:0] node1603;
	wire [4-1:0] node1607;
	wire [4-1:0] node1609;
	wire [4-1:0] node1610;
	wire [4-1:0] node1614;
	wire [4-1:0] node1615;
	wire [4-1:0] node1616;
	wire [4-1:0] node1620;
	wire [4-1:0] node1622;
	wire [4-1:0] node1623;
	wire [4-1:0] node1626;
	wire [4-1:0] node1629;
	wire [4-1:0] node1630;
	wire [4-1:0] node1631;
	wire [4-1:0] node1632;
	wire [4-1:0] node1636;
	wire [4-1:0] node1637;
	wire [4-1:0] node1639;
	wire [4-1:0] node1641;
	wire [4-1:0] node1644;
	wire [4-1:0] node1645;
	wire [4-1:0] node1646;
	wire [4-1:0] node1650;
	wire [4-1:0] node1652;
	wire [4-1:0] node1655;
	wire [4-1:0] node1656;
	wire [4-1:0] node1657;
	wire [4-1:0] node1659;
	wire [4-1:0] node1661;
	wire [4-1:0] node1664;
	wire [4-1:0] node1665;
	wire [4-1:0] node1666;
	wire [4-1:0] node1669;
	wire [4-1:0] node1672;
	wire [4-1:0] node1673;
	wire [4-1:0] node1676;
	wire [4-1:0] node1679;
	wire [4-1:0] node1680;
	wire [4-1:0] node1681;
	wire [4-1:0] node1682;
	wire [4-1:0] node1686;
	wire [4-1:0] node1689;
	wire [4-1:0] node1690;
	wire [4-1:0] node1692;
	wire [4-1:0] node1695;
	wire [4-1:0] node1698;
	wire [4-1:0] node1699;
	wire [4-1:0] node1700;
	wire [4-1:0] node1701;
	wire [4-1:0] node1702;
	wire [4-1:0] node1703;
	wire [4-1:0] node1704;
	wire [4-1:0] node1708;
	wire [4-1:0] node1709;
	wire [4-1:0] node1711;
	wire [4-1:0] node1714;
	wire [4-1:0] node1715;
	wire [4-1:0] node1719;
	wire [4-1:0] node1720;
	wire [4-1:0] node1721;
	wire [4-1:0] node1723;
	wire [4-1:0] node1728;
	wire [4-1:0] node1729;
	wire [4-1:0] node1730;
	wire [4-1:0] node1731;
	wire [4-1:0] node1732;
	wire [4-1:0] node1736;
	wire [4-1:0] node1737;
	wire [4-1:0] node1741;
	wire [4-1:0] node1744;
	wire [4-1:0] node1745;
	wire [4-1:0] node1747;
	wire [4-1:0] node1749;
	wire [4-1:0] node1752;
	wire [4-1:0] node1753;
	wire [4-1:0] node1757;
	wire [4-1:0] node1758;
	wire [4-1:0] node1759;
	wire [4-1:0] node1760;
	wire [4-1:0] node1761;
	wire [4-1:0] node1766;
	wire [4-1:0] node1768;
	wire [4-1:0] node1769;
	wire [4-1:0] node1771;
	wire [4-1:0] node1774;
	wire [4-1:0] node1775;
	wire [4-1:0] node1779;
	wire [4-1:0] node1780;
	wire [4-1:0] node1782;
	wire [4-1:0] node1785;
	wire [4-1:0] node1786;
	wire [4-1:0] node1788;
	wire [4-1:0] node1791;
	wire [4-1:0] node1792;
	wire [4-1:0] node1794;
	wire [4-1:0] node1797;
	wire [4-1:0] node1799;
	wire [4-1:0] node1802;
	wire [4-1:0] node1803;
	wire [4-1:0] node1804;
	wire [4-1:0] node1805;
	wire [4-1:0] node1806;
	wire [4-1:0] node1809;
	wire [4-1:0] node1812;
	wire [4-1:0] node1813;
	wire [4-1:0] node1814;
	wire [4-1:0] node1816;
	wire [4-1:0] node1820;
	wire [4-1:0] node1821;
	wire [4-1:0] node1825;
	wire [4-1:0] node1826;
	wire [4-1:0] node1827;
	wire [4-1:0] node1828;
	wire [4-1:0] node1829;
	wire [4-1:0] node1833;
	wire [4-1:0] node1834;
	wire [4-1:0] node1838;
	wire [4-1:0] node1839;
	wire [4-1:0] node1840;
	wire [4-1:0] node1845;
	wire [4-1:0] node1846;
	wire [4-1:0] node1847;
	wire [4-1:0] node1849;
	wire [4-1:0] node1853;
	wire [4-1:0] node1855;
	wire [4-1:0] node1858;
	wire [4-1:0] node1859;
	wire [4-1:0] node1860;
	wire [4-1:0] node1861;
	wire [4-1:0] node1864;
	wire [4-1:0] node1866;
	wire [4-1:0] node1867;
	wire [4-1:0] node1870;
	wire [4-1:0] node1873;
	wire [4-1:0] node1874;
	wire [4-1:0] node1876;
	wire [4-1:0] node1877;
	wire [4-1:0] node1880;
	wire [4-1:0] node1883;
	wire [4-1:0] node1885;
	wire [4-1:0] node1888;
	wire [4-1:0] node1889;
	wire [4-1:0] node1890;
	wire [4-1:0] node1891;
	wire [4-1:0] node1892;
	wire [4-1:0] node1898;
	wire [4-1:0] node1899;
	wire [4-1:0] node1902;
	wire [4-1:0] node1905;
	wire [4-1:0] node1906;
	wire [4-1:0] node1907;
	wire [4-1:0] node1908;
	wire [4-1:0] node1909;
	wire [4-1:0] node1910;
	wire [4-1:0] node1911;
	wire [4-1:0] node1912;
	wire [4-1:0] node1913;
	wire [4-1:0] node1914;
	wire [4-1:0] node1917;
	wire [4-1:0] node1920;
	wire [4-1:0] node1922;
	wire [4-1:0] node1925;
	wire [4-1:0] node1926;
	wire [4-1:0] node1928;
	wire [4-1:0] node1931;
	wire [4-1:0] node1933;
	wire [4-1:0] node1934;
	wire [4-1:0] node1938;
	wire [4-1:0] node1939;
	wire [4-1:0] node1940;
	wire [4-1:0] node1943;
	wire [4-1:0] node1945;
	wire [4-1:0] node1946;
	wire [4-1:0] node1950;
	wire [4-1:0] node1951;
	wire [4-1:0] node1953;
	wire [4-1:0] node1956;
	wire [4-1:0] node1959;
	wire [4-1:0] node1960;
	wire [4-1:0] node1961;
	wire [4-1:0] node1962;
	wire [4-1:0] node1965;
	wire [4-1:0] node1966;
	wire [4-1:0] node1967;
	wire [4-1:0] node1970;
	wire [4-1:0] node1973;
	wire [4-1:0] node1974;
	wire [4-1:0] node1978;
	wire [4-1:0] node1979;
	wire [4-1:0] node1982;
	wire [4-1:0] node1983;
	wire [4-1:0] node1987;
	wire [4-1:0] node1988;
	wire [4-1:0] node1989;
	wire [4-1:0] node1990;
	wire [4-1:0] node1993;
	wire [4-1:0] node1995;
	wire [4-1:0] node1998;
	wire [4-1:0] node2001;
	wire [4-1:0] node2002;
	wire [4-1:0] node2003;
	wire [4-1:0] node2004;
	wire [4-1:0] node2009;
	wire [4-1:0] node2012;
	wire [4-1:0] node2013;
	wire [4-1:0] node2014;
	wire [4-1:0] node2015;
	wire [4-1:0] node2016;
	wire [4-1:0] node2017;
	wire [4-1:0] node2019;
	wire [4-1:0] node2023;
	wire [4-1:0] node2024;
	wire [4-1:0] node2027;
	wire [4-1:0] node2028;
	wire [4-1:0] node2032;
	wire [4-1:0] node2033;
	wire [4-1:0] node2036;
	wire [4-1:0] node2038;
	wire [4-1:0] node2040;
	wire [4-1:0] node2043;
	wire [4-1:0] node2044;
	wire [4-1:0] node2045;
	wire [4-1:0] node2046;
	wire [4-1:0] node2049;
	wire [4-1:0] node2050;
	wire [4-1:0] node2053;
	wire [4-1:0] node2056;
	wire [4-1:0] node2059;
	wire [4-1:0] node2060;
	wire [4-1:0] node2062;
	wire [4-1:0] node2065;
	wire [4-1:0] node2066;
	wire [4-1:0] node2068;
	wire [4-1:0] node2072;
	wire [4-1:0] node2073;
	wire [4-1:0] node2074;
	wire [4-1:0] node2075;
	wire [4-1:0] node2077;
	wire [4-1:0] node2078;
	wire [4-1:0] node2082;
	wire [4-1:0] node2083;
	wire [4-1:0] node2087;
	wire [4-1:0] node2088;
	wire [4-1:0] node2089;
	wire [4-1:0] node2093;
	wire [4-1:0] node2096;
	wire [4-1:0] node2097;
	wire [4-1:0] node2098;
	wire [4-1:0] node2099;
	wire [4-1:0] node2101;
	wire [4-1:0] node2105;
	wire [4-1:0] node2106;
	wire [4-1:0] node2110;
	wire [4-1:0] node2111;
	wire [4-1:0] node2112;
	wire [4-1:0] node2113;
	wire [4-1:0] node2116;
	wire [4-1:0] node2119;
	wire [4-1:0] node2120;
	wire [4-1:0] node2124;
	wire [4-1:0] node2125;
	wire [4-1:0] node2126;
	wire [4-1:0] node2131;
	wire [4-1:0] node2132;
	wire [4-1:0] node2133;
	wire [4-1:0] node2134;
	wire [4-1:0] node2135;
	wire [4-1:0] node2136;
	wire [4-1:0] node2138;
	wire [4-1:0] node2140;
	wire [4-1:0] node2143;
	wire [4-1:0] node2145;
	wire [4-1:0] node2146;
	wire [4-1:0] node2150;
	wire [4-1:0] node2151;
	wire [4-1:0] node2152;
	wire [4-1:0] node2153;
	wire [4-1:0] node2157;
	wire [4-1:0] node2158;
	wire [4-1:0] node2162;
	wire [4-1:0] node2163;
	wire [4-1:0] node2167;
	wire [4-1:0] node2168;
	wire [4-1:0] node2169;
	wire [4-1:0] node2170;
	wire [4-1:0] node2171;
	wire [4-1:0] node2175;
	wire [4-1:0] node2176;
	wire [4-1:0] node2179;
	wire [4-1:0] node2183;
	wire [4-1:0] node2184;
	wire [4-1:0] node2185;
	wire [4-1:0] node2187;
	wire [4-1:0] node2191;
	wire [4-1:0] node2193;
	wire [4-1:0] node2196;
	wire [4-1:0] node2197;
	wire [4-1:0] node2198;
	wire [4-1:0] node2199;
	wire [4-1:0] node2200;
	wire [4-1:0] node2202;
	wire [4-1:0] node2205;
	wire [4-1:0] node2209;
	wire [4-1:0] node2210;
	wire [4-1:0] node2213;
	wire [4-1:0] node2214;
	wire [4-1:0] node2217;
	wire [4-1:0] node2219;
	wire [4-1:0] node2222;
	wire [4-1:0] node2223;
	wire [4-1:0] node2224;
	wire [4-1:0] node2225;
	wire [4-1:0] node2226;
	wire [4-1:0] node2231;
	wire [4-1:0] node2232;
	wire [4-1:0] node2233;
	wire [4-1:0] node2238;
	wire [4-1:0] node2240;
	wire [4-1:0] node2241;
	wire [4-1:0] node2242;
	wire [4-1:0] node2246;
	wire [4-1:0] node2249;
	wire [4-1:0] node2250;
	wire [4-1:0] node2251;
	wire [4-1:0] node2252;
	wire [4-1:0] node2253;
	wire [4-1:0] node2254;
	wire [4-1:0] node2256;
	wire [4-1:0] node2260;
	wire [4-1:0] node2263;
	wire [4-1:0] node2264;
	wire [4-1:0] node2265;
	wire [4-1:0] node2266;
	wire [4-1:0] node2270;
	wire [4-1:0] node2271;
	wire [4-1:0] node2275;
	wire [4-1:0] node2276;
	wire [4-1:0] node2277;
	wire [4-1:0] node2280;
	wire [4-1:0] node2284;
	wire [4-1:0] node2285;
	wire [4-1:0] node2286;
	wire [4-1:0] node2289;
	wire [4-1:0] node2290;
	wire [4-1:0] node2291;
	wire [4-1:0] node2294;
	wire [4-1:0] node2298;
	wire [4-1:0] node2299;
	wire [4-1:0] node2300;
	wire [4-1:0] node2301;
	wire [4-1:0] node2305;
	wire [4-1:0] node2307;
	wire [4-1:0] node2310;
	wire [4-1:0] node2311;
	wire [4-1:0] node2314;
	wire [4-1:0] node2316;
	wire [4-1:0] node2319;
	wire [4-1:0] node2320;
	wire [4-1:0] node2321;
	wire [4-1:0] node2322;
	wire [4-1:0] node2325;
	wire [4-1:0] node2326;
	wire [4-1:0] node2327;
	wire [4-1:0] node2331;
	wire [4-1:0] node2332;
	wire [4-1:0] node2336;
	wire [4-1:0] node2337;
	wire [4-1:0] node2339;
	wire [4-1:0] node2342;
	wire [4-1:0] node2344;
	wire [4-1:0] node2347;
	wire [4-1:0] node2348;
	wire [4-1:0] node2349;
	wire [4-1:0] node2351;
	wire [4-1:0] node2354;
	wire [4-1:0] node2355;
	wire [4-1:0] node2357;
	wire [4-1:0] node2361;
	wire [4-1:0] node2362;
	wire [4-1:0] node2363;
	wire [4-1:0] node2364;
	wire [4-1:0] node2368;
	wire [4-1:0] node2371;
	wire [4-1:0] node2372;
	wire [4-1:0] node2376;
	wire [4-1:0] node2377;
	wire [4-1:0] node2378;
	wire [4-1:0] node2379;
	wire [4-1:0] node2380;
	wire [4-1:0] node2381;
	wire [4-1:0] node2382;
	wire [4-1:0] node2383;
	wire [4-1:0] node2385;
	wire [4-1:0] node2390;
	wire [4-1:0] node2391;
	wire [4-1:0] node2392;
	wire [4-1:0] node2394;
	wire [4-1:0] node2397;
	wire [4-1:0] node2400;
	wire [4-1:0] node2402;
	wire [4-1:0] node2403;
	wire [4-1:0] node2407;
	wire [4-1:0] node2408;
	wire [4-1:0] node2409;
	wire [4-1:0] node2410;
	wire [4-1:0] node2413;
	wire [4-1:0] node2415;
	wire [4-1:0] node2418;
	wire [4-1:0] node2420;
	wire [4-1:0] node2422;
	wire [4-1:0] node2425;
	wire [4-1:0] node2426;
	wire [4-1:0] node2428;
	wire [4-1:0] node2429;
	wire [4-1:0] node2432;
	wire [4-1:0] node2435;
	wire [4-1:0] node2436;
	wire [4-1:0] node2437;
	wire [4-1:0] node2441;
	wire [4-1:0] node2442;
	wire [4-1:0] node2446;
	wire [4-1:0] node2447;
	wire [4-1:0] node2448;
	wire [4-1:0] node2449;
	wire [4-1:0] node2451;
	wire [4-1:0] node2453;
	wire [4-1:0] node2457;
	wire [4-1:0] node2458;
	wire [4-1:0] node2461;
	wire [4-1:0] node2462;
	wire [4-1:0] node2466;
	wire [4-1:0] node2467;
	wire [4-1:0] node2468;
	wire [4-1:0] node2469;
	wire [4-1:0] node2473;
	wire [4-1:0] node2474;
	wire [4-1:0] node2476;
	wire [4-1:0] node2479;
	wire [4-1:0] node2481;
	wire [4-1:0] node2484;
	wire [4-1:0] node2486;
	wire [4-1:0] node2489;
	wire [4-1:0] node2490;
	wire [4-1:0] node2491;
	wire [4-1:0] node2492;
	wire [4-1:0] node2493;
	wire [4-1:0] node2495;
	wire [4-1:0] node2496;
	wire [4-1:0] node2500;
	wire [4-1:0] node2501;
	wire [4-1:0] node2503;
	wire [4-1:0] node2506;
	wire [4-1:0] node2508;
	wire [4-1:0] node2511;
	wire [4-1:0] node2512;
	wire [4-1:0] node2515;
	wire [4-1:0] node2516;
	wire [4-1:0] node2518;
	wire [4-1:0] node2522;
	wire [4-1:0] node2523;
	wire [4-1:0] node2524;
	wire [4-1:0] node2526;
	wire [4-1:0] node2527;
	wire [4-1:0] node2531;
	wire [4-1:0] node2534;
	wire [4-1:0] node2535;
	wire [4-1:0] node2536;
	wire [4-1:0] node2539;
	wire [4-1:0] node2542;
	wire [4-1:0] node2543;
	wire [4-1:0] node2544;
	wire [4-1:0] node2548;
	wire [4-1:0] node2550;
	wire [4-1:0] node2553;
	wire [4-1:0] node2554;
	wire [4-1:0] node2555;
	wire [4-1:0] node2556;
	wire [4-1:0] node2557;
	wire [4-1:0] node2559;
	wire [4-1:0] node2563;
	wire [4-1:0] node2564;
	wire [4-1:0] node2566;
	wire [4-1:0] node2569;
	wire [4-1:0] node2570;
	wire [4-1:0] node2574;
	wire [4-1:0] node2575;
	wire [4-1:0] node2578;
	wire [4-1:0] node2581;
	wire [4-1:0] node2582;
	wire [4-1:0] node2583;
	wire [4-1:0] node2584;
	wire [4-1:0] node2588;
	wire [4-1:0] node2589;
	wire [4-1:0] node2590;
	wire [4-1:0] node2594;
	wire [4-1:0] node2595;
	wire [4-1:0] node2599;
	wire [4-1:0] node2600;
	wire [4-1:0] node2602;
	wire [4-1:0] node2604;
	wire [4-1:0] node2607;
	wire [4-1:0] node2608;
	wire [4-1:0] node2610;
	wire [4-1:0] node2613;
	wire [4-1:0] node2615;
	wire [4-1:0] node2618;
	wire [4-1:0] node2619;
	wire [4-1:0] node2620;
	wire [4-1:0] node2621;
	wire [4-1:0] node2622;
	wire [4-1:0] node2623;
	wire [4-1:0] node2624;
	wire [4-1:0] node2625;
	wire [4-1:0] node2628;
	wire [4-1:0] node2633;
	wire [4-1:0] node2634;
	wire [4-1:0] node2635;
	wire [4-1:0] node2637;
	wire [4-1:0] node2640;
	wire [4-1:0] node2643;
	wire [4-1:0] node2645;
	wire [4-1:0] node2646;
	wire [4-1:0] node2649;
	wire [4-1:0] node2652;
	wire [4-1:0] node2653;
	wire [4-1:0] node2654;
	wire [4-1:0] node2655;
	wire [4-1:0] node2658;
	wire [4-1:0] node2660;
	wire [4-1:0] node2664;
	wire [4-1:0] node2666;
	wire [4-1:0] node2667;
	wire [4-1:0] node2668;
	wire [4-1:0] node2672;
	wire [4-1:0] node2673;
	wire [4-1:0] node2677;
	wire [4-1:0] node2678;
	wire [4-1:0] node2679;
	wire [4-1:0] node2680;
	wire [4-1:0] node2681;
	wire [4-1:0] node2685;
	wire [4-1:0] node2686;
	wire [4-1:0] node2689;
	wire [4-1:0] node2692;
	wire [4-1:0] node2693;
	wire [4-1:0] node2695;
	wire [4-1:0] node2697;
	wire [4-1:0] node2700;
	wire [4-1:0] node2701;
	wire [4-1:0] node2705;
	wire [4-1:0] node2706;
	wire [4-1:0] node2707;
	wire [4-1:0] node2708;
	wire [4-1:0] node2712;
	wire [4-1:0] node2714;
	wire [4-1:0] node2717;
	wire [4-1:0] node2718;
	wire [4-1:0] node2719;
	wire [4-1:0] node2722;
	wire [4-1:0] node2725;
	wire [4-1:0] node2726;
	wire [4-1:0] node2728;
	wire [4-1:0] node2731;
	wire [4-1:0] node2733;
	wire [4-1:0] node2736;
	wire [4-1:0] node2737;
	wire [4-1:0] node2738;
	wire [4-1:0] node2739;
	wire [4-1:0] node2740;
	wire [4-1:0] node2741;
	wire [4-1:0] node2743;
	wire [4-1:0] node2746;
	wire [4-1:0] node2748;
	wire [4-1:0] node2751;
	wire [4-1:0] node2752;
	wire [4-1:0] node2753;
	wire [4-1:0] node2756;
	wire [4-1:0] node2760;
	wire [4-1:0] node2761;
	wire [4-1:0] node2763;
	wire [4-1:0] node2764;
	wire [4-1:0] node2768;
	wire [4-1:0] node2770;
	wire [4-1:0] node2771;
	wire [4-1:0] node2775;
	wire [4-1:0] node2776;
	wire [4-1:0] node2777;
	wire [4-1:0] node2780;
	wire [4-1:0] node2782;
	wire [4-1:0] node2785;
	wire [4-1:0] node2786;
	wire [4-1:0] node2787;
	wire [4-1:0] node2788;
	wire [4-1:0] node2791;
	wire [4-1:0] node2796;
	wire [4-1:0] node2797;
	wire [4-1:0] node2798;
	wire [4-1:0] node2799;
	wire [4-1:0] node2800;
	wire [4-1:0] node2804;
	wire [4-1:0] node2807;
	wire [4-1:0] node2809;
	wire [4-1:0] node2811;
	wire [4-1:0] node2814;
	wire [4-1:0] node2815;
	wire [4-1:0] node2816;
	wire [4-1:0] node2817;
	wire [4-1:0] node2821;
	wire [4-1:0] node2822;
	wire [4-1:0] node2823;
	wire [4-1:0] node2828;
	wire [4-1:0] node2829;
	wire [4-1:0] node2831;
	wire [4-1:0] node2832;
	wire [4-1:0] node2836;
	wire [4-1:0] node2837;
	wire [4-1:0] node2838;
	wire [4-1:0] node2841;
	wire [4-1:0] node2844;
	wire [4-1:0] node2845;
	wire [4-1:0] node2849;
	wire [4-1:0] node2850;
	wire [4-1:0] node2851;
	wire [4-1:0] node2852;
	wire [4-1:0] node2853;
	wire [4-1:0] node2854;
	wire [4-1:0] node2855;
	wire [4-1:0] node2856;
	wire [4-1:0] node2858;
	wire [4-1:0] node2861;
	wire [4-1:0] node2862;
	wire [4-1:0] node2865;
	wire [4-1:0] node2867;
	wire [4-1:0] node2870;
	wire [4-1:0] node2871;
	wire [4-1:0] node2873;
	wire [4-1:0] node2875;
	wire [4-1:0] node2878;
	wire [4-1:0] node2879;
	wire [4-1:0] node2883;
	wire [4-1:0] node2884;
	wire [4-1:0] node2885;
	wire [4-1:0] node2886;
	wire [4-1:0] node2888;
	wire [4-1:0] node2893;
	wire [4-1:0] node2894;
	wire [4-1:0] node2895;
	wire [4-1:0] node2899;
	wire [4-1:0] node2902;
	wire [4-1:0] node2903;
	wire [4-1:0] node2904;
	wire [4-1:0] node2905;
	wire [4-1:0] node2906;
	wire [4-1:0] node2910;
	wire [4-1:0] node2911;
	wire [4-1:0] node2914;
	wire [4-1:0] node2915;
	wire [4-1:0] node2919;
	wire [4-1:0] node2920;
	wire [4-1:0] node2922;
	wire [4-1:0] node2924;
	wire [4-1:0] node2927;
	wire [4-1:0] node2930;
	wire [4-1:0] node2931;
	wire [4-1:0] node2932;
	wire [4-1:0] node2935;
	wire [4-1:0] node2936;
	wire [4-1:0] node2937;
	wire [4-1:0] node2942;
	wire [4-1:0] node2943;
	wire [4-1:0] node2945;
	wire [4-1:0] node2946;
	wire [4-1:0] node2950;
	wire [4-1:0] node2951;
	wire [4-1:0] node2952;
	wire [4-1:0] node2956;
	wire [4-1:0] node2957;
	wire [4-1:0] node2961;
	wire [4-1:0] node2962;
	wire [4-1:0] node2963;
	wire [4-1:0] node2964;
	wire [4-1:0] node2965;
	wire [4-1:0] node2967;
	wire [4-1:0] node2968;
	wire [4-1:0] node2971;
	wire [4-1:0] node2974;
	wire [4-1:0] node2976;
	wire [4-1:0] node2977;
	wire [4-1:0] node2980;
	wire [4-1:0] node2983;
	wire [4-1:0] node2984;
	wire [4-1:0] node2986;
	wire [4-1:0] node2988;
	wire [4-1:0] node2991;
	wire [4-1:0] node2992;
	wire [4-1:0] node2993;
	wire [4-1:0] node2998;
	wire [4-1:0] node2999;
	wire [4-1:0] node3000;
	wire [4-1:0] node3003;
	wire [4-1:0] node3004;
	wire [4-1:0] node3007;
	wire [4-1:0] node3010;
	wire [4-1:0] node3012;
	wire [4-1:0] node3013;
	wire [4-1:0] node3014;
	wire [4-1:0] node3017;
	wire [4-1:0] node3021;
	wire [4-1:0] node3022;
	wire [4-1:0] node3023;
	wire [4-1:0] node3025;
	wire [4-1:0] node3026;
	wire [4-1:0] node3028;
	wire [4-1:0] node3032;
	wire [4-1:0] node3034;
	wire [4-1:0] node3035;
	wire [4-1:0] node3036;
	wire [4-1:0] node3039;
	wire [4-1:0] node3042;
	wire [4-1:0] node3044;
	wire [4-1:0] node3047;
	wire [4-1:0] node3048;
	wire [4-1:0] node3049;
	wire [4-1:0] node3050;
	wire [4-1:0] node3052;
	wire [4-1:0] node3056;
	wire [4-1:0] node3057;
	wire [4-1:0] node3061;
	wire [4-1:0] node3063;
	wire [4-1:0] node3065;
	wire [4-1:0] node3066;
	wire [4-1:0] node3070;
	wire [4-1:0] node3071;
	wire [4-1:0] node3072;
	wire [4-1:0] node3073;
	wire [4-1:0] node3074;
	wire [4-1:0] node3075;
	wire [4-1:0] node3077;
	wire [4-1:0] node3079;
	wire [4-1:0] node3082;
	wire [4-1:0] node3083;
	wire [4-1:0] node3086;
	wire [4-1:0] node3089;
	wire [4-1:0] node3090;
	wire [4-1:0] node3091;
	wire [4-1:0] node3092;
	wire [4-1:0] node3097;
	wire [4-1:0] node3098;
	wire [4-1:0] node3099;
	wire [4-1:0] node3103;
	wire [4-1:0] node3106;
	wire [4-1:0] node3107;
	wire [4-1:0] node3108;
	wire [4-1:0] node3109;
	wire [4-1:0] node3112;
	wire [4-1:0] node3114;
	wire [4-1:0] node3118;
	wire [4-1:0] node3119;
	wire [4-1:0] node3121;
	wire [4-1:0] node3122;
	wire [4-1:0] node3126;
	wire [4-1:0] node3129;
	wire [4-1:0] node3130;
	wire [4-1:0] node3131;
	wire [4-1:0] node3132;
	wire [4-1:0] node3133;
	wire [4-1:0] node3135;
	wire [4-1:0] node3139;
	wire [4-1:0] node3140;
	wire [4-1:0] node3143;
	wire [4-1:0] node3146;
	wire [4-1:0] node3147;
	wire [4-1:0] node3149;
	wire [4-1:0] node3150;
	wire [4-1:0] node3154;
	wire [4-1:0] node3157;
	wire [4-1:0] node3158;
	wire [4-1:0] node3159;
	wire [4-1:0] node3160;
	wire [4-1:0] node3164;
	wire [4-1:0] node3167;
	wire [4-1:0] node3168;
	wire [4-1:0] node3169;
	wire [4-1:0] node3171;
	wire [4-1:0] node3174;
	wire [4-1:0] node3176;
	wire [4-1:0] node3179;
	wire [4-1:0] node3181;
	wire [4-1:0] node3182;
	wire [4-1:0] node3186;
	wire [4-1:0] node3187;
	wire [4-1:0] node3188;
	wire [4-1:0] node3189;
	wire [4-1:0] node3190;
	wire [4-1:0] node3191;
	wire [4-1:0] node3195;
	wire [4-1:0] node3198;
	wire [4-1:0] node3200;
	wire [4-1:0] node3201;
	wire [4-1:0] node3202;
	wire [4-1:0] node3205;
	wire [4-1:0] node3208;
	wire [4-1:0] node3211;
	wire [4-1:0] node3212;
	wire [4-1:0] node3213;
	wire [4-1:0] node3214;
	wire [4-1:0] node3218;
	wire [4-1:0] node3219;
	wire [4-1:0] node3223;
	wire [4-1:0] node3225;
	wire [4-1:0] node3227;
	wire [4-1:0] node3230;
	wire [4-1:0] node3231;
	wire [4-1:0] node3232;
	wire [4-1:0] node3233;
	wire [4-1:0] node3234;
	wire [4-1:0] node3237;
	wire [4-1:0] node3238;
	wire [4-1:0] node3242;
	wire [4-1:0] node3243;
	wire [4-1:0] node3244;
	wire [4-1:0] node3248;
	wire [4-1:0] node3250;
	wire [4-1:0] node3253;
	wire [4-1:0] node3254;
	wire [4-1:0] node3256;
	wire [4-1:0] node3259;
	wire [4-1:0] node3260;
	wire [4-1:0] node3263;
	wire [4-1:0] node3264;
	wire [4-1:0] node3268;
	wire [4-1:0] node3269;
	wire [4-1:0] node3270;
	wire [4-1:0] node3271;
	wire [4-1:0] node3274;
	wire [4-1:0] node3275;
	wire [4-1:0] node3279;
	wire [4-1:0] node3282;
	wire [4-1:0] node3284;
	wire [4-1:0] node3285;
	wire [4-1:0] node3287;
	wire [4-1:0] node3291;
	wire [4-1:0] node3292;
	wire [4-1:0] node3293;
	wire [4-1:0] node3294;
	wire [4-1:0] node3295;
	wire [4-1:0] node3296;
	wire [4-1:0] node3298;
	wire [4-1:0] node3301;
	wire [4-1:0] node3303;
	wire [4-1:0] node3305;
	wire [4-1:0] node3306;
	wire [4-1:0] node3310;
	wire [4-1:0] node3311;
	wire [4-1:0] node3312;
	wire [4-1:0] node3314;
	wire [4-1:0] node3318;
	wire [4-1:0] node3319;
	wire [4-1:0] node3322;
	wire [4-1:0] node3325;
	wire [4-1:0] node3326;
	wire [4-1:0] node3327;
	wire [4-1:0] node3328;
	wire [4-1:0] node3330;
	wire [4-1:0] node3332;
	wire [4-1:0] node3335;
	wire [4-1:0] node3336;
	wire [4-1:0] node3339;
	wire [4-1:0] node3342;
	wire [4-1:0] node3343;
	wire [4-1:0] node3344;
	wire [4-1:0] node3347;
	wire [4-1:0] node3350;
	wire [4-1:0] node3351;
	wire [4-1:0] node3353;
	wire [4-1:0] node3356;
	wire [4-1:0] node3358;
	wire [4-1:0] node3361;
	wire [4-1:0] node3362;
	wire [4-1:0] node3363;
	wire [4-1:0] node3364;
	wire [4-1:0] node3368;
	wire [4-1:0] node3371;
	wire [4-1:0] node3372;
	wire [4-1:0] node3373;
	wire [4-1:0] node3375;
	wire [4-1:0] node3378;
	wire [4-1:0] node3379;
	wire [4-1:0] node3383;
	wire [4-1:0] node3386;
	wire [4-1:0] node3387;
	wire [4-1:0] node3388;
	wire [4-1:0] node3389;
	wire [4-1:0] node3391;
	wire [4-1:0] node3392;
	wire [4-1:0] node3396;
	wire [4-1:0] node3397;
	wire [4-1:0] node3398;
	wire [4-1:0] node3399;
	wire [4-1:0] node3403;
	wire [4-1:0] node3406;
	wire [4-1:0] node3408;
	wire [4-1:0] node3409;
	wire [4-1:0] node3413;
	wire [4-1:0] node3414;
	wire [4-1:0] node3415;
	wire [4-1:0] node3417;
	wire [4-1:0] node3418;
	wire [4-1:0] node3421;
	wire [4-1:0] node3424;
	wire [4-1:0] node3425;
	wire [4-1:0] node3429;
	wire [4-1:0] node3430;
	wire [4-1:0] node3432;
	wire [4-1:0] node3435;
	wire [4-1:0] node3438;
	wire [4-1:0] node3439;
	wire [4-1:0] node3440;
	wire [4-1:0] node3441;
	wire [4-1:0] node3442;
	wire [4-1:0] node3446;
	wire [4-1:0] node3448;
	wire [4-1:0] node3449;
	wire [4-1:0] node3453;
	wire [4-1:0] node3454;
	wire [4-1:0] node3457;
	wire [4-1:0] node3460;
	wire [4-1:0] node3461;
	wire [4-1:0] node3462;
	wire [4-1:0] node3463;
	wire [4-1:0] node3464;
	wire [4-1:0] node3470;
	wire [4-1:0] node3471;
	wire [4-1:0] node3472;
	wire [4-1:0] node3473;
	wire [4-1:0] node3478;
	wire [4-1:0] node3479;
	wire [4-1:0] node3483;
	wire [4-1:0] node3484;
	wire [4-1:0] node3485;
	wire [4-1:0] node3486;
	wire [4-1:0] node3487;
	wire [4-1:0] node3488;
	wire [4-1:0] node3490;
	wire [4-1:0] node3491;
	wire [4-1:0] node3496;
	wire [4-1:0] node3497;
	wire [4-1:0] node3499;
	wire [4-1:0] node3502;
	wire [4-1:0] node3503;
	wire [4-1:0] node3505;
	wire [4-1:0] node3508;
	wire [4-1:0] node3511;
	wire [4-1:0] node3512;
	wire [4-1:0] node3513;
	wire [4-1:0] node3515;
	wire [4-1:0] node3518;
	wire [4-1:0] node3519;
	wire [4-1:0] node3523;
	wire [4-1:0] node3524;
	wire [4-1:0] node3525;
	wire [4-1:0] node3526;
	wire [4-1:0] node3531;
	wire [4-1:0] node3532;
	wire [4-1:0] node3536;
	wire [4-1:0] node3537;
	wire [4-1:0] node3538;
	wire [4-1:0] node3539;
	wire [4-1:0] node3541;
	wire [4-1:0] node3544;
	wire [4-1:0] node3546;
	wire [4-1:0] node3547;
	wire [4-1:0] node3550;
	wire [4-1:0] node3553;
	wire [4-1:0] node3554;
	wire [4-1:0] node3556;
	wire [4-1:0] node3559;
	wire [4-1:0] node3560;
	wire [4-1:0] node3561;
	wire [4-1:0] node3565;
	wire [4-1:0] node3566;
	wire [4-1:0] node3570;
	wire [4-1:0] node3571;
	wire [4-1:0] node3572;
	wire [4-1:0] node3573;
	wire [4-1:0] node3574;
	wire [4-1:0] node3578;
	wire [4-1:0] node3580;
	wire [4-1:0] node3583;
	wire [4-1:0] node3584;
	wire [4-1:0] node3585;
	wire [4-1:0] node3588;
	wire [4-1:0] node3591;
	wire [4-1:0] node3592;
	wire [4-1:0] node3595;
	wire [4-1:0] node3598;
	wire [4-1:0] node3599;
	wire [4-1:0] node3600;
	wire [4-1:0] node3601;
	wire [4-1:0] node3605;
	wire [4-1:0] node3606;
	wire [4-1:0] node3610;
	wire [4-1:0] node3611;
	wire [4-1:0] node3613;
	wire [4-1:0] node3616;
	wire [4-1:0] node3617;
	wire [4-1:0] node3620;
	wire [4-1:0] node3623;
	wire [4-1:0] node3624;
	wire [4-1:0] node3625;
	wire [4-1:0] node3626;
	wire [4-1:0] node3627;
	wire [4-1:0] node3628;
	wire [4-1:0] node3630;
	wire [4-1:0] node3634;
	wire [4-1:0] node3636;
	wire [4-1:0] node3639;
	wire [4-1:0] node3640;
	wire [4-1:0] node3643;
	wire [4-1:0] node3644;
	wire [4-1:0] node3646;
	wire [4-1:0] node3649;
	wire [4-1:0] node3652;
	wire [4-1:0] node3653;
	wire [4-1:0] node3654;
	wire [4-1:0] node3655;
	wire [4-1:0] node3660;
	wire [4-1:0] node3661;
	wire [4-1:0] node3662;
	wire [4-1:0] node3667;
	wire [4-1:0] node3668;
	wire [4-1:0] node3669;
	wire [4-1:0] node3670;
	wire [4-1:0] node3671;
	wire [4-1:0] node3676;
	wire [4-1:0] node3677;
	wire [4-1:0] node3678;
	wire [4-1:0] node3679;
	wire [4-1:0] node3682;
	wire [4-1:0] node3686;
	wire [4-1:0] node3687;
	wire [4-1:0] node3688;
	wire [4-1:0] node3693;
	wire [4-1:0] node3694;
	wire [4-1:0] node3695;
	wire [4-1:0] node3698;
	wire [4-1:0] node3699;
	wire [4-1:0] node3703;
	wire [4-1:0] node3705;
	wire [4-1:0] node3708;
	wire [4-1:0] node3709;
	wire [4-1:0] node3710;
	wire [4-1:0] node3711;
	wire [4-1:0] node3712;
	wire [4-1:0] node3713;
	wire [4-1:0] node3714;
	wire [4-1:0] node3715;
	wire [4-1:0] node3716;
	wire [4-1:0] node3717;
	wire [4-1:0] node3719;
	wire [4-1:0] node3722;
	wire [4-1:0] node3723;
	wire [4-1:0] node3727;
	wire [4-1:0] node3728;
	wire [4-1:0] node3730;
	wire [4-1:0] node3734;
	wire [4-1:0] node3735;
	wire [4-1:0] node3736;
	wire [4-1:0] node3740;
	wire [4-1:0] node3741;
	wire [4-1:0] node3743;
	wire [4-1:0] node3744;
	wire [4-1:0] node3749;
	wire [4-1:0] node3750;
	wire [4-1:0] node3751;
	wire [4-1:0] node3752;
	wire [4-1:0] node3755;
	wire [4-1:0] node3756;
	wire [4-1:0] node3757;
	wire [4-1:0] node3762;
	wire [4-1:0] node3763;
	wire [4-1:0] node3764;
	wire [4-1:0] node3767;
	wire [4-1:0] node3768;
	wire [4-1:0] node3772;
	wire [4-1:0] node3773;
	wire [4-1:0] node3776;
	wire [4-1:0] node3778;
	wire [4-1:0] node3781;
	wire [4-1:0] node3782;
	wire [4-1:0] node3783;
	wire [4-1:0] node3784;
	wire [4-1:0] node3788;
	wire [4-1:0] node3790;
	wire [4-1:0] node3793;
	wire [4-1:0] node3794;
	wire [4-1:0] node3797;
	wire [4-1:0] node3800;
	wire [4-1:0] node3801;
	wire [4-1:0] node3802;
	wire [4-1:0] node3803;
	wire [4-1:0] node3804;
	wire [4-1:0] node3805;
	wire [4-1:0] node3807;
	wire [4-1:0] node3810;
	wire [4-1:0] node3813;
	wire [4-1:0] node3814;
	wire [4-1:0] node3817;
	wire [4-1:0] node3819;
	wire [4-1:0] node3822;
	wire [4-1:0] node3823;
	wire [4-1:0] node3825;
	wire [4-1:0] node3827;
	wire [4-1:0] node3830;
	wire [4-1:0] node3831;
	wire [4-1:0] node3834;
	wire [4-1:0] node3837;
	wire [4-1:0] node3838;
	wire [4-1:0] node3839;
	wire [4-1:0] node3840;
	wire [4-1:0] node3843;
	wire [4-1:0] node3844;
	wire [4-1:0] node3848;
	wire [4-1:0] node3851;
	wire [4-1:0] node3852;
	wire [4-1:0] node3853;
	wire [4-1:0] node3855;
	wire [4-1:0] node3859;
	wire [4-1:0] node3861;
	wire [4-1:0] node3864;
	wire [4-1:0] node3865;
	wire [4-1:0] node3866;
	wire [4-1:0] node3867;
	wire [4-1:0] node3868;
	wire [4-1:0] node3872;
	wire [4-1:0] node3874;
	wire [4-1:0] node3877;
	wire [4-1:0] node3878;
	wire [4-1:0] node3879;
	wire [4-1:0] node3882;
	wire [4-1:0] node3885;
	wire [4-1:0] node3888;
	wire [4-1:0] node3889;
	wire [4-1:0] node3890;
	wire [4-1:0] node3891;
	wire [4-1:0] node3894;
	wire [4-1:0] node3895;
	wire [4-1:0] node3899;
	wire [4-1:0] node3901;
	wire [4-1:0] node3902;
	wire [4-1:0] node3905;
	wire [4-1:0] node3908;
	wire [4-1:0] node3909;
	wire [4-1:0] node3910;
	wire [4-1:0] node3914;
	wire [4-1:0] node3915;
	wire [4-1:0] node3918;
	wire [4-1:0] node3921;
	wire [4-1:0] node3922;
	wire [4-1:0] node3923;
	wire [4-1:0] node3924;
	wire [4-1:0] node3925;
	wire [4-1:0] node3926;
	wire [4-1:0] node3927;
	wire [4-1:0] node3931;
	wire [4-1:0] node3932;
	wire [4-1:0] node3933;
	wire [4-1:0] node3936;
	wire [4-1:0] node3940;
	wire [4-1:0] node3942;
	wire [4-1:0] node3943;
	wire [4-1:0] node3944;
	wire [4-1:0] node3949;
	wire [4-1:0] node3950;
	wire [4-1:0] node3952;
	wire [4-1:0] node3954;
	wire [4-1:0] node3956;
	wire [4-1:0] node3959;
	wire [4-1:0] node3960;
	wire [4-1:0] node3962;
	wire [4-1:0] node3965;
	wire [4-1:0] node3966;
	wire [4-1:0] node3969;
	wire [4-1:0] node3972;
	wire [4-1:0] node3973;
	wire [4-1:0] node3974;
	wire [4-1:0] node3975;
	wire [4-1:0] node3977;
	wire [4-1:0] node3980;
	wire [4-1:0] node3981;
	wire [4-1:0] node3982;
	wire [4-1:0] node3986;
	wire [4-1:0] node3989;
	wire [4-1:0] node3992;
	wire [4-1:0] node3993;
	wire [4-1:0] node3994;
	wire [4-1:0] node3995;
	wire [4-1:0] node3997;
	wire [4-1:0] node4000;
	wire [4-1:0] node4004;
	wire [4-1:0] node4005;
	wire [4-1:0] node4007;
	wire [4-1:0] node4010;
	wire [4-1:0] node4012;
	wire [4-1:0] node4015;
	wire [4-1:0] node4016;
	wire [4-1:0] node4017;
	wire [4-1:0] node4018;
	wire [4-1:0] node4019;
	wire [4-1:0] node4021;
	wire [4-1:0] node4024;
	wire [4-1:0] node4027;
	wire [4-1:0] node4028;
	wire [4-1:0] node4029;
	wire [4-1:0] node4031;
	wire [4-1:0] node4034;
	wire [4-1:0] node4037;
	wire [4-1:0] node4038;
	wire [4-1:0] node4042;
	wire [4-1:0] node4043;
	wire [4-1:0] node4044;
	wire [4-1:0] node4045;
	wire [4-1:0] node4046;
	wire [4-1:0] node4050;
	wire [4-1:0] node4053;
	wire [4-1:0] node4055;
	wire [4-1:0] node4056;
	wire [4-1:0] node4060;
	wire [4-1:0] node4061;
	wire [4-1:0] node4062;
	wire [4-1:0] node4065;
	wire [4-1:0] node4066;
	wire [4-1:0] node4070;
	wire [4-1:0] node4072;
	wire [4-1:0] node4074;
	wire [4-1:0] node4077;
	wire [4-1:0] node4078;
	wire [4-1:0] node4079;
	wire [4-1:0] node4080;
	wire [4-1:0] node4082;
	wire [4-1:0] node4084;
	wire [4-1:0] node4088;
	wire [4-1:0] node4089;
	wire [4-1:0] node4091;
	wire [4-1:0] node4092;
	wire [4-1:0] node4095;
	wire [4-1:0] node4098;
	wire [4-1:0] node4099;
	wire [4-1:0] node4101;
	wire [4-1:0] node4104;
	wire [4-1:0] node4105;
	wire [4-1:0] node4108;
	wire [4-1:0] node4111;
	wire [4-1:0] node4112;
	wire [4-1:0] node4113;
	wire [4-1:0] node4114;
	wire [4-1:0] node4115;
	wire [4-1:0] node4119;
	wire [4-1:0] node4122;
	wire [4-1:0] node4123;
	wire [4-1:0] node4127;
	wire [4-1:0] node4128;
	wire [4-1:0] node4129;
	wire [4-1:0] node4130;
	wire [4-1:0] node4133;
	wire [4-1:0] node4136;
	wire [4-1:0] node4137;
	wire [4-1:0] node4141;
	wire [4-1:0] node4142;
	wire [4-1:0] node4144;
	wire [4-1:0] node4148;
	wire [4-1:0] node4149;
	wire [4-1:0] node4150;
	wire [4-1:0] node4151;
	wire [4-1:0] node4152;
	wire [4-1:0] node4153;
	wire [4-1:0] node4156;
	wire [4-1:0] node4157;
	wire [4-1:0] node4160;
	wire [4-1:0] node4161;
	wire [4-1:0] node4164;
	wire [4-1:0] node4165;
	wire [4-1:0] node4169;
	wire [4-1:0] node4170;
	wire [4-1:0] node4171;
	wire [4-1:0] node4174;
	wire [4-1:0] node4175;
	wire [4-1:0] node4177;
	wire [4-1:0] node4180;
	wire [4-1:0] node4183;
	wire [4-1:0] node4184;
	wire [4-1:0] node4186;
	wire [4-1:0] node4189;
	wire [4-1:0] node4191;
	wire [4-1:0] node4192;
	wire [4-1:0] node4196;
	wire [4-1:0] node4197;
	wire [4-1:0] node4198;
	wire [4-1:0] node4200;
	wire [4-1:0] node4201;
	wire [4-1:0] node4205;
	wire [4-1:0] node4206;
	wire [4-1:0] node4207;
	wire [4-1:0] node4209;
	wire [4-1:0] node4213;
	wire [4-1:0] node4214;
	wire [4-1:0] node4217;
	wire [4-1:0] node4218;
	wire [4-1:0] node4222;
	wire [4-1:0] node4223;
	wire [4-1:0] node4224;
	wire [4-1:0] node4226;
	wire [4-1:0] node4227;
	wire [4-1:0] node4231;
	wire [4-1:0] node4232;
	wire [4-1:0] node4234;
	wire [4-1:0] node4237;
	wire [4-1:0] node4240;
	wire [4-1:0] node4241;
	wire [4-1:0] node4244;
	wire [4-1:0] node4247;
	wire [4-1:0] node4248;
	wire [4-1:0] node4249;
	wire [4-1:0] node4251;
	wire [4-1:0] node4253;
	wire [4-1:0] node4255;
	wire [4-1:0] node4257;
	wire [4-1:0] node4260;
	wire [4-1:0] node4261;
	wire [4-1:0] node4263;
	wire [4-1:0] node4264;
	wire [4-1:0] node4267;
	wire [4-1:0] node4270;
	wire [4-1:0] node4271;
	wire [4-1:0] node4272;
	wire [4-1:0] node4273;
	wire [4-1:0] node4277;
	wire [4-1:0] node4280;
	wire [4-1:0] node4281;
	wire [4-1:0] node4283;
	wire [4-1:0] node4287;
	wire [4-1:0] node4288;
	wire [4-1:0] node4289;
	wire [4-1:0] node4290;
	wire [4-1:0] node4291;
	wire [4-1:0] node4294;
	wire [4-1:0] node4295;
	wire [4-1:0] node4299;
	wire [4-1:0] node4301;
	wire [4-1:0] node4303;
	wire [4-1:0] node4306;
	wire [4-1:0] node4307;
	wire [4-1:0] node4308;
	wire [4-1:0] node4310;
	wire [4-1:0] node4313;
	wire [4-1:0] node4317;
	wire [4-1:0] node4318;
	wire [4-1:0] node4319;
	wire [4-1:0] node4320;
	wire [4-1:0] node4323;
	wire [4-1:0] node4327;
	wire [4-1:0] node4328;
	wire [4-1:0] node4329;
	wire [4-1:0] node4332;
	wire [4-1:0] node4333;
	wire [4-1:0] node4337;
	wire [4-1:0] node4338;
	wire [4-1:0] node4342;
	wire [4-1:0] node4343;
	wire [4-1:0] node4344;
	wire [4-1:0] node4345;
	wire [4-1:0] node4346;
	wire [4-1:0] node4348;
	wire [4-1:0] node4349;
	wire [4-1:0] node4350;
	wire [4-1:0] node4354;
	wire [4-1:0] node4358;
	wire [4-1:0] node4359;
	wire [4-1:0] node4360;
	wire [4-1:0] node4361;
	wire [4-1:0] node4363;
	wire [4-1:0] node4367;
	wire [4-1:0] node4369;
	wire [4-1:0] node4371;
	wire [4-1:0] node4374;
	wire [4-1:0] node4375;
	wire [4-1:0] node4376;
	wire [4-1:0] node4380;
	wire [4-1:0] node4381;
	wire [4-1:0] node4382;
	wire [4-1:0] node4387;
	wire [4-1:0] node4388;
	wire [4-1:0] node4389;
	wire [4-1:0] node4390;
	wire [4-1:0] node4391;
	wire [4-1:0] node4392;
	wire [4-1:0] node4397;
	wire [4-1:0] node4399;
	wire [4-1:0] node4400;
	wire [4-1:0] node4403;
	wire [4-1:0] node4406;
	wire [4-1:0] node4407;
	wire [4-1:0] node4408;
	wire [4-1:0] node4409;
	wire [4-1:0] node4413;
	wire [4-1:0] node4416;
	wire [4-1:0] node4417;
	wire [4-1:0] node4419;
	wire [4-1:0] node4423;
	wire [4-1:0] node4424;
	wire [4-1:0] node4425;
	wire [4-1:0] node4427;
	wire [4-1:0] node4430;
	wire [4-1:0] node4432;
	wire [4-1:0] node4433;
	wire [4-1:0] node4436;
	wire [4-1:0] node4439;
	wire [4-1:0] node4440;
	wire [4-1:0] node4442;
	wire [4-1:0] node4443;
	wire [4-1:0] node4446;
	wire [4-1:0] node4450;
	wire [4-1:0] node4451;
	wire [4-1:0] node4452;
	wire [4-1:0] node4453;
	wire [4-1:0] node4454;
	wire [4-1:0] node4456;
	wire [4-1:0] node4459;
	wire [4-1:0] node4460;
	wire [4-1:0] node4463;
	wire [4-1:0] node4465;
	wire [4-1:0] node4468;
	wire [4-1:0] node4469;
	wire [4-1:0] node4472;
	wire [4-1:0] node4475;
	wire [4-1:0] node4476;
	wire [4-1:0] node4477;
	wire [4-1:0] node4479;
	wire [4-1:0] node4481;
	wire [4-1:0] node4484;
	wire [4-1:0] node4487;
	wire [4-1:0] node4488;
	wire [4-1:0] node4489;
	wire [4-1:0] node4490;
	wire [4-1:0] node4493;
	wire [4-1:0] node4497;
	wire [4-1:0] node4498;
	wire [4-1:0] node4502;
	wire [4-1:0] node4503;
	wire [4-1:0] node4504;
	wire [4-1:0] node4505;
	wire [4-1:0] node4506;
	wire [4-1:0] node4508;
	wire [4-1:0] node4511;
	wire [4-1:0] node4512;
	wire [4-1:0] node4516;
	wire [4-1:0] node4519;
	wire [4-1:0] node4522;
	wire [4-1:0] node4523;
	wire [4-1:0] node4524;
	wire [4-1:0] node4525;
	wire [4-1:0] node4526;
	wire [4-1:0] node4530;
	wire [4-1:0] node4531;
	wire [4-1:0] node4534;
	wire [4-1:0] node4537;
	wire [4-1:0] node4539;
	wire [4-1:0] node4541;
	wire [4-1:0] node4544;
	wire [4-1:0] node4545;
	wire [4-1:0] node4547;
	wire [4-1:0] node4548;
	wire [4-1:0] node4552;
	wire [4-1:0] node4555;
	wire [4-1:0] node4556;
	wire [4-1:0] node4557;
	wire [4-1:0] node4558;
	wire [4-1:0] node4559;
	wire [4-1:0] node4560;
	wire [4-1:0] node4561;
	wire [4-1:0] node4564;
	wire [4-1:0] node4565;
	wire [4-1:0] node4567;
	wire [4-1:0] node4570;
	wire [4-1:0] node4573;
	wire [4-1:0] node4574;
	wire [4-1:0] node4575;
	wire [4-1:0] node4577;
	wire [4-1:0] node4580;
	wire [4-1:0] node4583;
	wire [4-1:0] node4584;
	wire [4-1:0] node4585;
	wire [4-1:0] node4589;
	wire [4-1:0] node4590;
	wire [4-1:0] node4594;
	wire [4-1:0] node4595;
	wire [4-1:0] node4596;
	wire [4-1:0] node4598;
	wire [4-1:0] node4600;
	wire [4-1:0] node4601;
	wire [4-1:0] node4605;
	wire [4-1:0] node4606;
	wire [4-1:0] node4607;
	wire [4-1:0] node4608;
	wire [4-1:0] node4612;
	wire [4-1:0] node4615;
	wire [4-1:0] node4617;
	wire [4-1:0] node4620;
	wire [4-1:0] node4621;
	wire [4-1:0] node4622;
	wire [4-1:0] node4623;
	wire [4-1:0] node4626;
	wire [4-1:0] node4627;
	wire [4-1:0] node4632;
	wire [4-1:0] node4633;
	wire [4-1:0] node4636;
	wire [4-1:0] node4637;
	wire [4-1:0] node4638;
	wire [4-1:0] node4643;
	wire [4-1:0] node4644;
	wire [4-1:0] node4645;
	wire [4-1:0] node4646;
	wire [4-1:0] node4647;
	wire [4-1:0] node4648;
	wire [4-1:0] node4649;
	wire [4-1:0] node4652;
	wire [4-1:0] node4656;
	wire [4-1:0] node4657;
	wire [4-1:0] node4658;
	wire [4-1:0] node4661;
	wire [4-1:0] node4665;
	wire [4-1:0] node4666;
	wire [4-1:0] node4668;
	wire [4-1:0] node4670;
	wire [4-1:0] node4673;
	wire [4-1:0] node4676;
	wire [4-1:0] node4677;
	wire [4-1:0] node4678;
	wire [4-1:0] node4681;
	wire [4-1:0] node4682;
	wire [4-1:0] node4685;
	wire [4-1:0] node4688;
	wire [4-1:0] node4689;
	wire [4-1:0] node4691;
	wire [4-1:0] node4693;
	wire [4-1:0] node4696;
	wire [4-1:0] node4697;
	wire [4-1:0] node4700;
	wire [4-1:0] node4701;
	wire [4-1:0] node4705;
	wire [4-1:0] node4706;
	wire [4-1:0] node4707;
	wire [4-1:0] node4708;
	wire [4-1:0] node4709;
	wire [4-1:0] node4711;
	wire [4-1:0] node4714;
	wire [4-1:0] node4715;
	wire [4-1:0] node4719;
	wire [4-1:0] node4722;
	wire [4-1:0] node4723;
	wire [4-1:0] node4724;
	wire [4-1:0] node4726;
	wire [4-1:0] node4729;
	wire [4-1:0] node4730;
	wire [4-1:0] node4734;
	wire [4-1:0] node4736;
	wire [4-1:0] node4739;
	wire [4-1:0] node4740;
	wire [4-1:0] node4742;
	wire [4-1:0] node4743;
	wire [4-1:0] node4745;
	wire [4-1:0] node4749;
	wire [4-1:0] node4750;
	wire [4-1:0] node4751;
	wire [4-1:0] node4755;
	wire [4-1:0] node4756;
	wire [4-1:0] node4759;
	wire [4-1:0] node4762;
	wire [4-1:0] node4763;
	wire [4-1:0] node4764;
	wire [4-1:0] node4765;
	wire [4-1:0] node4766;
	wire [4-1:0] node4767;
	wire [4-1:0] node4769;
	wire [4-1:0] node4772;
	wire [4-1:0] node4773;
	wire [4-1:0] node4775;
	wire [4-1:0] node4778;
	wire [4-1:0] node4780;
	wire [4-1:0] node4783;
	wire [4-1:0] node4784;
	wire [4-1:0] node4785;
	wire [4-1:0] node4786;
	wire [4-1:0] node4790;
	wire [4-1:0] node4794;
	wire [4-1:0] node4795;
	wire [4-1:0] node4796;
	wire [4-1:0] node4797;
	wire [4-1:0] node4800;
	wire [4-1:0] node4803;
	wire [4-1:0] node4804;
	wire [4-1:0] node4805;
	wire [4-1:0] node4808;
	wire [4-1:0] node4812;
	wire [4-1:0] node4813;
	wire [4-1:0] node4816;
	wire [4-1:0] node4817;
	wire [4-1:0] node4818;
	wire [4-1:0] node4823;
	wire [4-1:0] node4824;
	wire [4-1:0] node4825;
	wire [4-1:0] node4826;
	wire [4-1:0] node4827;
	wire [4-1:0] node4828;
	wire [4-1:0] node4831;
	wire [4-1:0] node4834;
	wire [4-1:0] node4837;
	wire [4-1:0] node4838;
	wire [4-1:0] node4842;
	wire [4-1:0] node4843;
	wire [4-1:0] node4845;
	wire [4-1:0] node4846;
	wire [4-1:0] node4850;
	wire [4-1:0] node4851;
	wire [4-1:0] node4853;
	wire [4-1:0] node4856;
	wire [4-1:0] node4858;
	wire [4-1:0] node4861;
	wire [4-1:0] node4862;
	wire [4-1:0] node4863;
	wire [4-1:0] node4866;
	wire [4-1:0] node4867;
	wire [4-1:0] node4869;
	wire [4-1:0] node4872;
	wire [4-1:0] node4873;
	wire [4-1:0] node4877;
	wire [4-1:0] node4878;
	wire [4-1:0] node4880;
	wire [4-1:0] node4883;
	wire [4-1:0] node4884;
	wire [4-1:0] node4887;
	wire [4-1:0] node4890;
	wire [4-1:0] node4891;
	wire [4-1:0] node4892;
	wire [4-1:0] node4893;
	wire [4-1:0] node4894;
	wire [4-1:0] node4895;
	wire [4-1:0] node4896;
	wire [4-1:0] node4900;
	wire [4-1:0] node4901;
	wire [4-1:0] node4904;
	wire [4-1:0] node4908;
	wire [4-1:0] node4909;
	wire [4-1:0] node4910;
	wire [4-1:0] node4913;
	wire [4-1:0] node4914;
	wire [4-1:0] node4918;
	wire [4-1:0] node4919;
	wire [4-1:0] node4923;
	wire [4-1:0] node4924;
	wire [4-1:0] node4925;
	wire [4-1:0] node4927;
	wire [4-1:0] node4931;
	wire [4-1:0] node4932;
	wire [4-1:0] node4933;
	wire [4-1:0] node4934;
	wire [4-1:0] node4937;
	wire [4-1:0] node4940;
	wire [4-1:0] node4941;
	wire [4-1:0] node4944;
	wire [4-1:0] node4947;
	wire [4-1:0] node4948;
	wire [4-1:0] node4950;
	wire [4-1:0] node4953;
	wire [4-1:0] node4954;
	wire [4-1:0] node4958;
	wire [4-1:0] node4959;
	wire [4-1:0] node4960;
	wire [4-1:0] node4961;
	wire [4-1:0] node4962;
	wire [4-1:0] node4966;
	wire [4-1:0] node4969;
	wire [4-1:0] node4970;
	wire [4-1:0] node4972;
	wire [4-1:0] node4975;
	wire [4-1:0] node4978;
	wire [4-1:0] node4979;
	wire [4-1:0] node4980;
	wire [4-1:0] node4982;
	wire [4-1:0] node4985;
	wire [4-1:0] node4986;
	wire [4-1:0] node4989;
	wire [4-1:0] node4992;
	wire [4-1:0] node4993;
	wire [4-1:0] node4994;
	wire [4-1:0] node4996;
	wire [4-1:0] node5000;
	wire [4-1:0] node5003;
	wire [4-1:0] node5004;
	wire [4-1:0] node5005;
	wire [4-1:0] node5006;
	wire [4-1:0] node5007;
	wire [4-1:0] node5008;
	wire [4-1:0] node5009;
	wire [4-1:0] node5012;
	wire [4-1:0] node5014;
	wire [4-1:0] node5017;
	wire [4-1:0] node5018;
	wire [4-1:0] node5021;
	wire [4-1:0] node5023;
	wire [4-1:0] node5026;
	wire [4-1:0] node5027;
	wire [4-1:0] node5028;
	wire [4-1:0] node5029;
	wire [4-1:0] node5033;
	wire [4-1:0] node5034;
	wire [4-1:0] node5038;
	wire [4-1:0] node5039;
	wire [4-1:0] node5040;
	wire [4-1:0] node5044;
	wire [4-1:0] node5045;
	wire [4-1:0] node5046;
	wire [4-1:0] node5049;
	wire [4-1:0] node5052;
	wire [4-1:0] node5055;
	wire [4-1:0] node5056;
	wire [4-1:0] node5057;
	wire [4-1:0] node5058;
	wire [4-1:0] node5059;
	wire [4-1:0] node5062;
	wire [4-1:0] node5063;
	wire [4-1:0] node5066;
	wire [4-1:0] node5069;
	wire [4-1:0] node5070;
	wire [4-1:0] node5071;
	wire [4-1:0] node5076;
	wire [4-1:0] node5078;
	wire [4-1:0] node5081;
	wire [4-1:0] node5082;
	wire [4-1:0] node5083;
	wire [4-1:0] node5084;
	wire [4-1:0] node5088;
	wire [4-1:0] node5090;
	wire [4-1:0] node5093;
	wire [4-1:0] node5094;
	wire [4-1:0] node5096;
	wire [4-1:0] node5099;
	wire [4-1:0] node5100;
	wire [4-1:0] node5104;
	wire [4-1:0] node5105;
	wire [4-1:0] node5106;
	wire [4-1:0] node5107;
	wire [4-1:0] node5108;
	wire [4-1:0] node5109;
	wire [4-1:0] node5114;
	wire [4-1:0] node5115;
	wire [4-1:0] node5116;
	wire [4-1:0] node5119;
	wire [4-1:0] node5120;
	wire [4-1:0] node5124;
	wire [4-1:0] node5126;
	wire [4-1:0] node5127;
	wire [4-1:0] node5130;
	wire [4-1:0] node5133;
	wire [4-1:0] node5134;
	wire [4-1:0] node5136;
	wire [4-1:0] node5137;
	wire [4-1:0] node5140;
	wire [4-1:0] node5141;
	wire [4-1:0] node5145;
	wire [4-1:0] node5146;
	wire [4-1:0] node5147;
	wire [4-1:0] node5151;
	wire [4-1:0] node5152;
	wire [4-1:0] node5156;
	wire [4-1:0] node5157;
	wire [4-1:0] node5158;
	wire [4-1:0] node5159;
	wire [4-1:0] node5160;
	wire [4-1:0] node5162;
	wire [4-1:0] node5165;
	wire [4-1:0] node5166;
	wire [4-1:0] node5169;
	wire [4-1:0] node5172;
	wire [4-1:0] node5173;
	wire [4-1:0] node5176;
	wire [4-1:0] node5177;
	wire [4-1:0] node5181;
	wire [4-1:0] node5182;
	wire [4-1:0] node5183;
	wire [4-1:0] node5184;
	wire [4-1:0] node5187;
	wire [4-1:0] node5190;
	wire [4-1:0] node5193;
	wire [4-1:0] node5194;
	wire [4-1:0] node5195;
	wire [4-1:0] node5198;
	wire [4-1:0] node5202;
	wire [4-1:0] node5203;
	wire [4-1:0] node5204;
	wire [4-1:0] node5206;
	wire [4-1:0] node5209;
	wire [4-1:0] node5211;
	wire [4-1:0] node5213;
	wire [4-1:0] node5216;
	wire [4-1:0] node5218;
	wire [4-1:0] node5220;
	wire [4-1:0] node5223;
	wire [4-1:0] node5224;
	wire [4-1:0] node5225;
	wire [4-1:0] node5226;
	wire [4-1:0] node5227;
	wire [4-1:0] node5228;
	wire [4-1:0] node5229;
	wire [4-1:0] node5233;
	wire [4-1:0] node5234;
	wire [4-1:0] node5235;
	wire [4-1:0] node5240;
	wire [4-1:0] node5241;
	wire [4-1:0] node5243;
	wire [4-1:0] node5246;
	wire [4-1:0] node5247;
	wire [4-1:0] node5250;
	wire [4-1:0] node5252;
	wire [4-1:0] node5255;
	wire [4-1:0] node5256;
	wire [4-1:0] node5257;
	wire [4-1:0] node5259;
	wire [4-1:0] node5261;
	wire [4-1:0] node5264;
	wire [4-1:0] node5265;
	wire [4-1:0] node5266;
	wire [4-1:0] node5269;
	wire [4-1:0] node5272;
	wire [4-1:0] node5273;
	wire [4-1:0] node5277;
	wire [4-1:0] node5279;
	wire [4-1:0] node5280;
	wire [4-1:0] node5283;
	wire [4-1:0] node5284;
	wire [4-1:0] node5287;
	wire [4-1:0] node5290;
	wire [4-1:0] node5291;
	wire [4-1:0] node5292;
	wire [4-1:0] node5293;
	wire [4-1:0] node5294;
	wire [4-1:0] node5297;
	wire [4-1:0] node5298;
	wire [4-1:0] node5301;
	wire [4-1:0] node5304;
	wire [4-1:0] node5306;
	wire [4-1:0] node5309;
	wire [4-1:0] node5310;
	wire [4-1:0] node5311;
	wire [4-1:0] node5313;
	wire [4-1:0] node5316;
	wire [4-1:0] node5317;
	wire [4-1:0] node5320;
	wire [4-1:0] node5323;
	wire [4-1:0] node5324;
	wire [4-1:0] node5325;
	wire [4-1:0] node5330;
	wire [4-1:0] node5331;
	wire [4-1:0] node5332;
	wire [4-1:0] node5335;
	wire [4-1:0] node5336;
	wire [4-1:0] node5339;
	wire [4-1:0] node5342;
	wire [4-1:0] node5343;
	wire [4-1:0] node5344;
	wire [4-1:0] node5348;
	wire [4-1:0] node5349;
	wire [4-1:0] node5352;
	wire [4-1:0] node5355;
	wire [4-1:0] node5356;
	wire [4-1:0] node5357;
	wire [4-1:0] node5358;
	wire [4-1:0] node5359;
	wire [4-1:0] node5361;
	wire [4-1:0] node5362;
	wire [4-1:0] node5367;
	wire [4-1:0] node5369;
	wire [4-1:0] node5370;
	wire [4-1:0] node5372;
	wire [4-1:0] node5376;
	wire [4-1:0] node5377;
	wire [4-1:0] node5378;
	wire [4-1:0] node5380;
	wire [4-1:0] node5384;
	wire [4-1:0] node5385;
	wire [4-1:0] node5386;
	wire [4-1:0] node5388;
	wire [4-1:0] node5391;
	wire [4-1:0] node5394;
	wire [4-1:0] node5395;
	wire [4-1:0] node5397;
	wire [4-1:0] node5400;
	wire [4-1:0] node5401;
	wire [4-1:0] node5405;
	wire [4-1:0] node5406;
	wire [4-1:0] node5407;
	wire [4-1:0] node5408;
	wire [4-1:0] node5409;
	wire [4-1:0] node5411;
	wire [4-1:0] node5414;
	wire [4-1:0] node5415;
	wire [4-1:0] node5420;
	wire [4-1:0] node5421;
	wire [4-1:0] node5422;
	wire [4-1:0] node5423;
	wire [4-1:0] node5426;
	wire [4-1:0] node5430;
	wire [4-1:0] node5432;
	wire [4-1:0] node5435;
	wire [4-1:0] node5436;
	wire [4-1:0] node5437;
	wire [4-1:0] node5439;
	wire [4-1:0] node5442;
	wire [4-1:0] node5443;
	wire [4-1:0] node5447;
	wire [4-1:0] node5448;
	wire [4-1:0] node5451;
	wire [4-1:0] node5453;
	wire [4-1:0] node5455;
	wire [4-1:0] node5458;
	wire [4-1:0] node5459;
	wire [4-1:0] node5460;
	wire [4-1:0] node5461;
	wire [4-1:0] node5462;
	wire [4-1:0] node5463;
	wire [4-1:0] node5464;
	wire [4-1:0] node5465;
	wire [4-1:0] node5466;
	wire [4-1:0] node5468;
	wire [4-1:0] node5471;
	wire [4-1:0] node5472;
	wire [4-1:0] node5475;
	wire [4-1:0] node5478;
	wire [4-1:0] node5479;
	wire [4-1:0] node5480;
	wire [4-1:0] node5482;
	wire [4-1:0] node5486;
	wire [4-1:0] node5487;
	wire [4-1:0] node5488;
	wire [4-1:0] node5493;
	wire [4-1:0] node5494;
	wire [4-1:0] node5495;
	wire [4-1:0] node5497;
	wire [4-1:0] node5500;
	wire [4-1:0] node5501;
	wire [4-1:0] node5504;
	wire [4-1:0] node5505;
	wire [4-1:0] node5508;
	wire [4-1:0] node5511;
	wire [4-1:0] node5512;
	wire [4-1:0] node5514;
	wire [4-1:0] node5516;
	wire [4-1:0] node5519;
	wire [4-1:0] node5520;
	wire [4-1:0] node5524;
	wire [4-1:0] node5525;
	wire [4-1:0] node5526;
	wire [4-1:0] node5527;
	wire [4-1:0] node5529;
	wire [4-1:0] node5530;
	wire [4-1:0] node5534;
	wire [4-1:0] node5536;
	wire [4-1:0] node5539;
	wire [4-1:0] node5540;
	wire [4-1:0] node5541;
	wire [4-1:0] node5545;
	wire [4-1:0] node5548;
	wire [4-1:0] node5549;
	wire [4-1:0] node5551;
	wire [4-1:0] node5552;
	wire [4-1:0] node5553;
	wire [4-1:0] node5557;
	wire [4-1:0] node5559;
	wire [4-1:0] node5562;
	wire [4-1:0] node5563;
	wire [4-1:0] node5564;
	wire [4-1:0] node5566;
	wire [4-1:0] node5570;
	wire [4-1:0] node5571;
	wire [4-1:0] node5575;
	wire [4-1:0] node5576;
	wire [4-1:0] node5577;
	wire [4-1:0] node5578;
	wire [4-1:0] node5579;
	wire [4-1:0] node5580;
	wire [4-1:0] node5581;
	wire [4-1:0] node5586;
	wire [4-1:0] node5588;
	wire [4-1:0] node5591;
	wire [4-1:0] node5592;
	wire [4-1:0] node5595;
	wire [4-1:0] node5596;
	wire [4-1:0] node5598;
	wire [4-1:0] node5601;
	wire [4-1:0] node5604;
	wire [4-1:0] node5605;
	wire [4-1:0] node5606;
	wire [4-1:0] node5607;
	wire [4-1:0] node5611;
	wire [4-1:0] node5614;
	wire [4-1:0] node5615;
	wire [4-1:0] node5616;
	wire [4-1:0] node5617;
	wire [4-1:0] node5623;
	wire [4-1:0] node5624;
	wire [4-1:0] node5625;
	wire [4-1:0] node5626;
	wire [4-1:0] node5630;
	wire [4-1:0] node5631;
	wire [4-1:0] node5633;
	wire [4-1:0] node5636;
	wire [4-1:0] node5638;
	wire [4-1:0] node5639;
	wire [4-1:0] node5643;
	wire [4-1:0] node5644;
	wire [4-1:0] node5645;
	wire [4-1:0] node5647;
	wire [4-1:0] node5651;
	wire [4-1:0] node5652;
	wire [4-1:0] node5655;
	wire [4-1:0] node5658;
	wire [4-1:0] node5659;
	wire [4-1:0] node5660;
	wire [4-1:0] node5661;
	wire [4-1:0] node5662;
	wire [4-1:0] node5663;
	wire [4-1:0] node5665;
	wire [4-1:0] node5667;
	wire [4-1:0] node5670;
	wire [4-1:0] node5671;
	wire [4-1:0] node5672;
	wire [4-1:0] node5677;
	wire [4-1:0] node5678;
	wire [4-1:0] node5679;
	wire [4-1:0] node5681;
	wire [4-1:0] node5684;
	wire [4-1:0] node5685;
	wire [4-1:0] node5690;
	wire [4-1:0] node5691;
	wire [4-1:0] node5692;
	wire [4-1:0] node5693;
	wire [4-1:0] node5694;
	wire [4-1:0] node5697;
	wire [4-1:0] node5701;
	wire [4-1:0] node5703;
	wire [4-1:0] node5704;
	wire [4-1:0] node5708;
	wire [4-1:0] node5709;
	wire [4-1:0] node5710;
	wire [4-1:0] node5714;
	wire [4-1:0] node5717;
	wire [4-1:0] node5718;
	wire [4-1:0] node5719;
	wire [4-1:0] node5720;
	wire [4-1:0] node5721;
	wire [4-1:0] node5722;
	wire [4-1:0] node5727;
	wire [4-1:0] node5729;
	wire [4-1:0] node5732;
	wire [4-1:0] node5733;
	wire [4-1:0] node5735;
	wire [4-1:0] node5739;
	wire [4-1:0] node5740;
	wire [4-1:0] node5741;
	wire [4-1:0] node5744;
	wire [4-1:0] node5746;
	wire [4-1:0] node5747;
	wire [4-1:0] node5750;
	wire [4-1:0] node5753;
	wire [4-1:0] node5754;
	wire [4-1:0] node5756;
	wire [4-1:0] node5759;
	wire [4-1:0] node5760;
	wire [4-1:0] node5761;
	wire [4-1:0] node5764;
	wire [4-1:0] node5767;
	wire [4-1:0] node5768;
	wire [4-1:0] node5772;
	wire [4-1:0] node5773;
	wire [4-1:0] node5774;
	wire [4-1:0] node5775;
	wire [4-1:0] node5776;
	wire [4-1:0] node5778;
	wire [4-1:0] node5781;
	wire [4-1:0] node5782;
	wire [4-1:0] node5783;
	wire [4-1:0] node5788;
	wire [4-1:0] node5789;
	wire [4-1:0] node5790;
	wire [4-1:0] node5791;
	wire [4-1:0] node5794;
	wire [4-1:0] node5798;
	wire [4-1:0] node5799;
	wire [4-1:0] node5801;
	wire [4-1:0] node5804;
	wire [4-1:0] node5806;
	wire [4-1:0] node5809;
	wire [4-1:0] node5810;
	wire [4-1:0] node5811;
	wire [4-1:0] node5812;
	wire [4-1:0] node5814;
	wire [4-1:0] node5818;
	wire [4-1:0] node5820;
	wire [4-1:0] node5822;
	wire [4-1:0] node5825;
	wire [4-1:0] node5826;
	wire [4-1:0] node5827;
	wire [4-1:0] node5831;
	wire [4-1:0] node5832;
	wire [4-1:0] node5833;
	wire [4-1:0] node5837;
	wire [4-1:0] node5840;
	wire [4-1:0] node5841;
	wire [4-1:0] node5842;
	wire [4-1:0] node5843;
	wire [4-1:0] node5845;
	wire [4-1:0] node5848;
	wire [4-1:0] node5849;
	wire [4-1:0] node5851;
	wire [4-1:0] node5854;
	wire [4-1:0] node5857;
	wire [4-1:0] node5858;
	wire [4-1:0] node5859;
	wire [4-1:0] node5863;
	wire [4-1:0] node5866;
	wire [4-1:0] node5867;
	wire [4-1:0] node5868;
	wire [4-1:0] node5869;
	wire [4-1:0] node5871;
	wire [4-1:0] node5874;
	wire [4-1:0] node5878;
	wire [4-1:0] node5879;
	wire [4-1:0] node5880;
	wire [4-1:0] node5884;
	wire [4-1:0] node5885;
	wire [4-1:0] node5886;
	wire [4-1:0] node5890;
	wire [4-1:0] node5891;
	wire [4-1:0] node5895;
	wire [4-1:0] node5896;
	wire [4-1:0] node5897;
	wire [4-1:0] node5898;
	wire [4-1:0] node5899;
	wire [4-1:0] node5900;
	wire [4-1:0] node5901;
	wire [4-1:0] node5902;
	wire [4-1:0] node5906;
	wire [4-1:0] node5907;
	wire [4-1:0] node5908;
	wire [4-1:0] node5913;
	wire [4-1:0] node5914;
	wire [4-1:0] node5915;
	wire [4-1:0] node5919;
	wire [4-1:0] node5921;
	wire [4-1:0] node5924;
	wire [4-1:0] node5925;
	wire [4-1:0] node5926;
	wire [4-1:0] node5927;
	wire [4-1:0] node5930;
	wire [4-1:0] node5931;
	wire [4-1:0] node5935;
	wire [4-1:0] node5938;
	wire [4-1:0] node5939;
	wire [4-1:0] node5942;
	wire [4-1:0] node5944;
	wire [4-1:0] node5946;
	wire [4-1:0] node5949;
	wire [4-1:0] node5950;
	wire [4-1:0] node5951;
	wire [4-1:0] node5952;
	wire [4-1:0] node5953;
	wire [4-1:0] node5954;
	wire [4-1:0] node5957;
	wire [4-1:0] node5960;
	wire [4-1:0] node5963;
	wire [4-1:0] node5964;
	wire [4-1:0] node5965;
	wire [4-1:0] node5969;
	wire [4-1:0] node5972;
	wire [4-1:0] node5973;
	wire [4-1:0] node5974;
	wire [4-1:0] node5976;
	wire [4-1:0] node5979;
	wire [4-1:0] node5982;
	wire [4-1:0] node5984;
	wire [4-1:0] node5987;
	wire [4-1:0] node5988;
	wire [4-1:0] node5989;
	wire [4-1:0] node5990;
	wire [4-1:0] node5991;
	wire [4-1:0] node5997;
	wire [4-1:0] node5998;
	wire [4-1:0] node5999;
	wire [4-1:0] node6003;
	wire [4-1:0] node6004;
	wire [4-1:0] node6005;
	wire [4-1:0] node6009;
	wire [4-1:0] node6011;
	wire [4-1:0] node6014;
	wire [4-1:0] node6015;
	wire [4-1:0] node6016;
	wire [4-1:0] node6017;
	wire [4-1:0] node6018;
	wire [4-1:0] node6019;
	wire [4-1:0] node6022;
	wire [4-1:0] node6025;
	wire [4-1:0] node6026;
	wire [4-1:0] node6028;
	wire [4-1:0] node6032;
	wire [4-1:0] node6033;
	wire [4-1:0] node6035;
	wire [4-1:0] node6038;
	wire [4-1:0] node6039;
	wire [4-1:0] node6040;
	wire [4-1:0] node6043;
	wire [4-1:0] node6046;
	wire [4-1:0] node6049;
	wire [4-1:0] node6050;
	wire [4-1:0] node6051;
	wire [4-1:0] node6052;
	wire [4-1:0] node6057;
	wire [4-1:0] node6058;
	wire [4-1:0] node6061;
	wire [4-1:0] node6062;
	wire [4-1:0] node6064;
	wire [4-1:0] node6068;
	wire [4-1:0] node6069;
	wire [4-1:0] node6070;
	wire [4-1:0] node6071;
	wire [4-1:0] node6072;
	wire [4-1:0] node6076;
	wire [4-1:0] node6077;
	wire [4-1:0] node6078;
	wire [4-1:0] node6082;
	wire [4-1:0] node6083;
	wire [4-1:0] node6086;
	wire [4-1:0] node6089;
	wire [4-1:0] node6090;
	wire [4-1:0] node6091;
	wire [4-1:0] node6096;
	wire [4-1:0] node6097;
	wire [4-1:0] node6098;
	wire [4-1:0] node6099;
	wire [4-1:0] node6103;
	wire [4-1:0] node6105;
	wire [4-1:0] node6106;
	wire [4-1:0] node6110;
	wire [4-1:0] node6111;
	wire [4-1:0] node6112;
	wire [4-1:0] node6113;
	wire [4-1:0] node6116;
	wire [4-1:0] node6119;
	wire [4-1:0] node6121;
	wire [4-1:0] node6125;
	wire [4-1:0] node6126;
	wire [4-1:0] node6127;
	wire [4-1:0] node6128;
	wire [4-1:0] node6129;
	wire [4-1:0] node6130;
	wire [4-1:0] node6133;
	wire [4-1:0] node6135;
	wire [4-1:0] node6136;
	wire [4-1:0] node6140;
	wire [4-1:0] node6141;
	wire [4-1:0] node6142;
	wire [4-1:0] node6144;
	wire [4-1:0] node6147;
	wire [4-1:0] node6148;
	wire [4-1:0] node6152;
	wire [4-1:0] node6153;
	wire [4-1:0] node6154;
	wire [4-1:0] node6157;
	wire [4-1:0] node6160;
	wire [4-1:0] node6163;
	wire [4-1:0] node6164;
	wire [4-1:0] node6165;
	wire [4-1:0] node6168;
	wire [4-1:0] node6169;
	wire [4-1:0] node6171;
	wire [4-1:0] node6174;
	wire [4-1:0] node6175;
	wire [4-1:0] node6179;
	wire [4-1:0] node6180;
	wire [4-1:0] node6181;
	wire [4-1:0] node6185;
	wire [4-1:0] node6186;
	wire [4-1:0] node6188;
	wire [4-1:0] node6191;
	wire [4-1:0] node6193;
	wire [4-1:0] node6196;
	wire [4-1:0] node6197;
	wire [4-1:0] node6198;
	wire [4-1:0] node6199;
	wire [4-1:0] node6200;
	wire [4-1:0] node6203;
	wire [4-1:0] node6204;
	wire [4-1:0] node6208;
	wire [4-1:0] node6209;
	wire [4-1:0] node6212;
	wire [4-1:0] node6214;
	wire [4-1:0] node6217;
	wire [4-1:0] node6218;
	wire [4-1:0] node6220;
	wire [4-1:0] node6221;
	wire [4-1:0] node6224;
	wire [4-1:0] node6227;
	wire [4-1:0] node6229;
	wire [4-1:0] node6232;
	wire [4-1:0] node6233;
	wire [4-1:0] node6234;
	wire [4-1:0] node6237;
	wire [4-1:0] node6238;
	wire [4-1:0] node6239;
	wire [4-1:0] node6244;
	wire [4-1:0] node6245;
	wire [4-1:0] node6246;
	wire [4-1:0] node6249;
	wire [4-1:0] node6251;
	wire [4-1:0] node6254;
	wire [4-1:0] node6256;
	wire [4-1:0] node6257;
	wire [4-1:0] node6261;
	wire [4-1:0] node6262;
	wire [4-1:0] node6263;
	wire [4-1:0] node6264;
	wire [4-1:0] node6265;
	wire [4-1:0] node6267;
	wire [4-1:0] node6268;
	wire [4-1:0] node6272;
	wire [4-1:0] node6273;
	wire [4-1:0] node6274;
	wire [4-1:0] node6279;
	wire [4-1:0] node6280;
	wire [4-1:0] node6283;
	wire [4-1:0] node6284;
	wire [4-1:0] node6285;
	wire [4-1:0] node6289;
	wire [4-1:0] node6290;
	wire [4-1:0] node6293;
	wire [4-1:0] node6296;
	wire [4-1:0] node6297;
	wire [4-1:0] node6299;
	wire [4-1:0] node6301;
	wire [4-1:0] node6304;
	wire [4-1:0] node6305;
	wire [4-1:0] node6307;
	wire [4-1:0] node6308;
	wire [4-1:0] node6312;
	wire [4-1:0] node6313;
	wire [4-1:0] node6317;
	wire [4-1:0] node6318;
	wire [4-1:0] node6319;
	wire [4-1:0] node6320;
	wire [4-1:0] node6322;
	wire [4-1:0] node6325;
	wire [4-1:0] node6326;
	wire [4-1:0] node6329;
	wire [4-1:0] node6332;
	wire [4-1:0] node6333;
	wire [4-1:0] node6334;
	wire [4-1:0] node6335;
	wire [4-1:0] node6339;
	wire [4-1:0] node6340;
	wire [4-1:0] node6344;
	wire [4-1:0] node6345;
	wire [4-1:0] node6349;
	wire [4-1:0] node6350;
	wire [4-1:0] node6351;
	wire [4-1:0] node6352;
	wire [4-1:0] node6356;
	wire [4-1:0] node6359;
	wire [4-1:0] node6360;
	wire [4-1:0] node6361;
	wire [4-1:0] node6363;
	wire [4-1:0] node6366;
	wire [4-1:0] node6369;
	wire [4-1:0] node6371;
	wire [4-1:0] node6374;
	wire [4-1:0] node6375;
	wire [4-1:0] node6376;
	wire [4-1:0] node6377;
	wire [4-1:0] node6378;
	wire [4-1:0] node6379;
	wire [4-1:0] node6380;
	wire [4-1:0] node6381;
	wire [4-1:0] node6384;
	wire [4-1:0] node6386;
	wire [4-1:0] node6389;
	wire [4-1:0] node6390;
	wire [4-1:0] node6392;
	wire [4-1:0] node6393;
	wire [4-1:0] node6396;
	wire [4-1:0] node6399;
	wire [4-1:0] node6401;
	wire [4-1:0] node6404;
	wire [4-1:0] node6405;
	wire [4-1:0] node6406;
	wire [4-1:0] node6408;
	wire [4-1:0] node6411;
	wire [4-1:0] node6414;
	wire [4-1:0] node6415;
	wire [4-1:0] node6416;
	wire [4-1:0] node6417;
	wire [4-1:0] node6421;
	wire [4-1:0] node6423;
	wire [4-1:0] node6426;
	wire [4-1:0] node6427;
	wire [4-1:0] node6428;
	wire [4-1:0] node6432;
	wire [4-1:0] node6433;
	wire [4-1:0] node6437;
	wire [4-1:0] node6438;
	wire [4-1:0] node6439;
	wire [4-1:0] node6440;
	wire [4-1:0] node6443;
	wire [4-1:0] node6444;
	wire [4-1:0] node6447;
	wire [4-1:0] node6450;
	wire [4-1:0] node6451;
	wire [4-1:0] node6452;
	wire [4-1:0] node6455;
	wire [4-1:0] node6456;
	wire [4-1:0] node6461;
	wire [4-1:0] node6462;
	wire [4-1:0] node6463;
	wire [4-1:0] node6465;
	wire [4-1:0] node6467;
	wire [4-1:0] node6470;
	wire [4-1:0] node6471;
	wire [4-1:0] node6474;
	wire [4-1:0] node6475;
	wire [4-1:0] node6478;
	wire [4-1:0] node6481;
	wire [4-1:0] node6482;
	wire [4-1:0] node6483;
	wire [4-1:0] node6487;
	wire [4-1:0] node6490;
	wire [4-1:0] node6491;
	wire [4-1:0] node6492;
	wire [4-1:0] node6493;
	wire [4-1:0] node6494;
	wire [4-1:0] node6496;
	wire [4-1:0] node6499;
	wire [4-1:0] node6500;
	wire [4-1:0] node6504;
	wire [4-1:0] node6505;
	wire [4-1:0] node6507;
	wire [4-1:0] node6510;
	wire [4-1:0] node6511;
	wire [4-1:0] node6512;
	wire [4-1:0] node6516;
	wire [4-1:0] node6517;
	wire [4-1:0] node6521;
	wire [4-1:0] node6522;
	wire [4-1:0] node6523;
	wire [4-1:0] node6524;
	wire [4-1:0] node6526;
	wire [4-1:0] node6530;
	wire [4-1:0] node6532;
	wire [4-1:0] node6533;
	wire [4-1:0] node6537;
	wire [4-1:0] node6538;
	wire [4-1:0] node6539;
	wire [4-1:0] node6542;
	wire [4-1:0] node6545;
	wire [4-1:0] node6546;
	wire [4-1:0] node6550;
	wire [4-1:0] node6551;
	wire [4-1:0] node6552;
	wire [4-1:0] node6553;
	wire [4-1:0] node6556;
	wire [4-1:0] node6559;
	wire [4-1:0] node6560;
	wire [4-1:0] node6562;
	wire [4-1:0] node6563;
	wire [4-1:0] node6568;
	wire [4-1:0] node6569;
	wire [4-1:0] node6570;
	wire [4-1:0] node6573;
	wire [4-1:0] node6576;
	wire [4-1:0] node6577;
	wire [4-1:0] node6578;
	wire [4-1:0] node6582;
	wire [4-1:0] node6584;
	wire [4-1:0] node6587;
	wire [4-1:0] node6588;
	wire [4-1:0] node6589;
	wire [4-1:0] node6590;
	wire [4-1:0] node6591;
	wire [4-1:0] node6592;
	wire [4-1:0] node6594;
	wire [4-1:0] node6595;
	wire [4-1:0] node6599;
	wire [4-1:0] node6600;
	wire [4-1:0] node6603;
	wire [4-1:0] node6605;
	wire [4-1:0] node6608;
	wire [4-1:0] node6609;
	wire [4-1:0] node6611;
	wire [4-1:0] node6614;
	wire [4-1:0] node6615;
	wire [4-1:0] node6618;
	wire [4-1:0] node6621;
	wire [4-1:0] node6622;
	wire [4-1:0] node6623;
	wire [4-1:0] node6624;
	wire [4-1:0] node6626;
	wire [4-1:0] node6630;
	wire [4-1:0] node6632;
	wire [4-1:0] node6635;
	wire [4-1:0] node6636;
	wire [4-1:0] node6637;
	wire [4-1:0] node6640;
	wire [4-1:0] node6642;
	wire [4-1:0] node6645;
	wire [4-1:0] node6646;
	wire [4-1:0] node6649;
	wire [4-1:0] node6652;
	wire [4-1:0] node6653;
	wire [4-1:0] node6654;
	wire [4-1:0] node6656;
	wire [4-1:0] node6657;
	wire [4-1:0] node6659;
	wire [4-1:0] node6662;
	wire [4-1:0] node6665;
	wire [4-1:0] node6666;
	wire [4-1:0] node6667;
	wire [4-1:0] node6670;
	wire [4-1:0] node6672;
	wire [4-1:0] node6675;
	wire [4-1:0] node6678;
	wire [4-1:0] node6679;
	wire [4-1:0] node6680;
	wire [4-1:0] node6682;
	wire [4-1:0] node6685;
	wire [4-1:0] node6687;
	wire [4-1:0] node6689;
	wire [4-1:0] node6692;
	wire [4-1:0] node6693;
	wire [4-1:0] node6695;
	wire [4-1:0] node6698;
	wire [4-1:0] node6699;
	wire [4-1:0] node6700;
	wire [4-1:0] node6705;
	wire [4-1:0] node6706;
	wire [4-1:0] node6707;
	wire [4-1:0] node6708;
	wire [4-1:0] node6709;
	wire [4-1:0] node6712;
	wire [4-1:0] node6715;
	wire [4-1:0] node6716;
	wire [4-1:0] node6718;
	wire [4-1:0] node6720;
	wire [4-1:0] node6724;
	wire [4-1:0] node6725;
	wire [4-1:0] node6726;
	wire [4-1:0] node6727;
	wire [4-1:0] node6728;
	wire [4-1:0] node6733;
	wire [4-1:0] node6736;
	wire [4-1:0] node6737;
	wire [4-1:0] node6741;
	wire [4-1:0] node6742;
	wire [4-1:0] node6743;
	wire [4-1:0] node6745;
	wire [4-1:0] node6746;
	wire [4-1:0] node6750;
	wire [4-1:0] node6751;
	wire [4-1:0] node6752;
	wire [4-1:0] node6755;
	wire [4-1:0] node6758;
	wire [4-1:0] node6759;
	wire [4-1:0] node6760;
	wire [4-1:0] node6765;
	wire [4-1:0] node6766;
	wire [4-1:0] node6767;
	wire [4-1:0] node6768;
	wire [4-1:0] node6771;
	wire [4-1:0] node6774;
	wire [4-1:0] node6776;
	wire [4-1:0] node6779;
	wire [4-1:0] node6780;
	wire [4-1:0] node6784;
	wire [4-1:0] node6785;
	wire [4-1:0] node6786;
	wire [4-1:0] node6787;
	wire [4-1:0] node6788;
	wire [4-1:0] node6789;
	wire [4-1:0] node6790;
	wire [4-1:0] node6793;
	wire [4-1:0] node6796;
	wire [4-1:0] node6797;
	wire [4-1:0] node6798;
	wire [4-1:0] node6802;
	wire [4-1:0] node6805;
	wire [4-1:0] node6806;
	wire [4-1:0] node6807;
	wire [4-1:0] node6808;
	wire [4-1:0] node6811;
	wire [4-1:0] node6814;
	wire [4-1:0] node6815;
	wire [4-1:0] node6819;
	wire [4-1:0] node6820;
	wire [4-1:0] node6822;
	wire [4-1:0] node6823;
	wire [4-1:0] node6827;
	wire [4-1:0] node6828;
	wire [4-1:0] node6832;
	wire [4-1:0] node6833;
	wire [4-1:0] node6834;
	wire [4-1:0] node6835;
	wire [4-1:0] node6836;
	wire [4-1:0] node6839;
	wire [4-1:0] node6840;
	wire [4-1:0] node6843;
	wire [4-1:0] node6846;
	wire [4-1:0] node6847;
	wire [4-1:0] node6848;
	wire [4-1:0] node6852;
	wire [4-1:0] node6855;
	wire [4-1:0] node6856;
	wire [4-1:0] node6857;
	wire [4-1:0] node6860;
	wire [4-1:0] node6862;
	wire [4-1:0] node6865;
	wire [4-1:0] node6868;
	wire [4-1:0] node6869;
	wire [4-1:0] node6870;
	wire [4-1:0] node6871;
	wire [4-1:0] node6876;
	wire [4-1:0] node6877;
	wire [4-1:0] node6878;
	wire [4-1:0] node6880;
	wire [4-1:0] node6883;
	wire [4-1:0] node6887;
	wire [4-1:0] node6888;
	wire [4-1:0] node6889;
	wire [4-1:0] node6890;
	wire [4-1:0] node6891;
	wire [4-1:0] node6893;
	wire [4-1:0] node6896;
	wire [4-1:0] node6897;
	wire [4-1:0] node6898;
	wire [4-1:0] node6903;
	wire [4-1:0] node6904;
	wire [4-1:0] node6905;
	wire [4-1:0] node6908;
	wire [4-1:0] node6912;
	wire [4-1:0] node6913;
	wire [4-1:0] node6914;
	wire [4-1:0] node6916;
	wire [4-1:0] node6920;
	wire [4-1:0] node6921;
	wire [4-1:0] node6923;
	wire [4-1:0] node6927;
	wire [4-1:0] node6928;
	wire [4-1:0] node6929;
	wire [4-1:0] node6930;
	wire [4-1:0] node6933;
	wire [4-1:0] node6935;
	wire [4-1:0] node6938;
	wire [4-1:0] node6940;
	wire [4-1:0] node6941;
	wire [4-1:0] node6942;
	wire [4-1:0] node6946;
	wire [4-1:0] node6949;
	wire [4-1:0] node6950;
	wire [4-1:0] node6951;
	wire [4-1:0] node6952;
	wire [4-1:0] node6955;
	wire [4-1:0] node6958;
	wire [4-1:0] node6959;
	wire [4-1:0] node6963;
	wire [4-1:0] node6964;
	wire [4-1:0] node6967;
	wire [4-1:0] node6969;
	wire [4-1:0] node6971;
	wire [4-1:0] node6974;
	wire [4-1:0] node6975;
	wire [4-1:0] node6976;
	wire [4-1:0] node6977;
	wire [4-1:0] node6978;
	wire [4-1:0] node6979;
	wire [4-1:0] node6982;
	wire [4-1:0] node6984;
	wire [4-1:0] node6987;
	wire [4-1:0] node6988;
	wire [4-1:0] node6989;
	wire [4-1:0] node6992;
	wire [4-1:0] node6993;
	wire [4-1:0] node6997;
	wire [4-1:0] node6999;
	wire [4-1:0] node7002;
	wire [4-1:0] node7003;
	wire [4-1:0] node7004;
	wire [4-1:0] node7007;
	wire [4-1:0] node7010;
	wire [4-1:0] node7012;
	wire [4-1:0] node7014;
	wire [4-1:0] node7017;
	wire [4-1:0] node7018;
	wire [4-1:0] node7019;
	wire [4-1:0] node7020;
	wire [4-1:0] node7021;
	wire [4-1:0] node7023;
	wire [4-1:0] node7026;
	wire [4-1:0] node7028;
	wire [4-1:0] node7031;
	wire [4-1:0] node7032;
	wire [4-1:0] node7034;
	wire [4-1:0] node7037;
	wire [4-1:0] node7039;
	wire [4-1:0] node7042;
	wire [4-1:0] node7043;
	wire [4-1:0] node7044;
	wire [4-1:0] node7046;
	wire [4-1:0] node7049;
	wire [4-1:0] node7051;
	wire [4-1:0] node7054;
	wire [4-1:0] node7057;
	wire [4-1:0] node7058;
	wire [4-1:0] node7059;
	wire [4-1:0] node7060;
	wire [4-1:0] node7062;
	wire [4-1:0] node7065;
	wire [4-1:0] node7066;
	wire [4-1:0] node7069;
	wire [4-1:0] node7072;
	wire [4-1:0] node7075;
	wire [4-1:0] node7076;
	wire [4-1:0] node7079;
	wire [4-1:0] node7080;
	wire [4-1:0] node7083;
	wire [4-1:0] node7084;
	wire [4-1:0] node7088;
	wire [4-1:0] node7089;
	wire [4-1:0] node7090;
	wire [4-1:0] node7091;
	wire [4-1:0] node7092;
	wire [4-1:0] node7094;
	wire [4-1:0] node7097;
	wire [4-1:0] node7098;
	wire [4-1:0] node7102;
	wire [4-1:0] node7103;
	wire [4-1:0] node7105;
	wire [4-1:0] node7106;
	wire [4-1:0] node7110;
	wire [4-1:0] node7112;
	wire [4-1:0] node7115;
	wire [4-1:0] node7116;
	wire [4-1:0] node7119;
	wire [4-1:0] node7122;
	wire [4-1:0] node7123;
	wire [4-1:0] node7124;
	wire [4-1:0] node7125;
	wire [4-1:0] node7127;
	wire [4-1:0] node7131;
	wire [4-1:0] node7133;
	wire [4-1:0] node7134;
	wire [4-1:0] node7138;
	wire [4-1:0] node7139;
	wire [4-1:0] node7140;
	wire [4-1:0] node7142;
	wire [4-1:0] node7143;
	wire [4-1:0] node7146;
	wire [4-1:0] node7149;
	wire [4-1:0] node7150;
	wire [4-1:0] node7152;
	wire [4-1:0] node7156;
	wire [4-1:0] node7157;
	wire [4-1:0] node7158;
	wire [4-1:0] node7160;
	wire [4-1:0] node7165;
	wire [4-1:0] node7166;
	wire [4-1:0] node7167;
	wire [4-1:0] node7168;
	wire [4-1:0] node7169;
	wire [4-1:0] node7170;
	wire [4-1:0] node7171;
	wire [4-1:0] node7172;
	wire [4-1:0] node7173;
	wire [4-1:0] node7174;
	wire [4-1:0] node7175;
	wire [4-1:0] node7177;
	wire [4-1:0] node7180;
	wire [4-1:0] node7181;
	wire [4-1:0] node7185;
	wire [4-1:0] node7186;
	wire [4-1:0] node7188;
	wire [4-1:0] node7190;
	wire [4-1:0] node7193;
	wire [4-1:0] node7194;
	wire [4-1:0] node7196;
	wire [4-1:0] node7200;
	wire [4-1:0] node7201;
	wire [4-1:0] node7202;
	wire [4-1:0] node7203;
	wire [4-1:0] node7204;
	wire [4-1:0] node7209;
	wire [4-1:0] node7210;
	wire [4-1:0] node7211;
	wire [4-1:0] node7214;
	wire [4-1:0] node7217;
	wire [4-1:0] node7219;
	wire [4-1:0] node7222;
	wire [4-1:0] node7223;
	wire [4-1:0] node7225;
	wire [4-1:0] node7228;
	wire [4-1:0] node7230;
	wire [4-1:0] node7231;
	wire [4-1:0] node7234;
	wire [4-1:0] node7237;
	wire [4-1:0] node7238;
	wire [4-1:0] node7239;
	wire [4-1:0] node7240;
	wire [4-1:0] node7241;
	wire [4-1:0] node7243;
	wire [4-1:0] node7246;
	wire [4-1:0] node7248;
	wire [4-1:0] node7251;
	wire [4-1:0] node7252;
	wire [4-1:0] node7256;
	wire [4-1:0] node7257;
	wire [4-1:0] node7261;
	wire [4-1:0] node7262;
	wire [4-1:0] node7263;
	wire [4-1:0] node7264;
	wire [4-1:0] node7265;
	wire [4-1:0] node7268;
	wire [4-1:0] node7271;
	wire [4-1:0] node7272;
	wire [4-1:0] node7276;
	wire [4-1:0] node7278;
	wire [4-1:0] node7280;
	wire [4-1:0] node7283;
	wire [4-1:0] node7284;
	wire [4-1:0] node7286;
	wire [4-1:0] node7288;
	wire [4-1:0] node7291;
	wire [4-1:0] node7294;
	wire [4-1:0] node7295;
	wire [4-1:0] node7296;
	wire [4-1:0] node7297;
	wire [4-1:0] node7298;
	wire [4-1:0] node7299;
	wire [4-1:0] node7300;
	wire [4-1:0] node7303;
	wire [4-1:0] node7306;
	wire [4-1:0] node7308;
	wire [4-1:0] node7311;
	wire [4-1:0] node7312;
	wire [4-1:0] node7315;
	wire [4-1:0] node7316;
	wire [4-1:0] node7320;
	wire [4-1:0] node7321;
	wire [4-1:0] node7322;
	wire [4-1:0] node7324;
	wire [4-1:0] node7328;
	wire [4-1:0] node7330;
	wire [4-1:0] node7333;
	wire [4-1:0] node7334;
	wire [4-1:0] node7335;
	wire [4-1:0] node7336;
	wire [4-1:0] node7338;
	wire [4-1:0] node7341;
	wire [4-1:0] node7344;
	wire [4-1:0] node7346;
	wire [4-1:0] node7349;
	wire [4-1:0] node7350;
	wire [4-1:0] node7352;
	wire [4-1:0] node7354;
	wire [4-1:0] node7357;
	wire [4-1:0] node7358;
	wire [4-1:0] node7359;
	wire [4-1:0] node7363;
	wire [4-1:0] node7364;
	wire [4-1:0] node7368;
	wire [4-1:0] node7369;
	wire [4-1:0] node7370;
	wire [4-1:0] node7371;
	wire [4-1:0] node7372;
	wire [4-1:0] node7373;
	wire [4-1:0] node7377;
	wire [4-1:0] node7380;
	wire [4-1:0] node7381;
	wire [4-1:0] node7384;
	wire [4-1:0] node7387;
	wire [4-1:0] node7388;
	wire [4-1:0] node7389;
	wire [4-1:0] node7392;
	wire [4-1:0] node7394;
	wire [4-1:0] node7397;
	wire [4-1:0] node7398;
	wire [4-1:0] node7401;
	wire [4-1:0] node7404;
	wire [4-1:0] node7405;
	wire [4-1:0] node7406;
	wire [4-1:0] node7407;
	wire [4-1:0] node7410;
	wire [4-1:0] node7413;
	wire [4-1:0] node7414;
	wire [4-1:0] node7416;
	wire [4-1:0] node7420;
	wire [4-1:0] node7422;
	wire [4-1:0] node7424;
	wire [4-1:0] node7426;
	wire [4-1:0] node7429;
	wire [4-1:0] node7430;
	wire [4-1:0] node7431;
	wire [4-1:0] node7432;
	wire [4-1:0] node7433;
	wire [4-1:0] node7436;
	wire [4-1:0] node7437;
	wire [4-1:0] node7438;
	wire [4-1:0] node7443;
	wire [4-1:0] node7444;
	wire [4-1:0] node7445;
	wire [4-1:0] node7446;
	wire [4-1:0] node7450;
	wire [4-1:0] node7451;
	wire [4-1:0] node7453;
	wire [4-1:0] node7456;
	wire [4-1:0] node7457;
	wire [4-1:0] node7460;
	wire [4-1:0] node7463;
	wire [4-1:0] node7464;
	wire [4-1:0] node7466;
	wire [4-1:0] node7469;
	wire [4-1:0] node7471;
	wire [4-1:0] node7472;
	wire [4-1:0] node7476;
	wire [4-1:0] node7477;
	wire [4-1:0] node7478;
	wire [4-1:0] node7479;
	wire [4-1:0] node7481;
	wire [4-1:0] node7484;
	wire [4-1:0] node7485;
	wire [4-1:0] node7489;
	wire [4-1:0] node7490;
	wire [4-1:0] node7492;
	wire [4-1:0] node7493;
	wire [4-1:0] node7498;
	wire [4-1:0] node7499;
	wire [4-1:0] node7501;
	wire [4-1:0] node7502;
	wire [4-1:0] node7503;
	wire [4-1:0] node7506;
	wire [4-1:0] node7509;
	wire [4-1:0] node7512;
	wire [4-1:0] node7514;
	wire [4-1:0] node7515;
	wire [4-1:0] node7518;
	wire [4-1:0] node7521;
	wire [4-1:0] node7522;
	wire [4-1:0] node7523;
	wire [4-1:0] node7524;
	wire [4-1:0] node7525;
	wire [4-1:0] node7528;
	wire [4-1:0] node7529;
	wire [4-1:0] node7532;
	wire [4-1:0] node7533;
	wire [4-1:0] node7536;
	wire [4-1:0] node7539;
	wire [4-1:0] node7540;
	wire [4-1:0] node7541;
	wire [4-1:0] node7543;
	wire [4-1:0] node7546;
	wire [4-1:0] node7549;
	wire [4-1:0] node7551;
	wire [4-1:0] node7553;
	wire [4-1:0] node7556;
	wire [4-1:0] node7557;
	wire [4-1:0] node7558;
	wire [4-1:0] node7561;
	wire [4-1:0] node7562;
	wire [4-1:0] node7563;
	wire [4-1:0] node7567;
	wire [4-1:0] node7569;
	wire [4-1:0] node7572;
	wire [4-1:0] node7573;
	wire [4-1:0] node7574;
	wire [4-1:0] node7576;
	wire [4-1:0] node7579;
	wire [4-1:0] node7582;
	wire [4-1:0] node7584;
	wire [4-1:0] node7587;
	wire [4-1:0] node7588;
	wire [4-1:0] node7589;
	wire [4-1:0] node7591;
	wire [4-1:0] node7594;
	wire [4-1:0] node7596;
	wire [4-1:0] node7599;
	wire [4-1:0] node7600;
	wire [4-1:0] node7601;
	wire [4-1:0] node7604;
	wire [4-1:0] node7605;
	wire [4-1:0] node7607;
	wire [4-1:0] node7610;
	wire [4-1:0] node7611;
	wire [4-1:0] node7614;
	wire [4-1:0] node7617;
	wire [4-1:0] node7618;
	wire [4-1:0] node7620;
	wire [4-1:0] node7622;
	wire [4-1:0] node7625;
	wire [4-1:0] node7626;
	wire [4-1:0] node7629;
	wire [4-1:0] node7630;
	wire [4-1:0] node7634;
	wire [4-1:0] node7635;
	wire [4-1:0] node7636;
	wire [4-1:0] node7637;
	wire [4-1:0] node7638;
	wire [4-1:0] node7639;
	wire [4-1:0] node7640;
	wire [4-1:0] node7644;
	wire [4-1:0] node7646;
	wire [4-1:0] node7647;
	wire [4-1:0] node7649;
	wire [4-1:0] node7652;
	wire [4-1:0] node7654;
	wire [4-1:0] node7657;
	wire [4-1:0] node7658;
	wire [4-1:0] node7659;
	wire [4-1:0] node7660;
	wire [4-1:0] node7664;
	wire [4-1:0] node7665;
	wire [4-1:0] node7667;
	wire [4-1:0] node7670;
	wire [4-1:0] node7671;
	wire [4-1:0] node7675;
	wire [4-1:0] node7676;
	wire [4-1:0] node7678;
	wire [4-1:0] node7679;
	wire [4-1:0] node7682;
	wire [4-1:0] node7685;
	wire [4-1:0] node7686;
	wire [4-1:0] node7690;
	wire [4-1:0] node7691;
	wire [4-1:0] node7692;
	wire [4-1:0] node7693;
	wire [4-1:0] node7694;
	wire [4-1:0] node7695;
	wire [4-1:0] node7699;
	wire [4-1:0] node7702;
	wire [4-1:0] node7703;
	wire [4-1:0] node7704;
	wire [4-1:0] node7709;
	wire [4-1:0] node7710;
	wire [4-1:0] node7711;
	wire [4-1:0] node7714;
	wire [4-1:0] node7717;
	wire [4-1:0] node7720;
	wire [4-1:0] node7721;
	wire [4-1:0] node7722;
	wire [4-1:0] node7723;
	wire [4-1:0] node7725;
	wire [4-1:0] node7728;
	wire [4-1:0] node7730;
	wire [4-1:0] node7733;
	wire [4-1:0] node7734;
	wire [4-1:0] node7736;
	wire [4-1:0] node7739;
	wire [4-1:0] node7742;
	wire [4-1:0] node7743;
	wire [4-1:0] node7744;
	wire [4-1:0] node7747;
	wire [4-1:0] node7748;
	wire [4-1:0] node7751;
	wire [4-1:0] node7754;
	wire [4-1:0] node7755;
	wire [4-1:0] node7758;
	wire [4-1:0] node7760;
	wire [4-1:0] node7763;
	wire [4-1:0] node7764;
	wire [4-1:0] node7765;
	wire [4-1:0] node7766;
	wire [4-1:0] node7767;
	wire [4-1:0] node7770;
	wire [4-1:0] node7771;
	wire [4-1:0] node7775;
	wire [4-1:0] node7777;
	wire [4-1:0] node7780;
	wire [4-1:0] node7781;
	wire [4-1:0] node7782;
	wire [4-1:0] node7783;
	wire [4-1:0] node7785;
	wire [4-1:0] node7788;
	wire [4-1:0] node7791;
	wire [4-1:0] node7793;
	wire [4-1:0] node7795;
	wire [4-1:0] node7798;
	wire [4-1:0] node7799;
	wire [4-1:0] node7800;
	wire [4-1:0] node7802;
	wire [4-1:0] node7807;
	wire [4-1:0] node7808;
	wire [4-1:0] node7809;
	wire [4-1:0] node7810;
	wire [4-1:0] node7811;
	wire [4-1:0] node7814;
	wire [4-1:0] node7817;
	wire [4-1:0] node7819;
	wire [4-1:0] node7822;
	wire [4-1:0] node7823;
	wire [4-1:0] node7825;
	wire [4-1:0] node7828;
	wire [4-1:0] node7830;
	wire [4-1:0] node7833;
	wire [4-1:0] node7834;
	wire [4-1:0] node7835;
	wire [4-1:0] node7836;
	wire [4-1:0] node7840;
	wire [4-1:0] node7842;
	wire [4-1:0] node7845;
	wire [4-1:0] node7846;
	wire [4-1:0] node7847;
	wire [4-1:0] node7848;
	wire [4-1:0] node7853;
	wire [4-1:0] node7854;
	wire [4-1:0] node7855;
	wire [4-1:0] node7859;
	wire [4-1:0] node7862;
	wire [4-1:0] node7863;
	wire [4-1:0] node7864;
	wire [4-1:0] node7865;
	wire [4-1:0] node7866;
	wire [4-1:0] node7867;
	wire [4-1:0] node7869;
	wire [4-1:0] node7870;
	wire [4-1:0] node7873;
	wire [4-1:0] node7876;
	wire [4-1:0] node7878;
	wire [4-1:0] node7879;
	wire [4-1:0] node7882;
	wire [4-1:0] node7885;
	wire [4-1:0] node7887;
	wire [4-1:0] node7889;
	wire [4-1:0] node7890;
	wire [4-1:0] node7894;
	wire [4-1:0] node7895;
	wire [4-1:0] node7896;
	wire [4-1:0] node7897;
	wire [4-1:0] node7900;
	wire [4-1:0] node7904;
	wire [4-1:0] node7905;
	wire [4-1:0] node7906;
	wire [4-1:0] node7909;
	wire [4-1:0] node7910;
	wire [4-1:0] node7914;
	wire [4-1:0] node7915;
	wire [4-1:0] node7919;
	wire [4-1:0] node7920;
	wire [4-1:0] node7921;
	wire [4-1:0] node7922;
	wire [4-1:0] node7923;
	wire [4-1:0] node7927;
	wire [4-1:0] node7928;
	wire [4-1:0] node7930;
	wire [4-1:0] node7933;
	wire [4-1:0] node7936;
	wire [4-1:0] node7937;
	wire [4-1:0] node7941;
	wire [4-1:0] node7942;
	wire [4-1:0] node7943;
	wire [4-1:0] node7945;
	wire [4-1:0] node7949;
	wire [4-1:0] node7950;
	wire [4-1:0] node7951;
	wire [4-1:0] node7955;
	wire [4-1:0] node7957;
	wire [4-1:0] node7960;
	wire [4-1:0] node7961;
	wire [4-1:0] node7962;
	wire [4-1:0] node7963;
	wire [4-1:0] node7964;
	wire [4-1:0] node7965;
	wire [4-1:0] node7970;
	wire [4-1:0] node7971;
	wire [4-1:0] node7974;
	wire [4-1:0] node7976;
	wire [4-1:0] node7979;
	wire [4-1:0] node7981;
	wire [4-1:0] node7982;
	wire [4-1:0] node7984;
	wire [4-1:0] node7987;
	wire [4-1:0] node7988;
	wire [4-1:0] node7992;
	wire [4-1:0] node7993;
	wire [4-1:0] node7994;
	wire [4-1:0] node7995;
	wire [4-1:0] node7996;
	wire [4-1:0] node7998;
	wire [4-1:0] node8002;
	wire [4-1:0] node8003;
	wire [4-1:0] node8005;
	wire [4-1:0] node8009;
	wire [4-1:0] node8010;
	wire [4-1:0] node8013;
	wire [4-1:0] node8014;
	wire [4-1:0] node8017;
	wire [4-1:0] node8020;
	wire [4-1:0] node8021;
	wire [4-1:0] node8022;
	wire [4-1:0] node8023;
	wire [4-1:0] node8026;
	wire [4-1:0] node8028;
	wire [4-1:0] node8031;
	wire [4-1:0] node8032;
	wire [4-1:0] node8034;
	wire [4-1:0] node8038;
	wire [4-1:0] node8039;
	wire [4-1:0] node8041;
	wire [4-1:0] node8042;
	wire [4-1:0] node8045;
	wire [4-1:0] node8048;
	wire [4-1:0] node8049;
	wire [4-1:0] node8050;
	wire [4-1:0] node8053;
	wire [4-1:0] node8056;
	wire [4-1:0] node8059;
	wire [4-1:0] node8060;
	wire [4-1:0] node8061;
	wire [4-1:0] node8062;
	wire [4-1:0] node8063;
	wire [4-1:0] node8064;
	wire [4-1:0] node8065;
	wire [4-1:0] node8066;
	wire [4-1:0] node8068;
	wire [4-1:0] node8072;
	wire [4-1:0] node8073;
	wire [4-1:0] node8075;
	wire [4-1:0] node8078;
	wire [4-1:0] node8081;
	wire [4-1:0] node8082;
	wire [4-1:0] node8083;
	wire [4-1:0] node8085;
	wire [4-1:0] node8087;
	wire [4-1:0] node8091;
	wire [4-1:0] node8092;
	wire [4-1:0] node8094;
	wire [4-1:0] node8097;
	wire [4-1:0] node8100;
	wire [4-1:0] node8101;
	wire [4-1:0] node8102;
	wire [4-1:0] node8103;
	wire [4-1:0] node8104;
	wire [4-1:0] node8106;
	wire [4-1:0] node8110;
	wire [4-1:0] node8112;
	wire [4-1:0] node8115;
	wire [4-1:0] node8116;
	wire [4-1:0] node8118;
	wire [4-1:0] node8121;
	wire [4-1:0] node8122;
	wire [4-1:0] node8125;
	wire [4-1:0] node8126;
	wire [4-1:0] node8130;
	wire [4-1:0] node8131;
	wire [4-1:0] node8132;
	wire [4-1:0] node8135;
	wire [4-1:0] node8137;
	wire [4-1:0] node8140;
	wire [4-1:0] node8141;
	wire [4-1:0] node8143;
	wire [4-1:0] node8146;
	wire [4-1:0] node8147;
	wire [4-1:0] node8151;
	wire [4-1:0] node8152;
	wire [4-1:0] node8153;
	wire [4-1:0] node8154;
	wire [4-1:0] node8155;
	wire [4-1:0] node8156;
	wire [4-1:0] node8158;
	wire [4-1:0] node8161;
	wire [4-1:0] node8164;
	wire [4-1:0] node8165;
	wire [4-1:0] node8169;
	wire [4-1:0] node8171;
	wire [4-1:0] node8174;
	wire [4-1:0] node8175;
	wire [4-1:0] node8176;
	wire [4-1:0] node8178;
	wire [4-1:0] node8179;
	wire [4-1:0] node8182;
	wire [4-1:0] node8185;
	wire [4-1:0] node8187;
	wire [4-1:0] node8189;
	wire [4-1:0] node8192;
	wire [4-1:0] node8193;
	wire [4-1:0] node8196;
	wire [4-1:0] node8198;
	wire [4-1:0] node8200;
	wire [4-1:0] node8203;
	wire [4-1:0] node8204;
	wire [4-1:0] node8205;
	wire [4-1:0] node8206;
	wire [4-1:0] node8207;
	wire [4-1:0] node8211;
	wire [4-1:0] node8212;
	wire [4-1:0] node8213;
	wire [4-1:0] node8216;
	wire [4-1:0] node8220;
	wire [4-1:0] node8221;
	wire [4-1:0] node8222;
	wire [4-1:0] node8226;
	wire [4-1:0] node8228;
	wire [4-1:0] node8229;
	wire [4-1:0] node8232;
	wire [4-1:0] node8235;
	wire [4-1:0] node8236;
	wire [4-1:0] node8237;
	wire [4-1:0] node8240;
	wire [4-1:0] node8241;
	wire [4-1:0] node8245;
	wire [4-1:0] node8246;
	wire [4-1:0] node8248;
	wire [4-1:0] node8250;
	wire [4-1:0] node8253;
	wire [4-1:0] node8256;
	wire [4-1:0] node8257;
	wire [4-1:0] node8258;
	wire [4-1:0] node8259;
	wire [4-1:0] node8260;
	wire [4-1:0] node8261;
	wire [4-1:0] node8264;
	wire [4-1:0] node8265;
	wire [4-1:0] node8268;
	wire [4-1:0] node8271;
	wire [4-1:0] node8272;
	wire [4-1:0] node8273;
	wire [4-1:0] node8274;
	wire [4-1:0] node8277;
	wire [4-1:0] node8280;
	wire [4-1:0] node8283;
	wire [4-1:0] node8284;
	wire [4-1:0] node8285;
	wire [4-1:0] node8289;
	wire [4-1:0] node8291;
	wire [4-1:0] node8294;
	wire [4-1:0] node8295;
	wire [4-1:0] node8296;
	wire [4-1:0] node8298;
	wire [4-1:0] node8301;
	wire [4-1:0] node8302;
	wire [4-1:0] node8303;
	wire [4-1:0] node8306;
	wire [4-1:0] node8309;
	wire [4-1:0] node8310;
	wire [4-1:0] node8314;
	wire [4-1:0] node8315;
	wire [4-1:0] node8316;
	wire [4-1:0] node8320;
	wire [4-1:0] node8321;
	wire [4-1:0] node8325;
	wire [4-1:0] node8326;
	wire [4-1:0] node8327;
	wire [4-1:0] node8328;
	wire [4-1:0] node8331;
	wire [4-1:0] node8332;
	wire [4-1:0] node8333;
	wire [4-1:0] node8338;
	wire [4-1:0] node8340;
	wire [4-1:0] node8341;
	wire [4-1:0] node8342;
	wire [4-1:0] node8347;
	wire [4-1:0] node8348;
	wire [4-1:0] node8349;
	wire [4-1:0] node8351;
	wire [4-1:0] node8352;
	wire [4-1:0] node8356;
	wire [4-1:0] node8357;
	wire [4-1:0] node8358;
	wire [4-1:0] node8362;
	wire [4-1:0] node8365;
	wire [4-1:0] node8366;
	wire [4-1:0] node8369;
	wire [4-1:0] node8370;
	wire [4-1:0] node8373;
	wire [4-1:0] node8376;
	wire [4-1:0] node8377;
	wire [4-1:0] node8378;
	wire [4-1:0] node8379;
	wire [4-1:0] node8380;
	wire [4-1:0] node8381;
	wire [4-1:0] node8385;
	wire [4-1:0] node8387;
	wire [4-1:0] node8388;
	wire [4-1:0] node8392;
	wire [4-1:0] node8393;
	wire [4-1:0] node8395;
	wire [4-1:0] node8397;
	wire [4-1:0] node8400;
	wire [4-1:0] node8402;
	wire [4-1:0] node8404;
	wire [4-1:0] node8407;
	wire [4-1:0] node8408;
	wire [4-1:0] node8409;
	wire [4-1:0] node8411;
	wire [4-1:0] node8414;
	wire [4-1:0] node8417;
	wire [4-1:0] node8419;
	wire [4-1:0] node8420;
	wire [4-1:0] node8422;
	wire [4-1:0] node8425;
	wire [4-1:0] node8426;
	wire [4-1:0] node8430;
	wire [4-1:0] node8431;
	wire [4-1:0] node8432;
	wire [4-1:0] node8433;
	wire [4-1:0] node8434;
	wire [4-1:0] node8436;
	wire [4-1:0] node8440;
	wire [4-1:0] node8441;
	wire [4-1:0] node8445;
	wire [4-1:0] node8446;
	wire [4-1:0] node8447;
	wire [4-1:0] node8449;
	wire [4-1:0] node8452;
	wire [4-1:0] node8454;
	wire [4-1:0] node8457;
	wire [4-1:0] node8458;
	wire [4-1:0] node8461;
	wire [4-1:0] node8464;
	wire [4-1:0] node8465;
	wire [4-1:0] node8466;
	wire [4-1:0] node8468;
	wire [4-1:0] node8471;
	wire [4-1:0] node8472;
	wire [4-1:0] node8474;
	wire [4-1:0] node8477;
	wire [4-1:0] node8479;
	wire [4-1:0] node8482;
	wire [4-1:0] node8484;
	wire [4-1:0] node8487;
	wire [4-1:0] node8488;
	wire [4-1:0] node8489;
	wire [4-1:0] node8490;
	wire [4-1:0] node8491;
	wire [4-1:0] node8492;
	wire [4-1:0] node8493;
	wire [4-1:0] node8494;
	wire [4-1:0] node8498;
	wire [4-1:0] node8499;
	wire [4-1:0] node8503;
	wire [4-1:0] node8504;
	wire [4-1:0] node8505;
	wire [4-1:0] node8509;
	wire [4-1:0] node8510;
	wire [4-1:0] node8511;
	wire [4-1:0] node8515;
	wire [4-1:0] node8516;
	wire [4-1:0] node8520;
	wire [4-1:0] node8521;
	wire [4-1:0] node8523;
	wire [4-1:0] node8526;
	wire [4-1:0] node8528;
	wire [4-1:0] node8530;
	wire [4-1:0] node8531;
	wire [4-1:0] node8535;
	wire [4-1:0] node8536;
	wire [4-1:0] node8537;
	wire [4-1:0] node8538;
	wire [4-1:0] node8539;
	wire [4-1:0] node8543;
	wire [4-1:0] node8546;
	wire [4-1:0] node8548;
	wire [4-1:0] node8549;
	wire [4-1:0] node8552;
	wire [4-1:0] node8555;
	wire [4-1:0] node8556;
	wire [4-1:0] node8557;
	wire [4-1:0] node8560;
	wire [4-1:0] node8563;
	wire [4-1:0] node8564;
	wire [4-1:0] node8567;
	wire [4-1:0] node8569;
	wire [4-1:0] node8572;
	wire [4-1:0] node8573;
	wire [4-1:0] node8574;
	wire [4-1:0] node8575;
	wire [4-1:0] node8576;
	wire [4-1:0] node8579;
	wire [4-1:0] node8580;
	wire [4-1:0] node8582;
	wire [4-1:0] node8586;
	wire [4-1:0] node8587;
	wire [4-1:0] node8588;
	wire [4-1:0] node8592;
	wire [4-1:0] node8593;
	wire [4-1:0] node8597;
	wire [4-1:0] node8598;
	wire [4-1:0] node8600;
	wire [4-1:0] node8601;
	wire [4-1:0] node8605;
	wire [4-1:0] node8606;
	wire [4-1:0] node8610;
	wire [4-1:0] node8611;
	wire [4-1:0] node8612;
	wire [4-1:0] node8614;
	wire [4-1:0] node8616;
	wire [4-1:0] node8617;
	wire [4-1:0] node8620;
	wire [4-1:0] node8623;
	wire [4-1:0] node8625;
	wire [4-1:0] node8626;
	wire [4-1:0] node8629;
	wire [4-1:0] node8632;
	wire [4-1:0] node8633;
	wire [4-1:0] node8635;
	wire [4-1:0] node8636;
	wire [4-1:0] node8637;
	wire [4-1:0] node8641;
	wire [4-1:0] node8644;
	wire [4-1:0] node8646;
	wire [4-1:0] node8647;
	wire [4-1:0] node8648;
	wire [4-1:0] node8651;
	wire [4-1:0] node8655;
	wire [4-1:0] node8656;
	wire [4-1:0] node8657;
	wire [4-1:0] node8658;
	wire [4-1:0] node8659;
	wire [4-1:0] node8660;
	wire [4-1:0] node8661;
	wire [4-1:0] node8662;
	wire [4-1:0] node8666;
	wire [4-1:0] node8669;
	wire [4-1:0] node8670;
	wire [4-1:0] node8673;
	wire [4-1:0] node8675;
	wire [4-1:0] node8678;
	wire [4-1:0] node8679;
	wire [4-1:0] node8680;
	wire [4-1:0] node8682;
	wire [4-1:0] node8687;
	wire [4-1:0] node8688;
	wire [4-1:0] node8689;
	wire [4-1:0] node8691;
	wire [4-1:0] node8694;
	wire [4-1:0] node8696;
	wire [4-1:0] node8697;
	wire [4-1:0] node8700;
	wire [4-1:0] node8703;
	wire [4-1:0] node8705;
	wire [4-1:0] node8706;
	wire [4-1:0] node8707;
	wire [4-1:0] node8712;
	wire [4-1:0] node8713;
	wire [4-1:0] node8714;
	wire [4-1:0] node8715;
	wire [4-1:0] node8719;
	wire [4-1:0] node8721;
	wire [4-1:0] node8722;
	wire [4-1:0] node8723;
	wire [4-1:0] node8726;
	wire [4-1:0] node8730;
	wire [4-1:0] node8731;
	wire [4-1:0] node8732;
	wire [4-1:0] node8734;
	wire [4-1:0] node8735;
	wire [4-1:0] node8738;
	wire [4-1:0] node8742;
	wire [4-1:0] node8744;
	wire [4-1:0] node8745;
	wire [4-1:0] node8749;
	wire [4-1:0] node8750;
	wire [4-1:0] node8751;
	wire [4-1:0] node8752;
	wire [4-1:0] node8753;
	wire [4-1:0] node8754;
	wire [4-1:0] node8755;
	wire [4-1:0] node8760;
	wire [4-1:0] node8762;
	wire [4-1:0] node8765;
	wire [4-1:0] node8766;
	wire [4-1:0] node8767;
	wire [4-1:0] node8769;
	wire [4-1:0] node8772;
	wire [4-1:0] node8774;
	wire [4-1:0] node8777;
	wire [4-1:0] node8778;
	wire [4-1:0] node8781;
	wire [4-1:0] node8782;
	wire [4-1:0] node8786;
	wire [4-1:0] node8787;
	wire [4-1:0] node8788;
	wire [4-1:0] node8789;
	wire [4-1:0] node8791;
	wire [4-1:0] node8794;
	wire [4-1:0] node8797;
	wire [4-1:0] node8799;
	wire [4-1:0] node8800;
	wire [4-1:0] node8803;
	wire [4-1:0] node8806;
	wire [4-1:0] node8807;
	wire [4-1:0] node8809;
	wire [4-1:0] node8810;
	wire [4-1:0] node8814;
	wire [4-1:0] node8816;
	wire [4-1:0] node8817;
	wire [4-1:0] node8820;
	wire [4-1:0] node8823;
	wire [4-1:0] node8824;
	wire [4-1:0] node8825;
	wire [4-1:0] node8826;
	wire [4-1:0] node8827;
	wire [4-1:0] node8828;
	wire [4-1:0] node8831;
	wire [4-1:0] node8835;
	wire [4-1:0] node8837;
	wire [4-1:0] node8840;
	wire [4-1:0] node8842;
	wire [4-1:0] node8844;
	wire [4-1:0] node8847;
	wire [4-1:0] node8848;
	wire [4-1:0] node8849;
	wire [4-1:0] node8850;
	wire [4-1:0] node8853;
	wire [4-1:0] node8854;
	wire [4-1:0] node8859;
	wire [4-1:0] node8861;
	wire [4-1:0] node8862;
	wire [4-1:0] node8866;
	wire [4-1:0] node8867;
	wire [4-1:0] node8868;
	wire [4-1:0] node8869;
	wire [4-1:0] node8870;
	wire [4-1:0] node8871;
	wire [4-1:0] node8872;
	wire [4-1:0] node8873;
	wire [4-1:0] node8875;
	wire [4-1:0] node8877;
	wire [4-1:0] node8880;
	wire [4-1:0] node8882;
	wire [4-1:0] node8883;
	wire [4-1:0] node8886;
	wire [4-1:0] node8887;
	wire [4-1:0] node8891;
	wire [4-1:0] node8892;
	wire [4-1:0] node8893;
	wire [4-1:0] node8894;
	wire [4-1:0] node8897;
	wire [4-1:0] node8899;
	wire [4-1:0] node8902;
	wire [4-1:0] node8903;
	wire [4-1:0] node8905;
	wire [4-1:0] node8908;
	wire [4-1:0] node8910;
	wire [4-1:0] node8913;
	wire [4-1:0] node8914;
	wire [4-1:0] node8917;
	wire [4-1:0] node8918;
	wire [4-1:0] node8922;
	wire [4-1:0] node8923;
	wire [4-1:0] node8924;
	wire [4-1:0] node8925;
	wire [4-1:0] node8928;
	wire [4-1:0] node8930;
	wire [4-1:0] node8931;
	wire [4-1:0] node8935;
	wire [4-1:0] node8936;
	wire [4-1:0] node8939;
	wire [4-1:0] node8940;
	wire [4-1:0] node8942;
	wire [4-1:0] node8946;
	wire [4-1:0] node8947;
	wire [4-1:0] node8948;
	wire [4-1:0] node8949;
	wire [4-1:0] node8950;
	wire [4-1:0] node8954;
	wire [4-1:0] node8957;
	wire [4-1:0] node8958;
	wire [4-1:0] node8962;
	wire [4-1:0] node8963;
	wire [4-1:0] node8965;
	wire [4-1:0] node8967;
	wire [4-1:0] node8970;
	wire [4-1:0] node8973;
	wire [4-1:0] node8974;
	wire [4-1:0] node8975;
	wire [4-1:0] node8976;
	wire [4-1:0] node8977;
	wire [4-1:0] node8978;
	wire [4-1:0] node8981;
	wire [4-1:0] node8984;
	wire [4-1:0] node8985;
	wire [4-1:0] node8987;
	wire [4-1:0] node8991;
	wire [4-1:0] node8992;
	wire [4-1:0] node8994;
	wire [4-1:0] node8997;
	wire [4-1:0] node8998;
	wire [4-1:0] node9000;
	wire [4-1:0] node9004;
	wire [4-1:0] node9005;
	wire [4-1:0] node9007;
	wire [4-1:0] node9008;
	wire [4-1:0] node9011;
	wire [4-1:0] node9012;
	wire [4-1:0] node9016;
	wire [4-1:0] node9017;
	wire [4-1:0] node9019;
	wire [4-1:0] node9022;
	wire [4-1:0] node9023;
	wire [4-1:0] node9025;
	wire [4-1:0] node9028;
	wire [4-1:0] node9031;
	wire [4-1:0] node9032;
	wire [4-1:0] node9033;
	wire [4-1:0] node9034;
	wire [4-1:0] node9036;
	wire [4-1:0] node9039;
	wire [4-1:0] node9040;
	wire [4-1:0] node9042;
	wire [4-1:0] node9045;
	wire [4-1:0] node9047;
	wire [4-1:0] node9050;
	wire [4-1:0] node9051;
	wire [4-1:0] node9054;
	wire [4-1:0] node9056;
	wire [4-1:0] node9057;
	wire [4-1:0] node9060;
	wire [4-1:0] node9063;
	wire [4-1:0] node9064;
	wire [4-1:0] node9065;
	wire [4-1:0] node9066;
	wire [4-1:0] node9067;
	wire [4-1:0] node9070;
	wire [4-1:0] node9075;
	wire [4-1:0] node9076;
	wire [4-1:0] node9078;
	wire [4-1:0] node9081;
	wire [4-1:0] node9084;
	wire [4-1:0] node9085;
	wire [4-1:0] node9086;
	wire [4-1:0] node9087;
	wire [4-1:0] node9088;
	wire [4-1:0] node9089;
	wire [4-1:0] node9091;
	wire [4-1:0] node9092;
	wire [4-1:0] node9096;
	wire [4-1:0] node9099;
	wire [4-1:0] node9100;
	wire [4-1:0] node9103;
	wire [4-1:0] node9104;
	wire [4-1:0] node9107;
	wire [4-1:0] node9108;
	wire [4-1:0] node9111;
	wire [4-1:0] node9114;
	wire [4-1:0] node9115;
	wire [4-1:0] node9116;
	wire [4-1:0] node9118;
	wire [4-1:0] node9122;
	wire [4-1:0] node9123;
	wire [4-1:0] node9125;
	wire [4-1:0] node9127;
	wire [4-1:0] node9130;
	wire [4-1:0] node9131;
	wire [4-1:0] node9135;
	wire [4-1:0] node9136;
	wire [4-1:0] node9137;
	wire [4-1:0] node9138;
	wire [4-1:0] node9141;
	wire [4-1:0] node9144;
	wire [4-1:0] node9145;
	wire [4-1:0] node9146;
	wire [4-1:0] node9149;
	wire [4-1:0] node9152;
	wire [4-1:0] node9153;
	wire [4-1:0] node9154;
	wire [4-1:0] node9159;
	wire [4-1:0] node9160;
	wire [4-1:0] node9161;
	wire [4-1:0] node9162;
	wire [4-1:0] node9163;
	wire [4-1:0] node9167;
	wire [4-1:0] node9169;
	wire [4-1:0] node9172;
	wire [4-1:0] node9173;
	wire [4-1:0] node9175;
	wire [4-1:0] node9178;
	wire [4-1:0] node9179;
	wire [4-1:0] node9183;
	wire [4-1:0] node9184;
	wire [4-1:0] node9185;
	wire [4-1:0] node9189;
	wire [4-1:0] node9190;
	wire [4-1:0] node9193;
	wire [4-1:0] node9194;
	wire [4-1:0] node9198;
	wire [4-1:0] node9199;
	wire [4-1:0] node9200;
	wire [4-1:0] node9201;
	wire [4-1:0] node9202;
	wire [4-1:0] node9205;
	wire [4-1:0] node9206;
	wire [4-1:0] node9207;
	wire [4-1:0] node9210;
	wire [4-1:0] node9214;
	wire [4-1:0] node9216;
	wire [4-1:0] node9217;
	wire [4-1:0] node9219;
	wire [4-1:0] node9222;
	wire [4-1:0] node9225;
	wire [4-1:0] node9226;
	wire [4-1:0] node9228;
	wire [4-1:0] node9229;
	wire [4-1:0] node9230;
	wire [4-1:0] node9233;
	wire [4-1:0] node9236;
	wire [4-1:0] node9239;
	wire [4-1:0] node9240;
	wire [4-1:0] node9241;
	wire [4-1:0] node9243;
	wire [4-1:0] node9247;
	wire [4-1:0] node9248;
	wire [4-1:0] node9249;
	wire [4-1:0] node9253;
	wire [4-1:0] node9255;
	wire [4-1:0] node9258;
	wire [4-1:0] node9259;
	wire [4-1:0] node9260;
	wire [4-1:0] node9261;
	wire [4-1:0] node9265;
	wire [4-1:0] node9266;
	wire [4-1:0] node9267;
	wire [4-1:0] node9269;
	wire [4-1:0] node9273;
	wire [4-1:0] node9274;
	wire [4-1:0] node9276;
	wire [4-1:0] node9280;
	wire [4-1:0] node9281;
	wire [4-1:0] node9282;
	wire [4-1:0] node9283;
	wire [4-1:0] node9284;
	wire [4-1:0] node9287;
	wire [4-1:0] node9290;
	wire [4-1:0] node9293;
	wire [4-1:0] node9296;
	wire [4-1:0] node9297;
	wire [4-1:0] node9298;
	wire [4-1:0] node9302;
	wire [4-1:0] node9304;
	wire [4-1:0] node9307;
	wire [4-1:0] node9308;
	wire [4-1:0] node9309;
	wire [4-1:0] node9310;
	wire [4-1:0] node9311;
	wire [4-1:0] node9312;
	wire [4-1:0] node9313;
	wire [4-1:0] node9316;
	wire [4-1:0] node9318;
	wire [4-1:0] node9321;
	wire [4-1:0] node9322;
	wire [4-1:0] node9324;
	wire [4-1:0] node9327;
	wire [4-1:0] node9329;
	wire [4-1:0] node9332;
	wire [4-1:0] node9333;
	wire [4-1:0] node9334;
	wire [4-1:0] node9336;
	wire [4-1:0] node9339;
	wire [4-1:0] node9340;
	wire [4-1:0] node9344;
	wire [4-1:0] node9345;
	wire [4-1:0] node9346;
	wire [4-1:0] node9349;
	wire [4-1:0] node9350;
	wire [4-1:0] node9353;
	wire [4-1:0] node9356;
	wire [4-1:0] node9357;
	wire [4-1:0] node9360;
	wire [4-1:0] node9362;
	wire [4-1:0] node9365;
	wire [4-1:0] node9366;
	wire [4-1:0] node9367;
	wire [4-1:0] node9368;
	wire [4-1:0] node9369;
	wire [4-1:0] node9373;
	wire [4-1:0] node9375;
	wire [4-1:0] node9377;
	wire [4-1:0] node9380;
	wire [4-1:0] node9381;
	wire [4-1:0] node9382;
	wire [4-1:0] node9386;
	wire [4-1:0] node9388;
	wire [4-1:0] node9391;
	wire [4-1:0] node9392;
	wire [4-1:0] node9393;
	wire [4-1:0] node9395;
	wire [4-1:0] node9398;
	wire [4-1:0] node9399;
	wire [4-1:0] node9402;
	wire [4-1:0] node9403;
	wire [4-1:0] node9406;
	wire [4-1:0] node9409;
	wire [4-1:0] node9411;
	wire [4-1:0] node9412;
	wire [4-1:0] node9416;
	wire [4-1:0] node9417;
	wire [4-1:0] node9418;
	wire [4-1:0] node9419;
	wire [4-1:0] node9420;
	wire [4-1:0] node9423;
	wire [4-1:0] node9424;
	wire [4-1:0] node9426;
	wire [4-1:0] node9430;
	wire [4-1:0] node9431;
	wire [4-1:0] node9433;
	wire [4-1:0] node9436;
	wire [4-1:0] node9439;
	wire [4-1:0] node9440;
	wire [4-1:0] node9441;
	wire [4-1:0] node9443;
	wire [4-1:0] node9446;
	wire [4-1:0] node9448;
	wire [4-1:0] node9451;
	wire [4-1:0] node9452;
	wire [4-1:0] node9453;
	wire [4-1:0] node9455;
	wire [4-1:0] node9458;
	wire [4-1:0] node9459;
	wire [4-1:0] node9463;
	wire [4-1:0] node9464;
	wire [4-1:0] node9467;
	wire [4-1:0] node9470;
	wire [4-1:0] node9471;
	wire [4-1:0] node9472;
	wire [4-1:0] node9473;
	wire [4-1:0] node9476;
	wire [4-1:0] node9477;
	wire [4-1:0] node9478;
	wire [4-1:0] node9481;
	wire [4-1:0] node9484;
	wire [4-1:0] node9487;
	wire [4-1:0] node9488;
	wire [4-1:0] node9489;
	wire [4-1:0] node9493;
	wire [4-1:0] node9495;
	wire [4-1:0] node9498;
	wire [4-1:0] node9499;
	wire [4-1:0] node9500;
	wire [4-1:0] node9501;
	wire [4-1:0] node9503;
	wire [4-1:0] node9506;
	wire [4-1:0] node9509;
	wire [4-1:0] node9511;
	wire [4-1:0] node9512;
	wire [4-1:0] node9516;
	wire [4-1:0] node9517;
	wire [4-1:0] node9519;
	wire [4-1:0] node9522;
	wire [4-1:0] node9525;
	wire [4-1:0] node9526;
	wire [4-1:0] node9527;
	wire [4-1:0] node9528;
	wire [4-1:0] node9529;
	wire [4-1:0] node9530;
	wire [4-1:0] node9532;
	wire [4-1:0] node9535;
	wire [4-1:0] node9536;
	wire [4-1:0] node9540;
	wire [4-1:0] node9541;
	wire [4-1:0] node9542;
	wire [4-1:0] node9543;
	wire [4-1:0] node9547;
	wire [4-1:0] node9548;
	wire [4-1:0] node9551;
	wire [4-1:0] node9554;
	wire [4-1:0] node9556;
	wire [4-1:0] node9559;
	wire [4-1:0] node9560;
	wire [4-1:0] node9561;
	wire [4-1:0] node9564;
	wire [4-1:0] node9565;
	wire [4-1:0] node9568;
	wire [4-1:0] node9571;
	wire [4-1:0] node9572;
	wire [4-1:0] node9574;
	wire [4-1:0] node9577;
	wire [4-1:0] node9578;
	wire [4-1:0] node9579;
	wire [4-1:0] node9584;
	wire [4-1:0] node9585;
	wire [4-1:0] node9586;
	wire [4-1:0] node9587;
	wire [4-1:0] node9589;
	wire [4-1:0] node9592;
	wire [4-1:0] node9593;
	wire [4-1:0] node9595;
	wire [4-1:0] node9598;
	wire [4-1:0] node9599;
	wire [4-1:0] node9602;
	wire [4-1:0] node9605;
	wire [4-1:0] node9606;
	wire [4-1:0] node9607;
	wire [4-1:0] node9610;
	wire [4-1:0] node9611;
	wire [4-1:0] node9614;
	wire [4-1:0] node9617;
	wire [4-1:0] node9618;
	wire [4-1:0] node9619;
	wire [4-1:0] node9623;
	wire [4-1:0] node9624;
	wire [4-1:0] node9628;
	wire [4-1:0] node9629;
	wire [4-1:0] node9630;
	wire [4-1:0] node9632;
	wire [4-1:0] node9634;
	wire [4-1:0] node9637;
	wire [4-1:0] node9638;
	wire [4-1:0] node9641;
	wire [4-1:0] node9644;
	wire [4-1:0] node9645;
	wire [4-1:0] node9646;
	wire [4-1:0] node9649;
	wire [4-1:0] node9651;
	wire [4-1:0] node9654;
	wire [4-1:0] node9656;
	wire [4-1:0] node9657;
	wire [4-1:0] node9661;
	wire [4-1:0] node9662;
	wire [4-1:0] node9663;
	wire [4-1:0] node9664;
	wire [4-1:0] node9665;
	wire [4-1:0] node9667;
	wire [4-1:0] node9670;
	wire [4-1:0] node9672;
	wire [4-1:0] node9674;
	wire [4-1:0] node9677;
	wire [4-1:0] node9678;
	wire [4-1:0] node9681;
	wire [4-1:0] node9682;
	wire [4-1:0] node9686;
	wire [4-1:0] node9687;
	wire [4-1:0] node9689;
	wire [4-1:0] node9691;
	wire [4-1:0] node9694;
	wire [4-1:0] node9695;
	wire [4-1:0] node9698;
	wire [4-1:0] node9699;
	wire [4-1:0] node9700;
	wire [4-1:0] node9705;
	wire [4-1:0] node9706;
	wire [4-1:0] node9707;
	wire [4-1:0] node9708;
	wire [4-1:0] node9709;
	wire [4-1:0] node9712;
	wire [4-1:0] node9716;
	wire [4-1:0] node9717;
	wire [4-1:0] node9718;
	wire [4-1:0] node9721;
	wire [4-1:0] node9724;
	wire [4-1:0] node9727;
	wire [4-1:0] node9728;
	wire [4-1:0] node9729;
	wire [4-1:0] node9732;
	wire [4-1:0] node9735;
	wire [4-1:0] node9736;
	wire [4-1:0] node9737;
	wire [4-1:0] node9738;
	wire [4-1:0] node9741;
	wire [4-1:0] node9745;
	wire [4-1:0] node9748;
	wire [4-1:0] node9749;
	wire [4-1:0] node9750;
	wire [4-1:0] node9751;
	wire [4-1:0] node9752;
	wire [4-1:0] node9753;
	wire [4-1:0] node9754;
	wire [4-1:0] node9755;
	wire [4-1:0] node9756;
	wire [4-1:0] node9759;
	wire [4-1:0] node9762;
	wire [4-1:0] node9764;
	wire [4-1:0] node9767;
	wire [4-1:0] node9768;
	wire [4-1:0] node9769;
	wire [4-1:0] node9770;
	wire [4-1:0] node9774;
	wire [4-1:0] node9777;
	wire [4-1:0] node9778;
	wire [4-1:0] node9780;
	wire [4-1:0] node9783;
	wire [4-1:0] node9784;
	wire [4-1:0] node9788;
	wire [4-1:0] node9789;
	wire [4-1:0] node9790;
	wire [4-1:0] node9793;
	wire [4-1:0] node9795;
	wire [4-1:0] node9798;
	wire [4-1:0] node9799;
	wire [4-1:0] node9800;
	wire [4-1:0] node9803;
	wire [4-1:0] node9806;
	wire [4-1:0] node9807;
	wire [4-1:0] node9810;
	wire [4-1:0] node9812;
	wire [4-1:0] node9815;
	wire [4-1:0] node9816;
	wire [4-1:0] node9817;
	wire [4-1:0] node9818;
	wire [4-1:0] node9819;
	wire [4-1:0] node9823;
	wire [4-1:0] node9825;
	wire [4-1:0] node9828;
	wire [4-1:0] node9829;
	wire [4-1:0] node9832;
	wire [4-1:0] node9833;
	wire [4-1:0] node9834;
	wire [4-1:0] node9839;
	wire [4-1:0] node9840;
	wire [4-1:0] node9841;
	wire [4-1:0] node9842;
	wire [4-1:0] node9845;
	wire [4-1:0] node9847;
	wire [4-1:0] node9850;
	wire [4-1:0] node9853;
	wire [4-1:0] node9854;
	wire [4-1:0] node9856;
	wire [4-1:0] node9859;
	wire [4-1:0] node9862;
	wire [4-1:0] node9863;
	wire [4-1:0] node9864;
	wire [4-1:0] node9865;
	wire [4-1:0] node9866;
	wire [4-1:0] node9867;
	wire [4-1:0] node9871;
	wire [4-1:0] node9872;
	wire [4-1:0] node9876;
	wire [4-1:0] node9878;
	wire [4-1:0] node9879;
	wire [4-1:0] node9882;
	wire [4-1:0] node9883;
	wire [4-1:0] node9886;
	wire [4-1:0] node9889;
	wire [4-1:0] node9890;
	wire [4-1:0] node9891;
	wire [4-1:0] node9893;
	wire [4-1:0] node9895;
	wire [4-1:0] node9898;
	wire [4-1:0] node9901;
	wire [4-1:0] node9902;
	wire [4-1:0] node9903;
	wire [4-1:0] node9907;
	wire [4-1:0] node9908;
	wire [4-1:0] node9911;
	wire [4-1:0] node9912;
	wire [4-1:0] node9915;
	wire [4-1:0] node9918;
	wire [4-1:0] node9919;
	wire [4-1:0] node9920;
	wire [4-1:0] node9921;
	wire [4-1:0] node9924;
	wire [4-1:0] node9925;
	wire [4-1:0] node9928;
	wire [4-1:0] node9931;
	wire [4-1:0] node9932;
	wire [4-1:0] node9933;
	wire [4-1:0] node9937;
	wire [4-1:0] node9940;
	wire [4-1:0] node9941;
	wire [4-1:0] node9943;
	wire [4-1:0] node9946;
	wire [4-1:0] node9948;
	wire [4-1:0] node9951;
	wire [4-1:0] node9952;
	wire [4-1:0] node9953;
	wire [4-1:0] node9954;
	wire [4-1:0] node9955;
	wire [4-1:0] node9956;
	wire [4-1:0] node9959;
	wire [4-1:0] node9962;
	wire [4-1:0] node9963;
	wire [4-1:0] node9965;
	wire [4-1:0] node9968;
	wire [4-1:0] node9970;
	wire [4-1:0] node9971;
	wire [4-1:0] node9975;
	wire [4-1:0] node9976;
	wire [4-1:0] node9977;
	wire [4-1:0] node9978;
	wire [4-1:0] node9983;
	wire [4-1:0] node9984;
	wire [4-1:0] node9985;
	wire [4-1:0] node9986;
	wire [4-1:0] node9989;
	wire [4-1:0] node9993;
	wire [4-1:0] node9995;
	wire [4-1:0] node9997;
	wire [4-1:0] node10000;
	wire [4-1:0] node10001;
	wire [4-1:0] node10002;
	wire [4-1:0] node10003;
	wire [4-1:0] node10006;
	wire [4-1:0] node10009;
	wire [4-1:0] node10010;
	wire [4-1:0] node10011;
	wire [4-1:0] node10013;
	wire [4-1:0] node10017;
	wire [4-1:0] node10020;
	wire [4-1:0] node10021;
	wire [4-1:0] node10022;
	wire [4-1:0] node10024;
	wire [4-1:0] node10028;
	wire [4-1:0] node10029;
	wire [4-1:0] node10033;
	wire [4-1:0] node10034;
	wire [4-1:0] node10035;
	wire [4-1:0] node10036;
	wire [4-1:0] node10037;
	wire [4-1:0] node10041;
	wire [4-1:0] node10042;
	wire [4-1:0] node10043;
	wire [4-1:0] node10046;
	wire [4-1:0] node10049;
	wire [4-1:0] node10051;
	wire [4-1:0] node10054;
	wire [4-1:0] node10055;
	wire [4-1:0] node10056;
	wire [4-1:0] node10058;
	wire [4-1:0] node10061;
	wire [4-1:0] node10064;
	wire [4-1:0] node10065;
	wire [4-1:0] node10067;
	wire [4-1:0] node10070;
	wire [4-1:0] node10072;
	wire [4-1:0] node10075;
	wire [4-1:0] node10076;
	wire [4-1:0] node10077;
	wire [4-1:0] node10078;
	wire [4-1:0] node10079;
	wire [4-1:0] node10083;
	wire [4-1:0] node10085;
	wire [4-1:0] node10087;
	wire [4-1:0] node10090;
	wire [4-1:0] node10091;
	wire [4-1:0] node10092;
	wire [4-1:0] node10097;
	wire [4-1:0] node10098;
	wire [4-1:0] node10099;
	wire [4-1:0] node10104;
	wire [4-1:0] node10105;
	wire [4-1:0] node10106;
	wire [4-1:0] node10107;
	wire [4-1:0] node10108;
	wire [4-1:0] node10109;
	wire [4-1:0] node10110;
	wire [4-1:0] node10112;
	wire [4-1:0] node10115;
	wire [4-1:0] node10118;
	wire [4-1:0] node10119;
	wire [4-1:0] node10122;
	wire [4-1:0] node10125;
	wire [4-1:0] node10126;
	wire [4-1:0] node10129;
	wire [4-1:0] node10130;
	wire [4-1:0] node10132;
	wire [4-1:0] node10135;
	wire [4-1:0] node10138;
	wire [4-1:0] node10139;
	wire [4-1:0] node10140;
	wire [4-1:0] node10143;
	wire [4-1:0] node10144;
	wire [4-1:0] node10147;
	wire [4-1:0] node10150;
	wire [4-1:0] node10151;
	wire [4-1:0] node10152;
	wire [4-1:0] node10153;
	wire [4-1:0] node10154;
	wire [4-1:0] node10157;
	wire [4-1:0] node10160;
	wire [4-1:0] node10162;
	wire [4-1:0] node10165;
	wire [4-1:0] node10166;
	wire [4-1:0] node10170;
	wire [4-1:0] node10172;
	wire [4-1:0] node10173;
	wire [4-1:0] node10177;
	wire [4-1:0] node10178;
	wire [4-1:0] node10179;
	wire [4-1:0] node10180;
	wire [4-1:0] node10181;
	wire [4-1:0] node10184;
	wire [4-1:0] node10185;
	wire [4-1:0] node10189;
	wire [4-1:0] node10190;
	wire [4-1:0] node10192;
	wire [4-1:0] node10195;
	wire [4-1:0] node10196;
	wire [4-1:0] node10200;
	wire [4-1:0] node10201;
	wire [4-1:0] node10202;
	wire [4-1:0] node10203;
	wire [4-1:0] node10204;
	wire [4-1:0] node10209;
	wire [4-1:0] node10210;
	wire [4-1:0] node10214;
	wire [4-1:0] node10215;
	wire [4-1:0] node10216;
	wire [4-1:0] node10219;
	wire [4-1:0] node10222;
	wire [4-1:0] node10223;
	wire [4-1:0] node10227;
	wire [4-1:0] node10228;
	wire [4-1:0] node10229;
	wire [4-1:0] node10230;
	wire [4-1:0] node10231;
	wire [4-1:0] node10234;
	wire [4-1:0] node10237;
	wire [4-1:0] node10240;
	wire [4-1:0] node10241;
	wire [4-1:0] node10243;
	wire [4-1:0] node10246;
	wire [4-1:0] node10248;
	wire [4-1:0] node10251;
	wire [4-1:0] node10252;
	wire [4-1:0] node10253;
	wire [4-1:0] node10254;
	wire [4-1:0] node10257;
	wire [4-1:0] node10259;
	wire [4-1:0] node10262;
	wire [4-1:0] node10263;
	wire [4-1:0] node10265;
	wire [4-1:0] node10269;
	wire [4-1:0] node10270;
	wire [4-1:0] node10272;
	wire [4-1:0] node10275;
	wire [4-1:0] node10278;
	wire [4-1:0] node10279;
	wire [4-1:0] node10280;
	wire [4-1:0] node10281;
	wire [4-1:0] node10282;
	wire [4-1:0] node10283;
	wire [4-1:0] node10284;
	wire [4-1:0] node10288;
	wire [4-1:0] node10291;
	wire [4-1:0] node10292;
	wire [4-1:0] node10294;
	wire [4-1:0] node10297;
	wire [4-1:0] node10298;
	wire [4-1:0] node10301;
	wire [4-1:0] node10304;
	wire [4-1:0] node10305;
	wire [4-1:0] node10306;
	wire [4-1:0] node10307;
	wire [4-1:0] node10309;
	wire [4-1:0] node10313;
	wire [4-1:0] node10315;
	wire [4-1:0] node10318;
	wire [4-1:0] node10319;
	wire [4-1:0] node10321;
	wire [4-1:0] node10323;
	wire [4-1:0] node10326;
	wire [4-1:0] node10329;
	wire [4-1:0] node10330;
	wire [4-1:0] node10331;
	wire [4-1:0] node10332;
	wire [4-1:0] node10335;
	wire [4-1:0] node10336;
	wire [4-1:0] node10338;
	wire [4-1:0] node10341;
	wire [4-1:0] node10343;
	wire [4-1:0] node10346;
	wire [4-1:0] node10348;
	wire [4-1:0] node10351;
	wire [4-1:0] node10352;
	wire [4-1:0] node10353;
	wire [4-1:0] node10354;
	wire [4-1:0] node10358;
	wire [4-1:0] node10360;
	wire [4-1:0] node10362;
	wire [4-1:0] node10365;
	wire [4-1:0] node10366;
	wire [4-1:0] node10367;
	wire [4-1:0] node10368;
	wire [4-1:0] node10372;
	wire [4-1:0] node10373;
	wire [4-1:0] node10376;
	wire [4-1:0] node10379;
	wire [4-1:0] node10382;
	wire [4-1:0] node10383;
	wire [4-1:0] node10384;
	wire [4-1:0] node10385;
	wire [4-1:0] node10386;
	wire [4-1:0] node10389;
	wire [4-1:0] node10392;
	wire [4-1:0] node10394;
	wire [4-1:0] node10397;
	wire [4-1:0] node10398;
	wire [4-1:0] node10399;
	wire [4-1:0] node10400;
	wire [4-1:0] node10401;
	wire [4-1:0] node10405;
	wire [4-1:0] node10407;
	wire [4-1:0] node10411;
	wire [4-1:0] node10412;
	wire [4-1:0] node10415;
	wire [4-1:0] node10418;
	wire [4-1:0] node10419;
	wire [4-1:0] node10420;
	wire [4-1:0] node10421;
	wire [4-1:0] node10423;
	wire [4-1:0] node10426;
	wire [4-1:0] node10427;
	wire [4-1:0] node10431;
	wire [4-1:0] node10432;
	wire [4-1:0] node10433;
	wire [4-1:0] node10436;
	wire [4-1:0] node10439;
	wire [4-1:0] node10442;
	wire [4-1:0] node10443;
	wire [4-1:0] node10444;
	wire [4-1:0] node10445;
	wire [4-1:0] node10449;
	wire [4-1:0] node10450;
	wire [4-1:0] node10454;
	wire [4-1:0] node10455;
	wire [4-1:0] node10456;
	wire [4-1:0] node10459;
	wire [4-1:0] node10463;
	wire [4-1:0] node10464;
	wire [4-1:0] node10465;
	wire [4-1:0] node10466;
	wire [4-1:0] node10467;
	wire [4-1:0] node10468;
	wire [4-1:0] node10469;
	wire [4-1:0] node10470;
	wire [4-1:0] node10471;
	wire [4-1:0] node10472;
	wire [4-1:0] node10475;
	wire [4-1:0] node10476;
	wire [4-1:0] node10480;
	wire [4-1:0] node10481;
	wire [4-1:0] node10482;
	wire [4-1:0] node10486;
	wire [4-1:0] node10487;
	wire [4-1:0] node10488;
	wire [4-1:0] node10492;
	wire [4-1:0] node10495;
	wire [4-1:0] node10496;
	wire [4-1:0] node10497;
	wire [4-1:0] node10498;
	wire [4-1:0] node10499;
	wire [4-1:0] node10503;
	wire [4-1:0] node10505;
	wire [4-1:0] node10508;
	wire [4-1:0] node10511;
	wire [4-1:0] node10513;
	wire [4-1:0] node10514;
	wire [4-1:0] node10515;
	wire [4-1:0] node10518;
	wire [4-1:0] node10521;
	wire [4-1:0] node10522;
	wire [4-1:0] node10526;
	wire [4-1:0] node10527;
	wire [4-1:0] node10528;
	wire [4-1:0] node10529;
	wire [4-1:0] node10531;
	wire [4-1:0] node10534;
	wire [4-1:0] node10536;
	wire [4-1:0] node10537;
	wire [4-1:0] node10541;
	wire [4-1:0] node10542;
	wire [4-1:0] node10545;
	wire [4-1:0] node10546;
	wire [4-1:0] node10547;
	wire [4-1:0] node10550;
	wire [4-1:0] node10553;
	wire [4-1:0] node10554;
	wire [4-1:0] node10558;
	wire [4-1:0] node10559;
	wire [4-1:0] node10560;
	wire [4-1:0] node10562;
	wire [4-1:0] node10565;
	wire [4-1:0] node10567;
	wire [4-1:0] node10568;
	wire [4-1:0] node10572;
	wire [4-1:0] node10573;
	wire [4-1:0] node10575;
	wire [4-1:0] node10578;
	wire [4-1:0] node10580;
	wire [4-1:0] node10581;
	wire [4-1:0] node10585;
	wire [4-1:0] node10586;
	wire [4-1:0] node10587;
	wire [4-1:0] node10588;
	wire [4-1:0] node10589;
	wire [4-1:0] node10590;
	wire [4-1:0] node10592;
	wire [4-1:0] node10595;
	wire [4-1:0] node10596;
	wire [4-1:0] node10601;
	wire [4-1:0] node10603;
	wire [4-1:0] node10606;
	wire [4-1:0] node10607;
	wire [4-1:0] node10608;
	wire [4-1:0] node10609;
	wire [4-1:0] node10612;
	wire [4-1:0] node10616;
	wire [4-1:0] node10617;
	wire [4-1:0] node10618;
	wire [4-1:0] node10621;
	wire [4-1:0] node10622;
	wire [4-1:0] node10626;
	wire [4-1:0] node10628;
	wire [4-1:0] node10629;
	wire [4-1:0] node10633;
	wire [4-1:0] node10634;
	wire [4-1:0] node10635;
	wire [4-1:0] node10636;
	wire [4-1:0] node10637;
	wire [4-1:0] node10638;
	wire [4-1:0] node10643;
	wire [4-1:0] node10644;
	wire [4-1:0] node10646;
	wire [4-1:0] node10650;
	wire [4-1:0] node10651;
	wire [4-1:0] node10652;
	wire [4-1:0] node10653;
	wire [4-1:0] node10656;
	wire [4-1:0] node10659;
	wire [4-1:0] node10662;
	wire [4-1:0] node10663;
	wire [4-1:0] node10664;
	wire [4-1:0] node10667;
	wire [4-1:0] node10670;
	wire [4-1:0] node10672;
	wire [4-1:0] node10675;
	wire [4-1:0] node10676;
	wire [4-1:0] node10677;
	wire [4-1:0] node10678;
	wire [4-1:0] node10682;
	wire [4-1:0] node10683;
	wire [4-1:0] node10684;
	wire [4-1:0] node10689;
	wire [4-1:0] node10690;
	wire [4-1:0] node10691;
	wire [4-1:0] node10694;
	wire [4-1:0] node10697;
	wire [4-1:0] node10700;
	wire [4-1:0] node10701;
	wire [4-1:0] node10702;
	wire [4-1:0] node10703;
	wire [4-1:0] node10704;
	wire [4-1:0] node10705;
	wire [4-1:0] node10708;
	wire [4-1:0] node10711;
	wire [4-1:0] node10712;
	wire [4-1:0] node10714;
	wire [4-1:0] node10717;
	wire [4-1:0] node10718;
	wire [4-1:0] node10722;
	wire [4-1:0] node10723;
	wire [4-1:0] node10724;
	wire [4-1:0] node10726;
	wire [4-1:0] node10728;
	wire [4-1:0] node10731;
	wire [4-1:0] node10734;
	wire [4-1:0] node10735;
	wire [4-1:0] node10736;
	wire [4-1:0] node10739;
	wire [4-1:0] node10740;
	wire [4-1:0] node10744;
	wire [4-1:0] node10745;
	wire [4-1:0] node10749;
	wire [4-1:0] node10750;
	wire [4-1:0] node10751;
	wire [4-1:0] node10753;
	wire [4-1:0] node10756;
	wire [4-1:0] node10758;
	wire [4-1:0] node10759;
	wire [4-1:0] node10762;
	wire [4-1:0] node10765;
	wire [4-1:0] node10766;
	wire [4-1:0] node10767;
	wire [4-1:0] node10769;
	wire [4-1:0] node10773;
	wire [4-1:0] node10774;
	wire [4-1:0] node10775;
	wire [4-1:0] node10779;
	wire [4-1:0] node10781;
	wire [4-1:0] node10783;
	wire [4-1:0] node10786;
	wire [4-1:0] node10787;
	wire [4-1:0] node10788;
	wire [4-1:0] node10789;
	wire [4-1:0] node10790;
	wire [4-1:0] node10793;
	wire [4-1:0] node10794;
	wire [4-1:0] node10798;
	wire [4-1:0] node10799;
	wire [4-1:0] node10801;
	wire [4-1:0] node10804;
	wire [4-1:0] node10805;
	wire [4-1:0] node10806;
	wire [4-1:0] node10810;
	wire [4-1:0] node10813;
	wire [4-1:0] node10814;
	wire [4-1:0] node10815;
	wire [4-1:0] node10817;
	wire [4-1:0] node10820;
	wire [4-1:0] node10821;
	wire [4-1:0] node10825;
	wire [4-1:0] node10826;
	wire [4-1:0] node10828;
	wire [4-1:0] node10829;
	wire [4-1:0] node10832;
	wire [4-1:0] node10835;
	wire [4-1:0] node10837;
	wire [4-1:0] node10839;
	wire [4-1:0] node10842;
	wire [4-1:0] node10843;
	wire [4-1:0] node10844;
	wire [4-1:0] node10845;
	wire [4-1:0] node10847;
	wire [4-1:0] node10848;
	wire [4-1:0] node10852;
	wire [4-1:0] node10855;
	wire [4-1:0] node10856;
	wire [4-1:0] node10858;
	wire [4-1:0] node10861;
	wire [4-1:0] node10862;
	wire [4-1:0] node10864;
	wire [4-1:0] node10868;
	wire [4-1:0] node10869;
	wire [4-1:0] node10870;
	wire [4-1:0] node10871;
	wire [4-1:0] node10874;
	wire [4-1:0] node10875;
	wire [4-1:0] node10878;
	wire [4-1:0] node10882;
	wire [4-1:0] node10883;
	wire [4-1:0] node10886;
	wire [4-1:0] node10887;
	wire [4-1:0] node10891;
	wire [4-1:0] node10892;
	wire [4-1:0] node10893;
	wire [4-1:0] node10894;
	wire [4-1:0] node10895;
	wire [4-1:0] node10898;
	wire [4-1:0] node10899;
	wire [4-1:0] node10901;
	wire [4-1:0] node10904;
	wire [4-1:0] node10905;
	wire [4-1:0] node10909;
	wire [4-1:0] node10910;
	wire [4-1:0] node10911;
	wire [4-1:0] node10912;
	wire [4-1:0] node10915;
	wire [4-1:0] node10918;
	wire [4-1:0] node10919;
	wire [4-1:0] node10921;
	wire [4-1:0] node10922;
	wire [4-1:0] node10925;
	wire [4-1:0] node10928;
	wire [4-1:0] node10930;
	wire [4-1:0] node10933;
	wire [4-1:0] node10934;
	wire [4-1:0] node10935;
	wire [4-1:0] node10939;
	wire [4-1:0] node10941;
	wire [4-1:0] node10944;
	wire [4-1:0] node10945;
	wire [4-1:0] node10946;
	wire [4-1:0] node10949;
	wire [4-1:0] node10950;
	wire [4-1:0] node10952;
	wire [4-1:0] node10955;
	wire [4-1:0] node10956;
	wire [4-1:0] node10960;
	wire [4-1:0] node10961;
	wire [4-1:0] node10962;
	wire [4-1:0] node10963;
	wire [4-1:0] node10965;
	wire [4-1:0] node10968;
	wire [4-1:0] node10971;
	wire [4-1:0] node10972;
	wire [4-1:0] node10974;
	wire [4-1:0] node10977;
	wire [4-1:0] node10980;
	wire [4-1:0] node10981;
	wire [4-1:0] node10982;
	wire [4-1:0] node10986;
	wire [4-1:0] node10988;
	wire [4-1:0] node10991;
	wire [4-1:0] node10992;
	wire [4-1:0] node10993;
	wire [4-1:0] node10994;
	wire [4-1:0] node10995;
	wire [4-1:0] node10996;
	wire [4-1:0] node10997;
	wire [4-1:0] node11001;
	wire [4-1:0] node11002;
	wire [4-1:0] node11003;
	wire [4-1:0] node11008;
	wire [4-1:0] node11009;
	wire [4-1:0] node11010;
	wire [4-1:0] node11013;
	wire [4-1:0] node11016;
	wire [4-1:0] node11017;
	wire [4-1:0] node11020;
	wire [4-1:0] node11021;
	wire [4-1:0] node11025;
	wire [4-1:0] node11026;
	wire [4-1:0] node11028;
	wire [4-1:0] node11030;
	wire [4-1:0] node11033;
	wire [4-1:0] node11034;
	wire [4-1:0] node11035;
	wire [4-1:0] node11036;
	wire [4-1:0] node11040;
	wire [4-1:0] node11044;
	wire [4-1:0] node11045;
	wire [4-1:0] node11046;
	wire [4-1:0] node11047;
	wire [4-1:0] node11050;
	wire [4-1:0] node11053;
	wire [4-1:0] node11054;
	wire [4-1:0] node11056;
	wire [4-1:0] node11059;
	wire [4-1:0] node11062;
	wire [4-1:0] node11063;
	wire [4-1:0] node11064;
	wire [4-1:0] node11067;
	wire [4-1:0] node11068;
	wire [4-1:0] node11070;
	wire [4-1:0] node11074;
	wire [4-1:0] node11075;
	wire [4-1:0] node11077;
	wire [4-1:0] node11080;
	wire [4-1:0] node11082;
	wire [4-1:0] node11085;
	wire [4-1:0] node11086;
	wire [4-1:0] node11087;
	wire [4-1:0] node11088;
	wire [4-1:0] node11089;
	wire [4-1:0] node11092;
	wire [4-1:0] node11093;
	wire [4-1:0] node11096;
	wire [4-1:0] node11098;
	wire [4-1:0] node11101;
	wire [4-1:0] node11103;
	wire [4-1:0] node11105;
	wire [4-1:0] node11108;
	wire [4-1:0] node11109;
	wire [4-1:0] node11110;
	wire [4-1:0] node11112;
	wire [4-1:0] node11113;
	wire [4-1:0] node11116;
	wire [4-1:0] node11119;
	wire [4-1:0] node11120;
	wire [4-1:0] node11122;
	wire [4-1:0] node11125;
	wire [4-1:0] node11128;
	wire [4-1:0] node11129;
	wire [4-1:0] node11132;
	wire [4-1:0] node11135;
	wire [4-1:0] node11136;
	wire [4-1:0] node11137;
	wire [4-1:0] node11138;
	wire [4-1:0] node11141;
	wire [4-1:0] node11144;
	wire [4-1:0] node11145;
	wire [4-1:0] node11146;
	wire [4-1:0] node11150;
	wire [4-1:0] node11151;
	wire [4-1:0] node11155;
	wire [4-1:0] node11156;
	wire [4-1:0] node11158;
	wire [4-1:0] node11161;
	wire [4-1:0] node11163;
	wire [4-1:0] node11166;
	wire [4-1:0] node11167;
	wire [4-1:0] node11168;
	wire [4-1:0] node11169;
	wire [4-1:0] node11170;
	wire [4-1:0] node11171;
	wire [4-1:0] node11172;
	wire [4-1:0] node11173;
	wire [4-1:0] node11174;
	wire [4-1:0] node11175;
	wire [4-1:0] node11178;
	wire [4-1:0] node11182;
	wire [4-1:0] node11184;
	wire [4-1:0] node11185;
	wire [4-1:0] node11189;
	wire [4-1:0] node11190;
	wire [4-1:0] node11193;
	wire [4-1:0] node11196;
	wire [4-1:0] node11197;
	wire [4-1:0] node11198;
	wire [4-1:0] node11199;
	wire [4-1:0] node11200;
	wire [4-1:0] node11203;
	wire [4-1:0] node11206;
	wire [4-1:0] node11207;
	wire [4-1:0] node11210;
	wire [4-1:0] node11213;
	wire [4-1:0] node11215;
	wire [4-1:0] node11216;
	wire [4-1:0] node11220;
	wire [4-1:0] node11221;
	wire [4-1:0] node11222;
	wire [4-1:0] node11223;
	wire [4-1:0] node11227;
	wire [4-1:0] node11228;
	wire [4-1:0] node11232;
	wire [4-1:0] node11233;
	wire [4-1:0] node11236;
	wire [4-1:0] node11239;
	wire [4-1:0] node11240;
	wire [4-1:0] node11241;
	wire [4-1:0] node11242;
	wire [4-1:0] node11243;
	wire [4-1:0] node11245;
	wire [4-1:0] node11249;
	wire [4-1:0] node11251;
	wire [4-1:0] node11254;
	wire [4-1:0] node11255;
	wire [4-1:0] node11257;
	wire [4-1:0] node11260;
	wire [4-1:0] node11262;
	wire [4-1:0] node11265;
	wire [4-1:0] node11266;
	wire [4-1:0] node11267;
	wire [4-1:0] node11268;
	wire [4-1:0] node11272;
	wire [4-1:0] node11275;
	wire [4-1:0] node11277;
	wire [4-1:0] node11278;
	wire [4-1:0] node11279;
	wire [4-1:0] node11283;
	wire [4-1:0] node11284;
	wire [4-1:0] node11288;
	wire [4-1:0] node11289;
	wire [4-1:0] node11290;
	wire [4-1:0] node11291;
	wire [4-1:0] node11292;
	wire [4-1:0] node11293;
	wire [4-1:0] node11297;
	wire [4-1:0] node11298;
	wire [4-1:0] node11301;
	wire [4-1:0] node11304;
	wire [4-1:0] node11305;
	wire [4-1:0] node11306;
	wire [4-1:0] node11308;
	wire [4-1:0] node11312;
	wire [4-1:0] node11313;
	wire [4-1:0] node11316;
	wire [4-1:0] node11319;
	wire [4-1:0] node11320;
	wire [4-1:0] node11321;
	wire [4-1:0] node11323;
	wire [4-1:0] node11325;
	wire [4-1:0] node11328;
	wire [4-1:0] node11331;
	wire [4-1:0] node11332;
	wire [4-1:0] node11334;
	wire [4-1:0] node11335;
	wire [4-1:0] node11338;
	wire [4-1:0] node11341;
	wire [4-1:0] node11343;
	wire [4-1:0] node11346;
	wire [4-1:0] node11347;
	wire [4-1:0] node11348;
	wire [4-1:0] node11350;
	wire [4-1:0] node11352;
	wire [4-1:0] node11354;
	wire [4-1:0] node11357;
	wire [4-1:0] node11358;
	wire [4-1:0] node11359;
	wire [4-1:0] node11361;
	wire [4-1:0] node11365;
	wire [4-1:0] node11366;
	wire [4-1:0] node11370;
	wire [4-1:0] node11371;
	wire [4-1:0] node11372;
	wire [4-1:0] node11375;
	wire [4-1:0] node11377;
	wire [4-1:0] node11378;
	wire [4-1:0] node11381;
	wire [4-1:0] node11384;
	wire [4-1:0] node11385;
	wire [4-1:0] node11389;
	wire [4-1:0] node11390;
	wire [4-1:0] node11391;
	wire [4-1:0] node11392;
	wire [4-1:0] node11393;
	wire [4-1:0] node11395;
	wire [4-1:0] node11396;
	wire [4-1:0] node11397;
	wire [4-1:0] node11401;
	wire [4-1:0] node11404;
	wire [4-1:0] node11405;
	wire [4-1:0] node11406;
	wire [4-1:0] node11407;
	wire [4-1:0] node11411;
	wire [4-1:0] node11414;
	wire [4-1:0] node11415;
	wire [4-1:0] node11418;
	wire [4-1:0] node11420;
	wire [4-1:0] node11423;
	wire [4-1:0] node11424;
	wire [4-1:0] node11425;
	wire [4-1:0] node11428;
	wire [4-1:0] node11429;
	wire [4-1:0] node11430;
	wire [4-1:0] node11433;
	wire [4-1:0] node11436;
	wire [4-1:0] node11437;
	wire [4-1:0] node11441;
	wire [4-1:0] node11442;
	wire [4-1:0] node11443;
	wire [4-1:0] node11444;
	wire [4-1:0] node11448;
	wire [4-1:0] node11449;
	wire [4-1:0] node11452;
	wire [4-1:0] node11455;
	wire [4-1:0] node11456;
	wire [4-1:0] node11458;
	wire [4-1:0] node11461;
	wire [4-1:0] node11462;
	wire [4-1:0] node11466;
	wire [4-1:0] node11467;
	wire [4-1:0] node11468;
	wire [4-1:0] node11470;
	wire [4-1:0] node11473;
	wire [4-1:0] node11474;
	wire [4-1:0] node11475;
	wire [4-1:0] node11476;
	wire [4-1:0] node11479;
	wire [4-1:0] node11484;
	wire [4-1:0] node11485;
	wire [4-1:0] node11486;
	wire [4-1:0] node11488;
	wire [4-1:0] node11493;
	wire [4-1:0] node11494;
	wire [4-1:0] node11495;
	wire [4-1:0] node11496;
	wire [4-1:0] node11497;
	wire [4-1:0] node11498;
	wire [4-1:0] node11502;
	wire [4-1:0] node11503;
	wire [4-1:0] node11507;
	wire [4-1:0] node11508;
	wire [4-1:0] node11509;
	wire [4-1:0] node11510;
	wire [4-1:0] node11513;
	wire [4-1:0] node11516;
	wire [4-1:0] node11518;
	wire [4-1:0] node11521;
	wire [4-1:0] node11522;
	wire [4-1:0] node11526;
	wire [4-1:0] node11527;
	wire [4-1:0] node11528;
	wire [4-1:0] node11529;
	wire [4-1:0] node11532;
	wire [4-1:0] node11533;
	wire [4-1:0] node11536;
	wire [4-1:0] node11539;
	wire [4-1:0] node11540;
	wire [4-1:0] node11544;
	wire [4-1:0] node11545;
	wire [4-1:0] node11546;
	wire [4-1:0] node11549;
	wire [4-1:0] node11552;
	wire [4-1:0] node11554;
	wire [4-1:0] node11557;
	wire [4-1:0] node11558;
	wire [4-1:0] node11559;
	wire [4-1:0] node11560;
	wire [4-1:0] node11561;
	wire [4-1:0] node11564;
	wire [4-1:0] node11567;
	wire [4-1:0] node11568;
	wire [4-1:0] node11572;
	wire [4-1:0] node11573;
	wire [4-1:0] node11574;
	wire [4-1:0] node11577;
	wire [4-1:0] node11581;
	wire [4-1:0] node11582;
	wire [4-1:0] node11583;
	wire [4-1:0] node11584;
	wire [4-1:0] node11586;
	wire [4-1:0] node11589;
	wire [4-1:0] node11592;
	wire [4-1:0] node11593;
	wire [4-1:0] node11594;
	wire [4-1:0] node11597;
	wire [4-1:0] node11601;
	wire [4-1:0] node11602;
	wire [4-1:0] node11603;
	wire [4-1:0] node11606;
	wire [4-1:0] node11610;
	wire [4-1:0] node11611;
	wire [4-1:0] node11612;
	wire [4-1:0] node11613;
	wire [4-1:0] node11614;
	wire [4-1:0] node11615;
	wire [4-1:0] node11616;
	wire [4-1:0] node11617;
	wire [4-1:0] node11618;
	wire [4-1:0] node11622;
	wire [4-1:0] node11625;
	wire [4-1:0] node11626;
	wire [4-1:0] node11627;
	wire [4-1:0] node11632;
	wire [4-1:0] node11633;
	wire [4-1:0] node11634;
	wire [4-1:0] node11636;
	wire [4-1:0] node11639;
	wire [4-1:0] node11640;
	wire [4-1:0] node11644;
	wire [4-1:0] node11645;
	wire [4-1:0] node11648;
	wire [4-1:0] node11651;
	wire [4-1:0] node11652;
	wire [4-1:0] node11653;
	wire [4-1:0] node11654;
	wire [4-1:0] node11658;
	wire [4-1:0] node11659;
	wire [4-1:0] node11661;
	wire [4-1:0] node11665;
	wire [4-1:0] node11666;
	wire [4-1:0] node11669;
	wire [4-1:0] node11670;
	wire [4-1:0] node11674;
	wire [4-1:0] node11675;
	wire [4-1:0] node11676;
	wire [4-1:0] node11677;
	wire [4-1:0] node11678;
	wire [4-1:0] node11679;
	wire [4-1:0] node11683;
	wire [4-1:0] node11686;
	wire [4-1:0] node11689;
	wire [4-1:0] node11690;
	wire [4-1:0] node11691;
	wire [4-1:0] node11692;
	wire [4-1:0] node11697;
	wire [4-1:0] node11698;
	wire [4-1:0] node11699;
	wire [4-1:0] node11703;
	wire [4-1:0] node11706;
	wire [4-1:0] node11707;
	wire [4-1:0] node11708;
	wire [4-1:0] node11710;
	wire [4-1:0] node11713;
	wire [4-1:0] node11715;
	wire [4-1:0] node11716;
	wire [4-1:0] node11719;
	wire [4-1:0] node11722;
	wire [4-1:0] node11723;
	wire [4-1:0] node11725;
	wire [4-1:0] node11728;
	wire [4-1:0] node11730;
	wire [4-1:0] node11733;
	wire [4-1:0] node11734;
	wire [4-1:0] node11735;
	wire [4-1:0] node11736;
	wire [4-1:0] node11737;
	wire [4-1:0] node11738;
	wire [4-1:0] node11739;
	wire [4-1:0] node11744;
	wire [4-1:0] node11745;
	wire [4-1:0] node11749;
	wire [4-1:0] node11750;
	wire [4-1:0] node11752;
	wire [4-1:0] node11755;
	wire [4-1:0] node11757;
	wire [4-1:0] node11759;
	wire [4-1:0] node11762;
	wire [4-1:0] node11763;
	wire [4-1:0] node11764;
	wire [4-1:0] node11765;
	wire [4-1:0] node11769;
	wire [4-1:0] node11770;
	wire [4-1:0] node11773;
	wire [4-1:0] node11776;
	wire [4-1:0] node11777;
	wire [4-1:0] node11778;
	wire [4-1:0] node11779;
	wire [4-1:0] node11784;
	wire [4-1:0] node11785;
	wire [4-1:0] node11787;
	wire [4-1:0] node11791;
	wire [4-1:0] node11792;
	wire [4-1:0] node11793;
	wire [4-1:0] node11794;
	wire [4-1:0] node11797;
	wire [4-1:0] node11798;
	wire [4-1:0] node11801;
	wire [4-1:0] node11802;
	wire [4-1:0] node11806;
	wire [4-1:0] node11807;
	wire [4-1:0] node11809;
	wire [4-1:0] node11812;
	wire [4-1:0] node11813;
	wire [4-1:0] node11817;
	wire [4-1:0] node11818;
	wire [4-1:0] node11819;
	wire [4-1:0] node11820;
	wire [4-1:0] node11822;
	wire [4-1:0] node11825;
	wire [4-1:0] node11828;
	wire [4-1:0] node11830;
	wire [4-1:0] node11831;
	wire [4-1:0] node11834;
	wire [4-1:0] node11837;
	wire [4-1:0] node11838;
	wire [4-1:0] node11839;
	wire [4-1:0] node11842;
	wire [4-1:0] node11843;
	wire [4-1:0] node11846;
	wire [4-1:0] node11849;
	wire [4-1:0] node11850;
	wire [4-1:0] node11854;
	wire [4-1:0] node11855;
	wire [4-1:0] node11856;
	wire [4-1:0] node11857;
	wire [4-1:0] node11858;
	wire [4-1:0] node11859;
	wire [4-1:0] node11860;
	wire [4-1:0] node11863;
	wire [4-1:0] node11865;
	wire [4-1:0] node11868;
	wire [4-1:0] node11871;
	wire [4-1:0] node11872;
	wire [4-1:0] node11873;
	wire [4-1:0] node11875;
	wire [4-1:0] node11878;
	wire [4-1:0] node11881;
	wire [4-1:0] node11883;
	wire [4-1:0] node11884;
	wire [4-1:0] node11888;
	wire [4-1:0] node11889;
	wire [4-1:0] node11891;
	wire [4-1:0] node11892;
	wire [4-1:0] node11894;
	wire [4-1:0] node11897;
	wire [4-1:0] node11900;
	wire [4-1:0] node11901;
	wire [4-1:0] node11903;
	wire [4-1:0] node11905;
	wire [4-1:0] node11908;
	wire [4-1:0] node11911;
	wire [4-1:0] node11912;
	wire [4-1:0] node11913;
	wire [4-1:0] node11916;
	wire [4-1:0] node11917;
	wire [4-1:0] node11918;
	wire [4-1:0] node11920;
	wire [4-1:0] node11923;
	wire [4-1:0] node11926;
	wire [4-1:0] node11927;
	wire [4-1:0] node11930;
	wire [4-1:0] node11933;
	wire [4-1:0] node11934;
	wire [4-1:0] node11935;
	wire [4-1:0] node11936;
	wire [4-1:0] node11938;
	wire [4-1:0] node11941;
	wire [4-1:0] node11943;
	wire [4-1:0] node11946;
	wire [4-1:0] node11947;
	wire [4-1:0] node11951;
	wire [4-1:0] node11952;
	wire [4-1:0] node11954;
	wire [4-1:0] node11957;
	wire [4-1:0] node11958;
	wire [4-1:0] node11961;
	wire [4-1:0] node11964;
	wire [4-1:0] node11965;
	wire [4-1:0] node11966;
	wire [4-1:0] node11967;
	wire [4-1:0] node11968;
	wire [4-1:0] node11971;
	wire [4-1:0] node11974;
	wire [4-1:0] node11975;
	wire [4-1:0] node11978;
	wire [4-1:0] node11980;
	wire [4-1:0] node11981;
	wire [4-1:0] node11985;
	wire [4-1:0] node11986;
	wire [4-1:0] node11987;
	wire [4-1:0] node11989;
	wire [4-1:0] node11993;
	wire [4-1:0] node11994;
	wire [4-1:0] node11996;
	wire [4-1:0] node11997;
	wire [4-1:0] node12002;
	wire [4-1:0] node12003;
	wire [4-1:0] node12004;
	wire [4-1:0] node12006;
	wire [4-1:0] node12008;
	wire [4-1:0] node12009;
	wire [4-1:0] node12013;
	wire [4-1:0] node12014;
	wire [4-1:0] node12015;
	wire [4-1:0] node12019;
	wire [4-1:0] node12020;
	wire [4-1:0] node12023;
	wire [4-1:0] node12026;
	wire [4-1:0] node12027;
	wire [4-1:0] node12028;
	wire [4-1:0] node12029;
	wire [4-1:0] node12030;
	wire [4-1:0] node12033;
	wire [4-1:0] node12037;
	wire [4-1:0] node12038;
	wire [4-1:0] node12039;
	wire [4-1:0] node12042;
	wire [4-1:0] node12046;
	wire [4-1:0] node12049;
	wire [4-1:0] node12050;
	wire [4-1:0] node12051;
	wire [4-1:0] node12052;
	wire [4-1:0] node12053;
	wire [4-1:0] node12054;
	wire [4-1:0] node12055;
	wire [4-1:0] node12056;
	wire [4-1:0] node12059;
	wire [4-1:0] node12061;
	wire [4-1:0] node12064;
	wire [4-1:0] node12065;
	wire [4-1:0] node12066;
	wire [4-1:0] node12067;
	wire [4-1:0] node12068;
	wire [4-1:0] node12072;
	wire [4-1:0] node12075;
	wire [4-1:0] node12077;
	wire [4-1:0] node12080;
	wire [4-1:0] node12081;
	wire [4-1:0] node12084;
	wire [4-1:0] node12087;
	wire [4-1:0] node12088;
	wire [4-1:0] node12089;
	wire [4-1:0] node12091;
	wire [4-1:0] node12095;
	wire [4-1:0] node12096;
	wire [4-1:0] node12099;
	wire [4-1:0] node12100;
	wire [4-1:0] node12101;
	wire [4-1:0] node12104;
	wire [4-1:0] node12107;
	wire [4-1:0] node12109;
	wire [4-1:0] node12111;
	wire [4-1:0] node12114;
	wire [4-1:0] node12115;
	wire [4-1:0] node12116;
	wire [4-1:0] node12117;
	wire [4-1:0] node12118;
	wire [4-1:0] node12121;
	wire [4-1:0] node12124;
	wire [4-1:0] node12126;
	wire [4-1:0] node12129;
	wire [4-1:0] node12130;
	wire [4-1:0] node12132;
	wire [4-1:0] node12133;
	wire [4-1:0] node12134;
	wire [4-1:0] node12138;
	wire [4-1:0] node12139;
	wire [4-1:0] node12143;
	wire [4-1:0] node12144;
	wire [4-1:0] node12147;
	wire [4-1:0] node12150;
	wire [4-1:0] node12151;
	wire [4-1:0] node12152;
	wire [4-1:0] node12154;
	wire [4-1:0] node12158;
	wire [4-1:0] node12159;
	wire [4-1:0] node12161;
	wire [4-1:0] node12164;
	wire [4-1:0] node12166;
	wire [4-1:0] node12168;
	wire [4-1:0] node12169;
	wire [4-1:0] node12173;
	wire [4-1:0] node12174;
	wire [4-1:0] node12175;
	wire [4-1:0] node12176;
	wire [4-1:0] node12177;
	wire [4-1:0] node12179;
	wire [4-1:0] node12182;
	wire [4-1:0] node12184;
	wire [4-1:0] node12185;
	wire [4-1:0] node12186;
	wire [4-1:0] node12191;
	wire [4-1:0] node12192;
	wire [4-1:0] node12194;
	wire [4-1:0] node12198;
	wire [4-1:0] node12199;
	wire [4-1:0] node12200;
	wire [4-1:0] node12201;
	wire [4-1:0] node12202;
	wire [4-1:0] node12206;
	wire [4-1:0] node12208;
	wire [4-1:0] node12209;
	wire [4-1:0] node12213;
	wire [4-1:0] node12214;
	wire [4-1:0] node12217;
	wire [4-1:0] node12220;
	wire [4-1:0] node12221;
	wire [4-1:0] node12222;
	wire [4-1:0] node12226;
	wire [4-1:0] node12227;
	wire [4-1:0] node12230;
	wire [4-1:0] node12233;
	wire [4-1:0] node12234;
	wire [4-1:0] node12235;
	wire [4-1:0] node12236;
	wire [4-1:0] node12237;
	wire [4-1:0] node12240;
	wire [4-1:0] node12241;
	wire [4-1:0] node12242;
	wire [4-1:0] node12246;
	wire [4-1:0] node12248;
	wire [4-1:0] node12251;
	wire [4-1:0] node12252;
	wire [4-1:0] node12254;
	wire [4-1:0] node12258;
	wire [4-1:0] node12259;
	wire [4-1:0] node12260;
	wire [4-1:0] node12262;
	wire [4-1:0] node12266;
	wire [4-1:0] node12267;
	wire [4-1:0] node12268;
	wire [4-1:0] node12272;
	wire [4-1:0] node12275;
	wire [4-1:0] node12276;
	wire [4-1:0] node12277;
	wire [4-1:0] node12280;
	wire [4-1:0] node12281;
	wire [4-1:0] node12282;
	wire [4-1:0] node12283;
	wire [4-1:0] node12286;
	wire [4-1:0] node12290;
	wire [4-1:0] node12291;
	wire [4-1:0] node12294;
	wire [4-1:0] node12297;
	wire [4-1:0] node12298;
	wire [4-1:0] node12299;
	wire [4-1:0] node12304;
	wire [4-1:0] node12305;
	wire [4-1:0] node12306;
	wire [4-1:0] node12307;
	wire [4-1:0] node12308;
	wire [4-1:0] node12309;
	wire [4-1:0] node12312;
	wire [4-1:0] node12315;
	wire [4-1:0] node12316;
	wire [4-1:0] node12318;
	wire [4-1:0] node12321;
	wire [4-1:0] node12322;
	wire [4-1:0] node12326;
	wire [4-1:0] node12327;
	wire [4-1:0] node12329;
	wire [4-1:0] node12332;
	wire [4-1:0] node12333;
	wire [4-1:0] node12337;
	wire [4-1:0] node12338;
	wire [4-1:0] node12339;
	wire [4-1:0] node12342;
	wire [4-1:0] node12343;
	wire [4-1:0] node12345;
	wire [4-1:0] node12346;
	wire [4-1:0] node12349;
	wire [4-1:0] node12352;
	wire [4-1:0] node12354;
	wire [4-1:0] node12357;
	wire [4-1:0] node12358;
	wire [4-1:0] node12362;
	wire [4-1:0] node12363;
	wire [4-1:0] node12364;
	wire [4-1:0] node12365;
	wire [4-1:0] node12366;
	wire [4-1:0] node12370;
	wire [4-1:0] node12371;
	wire [4-1:0] node12375;
	wire [4-1:0] node12376;
	wire [4-1:0] node12377;
	wire [4-1:0] node12380;
	wire [4-1:0] node12383;
	wire [4-1:0] node12386;
	wire [4-1:0] node12387;
	wire [4-1:0] node12388;
	wire [4-1:0] node12389;
	wire [4-1:0] node12392;
	wire [4-1:0] node12395;
	wire [4-1:0] node12396;
	wire [4-1:0] node12399;
	wire [4-1:0] node12402;
	wire [4-1:0] node12403;
	wire [4-1:0] node12404;
	wire [4-1:0] node12407;
	wire [4-1:0] node12410;
	wire [4-1:0] node12413;
	wire [4-1:0] node12414;
	wire [4-1:0] node12415;
	wire [4-1:0] node12416;
	wire [4-1:0] node12417;
	wire [4-1:0] node12418;
	wire [4-1:0] node12419;
	wire [4-1:0] node12421;
	wire [4-1:0] node12424;
	wire [4-1:0] node12426;
	wire [4-1:0] node12429;
	wire [4-1:0] node12430;
	wire [4-1:0] node12432;
	wire [4-1:0] node12435;
	wire [4-1:0] node12437;
	wire [4-1:0] node12440;
	wire [4-1:0] node12441;
	wire [4-1:0] node12442;
	wire [4-1:0] node12443;
	wire [4-1:0] node12446;
	wire [4-1:0] node12449;
	wire [4-1:0] node12450;
	wire [4-1:0] node12451;
	wire [4-1:0] node12452;
	wire [4-1:0] node12455;
	wire [4-1:0] node12460;
	wire [4-1:0] node12461;
	wire [4-1:0] node12462;
	wire [4-1:0] node12465;
	wire [4-1:0] node12468;
	wire [4-1:0] node12470;
	wire [4-1:0] node12471;
	wire [4-1:0] node12475;
	wire [4-1:0] node12476;
	wire [4-1:0] node12477;
	wire [4-1:0] node12479;
	wire [4-1:0] node12482;
	wire [4-1:0] node12484;
	wire [4-1:0] node12487;
	wire [4-1:0] node12488;
	wire [4-1:0] node12489;
	wire [4-1:0] node12493;
	wire [4-1:0] node12495;
	wire [4-1:0] node12498;
	wire [4-1:0] node12499;
	wire [4-1:0] node12500;
	wire [4-1:0] node12501;
	wire [4-1:0] node12504;
	wire [4-1:0] node12507;
	wire [4-1:0] node12508;
	wire [4-1:0] node12511;
	wire [4-1:0] node12514;
	wire [4-1:0] node12515;
	wire [4-1:0] node12518;
	wire [4-1:0] node12521;
	wire [4-1:0] node12522;
	wire [4-1:0] node12523;
	wire [4-1:0] node12524;
	wire [4-1:0] node12525;
	wire [4-1:0] node12526;
	wire [4-1:0] node12528;
	wire [4-1:0] node12529;
	wire [4-1:0] node12533;
	wire [4-1:0] node12534;
	wire [4-1:0] node12536;
	wire [4-1:0] node12537;
	wire [4-1:0] node12540;
	wire [4-1:0] node12543;
	wire [4-1:0] node12544;
	wire [4-1:0] node12547;
	wire [4-1:0] node12550;
	wire [4-1:0] node12551;
	wire [4-1:0] node12552;
	wire [4-1:0] node12554;
	wire [4-1:0] node12557;
	wire [4-1:0] node12558;
	wire [4-1:0] node12559;
	wire [4-1:0] node12564;
	wire [4-1:0] node12565;
	wire [4-1:0] node12566;
	wire [4-1:0] node12568;
	wire [4-1:0] node12571;
	wire [4-1:0] node12572;
	wire [4-1:0] node12576;
	wire [4-1:0] node12578;
	wire [4-1:0] node12580;
	wire [4-1:0] node12583;
	wire [4-1:0] node12584;
	wire [4-1:0] node12585;
	wire [4-1:0] node12586;
	wire [4-1:0] node12587;
	wire [4-1:0] node12591;
	wire [4-1:0] node12592;
	wire [4-1:0] node12596;
	wire [4-1:0] node12597;
	wire [4-1:0] node12598;
	wire [4-1:0] node12603;
	wire [4-1:0] node12604;
	wire [4-1:0] node12606;
	wire [4-1:0] node12607;
	wire [4-1:0] node12610;
	wire [4-1:0] node12613;
	wire [4-1:0] node12615;
	wire [4-1:0] node12616;
	wire [4-1:0] node12618;
	wire [4-1:0] node12622;
	wire [4-1:0] node12623;
	wire [4-1:0] node12626;
	wire [4-1:0] node12629;
	wire [4-1:0] node12630;
	wire [4-1:0] node12631;
	wire [4-1:0] node12632;
	wire [4-1:0] node12633;
	wire [4-1:0] node12637;
	wire [4-1:0] node12638;
	wire [4-1:0] node12643;
	wire [4-1:0] node12644;
	wire [4-1:0] node12645;
	wire [4-1:0] node12646;
	wire [4-1:0] node12650;
	wire [4-1:0] node12651;
	wire [4-1:0] node12656;
	wire [4-1:0] node12657;
	wire [4-1:0] node12658;
	wire [4-1:0] node12659;
	wire [4-1:0] node12660;
	wire [4-1:0] node12661;
	wire [4-1:0] node12662;
	wire [4-1:0] node12663;
	wire [4-1:0] node12664;
	wire [4-1:0] node12665;
	wire [4-1:0] node12666;
	wire [4-1:0] node12667;
	wire [4-1:0] node12668;
	wire [4-1:0] node12670;
	wire [4-1:0] node12674;
	wire [4-1:0] node12676;
	wire [4-1:0] node12677;
	wire [4-1:0] node12680;
	wire [4-1:0] node12683;
	wire [4-1:0] node12684;
	wire [4-1:0] node12685;
	wire [4-1:0] node12689;
	wire [4-1:0] node12690;
	wire [4-1:0] node12694;
	wire [4-1:0] node12695;
	wire [4-1:0] node12696;
	wire [4-1:0] node12697;
	wire [4-1:0] node12699;
	wire [4-1:0] node12703;
	wire [4-1:0] node12706;
	wire [4-1:0] node12707;
	wire [4-1:0] node12708;
	wire [4-1:0] node12712;
	wire [4-1:0] node12715;
	wire [4-1:0] node12716;
	wire [4-1:0] node12717;
	wire [4-1:0] node12718;
	wire [4-1:0] node12720;
	wire [4-1:0] node12723;
	wire [4-1:0] node12724;
	wire [4-1:0] node12727;
	wire [4-1:0] node12730;
	wire [4-1:0] node12731;
	wire [4-1:0] node12732;
	wire [4-1:0] node12736;
	wire [4-1:0] node12738;
	wire [4-1:0] node12740;
	wire [4-1:0] node12743;
	wire [4-1:0] node12744;
	wire [4-1:0] node12745;
	wire [4-1:0] node12749;
	wire [4-1:0] node12751;
	wire [4-1:0] node12752;
	wire [4-1:0] node12753;
	wire [4-1:0] node12757;
	wire [4-1:0] node12760;
	wire [4-1:0] node12761;
	wire [4-1:0] node12762;
	wire [4-1:0] node12763;
	wire [4-1:0] node12764;
	wire [4-1:0] node12766;
	wire [4-1:0] node12769;
	wire [4-1:0] node12770;
	wire [4-1:0] node12774;
	wire [4-1:0] node12775;
	wire [4-1:0] node12778;
	wire [4-1:0] node12780;
	wire [4-1:0] node12782;
	wire [4-1:0] node12785;
	wire [4-1:0] node12786;
	wire [4-1:0] node12787;
	wire [4-1:0] node12788;
	wire [4-1:0] node12792;
	wire [4-1:0] node12793;
	wire [4-1:0] node12795;
	wire [4-1:0] node12799;
	wire [4-1:0] node12800;
	wire [4-1:0] node12803;
	wire [4-1:0] node12804;
	wire [4-1:0] node12805;
	wire [4-1:0] node12808;
	wire [4-1:0] node12812;
	wire [4-1:0] node12813;
	wire [4-1:0] node12814;
	wire [4-1:0] node12815;
	wire [4-1:0] node12816;
	wire [4-1:0] node12818;
	wire [4-1:0] node12822;
	wire [4-1:0] node12823;
	wire [4-1:0] node12827;
	wire [4-1:0] node12828;
	wire [4-1:0] node12829;
	wire [4-1:0] node12833;
	wire [4-1:0] node12834;
	wire [4-1:0] node12836;
	wire [4-1:0] node12840;
	wire [4-1:0] node12841;
	wire [4-1:0] node12842;
	wire [4-1:0] node12844;
	wire [4-1:0] node12848;
	wire [4-1:0] node12849;
	wire [4-1:0] node12851;
	wire [4-1:0] node12852;
	wire [4-1:0] node12856;
	wire [4-1:0] node12857;
	wire [4-1:0] node12858;
	wire [4-1:0] node12861;
	wire [4-1:0] node12865;
	wire [4-1:0] node12866;
	wire [4-1:0] node12867;
	wire [4-1:0] node12868;
	wire [4-1:0] node12869;
	wire [4-1:0] node12871;
	wire [4-1:0] node12873;
	wire [4-1:0] node12876;
	wire [4-1:0] node12877;
	wire [4-1:0] node12878;
	wire [4-1:0] node12879;
	wire [4-1:0] node12882;
	wire [4-1:0] node12885;
	wire [4-1:0] node12886;
	wire [4-1:0] node12890;
	wire [4-1:0] node12892;
	wire [4-1:0] node12895;
	wire [4-1:0] node12896;
	wire [4-1:0] node12897;
	wire [4-1:0] node12899;
	wire [4-1:0] node12900;
	wire [4-1:0] node12905;
	wire [4-1:0] node12906;
	wire [4-1:0] node12907;
	wire [4-1:0] node12908;
	wire [4-1:0] node12913;
	wire [4-1:0] node12915;
	wire [4-1:0] node12916;
	wire [4-1:0] node12920;
	wire [4-1:0] node12921;
	wire [4-1:0] node12922;
	wire [4-1:0] node12923;
	wire [4-1:0] node12926;
	wire [4-1:0] node12928;
	wire [4-1:0] node12929;
	wire [4-1:0] node12932;
	wire [4-1:0] node12935;
	wire [4-1:0] node12936;
	wire [4-1:0] node12937;
	wire [4-1:0] node12940;
	wire [4-1:0] node12943;
	wire [4-1:0] node12946;
	wire [4-1:0] node12947;
	wire [4-1:0] node12948;
	wire [4-1:0] node12950;
	wire [4-1:0] node12951;
	wire [4-1:0] node12956;
	wire [4-1:0] node12958;
	wire [4-1:0] node12960;
	wire [4-1:0] node12963;
	wire [4-1:0] node12964;
	wire [4-1:0] node12965;
	wire [4-1:0] node12966;
	wire [4-1:0] node12967;
	wire [4-1:0] node12969;
	wire [4-1:0] node12970;
	wire [4-1:0] node12974;
	wire [4-1:0] node12975;
	wire [4-1:0] node12977;
	wire [4-1:0] node12981;
	wire [4-1:0] node12982;
	wire [4-1:0] node12985;
	wire [4-1:0] node12987;
	wire [4-1:0] node12989;
	wire [4-1:0] node12992;
	wire [4-1:0] node12993;
	wire [4-1:0] node12994;
	wire [4-1:0] node12995;
	wire [4-1:0] node12998;
	wire [4-1:0] node12999;
	wire [4-1:0] node13002;
	wire [4-1:0] node13005;
	wire [4-1:0] node13007;
	wire [4-1:0] node13008;
	wire [4-1:0] node13011;
	wire [4-1:0] node13014;
	wire [4-1:0] node13015;
	wire [4-1:0] node13016;
	wire [4-1:0] node13017;
	wire [4-1:0] node13020;
	wire [4-1:0] node13023;
	wire [4-1:0] node13026;
	wire [4-1:0] node13028;
	wire [4-1:0] node13031;
	wire [4-1:0] node13032;
	wire [4-1:0] node13033;
	wire [4-1:0] node13034;
	wire [4-1:0] node13035;
	wire [4-1:0] node13037;
	wire [4-1:0] node13040;
	wire [4-1:0] node13042;
	wire [4-1:0] node13045;
	wire [4-1:0] node13046;
	wire [4-1:0] node13050;
	wire [4-1:0] node13052;
	wire [4-1:0] node13054;
	wire [4-1:0] node13057;
	wire [4-1:0] node13058;
	wire [4-1:0] node13059;
	wire [4-1:0] node13061;
	wire [4-1:0] node13064;
	wire [4-1:0] node13066;
	wire [4-1:0] node13067;
	wire [4-1:0] node13070;
	wire [4-1:0] node13073;
	wire [4-1:0] node13074;
	wire [4-1:0] node13076;
	wire [4-1:0] node13079;
	wire [4-1:0] node13080;
	wire [4-1:0] node13083;
	wire [4-1:0] node13084;
	wire [4-1:0] node13087;
	wire [4-1:0] node13090;
	wire [4-1:0] node13091;
	wire [4-1:0] node13092;
	wire [4-1:0] node13093;
	wire [4-1:0] node13094;
	wire [4-1:0] node13095;
	wire [4-1:0] node13096;
	wire [4-1:0] node13097;
	wire [4-1:0] node13101;
	wire [4-1:0] node13102;
	wire [4-1:0] node13106;
	wire [4-1:0] node13107;
	wire [4-1:0] node13111;
	wire [4-1:0] node13112;
	wire [4-1:0] node13113;
	wire [4-1:0] node13117;
	wire [4-1:0] node13118;
	wire [4-1:0] node13120;
	wire [4-1:0] node13123;
	wire [4-1:0] node13124;
	wire [4-1:0] node13126;
	wire [4-1:0] node13130;
	wire [4-1:0] node13131;
	wire [4-1:0] node13132;
	wire [4-1:0] node13133;
	wire [4-1:0] node13134;
	wire [4-1:0] node13135;
	wire [4-1:0] node13138;
	wire [4-1:0] node13141;
	wire [4-1:0] node13144;
	wire [4-1:0] node13146;
	wire [4-1:0] node13147;
	wire [4-1:0] node13151;
	wire [4-1:0] node13152;
	wire [4-1:0] node13153;
	wire [4-1:0] node13158;
	wire [4-1:0] node13159;
	wire [4-1:0] node13160;
	wire [4-1:0] node13161;
	wire [4-1:0] node13162;
	wire [4-1:0] node13165;
	wire [4-1:0] node13169;
	wire [4-1:0] node13172;
	wire [4-1:0] node13173;
	wire [4-1:0] node13176;
	wire [4-1:0] node13179;
	wire [4-1:0] node13180;
	wire [4-1:0] node13181;
	wire [4-1:0] node13182;
	wire [4-1:0] node13184;
	wire [4-1:0] node13185;
	wire [4-1:0] node13186;
	wire [4-1:0] node13190;
	wire [4-1:0] node13192;
	wire [4-1:0] node13195;
	wire [4-1:0] node13196;
	wire [4-1:0] node13199;
	wire [4-1:0] node13200;
	wire [4-1:0] node13201;
	wire [4-1:0] node13206;
	wire [4-1:0] node13207;
	wire [4-1:0] node13208;
	wire [4-1:0] node13211;
	wire [4-1:0] node13212;
	wire [4-1:0] node13213;
	wire [4-1:0] node13218;
	wire [4-1:0] node13219;
	wire [4-1:0] node13220;
	wire [4-1:0] node13223;
	wire [4-1:0] node13224;
	wire [4-1:0] node13228;
	wire [4-1:0] node13229;
	wire [4-1:0] node13233;
	wire [4-1:0] node13234;
	wire [4-1:0] node13235;
	wire [4-1:0] node13236;
	wire [4-1:0] node13237;
	wire [4-1:0] node13239;
	wire [4-1:0] node13243;
	wire [4-1:0] node13244;
	wire [4-1:0] node13245;
	wire [4-1:0] node13249;
	wire [4-1:0] node13251;
	wire [4-1:0] node13254;
	wire [4-1:0] node13255;
	wire [4-1:0] node13256;
	wire [4-1:0] node13257;
	wire [4-1:0] node13260;
	wire [4-1:0] node13264;
	wire [4-1:0] node13266;
	wire [4-1:0] node13268;
	wire [4-1:0] node13271;
	wire [4-1:0] node13272;
	wire [4-1:0] node13273;
	wire [4-1:0] node13275;
	wire [4-1:0] node13278;
	wire [4-1:0] node13281;
	wire [4-1:0] node13282;
	wire [4-1:0] node13284;
	wire [4-1:0] node13286;
	wire [4-1:0] node13289;
	wire [4-1:0] node13290;
	wire [4-1:0] node13291;
	wire [4-1:0] node13296;
	wire [4-1:0] node13297;
	wire [4-1:0] node13298;
	wire [4-1:0] node13299;
	wire [4-1:0] node13300;
	wire [4-1:0] node13301;
	wire [4-1:0] node13302;
	wire [4-1:0] node13305;
	wire [4-1:0] node13307;
	wire [4-1:0] node13310;
	wire [4-1:0] node13311;
	wire [4-1:0] node13313;
	wire [4-1:0] node13316;
	wire [4-1:0] node13319;
	wire [4-1:0] node13320;
	wire [4-1:0] node13322;
	wire [4-1:0] node13325;
	wire [4-1:0] node13326;
	wire [4-1:0] node13329;
	wire [4-1:0] node13332;
	wire [4-1:0] node13333;
	wire [4-1:0] node13335;
	wire [4-1:0] node13337;
	wire [4-1:0] node13340;
	wire [4-1:0] node13341;
	wire [4-1:0] node13343;
	wire [4-1:0] node13347;
	wire [4-1:0] node13348;
	wire [4-1:0] node13349;
	wire [4-1:0] node13350;
	wire [4-1:0] node13351;
	wire [4-1:0] node13355;
	wire [4-1:0] node13356;
	wire [4-1:0] node13360;
	wire [4-1:0] node13361;
	wire [4-1:0] node13362;
	wire [4-1:0] node13363;
	wire [4-1:0] node13368;
	wire [4-1:0] node13369;
	wire [4-1:0] node13370;
	wire [4-1:0] node13374;
	wire [4-1:0] node13377;
	wire [4-1:0] node13378;
	wire [4-1:0] node13379;
	wire [4-1:0] node13382;
	wire [4-1:0] node13384;
	wire [4-1:0] node13387;
	wire [4-1:0] node13388;
	wire [4-1:0] node13389;
	wire [4-1:0] node13391;
	wire [4-1:0] node13394;
	wire [4-1:0] node13397;
	wire [4-1:0] node13398;
	wire [4-1:0] node13401;
	wire [4-1:0] node13402;
	wire [4-1:0] node13406;
	wire [4-1:0] node13407;
	wire [4-1:0] node13408;
	wire [4-1:0] node13409;
	wire [4-1:0] node13410;
	wire [4-1:0] node13413;
	wire [4-1:0] node13414;
	wire [4-1:0] node13415;
	wire [4-1:0] node13419;
	wire [4-1:0] node13420;
	wire [4-1:0] node13424;
	wire [4-1:0] node13425;
	wire [4-1:0] node13426;
	wire [4-1:0] node13427;
	wire [4-1:0] node13430;
	wire [4-1:0] node13433;
	wire [4-1:0] node13436;
	wire [4-1:0] node13437;
	wire [4-1:0] node13438;
	wire [4-1:0] node13441;
	wire [4-1:0] node13444;
	wire [4-1:0] node13446;
	wire [4-1:0] node13449;
	wire [4-1:0] node13450;
	wire [4-1:0] node13451;
	wire [4-1:0] node13452;
	wire [4-1:0] node13455;
	wire [4-1:0] node13456;
	wire [4-1:0] node13460;
	wire [4-1:0] node13461;
	wire [4-1:0] node13464;
	wire [4-1:0] node13467;
	wire [4-1:0] node13468;
	wire [4-1:0] node13469;
	wire [4-1:0] node13471;
	wire [4-1:0] node13474;
	wire [4-1:0] node13476;
	wire [4-1:0] node13479;
	wire [4-1:0] node13480;
	wire [4-1:0] node13483;
	wire [4-1:0] node13484;
	wire [4-1:0] node13487;
	wire [4-1:0] node13490;
	wire [4-1:0] node13491;
	wire [4-1:0] node13492;
	wire [4-1:0] node13493;
	wire [4-1:0] node13494;
	wire [4-1:0] node13498;
	wire [4-1:0] node13501;
	wire [4-1:0] node13502;
	wire [4-1:0] node13503;
	wire [4-1:0] node13506;
	wire [4-1:0] node13509;
	wire [4-1:0] node13510;
	wire [4-1:0] node13512;
	wire [4-1:0] node13515;
	wire [4-1:0] node13516;
	wire [4-1:0] node13520;
	wire [4-1:0] node13521;
	wire [4-1:0] node13522;
	wire [4-1:0] node13523;
	wire [4-1:0] node13524;
	wire [4-1:0] node13527;
	wire [4-1:0] node13530;
	wire [4-1:0] node13532;
	wire [4-1:0] node13535;
	wire [4-1:0] node13536;
	wire [4-1:0] node13538;
	wire [4-1:0] node13541;
	wire [4-1:0] node13542;
	wire [4-1:0] node13546;
	wire [4-1:0] node13549;
	wire [4-1:0] node13550;
	wire [4-1:0] node13551;
	wire [4-1:0] node13552;
	wire [4-1:0] node13553;
	wire [4-1:0] node13554;
	wire [4-1:0] node13555;
	wire [4-1:0] node13556;
	wire [4-1:0] node13557;
	wire [4-1:0] node13559;
	wire [4-1:0] node13563;
	wire [4-1:0] node13564;
	wire [4-1:0] node13566;
	wire [4-1:0] node13570;
	wire [4-1:0] node13571;
	wire [4-1:0] node13573;
	wire [4-1:0] node13574;
	wire [4-1:0] node13578;
	wire [4-1:0] node13581;
	wire [4-1:0] node13582;
	wire [4-1:0] node13583;
	wire [4-1:0] node13585;
	wire [4-1:0] node13588;
	wire [4-1:0] node13589;
	wire [4-1:0] node13591;
	wire [4-1:0] node13595;
	wire [4-1:0] node13596;
	wire [4-1:0] node13597;
	wire [4-1:0] node13602;
	wire [4-1:0] node13603;
	wire [4-1:0] node13604;
	wire [4-1:0] node13605;
	wire [4-1:0] node13606;
	wire [4-1:0] node13609;
	wire [4-1:0] node13613;
	wire [4-1:0] node13614;
	wire [4-1:0] node13615;
	wire [4-1:0] node13616;
	wire [4-1:0] node13620;
	wire [4-1:0] node13621;
	wire [4-1:0] node13625;
	wire [4-1:0] node13626;
	wire [4-1:0] node13627;
	wire [4-1:0] node13632;
	wire [4-1:0] node13633;
	wire [4-1:0] node13634;
	wire [4-1:0] node13636;
	wire [4-1:0] node13637;
	wire [4-1:0] node13641;
	wire [4-1:0] node13643;
	wire [4-1:0] node13645;
	wire [4-1:0] node13648;
	wire [4-1:0] node13649;
	wire [4-1:0] node13650;
	wire [4-1:0] node13653;
	wire [4-1:0] node13656;
	wire [4-1:0] node13657;
	wire [4-1:0] node13661;
	wire [4-1:0] node13662;
	wire [4-1:0] node13663;
	wire [4-1:0] node13664;
	wire [4-1:0] node13665;
	wire [4-1:0] node13666;
	wire [4-1:0] node13669;
	wire [4-1:0] node13673;
	wire [4-1:0] node13674;
	wire [4-1:0] node13677;
	wire [4-1:0] node13678;
	wire [4-1:0] node13682;
	wire [4-1:0] node13683;
	wire [4-1:0] node13684;
	wire [4-1:0] node13685;
	wire [4-1:0] node13690;
	wire [4-1:0] node13691;
	wire [4-1:0] node13692;
	wire [4-1:0] node13696;
	wire [4-1:0] node13698;
	wire [4-1:0] node13701;
	wire [4-1:0] node13702;
	wire [4-1:0] node13703;
	wire [4-1:0] node13704;
	wire [4-1:0] node13706;
	wire [4-1:0] node13708;
	wire [4-1:0] node13711;
	wire [4-1:0] node13712;
	wire [4-1:0] node13715;
	wire [4-1:0] node13716;
	wire [4-1:0] node13720;
	wire [4-1:0] node13721;
	wire [4-1:0] node13722;
	wire [4-1:0] node13724;
	wire [4-1:0] node13727;
	wire [4-1:0] node13730;
	wire [4-1:0] node13731;
	wire [4-1:0] node13735;
	wire [4-1:0] node13736;
	wire [4-1:0] node13738;
	wire [4-1:0] node13740;
	wire [4-1:0] node13743;
	wire [4-1:0] node13744;
	wire [4-1:0] node13745;
	wire [4-1:0] node13746;
	wire [4-1:0] node13750;
	wire [4-1:0] node13751;
	wire [4-1:0] node13755;
	wire [4-1:0] node13757;
	wire [4-1:0] node13760;
	wire [4-1:0] node13761;
	wire [4-1:0] node13762;
	wire [4-1:0] node13763;
	wire [4-1:0] node13764;
	wire [4-1:0] node13765;
	wire [4-1:0] node13766;
	wire [4-1:0] node13768;
	wire [4-1:0] node13771;
	wire [4-1:0] node13772;
	wire [4-1:0] node13775;
	wire [4-1:0] node13778;
	wire [4-1:0] node13780;
	wire [4-1:0] node13783;
	wire [4-1:0] node13784;
	wire [4-1:0] node13785;
	wire [4-1:0] node13787;
	wire [4-1:0] node13790;
	wire [4-1:0] node13791;
	wire [4-1:0] node13795;
	wire [4-1:0] node13797;
	wire [4-1:0] node13799;
	wire [4-1:0] node13802;
	wire [4-1:0] node13803;
	wire [4-1:0] node13804;
	wire [4-1:0] node13805;
	wire [4-1:0] node13806;
	wire [4-1:0] node13810;
	wire [4-1:0] node13814;
	wire [4-1:0] node13815;
	wire [4-1:0] node13817;
	wire [4-1:0] node13818;
	wire [4-1:0] node13822;
	wire [4-1:0] node13824;
	wire [4-1:0] node13827;
	wire [4-1:0] node13828;
	wire [4-1:0] node13829;
	wire [4-1:0] node13830;
	wire [4-1:0] node13831;
	wire [4-1:0] node13835;
	wire [4-1:0] node13837;
	wire [4-1:0] node13840;
	wire [4-1:0] node13841;
	wire [4-1:0] node13844;
	wire [4-1:0] node13845;
	wire [4-1:0] node13848;
	wire [4-1:0] node13851;
	wire [4-1:0] node13852;
	wire [4-1:0] node13853;
	wire [4-1:0] node13854;
	wire [4-1:0] node13857;
	wire [4-1:0] node13858;
	wire [4-1:0] node13862;
	wire [4-1:0] node13863;
	wire [4-1:0] node13864;
	wire [4-1:0] node13868;
	wire [4-1:0] node13869;
	wire [4-1:0] node13872;
	wire [4-1:0] node13875;
	wire [4-1:0] node13876;
	wire [4-1:0] node13878;
	wire [4-1:0] node13881;
	wire [4-1:0] node13882;
	wire [4-1:0] node13883;
	wire [4-1:0] node13886;
	wire [4-1:0] node13889;
	wire [4-1:0] node13891;
	wire [4-1:0] node13894;
	wire [4-1:0] node13895;
	wire [4-1:0] node13896;
	wire [4-1:0] node13897;
	wire [4-1:0] node13899;
	wire [4-1:0] node13900;
	wire [4-1:0] node13901;
	wire [4-1:0] node13904;
	wire [4-1:0] node13907;
	wire [4-1:0] node13908;
	wire [4-1:0] node13912;
	wire [4-1:0] node13913;
	wire [4-1:0] node13915;
	wire [4-1:0] node13918;
	wire [4-1:0] node13920;
	wire [4-1:0] node13923;
	wire [4-1:0] node13924;
	wire [4-1:0] node13925;
	wire [4-1:0] node13926;
	wire [4-1:0] node13927;
	wire [4-1:0] node13931;
	wire [4-1:0] node13934;
	wire [4-1:0] node13936;
	wire [4-1:0] node13939;
	wire [4-1:0] node13940;
	wire [4-1:0] node13942;
	wire [4-1:0] node13945;
	wire [4-1:0] node13946;
	wire [4-1:0] node13949;
	wire [4-1:0] node13950;
	wire [4-1:0] node13954;
	wire [4-1:0] node13955;
	wire [4-1:0] node13956;
	wire [4-1:0] node13957;
	wire [4-1:0] node13958;
	wire [4-1:0] node13959;
	wire [4-1:0] node13964;
	wire [4-1:0] node13965;
	wire [4-1:0] node13966;
	wire [4-1:0] node13970;
	wire [4-1:0] node13971;
	wire [4-1:0] node13975;
	wire [4-1:0] node13976;
	wire [4-1:0] node13978;
	wire [4-1:0] node13981;
	wire [4-1:0] node13983;
	wire [4-1:0] node13985;
	wire [4-1:0] node13988;
	wire [4-1:0] node13989;
	wire [4-1:0] node13991;
	wire [4-1:0] node13992;
	wire [4-1:0] node13993;
	wire [4-1:0] node13996;
	wire [4-1:0] node14000;
	wire [4-1:0] node14001;
	wire [4-1:0] node14003;
	wire [4-1:0] node14004;
	wire [4-1:0] node14009;
	wire [4-1:0] node14010;
	wire [4-1:0] node14011;
	wire [4-1:0] node14012;
	wire [4-1:0] node14013;
	wire [4-1:0] node14014;
	wire [4-1:0] node14015;
	wire [4-1:0] node14016;
	wire [4-1:0] node14017;
	wire [4-1:0] node14021;
	wire [4-1:0] node14023;
	wire [4-1:0] node14026;
	wire [4-1:0] node14027;
	wire [4-1:0] node14029;
	wire [4-1:0] node14032;
	wire [4-1:0] node14033;
	wire [4-1:0] node14036;
	wire [4-1:0] node14039;
	wire [4-1:0] node14040;
	wire [4-1:0] node14041;
	wire [4-1:0] node14042;
	wire [4-1:0] node14046;
	wire [4-1:0] node14049;
	wire [4-1:0] node14050;
	wire [4-1:0] node14054;
	wire [4-1:0] node14055;
	wire [4-1:0] node14056;
	wire [4-1:0] node14057;
	wire [4-1:0] node14060;
	wire [4-1:0] node14062;
	wire [4-1:0] node14065;
	wire [4-1:0] node14067;
	wire [4-1:0] node14068;
	wire [4-1:0] node14071;
	wire [4-1:0] node14074;
	wire [4-1:0] node14075;
	wire [4-1:0] node14076;
	wire [4-1:0] node14077;
	wire [4-1:0] node14080;
	wire [4-1:0] node14084;
	wire [4-1:0] node14085;
	wire [4-1:0] node14088;
	wire [4-1:0] node14091;
	wire [4-1:0] node14092;
	wire [4-1:0] node14093;
	wire [4-1:0] node14094;
	wire [4-1:0] node14096;
	wire [4-1:0] node14100;
	wire [4-1:0] node14101;
	wire [4-1:0] node14102;
	wire [4-1:0] node14105;
	wire [4-1:0] node14106;
	wire [4-1:0] node14110;
	wire [4-1:0] node14113;
	wire [4-1:0] node14114;
	wire [4-1:0] node14115;
	wire [4-1:0] node14116;
	wire [4-1:0] node14118;
	wire [4-1:0] node14122;
	wire [4-1:0] node14123;
	wire [4-1:0] node14126;
	wire [4-1:0] node14129;
	wire [4-1:0] node14130;
	wire [4-1:0] node14131;
	wire [4-1:0] node14132;
	wire [4-1:0] node14137;
	wire [4-1:0] node14138;
	wire [4-1:0] node14139;
	wire [4-1:0] node14143;
	wire [4-1:0] node14145;
	wire [4-1:0] node14148;
	wire [4-1:0] node14149;
	wire [4-1:0] node14150;
	wire [4-1:0] node14151;
	wire [4-1:0] node14152;
	wire [4-1:0] node14153;
	wire [4-1:0] node14157;
	wire [4-1:0] node14159;
	wire [4-1:0] node14163;
	wire [4-1:0] node14164;
	wire [4-1:0] node14165;
	wire [4-1:0] node14166;
	wire [4-1:0] node14171;
	wire [4-1:0] node14172;
	wire [4-1:0] node14174;
	wire [4-1:0] node14177;
	wire [4-1:0] node14179;
	wire [4-1:0] node14182;
	wire [4-1:0] node14183;
	wire [4-1:0] node14184;
	wire [4-1:0] node14185;
	wire [4-1:0] node14188;
	wire [4-1:0] node14191;
	wire [4-1:0] node14192;
	wire [4-1:0] node14193;
	wire [4-1:0] node14198;
	wire [4-1:0] node14199;
	wire [4-1:0] node14200;
	wire [4-1:0] node14202;
	wire [4-1:0] node14205;
	wire [4-1:0] node14207;
	wire [4-1:0] node14210;
	wire [4-1:0] node14211;
	wire [4-1:0] node14212;
	wire [4-1:0] node14216;
	wire [4-1:0] node14218;
	wire [4-1:0] node14221;
	wire [4-1:0] node14222;
	wire [4-1:0] node14223;
	wire [4-1:0] node14224;
	wire [4-1:0] node14225;
	wire [4-1:0] node14226;
	wire [4-1:0] node14228;
	wire [4-1:0] node14230;
	wire [4-1:0] node14233;
	wire [4-1:0] node14234;
	wire [4-1:0] node14237;
	wire [4-1:0] node14238;
	wire [4-1:0] node14242;
	wire [4-1:0] node14243;
	wire [4-1:0] node14244;
	wire [4-1:0] node14245;
	wire [4-1:0] node14249;
	wire [4-1:0] node14252;
	wire [4-1:0] node14253;
	wire [4-1:0] node14254;
	wire [4-1:0] node14258;
	wire [4-1:0] node14260;
	wire [4-1:0] node14263;
	wire [4-1:0] node14264;
	wire [4-1:0] node14266;
	wire [4-1:0] node14267;
	wire [4-1:0] node14271;
	wire [4-1:0] node14272;
	wire [4-1:0] node14273;
	wire [4-1:0] node14276;
	wire [4-1:0] node14280;
	wire [4-1:0] node14281;
	wire [4-1:0] node14282;
	wire [4-1:0] node14284;
	wire [4-1:0] node14285;
	wire [4-1:0] node14288;
	wire [4-1:0] node14291;
	wire [4-1:0] node14292;
	wire [4-1:0] node14294;
	wire [4-1:0] node14297;
	wire [4-1:0] node14298;
	wire [4-1:0] node14300;
	wire [4-1:0] node14303;
	wire [4-1:0] node14305;
	wire [4-1:0] node14308;
	wire [4-1:0] node14309;
	wire [4-1:0] node14310;
	wire [4-1:0] node14311;
	wire [4-1:0] node14312;
	wire [4-1:0] node14316;
	wire [4-1:0] node14319;
	wire [4-1:0] node14320;
	wire [4-1:0] node14321;
	wire [4-1:0] node14324;
	wire [4-1:0] node14327;
	wire [4-1:0] node14328;
	wire [4-1:0] node14331;
	wire [4-1:0] node14334;
	wire [4-1:0] node14335;
	wire [4-1:0] node14339;
	wire [4-1:0] node14340;
	wire [4-1:0] node14341;
	wire [4-1:0] node14342;
	wire [4-1:0] node14343;
	wire [4-1:0] node14345;
	wire [4-1:0] node14348;
	wire [4-1:0] node14349;
	wire [4-1:0] node14350;
	wire [4-1:0] node14353;
	wire [4-1:0] node14356;
	wire [4-1:0] node14357;
	wire [4-1:0] node14361;
	wire [4-1:0] node14362;
	wire [4-1:0] node14364;
	wire [4-1:0] node14366;
	wire [4-1:0] node14369;
	wire [4-1:0] node14370;
	wire [4-1:0] node14372;
	wire [4-1:0] node14375;
	wire [4-1:0] node14376;
	wire [4-1:0] node14380;
	wire [4-1:0] node14381;
	wire [4-1:0] node14382;
	wire [4-1:0] node14384;
	wire [4-1:0] node14387;
	wire [4-1:0] node14388;
	wire [4-1:0] node14392;
	wire [4-1:0] node14393;
	wire [4-1:0] node14394;
	wire [4-1:0] node14398;
	wire [4-1:0] node14399;
	wire [4-1:0] node14400;
	wire [4-1:0] node14405;
	wire [4-1:0] node14406;
	wire [4-1:0] node14407;
	wire [4-1:0] node14408;
	wire [4-1:0] node14409;
	wire [4-1:0] node14412;
	wire [4-1:0] node14415;
	wire [4-1:0] node14416;
	wire [4-1:0] node14420;
	wire [4-1:0] node14421;
	wire [4-1:0] node14422;
	wire [4-1:0] node14423;
	wire [4-1:0] node14426;
	wire [4-1:0] node14429;
	wire [4-1:0] node14430;
	wire [4-1:0] node14433;
	wire [4-1:0] node14436;
	wire [4-1:0] node14437;
	wire [4-1:0] node14439;
	wire [4-1:0] node14443;
	wire [4-1:0] node14444;
	wire [4-1:0] node14446;
	wire [4-1:0] node14448;
	wire [4-1:0] node14450;
	wire [4-1:0] node14453;
	wire [4-1:0] node14454;
	wire [4-1:0] node14455;
	wire [4-1:0] node14456;
	wire [4-1:0] node14461;
	wire [4-1:0] node14462;
	wire [4-1:0] node14464;
	wire [4-1:0] node14467;
	wire [4-1:0] node14469;
	wire [4-1:0] node14472;
	wire [4-1:0] node14473;
	wire [4-1:0] node14474;
	wire [4-1:0] node14475;
	wire [4-1:0] node14476;
	wire [4-1:0] node14477;
	wire [4-1:0] node14478;
	wire [4-1:0] node14479;
	wire [4-1:0] node14480;
	wire [4-1:0] node14484;
	wire [4-1:0] node14485;
	wire [4-1:0] node14488;
	wire [4-1:0] node14490;
	wire [4-1:0] node14493;
	wire [4-1:0] node14494;
	wire [4-1:0] node14495;
	wire [4-1:0] node14497;
	wire [4-1:0] node14499;
	wire [4-1:0] node14502;
	wire [4-1:0] node14504;
	wire [4-1:0] node14506;
	wire [4-1:0] node14509;
	wire [4-1:0] node14510;
	wire [4-1:0] node14511;
	wire [4-1:0] node14512;
	wire [4-1:0] node14515;
	wire [4-1:0] node14519;
	wire [4-1:0] node14520;
	wire [4-1:0] node14521;
	wire [4-1:0] node14525;
	wire [4-1:0] node14527;
	wire [4-1:0] node14530;
	wire [4-1:0] node14531;
	wire [4-1:0] node14532;
	wire [4-1:0] node14533;
	wire [4-1:0] node14536;
	wire [4-1:0] node14537;
	wire [4-1:0] node14539;
	wire [4-1:0] node14542;
	wire [4-1:0] node14544;
	wire [4-1:0] node14547;
	wire [4-1:0] node14548;
	wire [4-1:0] node14549;
	wire [4-1:0] node14552;
	wire [4-1:0] node14555;
	wire [4-1:0] node14558;
	wire [4-1:0] node14559;
	wire [4-1:0] node14560;
	wire [4-1:0] node14561;
	wire [4-1:0] node14565;
	wire [4-1:0] node14567;
	wire [4-1:0] node14568;
	wire [4-1:0] node14572;
	wire [4-1:0] node14573;
	wire [4-1:0] node14574;
	wire [4-1:0] node14576;
	wire [4-1:0] node14579;
	wire [4-1:0] node14581;
	wire [4-1:0] node14584;
	wire [4-1:0] node14585;
	wire [4-1:0] node14589;
	wire [4-1:0] node14590;
	wire [4-1:0] node14591;
	wire [4-1:0] node14592;
	wire [4-1:0] node14593;
	wire [4-1:0] node14595;
	wire [4-1:0] node14598;
	wire [4-1:0] node14599;
	wire [4-1:0] node14601;
	wire [4-1:0] node14604;
	wire [4-1:0] node14606;
	wire [4-1:0] node14609;
	wire [4-1:0] node14610;
	wire [4-1:0] node14612;
	wire [4-1:0] node14613;
	wire [4-1:0] node14617;
	wire [4-1:0] node14618;
	wire [4-1:0] node14621;
	wire [4-1:0] node14624;
	wire [4-1:0] node14625;
	wire [4-1:0] node14626;
	wire [4-1:0] node14627;
	wire [4-1:0] node14630;
	wire [4-1:0] node14631;
	wire [4-1:0] node14634;
	wire [4-1:0] node14637;
	wire [4-1:0] node14638;
	wire [4-1:0] node14641;
	wire [4-1:0] node14644;
	wire [4-1:0] node14645;
	wire [4-1:0] node14646;
	wire [4-1:0] node14647;
	wire [4-1:0] node14650;
	wire [4-1:0] node14653;
	wire [4-1:0] node14655;
	wire [4-1:0] node14658;
	wire [4-1:0] node14659;
	wire [4-1:0] node14660;
	wire [4-1:0] node14663;
	wire [4-1:0] node14667;
	wire [4-1:0] node14668;
	wire [4-1:0] node14669;
	wire [4-1:0] node14670;
	wire [4-1:0] node14671;
	wire [4-1:0] node14672;
	wire [4-1:0] node14675;
	wire [4-1:0] node14678;
	wire [4-1:0] node14681;
	wire [4-1:0] node14682;
	wire [4-1:0] node14684;
	wire [4-1:0] node14688;
	wire [4-1:0] node14689;
	wire [4-1:0] node14690;
	wire [4-1:0] node14692;
	wire [4-1:0] node14695;
	wire [4-1:0] node14696;
	wire [4-1:0] node14700;
	wire [4-1:0] node14701;
	wire [4-1:0] node14705;
	wire [4-1:0] node14706;
	wire [4-1:0] node14708;
	wire [4-1:0] node14709;
	wire [4-1:0] node14712;
	wire [4-1:0] node14715;
	wire [4-1:0] node14716;
	wire [4-1:0] node14717;
	wire [4-1:0] node14721;
	wire [4-1:0] node14723;
	wire [4-1:0] node14726;
	wire [4-1:0] node14727;
	wire [4-1:0] node14728;
	wire [4-1:0] node14729;
	wire [4-1:0] node14730;
	wire [4-1:0] node14732;
	wire [4-1:0] node14733;
	wire [4-1:0] node14736;
	wire [4-1:0] node14739;
	wire [4-1:0] node14740;
	wire [4-1:0] node14741;
	wire [4-1:0] node14744;
	wire [4-1:0] node14746;
	wire [4-1:0] node14749;
	wire [4-1:0] node14752;
	wire [4-1:0] node14753;
	wire [4-1:0] node14754;
	wire [4-1:0] node14757;
	wire [4-1:0] node14758;
	wire [4-1:0] node14759;
	wire [4-1:0] node14764;
	wire [4-1:0] node14765;
	wire [4-1:0] node14766;
	wire [4-1:0] node14768;
	wire [4-1:0] node14772;
	wire [4-1:0] node14775;
	wire [4-1:0] node14776;
	wire [4-1:0] node14777;
	wire [4-1:0] node14778;
	wire [4-1:0] node14780;
	wire [4-1:0] node14783;
	wire [4-1:0] node14784;
	wire [4-1:0] node14785;
	wire [4-1:0] node14789;
	wire [4-1:0] node14790;
	wire [4-1:0] node14794;
	wire [4-1:0] node14795;
	wire [4-1:0] node14796;
	wire [4-1:0] node14799;
	wire [4-1:0] node14802;
	wire [4-1:0] node14803;
	wire [4-1:0] node14805;
	wire [4-1:0] node14808;
	wire [4-1:0] node14810;
	wire [4-1:0] node14813;
	wire [4-1:0] node14814;
	wire [4-1:0] node14815;
	wire [4-1:0] node14817;
	wire [4-1:0] node14818;
	wire [4-1:0] node14821;
	wire [4-1:0] node14824;
	wire [4-1:0] node14825;
	wire [4-1:0] node14829;
	wire [4-1:0] node14830;
	wire [4-1:0] node14832;
	wire [4-1:0] node14833;
	wire [4-1:0] node14836;
	wire [4-1:0] node14839;
	wire [4-1:0] node14840;
	wire [4-1:0] node14841;
	wire [4-1:0] node14844;
	wire [4-1:0] node14848;
	wire [4-1:0] node14849;
	wire [4-1:0] node14850;
	wire [4-1:0] node14851;
	wire [4-1:0] node14852;
	wire [4-1:0] node14854;
	wire [4-1:0] node14857;
	wire [4-1:0] node14858;
	wire [4-1:0] node14860;
	wire [4-1:0] node14864;
	wire [4-1:0] node14865;
	wire [4-1:0] node14868;
	wire [4-1:0] node14869;
	wire [4-1:0] node14872;
	wire [4-1:0] node14875;
	wire [4-1:0] node14876;
	wire [4-1:0] node14877;
	wire [4-1:0] node14878;
	wire [4-1:0] node14882;
	wire [4-1:0] node14883;
	wire [4-1:0] node14886;
	wire [4-1:0] node14887;
	wire [4-1:0] node14890;
	wire [4-1:0] node14893;
	wire [4-1:0] node14894;
	wire [4-1:0] node14896;
	wire [4-1:0] node14898;
	wire [4-1:0] node14901;
	wire [4-1:0] node14903;
	wire [4-1:0] node14904;
	wire [4-1:0] node14907;
	wire [4-1:0] node14910;
	wire [4-1:0] node14911;
	wire [4-1:0] node14912;
	wire [4-1:0] node14913;
	wire [4-1:0] node14914;
	wire [4-1:0] node14916;
	wire [4-1:0] node14919;
	wire [4-1:0] node14920;
	wire [4-1:0] node14924;
	wire [4-1:0] node14926;
	wire [4-1:0] node14929;
	wire [4-1:0] node14930;
	wire [4-1:0] node14933;
	wire [4-1:0] node14934;
	wire [4-1:0] node14935;
	wire [4-1:0] node14940;
	wire [4-1:0] node14941;
	wire [4-1:0] node14943;
	wire [4-1:0] node14944;
	wire [4-1:0] node14947;
	wire [4-1:0] node14948;
	wire [4-1:0] node14952;
	wire [4-1:0] node14953;
	wire [4-1:0] node14954;
	wire [4-1:0] node14955;
	wire [4-1:0] node14960;
	wire [4-1:0] node14961;
	wire [4-1:0] node14963;
	wire [4-1:0] node14966;
	wire [4-1:0] node14969;
	wire [4-1:0] node14970;
	wire [4-1:0] node14971;
	wire [4-1:0] node14972;
	wire [4-1:0] node14973;
	wire [4-1:0] node14974;
	wire [4-1:0] node14975;
	wire [4-1:0] node14977;
	wire [4-1:0] node14980;
	wire [4-1:0] node14981;
	wire [4-1:0] node14983;
	wire [4-1:0] node14987;
	wire [4-1:0] node14989;
	wire [4-1:0] node14992;
	wire [4-1:0] node14993;
	wire [4-1:0] node14994;
	wire [4-1:0] node14995;
	wire [4-1:0] node14997;
	wire [4-1:0] node15000;
	wire [4-1:0] node15003;
	wire [4-1:0] node15004;
	wire [4-1:0] node15005;
	wire [4-1:0] node15010;
	wire [4-1:0] node15011;
	wire [4-1:0] node15013;
	wire [4-1:0] node15016;
	wire [4-1:0] node15017;
	wire [4-1:0] node15018;
	wire [4-1:0] node15023;
	wire [4-1:0] node15024;
	wire [4-1:0] node15025;
	wire [4-1:0] node15026;
	wire [4-1:0] node15027;
	wire [4-1:0] node15029;
	wire [4-1:0] node15032;
	wire [4-1:0] node15035;
	wire [4-1:0] node15036;
	wire [4-1:0] node15037;
	wire [4-1:0] node15042;
	wire [4-1:0] node15043;
	wire [4-1:0] node15045;
	wire [4-1:0] node15047;
	wire [4-1:0] node15051;
	wire [4-1:0] node15052;
	wire [4-1:0] node15053;
	wire [4-1:0] node15054;
	wire [4-1:0] node15057;
	wire [4-1:0] node15058;
	wire [4-1:0] node15062;
	wire [4-1:0] node15063;
	wire [4-1:0] node15066;
	wire [4-1:0] node15068;
	wire [4-1:0] node15071;
	wire [4-1:0] node15072;
	wire [4-1:0] node15074;
	wire [4-1:0] node15076;
	wire [4-1:0] node15079;
	wire [4-1:0] node15081;
	wire [4-1:0] node15084;
	wire [4-1:0] node15085;
	wire [4-1:0] node15086;
	wire [4-1:0] node15087;
	wire [4-1:0] node15088;
	wire [4-1:0] node15089;
	wire [4-1:0] node15093;
	wire [4-1:0] node15095;
	wire [4-1:0] node15096;
	wire [4-1:0] node15100;
	wire [4-1:0] node15101;
	wire [4-1:0] node15103;
	wire [4-1:0] node15104;
	wire [4-1:0] node15108;
	wire [4-1:0] node15109;
	wire [4-1:0] node15113;
	wire [4-1:0] node15114;
	wire [4-1:0] node15115;
	wire [4-1:0] node15117;
	wire [4-1:0] node15118;
	wire [4-1:0] node15122;
	wire [4-1:0] node15125;
	wire [4-1:0] node15126;
	wire [4-1:0] node15127;
	wire [4-1:0] node15130;
	wire [4-1:0] node15133;
	wire [4-1:0] node15134;
	wire [4-1:0] node15135;
	wire [4-1:0] node15139;
	wire [4-1:0] node15140;
	wire [4-1:0] node15144;
	wire [4-1:0] node15145;
	wire [4-1:0] node15146;
	wire [4-1:0] node15147;
	wire [4-1:0] node15148;
	wire [4-1:0] node15152;
	wire [4-1:0] node15154;
	wire [4-1:0] node15157;
	wire [4-1:0] node15158;
	wire [4-1:0] node15160;
	wire [4-1:0] node15164;
	wire [4-1:0] node15165;
	wire [4-1:0] node15166;
	wire [4-1:0] node15167;
	wire [4-1:0] node15171;
	wire [4-1:0] node15174;
	wire [4-1:0] node15175;
	wire [4-1:0] node15176;
	wire [4-1:0] node15177;
	wire [4-1:0] node15181;
	wire [4-1:0] node15184;
	wire [4-1:0] node15186;
	wire [4-1:0] node15189;
	wire [4-1:0] node15190;
	wire [4-1:0] node15191;
	wire [4-1:0] node15192;
	wire [4-1:0] node15193;
	wire [4-1:0] node15194;
	wire [4-1:0] node15195;
	wire [4-1:0] node15196;
	wire [4-1:0] node15199;
	wire [4-1:0] node15202;
	wire [4-1:0] node15203;
	wire [4-1:0] node15207;
	wire [4-1:0] node15209;
	wire [4-1:0] node15210;
	wire [4-1:0] node15214;
	wire [4-1:0] node15215;
	wire [4-1:0] node15217;
	wire [4-1:0] node15220;
	wire [4-1:0] node15223;
	wire [4-1:0] node15224;
	wire [4-1:0] node15225;
	wire [4-1:0] node15226;
	wire [4-1:0] node15228;
	wire [4-1:0] node15231;
	wire [4-1:0] node15234;
	wire [4-1:0] node15235;
	wire [4-1:0] node15237;
	wire [4-1:0] node15240;
	wire [4-1:0] node15241;
	wire [4-1:0] node15244;
	wire [4-1:0] node15247;
	wire [4-1:0] node15248;
	wire [4-1:0] node15250;
	wire [4-1:0] node15254;
	wire [4-1:0] node15255;
	wire [4-1:0] node15256;
	wire [4-1:0] node15257;
	wire [4-1:0] node15258;
	wire [4-1:0] node15259;
	wire [4-1:0] node15262;
	wire [4-1:0] node15265;
	wire [4-1:0] node15267;
	wire [4-1:0] node15270;
	wire [4-1:0] node15273;
	wire [4-1:0] node15275;
	wire [4-1:0] node15276;
	wire [4-1:0] node15277;
	wire [4-1:0] node15280;
	wire [4-1:0] node15283;
	wire [4-1:0] node15286;
	wire [4-1:0] node15287;
	wire [4-1:0] node15288;
	wire [4-1:0] node15290;
	wire [4-1:0] node15293;
	wire [4-1:0] node15295;
	wire [4-1:0] node15298;
	wire [4-1:0] node15299;
	wire [4-1:0] node15300;
	wire [4-1:0] node15301;
	wire [4-1:0] node15306;
	wire [4-1:0] node15307;
	wire [4-1:0] node15310;
	wire [4-1:0] node15311;
	wire [4-1:0] node15315;
	wire [4-1:0] node15316;
	wire [4-1:0] node15317;
	wire [4-1:0] node15318;
	wire [4-1:0] node15319;
	wire [4-1:0] node15321;
	wire [4-1:0] node15324;
	wire [4-1:0] node15326;
	wire [4-1:0] node15328;
	wire [4-1:0] node15331;
	wire [4-1:0] node15332;
	wire [4-1:0] node15333;
	wire [4-1:0] node15336;
	wire [4-1:0] node15337;
	wire [4-1:0] node15341;
	wire [4-1:0] node15342;
	wire [4-1:0] node15345;
	wire [4-1:0] node15346;
	wire [4-1:0] node15349;
	wire [4-1:0] node15352;
	wire [4-1:0] node15353;
	wire [4-1:0] node15354;
	wire [4-1:0] node15356;
	wire [4-1:0] node15358;
	wire [4-1:0] node15361;
	wire [4-1:0] node15363;
	wire [4-1:0] node15364;
	wire [4-1:0] node15368;
	wire [4-1:0] node15370;
	wire [4-1:0] node15373;
	wire [4-1:0] node15374;
	wire [4-1:0] node15375;
	wire [4-1:0] node15376;
	wire [4-1:0] node15377;
	wire [4-1:0] node15379;
	wire [4-1:0] node15382;
	wire [4-1:0] node15385;
	wire [4-1:0] node15388;
	wire [4-1:0] node15389;
	wire [4-1:0] node15391;
	wire [4-1:0] node15394;
	wire [4-1:0] node15395;
	wire [4-1:0] node15398;
	wire [4-1:0] node15401;
	wire [4-1:0] node15402;
	wire [4-1:0] node15403;
	wire [4-1:0] node15404;
	wire [4-1:0] node15407;
	wire [4-1:0] node15409;
	wire [4-1:0] node15412;
	wire [4-1:0] node15415;
	wire [4-1:0] node15416;
	wire [4-1:0] node15420;
	wire [4-1:0] node15421;
	wire [4-1:0] node15422;
	wire [4-1:0] node15423;
	wire [4-1:0] node15424;
	wire [4-1:0] node15425;
	wire [4-1:0] node15426;
	wire [4-1:0] node15429;
	wire [4-1:0] node15430;
	wire [4-1:0] node15431;
	wire [4-1:0] node15433;
	wire [4-1:0] node15437;
	wire [4-1:0] node15438;
	wire [4-1:0] node15440;
	wire [4-1:0] node15443;
	wire [4-1:0] node15446;
	wire [4-1:0] node15447;
	wire [4-1:0] node15448;
	wire [4-1:0] node15449;
	wire [4-1:0] node15452;
	wire [4-1:0] node15453;
	wire [4-1:0] node15456;
	wire [4-1:0] node15459;
	wire [4-1:0] node15460;
	wire [4-1:0] node15461;
	wire [4-1:0] node15465;
	wire [4-1:0] node15468;
	wire [4-1:0] node15469;
	wire [4-1:0] node15470;
	wire [4-1:0] node15472;
	wire [4-1:0] node15475;
	wire [4-1:0] node15478;
	wire [4-1:0] node15479;
	wire [4-1:0] node15482;
	wire [4-1:0] node15483;
	wire [4-1:0] node15486;
	wire [4-1:0] node15489;
	wire [4-1:0] node15490;
	wire [4-1:0] node15491;
	wire [4-1:0] node15492;
	wire [4-1:0] node15493;
	wire [4-1:0] node15494;
	wire [4-1:0] node15498;
	wire [4-1:0] node15500;
	wire [4-1:0] node15503;
	wire [4-1:0] node15504;
	wire [4-1:0] node15507;
	wire [4-1:0] node15510;
	wire [4-1:0] node15511;
	wire [4-1:0] node15512;
	wire [4-1:0] node15516;
	wire [4-1:0] node15517;
	wire [4-1:0] node15518;
	wire [4-1:0] node15523;
	wire [4-1:0] node15524;
	wire [4-1:0] node15525;
	wire [4-1:0] node15527;
	wire [4-1:0] node15530;
	wire [4-1:0] node15531;
	wire [4-1:0] node15533;
	wire [4-1:0] node15536;
	wire [4-1:0] node15537;
	wire [4-1:0] node15540;
	wire [4-1:0] node15543;
	wire [4-1:0] node15545;
	wire [4-1:0] node15546;
	wire [4-1:0] node15550;
	wire [4-1:0] node15551;
	wire [4-1:0] node15552;
	wire [4-1:0] node15553;
	wire [4-1:0] node15554;
	wire [4-1:0] node15555;
	wire [4-1:0] node15556;
	wire [4-1:0] node15559;
	wire [4-1:0] node15563;
	wire [4-1:0] node15565;
	wire [4-1:0] node15568;
	wire [4-1:0] node15569;
	wire [4-1:0] node15570;
	wire [4-1:0] node15573;
	wire [4-1:0] node15574;
	wire [4-1:0] node15577;
	wire [4-1:0] node15580;
	wire [4-1:0] node15581;
	wire [4-1:0] node15582;
	wire [4-1:0] node15586;
	wire [4-1:0] node15587;
	wire [4-1:0] node15591;
	wire [4-1:0] node15592;
	wire [4-1:0] node15593;
	wire [4-1:0] node15597;
	wire [4-1:0] node15598;
	wire [4-1:0] node15600;
	wire [4-1:0] node15603;
	wire [4-1:0] node15604;
	wire [4-1:0] node15607;
	wire [4-1:0] node15610;
	wire [4-1:0] node15611;
	wire [4-1:0] node15612;
	wire [4-1:0] node15613;
	wire [4-1:0] node15615;
	wire [4-1:0] node15619;
	wire [4-1:0] node15620;
	wire [4-1:0] node15623;
	wire [4-1:0] node15624;
	wire [4-1:0] node15625;
	wire [4-1:0] node15629;
	wire [4-1:0] node15632;
	wire [4-1:0] node15633;
	wire [4-1:0] node15634;
	wire [4-1:0] node15635;
	wire [4-1:0] node15640;
	wire [4-1:0] node15641;
	wire [4-1:0] node15642;
	wire [4-1:0] node15643;
	wire [4-1:0] node15648;
	wire [4-1:0] node15649;
	wire [4-1:0] node15650;
	wire [4-1:0] node15655;
	wire [4-1:0] node15656;
	wire [4-1:0] node15657;
	wire [4-1:0] node15658;
	wire [4-1:0] node15659;
	wire [4-1:0] node15660;
	wire [4-1:0] node15662;
	wire [4-1:0] node15664;
	wire [4-1:0] node15667;
	wire [4-1:0] node15668;
	wire [4-1:0] node15669;
	wire [4-1:0] node15674;
	wire [4-1:0] node15675;
	wire [4-1:0] node15677;
	wire [4-1:0] node15680;
	wire [4-1:0] node15683;
	wire [4-1:0] node15684;
	wire [4-1:0] node15685;
	wire [4-1:0] node15686;
	wire [4-1:0] node15689;
	wire [4-1:0] node15691;
	wire [4-1:0] node15694;
	wire [4-1:0] node15695;
	wire [4-1:0] node15696;
	wire [4-1:0] node15700;
	wire [4-1:0] node15703;
	wire [4-1:0] node15704;
	wire [4-1:0] node15707;
	wire [4-1:0] node15708;
	wire [4-1:0] node15709;
	wire [4-1:0] node15714;
	wire [4-1:0] node15715;
	wire [4-1:0] node15716;
	wire [4-1:0] node15717;
	wire [4-1:0] node15720;
	wire [4-1:0] node15721;
	wire [4-1:0] node15722;
	wire [4-1:0] node15727;
	wire [4-1:0] node15728;
	wire [4-1:0] node15731;
	wire [4-1:0] node15733;
	wire [4-1:0] node15735;
	wire [4-1:0] node15738;
	wire [4-1:0] node15739;
	wire [4-1:0] node15740;
	wire [4-1:0] node15742;
	wire [4-1:0] node15744;
	wire [4-1:0] node15747;
	wire [4-1:0] node15750;
	wire [4-1:0] node15751;
	wire [4-1:0] node15753;
	wire [4-1:0] node15754;
	wire [4-1:0] node15757;
	wire [4-1:0] node15760;
	wire [4-1:0] node15762;
	wire [4-1:0] node15764;
	wire [4-1:0] node15767;
	wire [4-1:0] node15768;
	wire [4-1:0] node15769;
	wire [4-1:0] node15770;
	wire [4-1:0] node15771;
	wire [4-1:0] node15775;
	wire [4-1:0] node15776;
	wire [4-1:0] node15777;
	wire [4-1:0] node15779;
	wire [4-1:0] node15783;
	wire [4-1:0] node15785;
	wire [4-1:0] node15786;
	wire [4-1:0] node15789;
	wire [4-1:0] node15792;
	wire [4-1:0] node15793;
	wire [4-1:0] node15794;
	wire [4-1:0] node15795;
	wire [4-1:0] node15799;
	wire [4-1:0] node15800;
	wire [4-1:0] node15801;
	wire [4-1:0] node15805;
	wire [4-1:0] node15806;
	wire [4-1:0] node15809;
	wire [4-1:0] node15812;
	wire [4-1:0] node15813;
	wire [4-1:0] node15815;
	wire [4-1:0] node15817;
	wire [4-1:0] node15820;
	wire [4-1:0] node15821;
	wire [4-1:0] node15825;
	wire [4-1:0] node15826;
	wire [4-1:0] node15827;
	wire [4-1:0] node15828;
	wire [4-1:0] node15830;
	wire [4-1:0] node15831;
	wire [4-1:0] node15834;
	wire [4-1:0] node15837;
	wire [4-1:0] node15838;
	wire [4-1:0] node15839;
	wire [4-1:0] node15843;
	wire [4-1:0] node15845;
	wire [4-1:0] node15848;
	wire [4-1:0] node15849;
	wire [4-1:0] node15850;
	wire [4-1:0] node15851;
	wire [4-1:0] node15856;
	wire [4-1:0] node15857;
	wire [4-1:0] node15858;
	wire [4-1:0] node15862;
	wire [4-1:0] node15863;
	wire [4-1:0] node15867;
	wire [4-1:0] node15868;
	wire [4-1:0] node15869;
	wire [4-1:0] node15870;
	wire [4-1:0] node15871;
	wire [4-1:0] node15876;
	wire [4-1:0] node15877;
	wire [4-1:0] node15879;
	wire [4-1:0] node15883;
	wire [4-1:0] node15884;
	wire [4-1:0] node15885;
	wire [4-1:0] node15886;
	wire [4-1:0] node15891;
	wire [4-1:0] node15893;
	wire [4-1:0] node15896;
	wire [4-1:0] node15897;
	wire [4-1:0] node15898;
	wire [4-1:0] node15899;
	wire [4-1:0] node15900;
	wire [4-1:0] node15901;
	wire [4-1:0] node15902;
	wire [4-1:0] node15904;
	wire [4-1:0] node15906;
	wire [4-1:0] node15909;
	wire [4-1:0] node15910;
	wire [4-1:0] node15912;
	wire [4-1:0] node15915;
	wire [4-1:0] node15918;
	wire [4-1:0] node15919;
	wire [4-1:0] node15921;
	wire [4-1:0] node15924;
	wire [4-1:0] node15925;
	wire [4-1:0] node15927;
	wire [4-1:0] node15930;
	wire [4-1:0] node15931;
	wire [4-1:0] node15934;
	wire [4-1:0] node15937;
	wire [4-1:0] node15938;
	wire [4-1:0] node15939;
	wire [4-1:0] node15940;
	wire [4-1:0] node15941;
	wire [4-1:0] node15944;
	wire [4-1:0] node15948;
	wire [4-1:0] node15949;
	wire [4-1:0] node15952;
	wire [4-1:0] node15954;
	wire [4-1:0] node15957;
	wire [4-1:0] node15958;
	wire [4-1:0] node15961;
	wire [4-1:0] node15962;
	wire [4-1:0] node15963;
	wire [4-1:0] node15967;
	wire [4-1:0] node15969;
	wire [4-1:0] node15972;
	wire [4-1:0] node15973;
	wire [4-1:0] node15974;
	wire [4-1:0] node15975;
	wire [4-1:0] node15976;
	wire [4-1:0] node15980;
	wire [4-1:0] node15981;
	wire [4-1:0] node15983;
	wire [4-1:0] node15987;
	wire [4-1:0] node15988;
	wire [4-1:0] node15989;
	wire [4-1:0] node15994;
	wire [4-1:0] node15995;
	wire [4-1:0] node15996;
	wire [4-1:0] node15998;
	wire [4-1:0] node16001;
	wire [4-1:0] node16002;
	wire [4-1:0] node16003;
	wire [4-1:0] node16008;
	wire [4-1:0] node16010;
	wire [4-1:0] node16011;
	wire [4-1:0] node16012;
	wire [4-1:0] node16017;
	wire [4-1:0] node16018;
	wire [4-1:0] node16019;
	wire [4-1:0] node16020;
	wire [4-1:0] node16021;
	wire [4-1:0] node16022;
	wire [4-1:0] node16023;
	wire [4-1:0] node16026;
	wire [4-1:0] node16029;
	wire [4-1:0] node16033;
	wire [4-1:0] node16034;
	wire [4-1:0] node16035;
	wire [4-1:0] node16036;
	wire [4-1:0] node16039;
	wire [4-1:0] node16043;
	wire [4-1:0] node16044;
	wire [4-1:0] node16047;
	wire [4-1:0] node16048;
	wire [4-1:0] node16052;
	wire [4-1:0] node16053;
	wire [4-1:0] node16054;
	wire [4-1:0] node16055;
	wire [4-1:0] node16058;
	wire [4-1:0] node16060;
	wire [4-1:0] node16063;
	wire [4-1:0] node16065;
	wire [4-1:0] node16068;
	wire [4-1:0] node16070;
	wire [4-1:0] node16071;
	wire [4-1:0] node16073;
	wire [4-1:0] node16077;
	wire [4-1:0] node16078;
	wire [4-1:0] node16079;
	wire [4-1:0] node16080;
	wire [4-1:0] node16083;
	wire [4-1:0] node16084;
	wire [4-1:0] node16088;
	wire [4-1:0] node16089;
	wire [4-1:0] node16092;
	wire [4-1:0] node16095;
	wire [4-1:0] node16096;
	wire [4-1:0] node16097;
	wire [4-1:0] node16100;
	wire [4-1:0] node16102;
	wire [4-1:0] node16105;
	wire [4-1:0] node16106;
	wire [4-1:0] node16107;
	wire [4-1:0] node16108;
	wire [4-1:0] node16111;
	wire [4-1:0] node16115;
	wire [4-1:0] node16116;
	wire [4-1:0] node16120;
	wire [4-1:0] node16121;
	wire [4-1:0] node16122;
	wire [4-1:0] node16123;
	wire [4-1:0] node16124;
	wire [4-1:0] node16125;
	wire [4-1:0] node16126;
	wire [4-1:0] node16129;
	wire [4-1:0] node16130;
	wire [4-1:0] node16134;
	wire [4-1:0] node16137;
	wire [4-1:0] node16138;
	wire [4-1:0] node16139;
	wire [4-1:0] node16140;
	wire [4-1:0] node16143;
	wire [4-1:0] node16146;
	wire [4-1:0] node16149;
	wire [4-1:0] node16150;
	wire [4-1:0] node16151;
	wire [4-1:0] node16154;
	wire [4-1:0] node16157;
	wire [4-1:0] node16160;
	wire [4-1:0] node16161;
	wire [4-1:0] node16162;
	wire [4-1:0] node16165;
	wire [4-1:0] node16167;
	wire [4-1:0] node16170;
	wire [4-1:0] node16171;
	wire [4-1:0] node16172;
	wire [4-1:0] node16173;
	wire [4-1:0] node16177;
	wire [4-1:0] node16178;
	wire [4-1:0] node16182;
	wire [4-1:0] node16184;
	wire [4-1:0] node16187;
	wire [4-1:0] node16188;
	wire [4-1:0] node16189;
	wire [4-1:0] node16190;
	wire [4-1:0] node16191;
	wire [4-1:0] node16193;
	wire [4-1:0] node16197;
	wire [4-1:0] node16199;
	wire [4-1:0] node16201;
	wire [4-1:0] node16204;
	wire [4-1:0] node16205;
	wire [4-1:0] node16208;
	wire [4-1:0] node16211;
	wire [4-1:0] node16212;
	wire [4-1:0] node16213;
	wire [4-1:0] node16214;
	wire [4-1:0] node16216;
	wire [4-1:0] node16220;
	wire [4-1:0] node16221;
	wire [4-1:0] node16225;
	wire [4-1:0] node16226;
	wire [4-1:0] node16227;
	wire [4-1:0] node16228;
	wire [4-1:0] node16233;
	wire [4-1:0] node16236;
	wire [4-1:0] node16237;
	wire [4-1:0] node16238;
	wire [4-1:0] node16239;
	wire [4-1:0] node16240;
	wire [4-1:0] node16242;
	wire [4-1:0] node16245;
	wire [4-1:0] node16248;
	wire [4-1:0] node16249;
	wire [4-1:0] node16250;
	wire [4-1:0] node16251;
	wire [4-1:0] node16254;
	wire [4-1:0] node16257;
	wire [4-1:0] node16260;
	wire [4-1:0] node16263;
	wire [4-1:0] node16264;
	wire [4-1:0] node16266;
	wire [4-1:0] node16267;
	wire [4-1:0] node16268;
	wire [4-1:0] node16271;
	wire [4-1:0] node16275;
	wire [4-1:0] node16276;
	wire [4-1:0] node16278;
	wire [4-1:0] node16280;
	wire [4-1:0] node16283;
	wire [4-1:0] node16285;
	wire [4-1:0] node16288;
	wire [4-1:0] node16289;
	wire [4-1:0] node16290;
	wire [4-1:0] node16292;
	wire [4-1:0] node16293;
	wire [4-1:0] node16297;
	wire [4-1:0] node16298;
	wire [4-1:0] node16301;
	wire [4-1:0] node16302;
	wire [4-1:0] node16306;
	wire [4-1:0] node16307;
	wire [4-1:0] node16310;
	wire [4-1:0] node16311;
	wire [4-1:0] node16315;
	wire [4-1:0] node16316;
	wire [4-1:0] node16317;
	wire [4-1:0] node16318;
	wire [4-1:0] node16319;
	wire [4-1:0] node16320;
	wire [4-1:0] node16321;
	wire [4-1:0] node16322;
	wire [4-1:0] node16323;
	wire [4-1:0] node16324;
	wire [4-1:0] node16325;
	wire [4-1:0] node16328;
	wire [4-1:0] node16330;
	wire [4-1:0] node16333;
	wire [4-1:0] node16336;
	wire [4-1:0] node16337;
	wire [4-1:0] node16338;
	wire [4-1:0] node16342;
	wire [4-1:0] node16343;
	wire [4-1:0] node16344;
	wire [4-1:0] node16347;
	wire [4-1:0] node16350;
	wire [4-1:0] node16351;
	wire [4-1:0] node16354;
	wire [4-1:0] node16357;
	wire [4-1:0] node16358;
	wire [4-1:0] node16359;
	wire [4-1:0] node16360;
	wire [4-1:0] node16361;
	wire [4-1:0] node16364;
	wire [4-1:0] node16368;
	wire [4-1:0] node16370;
	wire [4-1:0] node16373;
	wire [4-1:0] node16374;
	wire [4-1:0] node16375;
	wire [4-1:0] node16378;
	wire [4-1:0] node16379;
	wire [4-1:0] node16382;
	wire [4-1:0] node16385;
	wire [4-1:0] node16386;
	wire [4-1:0] node16387;
	wire [4-1:0] node16392;
	wire [4-1:0] node16393;
	wire [4-1:0] node16394;
	wire [4-1:0] node16395;
	wire [4-1:0] node16397;
	wire [4-1:0] node16400;
	wire [4-1:0] node16401;
	wire [4-1:0] node16402;
	wire [4-1:0] node16406;
	wire [4-1:0] node16409;
	wire [4-1:0] node16410;
	wire [4-1:0] node16411;
	wire [4-1:0] node16412;
	wire [4-1:0] node16417;
	wire [4-1:0] node16419;
	wire [4-1:0] node16420;
	wire [4-1:0] node16424;
	wire [4-1:0] node16425;
	wire [4-1:0] node16426;
	wire [4-1:0] node16428;
	wire [4-1:0] node16431;
	wire [4-1:0] node16434;
	wire [4-1:0] node16435;
	wire [4-1:0] node16436;
	wire [4-1:0] node16439;
	wire [4-1:0] node16440;
	wire [4-1:0] node16444;
	wire [4-1:0] node16445;
	wire [4-1:0] node16449;
	wire [4-1:0] node16450;
	wire [4-1:0] node16451;
	wire [4-1:0] node16452;
	wire [4-1:0] node16454;
	wire [4-1:0] node16456;
	wire [4-1:0] node16459;
	wire [4-1:0] node16461;
	wire [4-1:0] node16463;
	wire [4-1:0] node16466;
	wire [4-1:0] node16467;
	wire [4-1:0] node16468;
	wire [4-1:0] node16469;
	wire [4-1:0] node16470;
	wire [4-1:0] node16473;
	wire [4-1:0] node16477;
	wire [4-1:0] node16478;
	wire [4-1:0] node16482;
	wire [4-1:0] node16483;
	wire [4-1:0] node16486;
	wire [4-1:0] node16487;
	wire [4-1:0] node16490;
	wire [4-1:0] node16493;
	wire [4-1:0] node16494;
	wire [4-1:0] node16495;
	wire [4-1:0] node16496;
	wire [4-1:0] node16497;
	wire [4-1:0] node16501;
	wire [4-1:0] node16503;
	wire [4-1:0] node16504;
	wire [4-1:0] node16507;
	wire [4-1:0] node16510;
	wire [4-1:0] node16511;
	wire [4-1:0] node16512;
	wire [4-1:0] node16515;
	wire [4-1:0] node16516;
	wire [4-1:0] node16520;
	wire [4-1:0] node16523;
	wire [4-1:0] node16524;
	wire [4-1:0] node16525;
	wire [4-1:0] node16527;
	wire [4-1:0] node16528;
	wire [4-1:0] node16532;
	wire [4-1:0] node16534;
	wire [4-1:0] node16537;
	wire [4-1:0] node16538;
	wire [4-1:0] node16539;
	wire [4-1:0] node16540;
	wire [4-1:0] node16545;
	wire [4-1:0] node16547;
	wire [4-1:0] node16550;
	wire [4-1:0] node16551;
	wire [4-1:0] node16552;
	wire [4-1:0] node16553;
	wire [4-1:0] node16554;
	wire [4-1:0] node16555;
	wire [4-1:0] node16557;
	wire [4-1:0] node16558;
	wire [4-1:0] node16562;
	wire [4-1:0] node16563;
	wire [4-1:0] node16566;
	wire [4-1:0] node16569;
	wire [4-1:0] node16570;
	wire [4-1:0] node16572;
	wire [4-1:0] node16574;
	wire [4-1:0] node16577;
	wire [4-1:0] node16579;
	wire [4-1:0] node16580;
	wire [4-1:0] node16584;
	wire [4-1:0] node16585;
	wire [4-1:0] node16586;
	wire [4-1:0] node16587;
	wire [4-1:0] node16589;
	wire [4-1:0] node16592;
	wire [4-1:0] node16595;
	wire [4-1:0] node16598;
	wire [4-1:0] node16599;
	wire [4-1:0] node16600;
	wire [4-1:0] node16601;
	wire [4-1:0] node16605;
	wire [4-1:0] node16608;
	wire [4-1:0] node16611;
	wire [4-1:0] node16612;
	wire [4-1:0] node16613;
	wire [4-1:0] node16614;
	wire [4-1:0] node16616;
	wire [4-1:0] node16619;
	wire [4-1:0] node16622;
	wire [4-1:0] node16623;
	wire [4-1:0] node16624;
	wire [4-1:0] node16625;
	wire [4-1:0] node16628;
	wire [4-1:0] node16631;
	wire [4-1:0] node16634;
	wire [4-1:0] node16635;
	wire [4-1:0] node16636;
	wire [4-1:0] node16641;
	wire [4-1:0] node16642;
	wire [4-1:0] node16643;
	wire [4-1:0] node16646;
	wire [4-1:0] node16647;
	wire [4-1:0] node16650;
	wire [4-1:0] node16653;
	wire [4-1:0] node16654;
	wire [4-1:0] node16655;
	wire [4-1:0] node16658;
	wire [4-1:0] node16661;
	wire [4-1:0] node16662;
	wire [4-1:0] node16663;
	wire [4-1:0] node16667;
	wire [4-1:0] node16670;
	wire [4-1:0] node16671;
	wire [4-1:0] node16672;
	wire [4-1:0] node16673;
	wire [4-1:0] node16675;
	wire [4-1:0] node16676;
	wire [4-1:0] node16678;
	wire [4-1:0] node16681;
	wire [4-1:0] node16682;
	wire [4-1:0] node16686;
	wire [4-1:0] node16687;
	wire [4-1:0] node16688;
	wire [4-1:0] node16691;
	wire [4-1:0] node16693;
	wire [4-1:0] node16696;
	wire [4-1:0] node16697;
	wire [4-1:0] node16699;
	wire [4-1:0] node16702;
	wire [4-1:0] node16703;
	wire [4-1:0] node16707;
	wire [4-1:0] node16708;
	wire [4-1:0] node16709;
	wire [4-1:0] node16710;
	wire [4-1:0] node16713;
	wire [4-1:0] node16714;
	wire [4-1:0] node16718;
	wire [4-1:0] node16719;
	wire [4-1:0] node16720;
	wire [4-1:0] node16724;
	wire [4-1:0] node16725;
	wire [4-1:0] node16728;
	wire [4-1:0] node16731;
	wire [4-1:0] node16732;
	wire [4-1:0] node16733;
	wire [4-1:0] node16736;
	wire [4-1:0] node16738;
	wire [4-1:0] node16741;
	wire [4-1:0] node16742;
	wire [4-1:0] node16745;
	wire [4-1:0] node16746;
	wire [4-1:0] node16749;
	wire [4-1:0] node16752;
	wire [4-1:0] node16753;
	wire [4-1:0] node16754;
	wire [4-1:0] node16755;
	wire [4-1:0] node16756;
	wire [4-1:0] node16759;
	wire [4-1:0] node16760;
	wire [4-1:0] node16764;
	wire [4-1:0] node16765;
	wire [4-1:0] node16766;
	wire [4-1:0] node16771;
	wire [4-1:0] node16772;
	wire [4-1:0] node16775;
	wire [4-1:0] node16777;
	wire [4-1:0] node16778;
	wire [4-1:0] node16781;
	wire [4-1:0] node16784;
	wire [4-1:0] node16785;
	wire [4-1:0] node16786;
	wire [4-1:0] node16787;
	wire [4-1:0] node16790;
	wire [4-1:0] node16793;
	wire [4-1:0] node16794;
	wire [4-1:0] node16796;
	wire [4-1:0] node16800;
	wire [4-1:0] node16801;
	wire [4-1:0] node16804;
	wire [4-1:0] node16807;
	wire [4-1:0] node16808;
	wire [4-1:0] node16809;
	wire [4-1:0] node16810;
	wire [4-1:0] node16811;
	wire [4-1:0] node16812;
	wire [4-1:0] node16813;
	wire [4-1:0] node16814;
	wire [4-1:0] node16816;
	wire [4-1:0] node16819;
	wire [4-1:0] node16823;
	wire [4-1:0] node16824;
	wire [4-1:0] node16825;
	wire [4-1:0] node16827;
	wire [4-1:0] node16831;
	wire [4-1:0] node16832;
	wire [4-1:0] node16835;
	wire [4-1:0] node16836;
	wire [4-1:0] node16840;
	wire [4-1:0] node16841;
	wire [4-1:0] node16842;
	wire [4-1:0] node16843;
	wire [4-1:0] node16846;
	wire [4-1:0] node16850;
	wire [4-1:0] node16851;
	wire [4-1:0] node16852;
	wire [4-1:0] node16854;
	wire [4-1:0] node16859;
	wire [4-1:0] node16860;
	wire [4-1:0] node16861;
	wire [4-1:0] node16863;
	wire [4-1:0] node16865;
	wire [4-1:0] node16868;
	wire [4-1:0] node16869;
	wire [4-1:0] node16872;
	wire [4-1:0] node16873;
	wire [4-1:0] node16874;
	wire [4-1:0] node16877;
	wire [4-1:0] node16880;
	wire [4-1:0] node16882;
	wire [4-1:0] node16885;
	wire [4-1:0] node16886;
	wire [4-1:0] node16887;
	wire [4-1:0] node16889;
	wire [4-1:0] node16892;
	wire [4-1:0] node16895;
	wire [4-1:0] node16896;
	wire [4-1:0] node16897;
	wire [4-1:0] node16898;
	wire [4-1:0] node16901;
	wire [4-1:0] node16904;
	wire [4-1:0] node16907;
	wire [4-1:0] node16909;
	wire [4-1:0] node16911;
	wire [4-1:0] node16914;
	wire [4-1:0] node16915;
	wire [4-1:0] node16916;
	wire [4-1:0] node16917;
	wire [4-1:0] node16918;
	wire [4-1:0] node16919;
	wire [4-1:0] node16922;
	wire [4-1:0] node16925;
	wire [4-1:0] node16926;
	wire [4-1:0] node16927;
	wire [4-1:0] node16930;
	wire [4-1:0] node16933;
	wire [4-1:0] node16934;
	wire [4-1:0] node16937;
	wire [4-1:0] node16940;
	wire [4-1:0] node16941;
	wire [4-1:0] node16942;
	wire [4-1:0] node16946;
	wire [4-1:0] node16947;
	wire [4-1:0] node16951;
	wire [4-1:0] node16952;
	wire [4-1:0] node16953;
	wire [4-1:0] node16956;
	wire [4-1:0] node16959;
	wire [4-1:0] node16960;
	wire [4-1:0] node16961;
	wire [4-1:0] node16965;
	wire [4-1:0] node16968;
	wire [4-1:0] node16969;
	wire [4-1:0] node16970;
	wire [4-1:0] node16972;
	wire [4-1:0] node16973;
	wire [4-1:0] node16975;
	wire [4-1:0] node16978;
	wire [4-1:0] node16981;
	wire [4-1:0] node16982;
	wire [4-1:0] node16985;
	wire [4-1:0] node16986;
	wire [4-1:0] node16989;
	wire [4-1:0] node16991;
	wire [4-1:0] node16994;
	wire [4-1:0] node16995;
	wire [4-1:0] node16997;
	wire [4-1:0] node17000;
	wire [4-1:0] node17001;
	wire [4-1:0] node17002;
	wire [4-1:0] node17005;
	wire [4-1:0] node17008;
	wire [4-1:0] node17009;
	wire [4-1:0] node17010;
	wire [4-1:0] node17015;
	wire [4-1:0] node17016;
	wire [4-1:0] node17017;
	wire [4-1:0] node17018;
	wire [4-1:0] node17019;
	wire [4-1:0] node17020;
	wire [4-1:0] node17021;
	wire [4-1:0] node17023;
	wire [4-1:0] node17027;
	wire [4-1:0] node17028;
	wire [4-1:0] node17032;
	wire [4-1:0] node17033;
	wire [4-1:0] node17035;
	wire [4-1:0] node17036;
	wire [4-1:0] node17041;
	wire [4-1:0] node17042;
	wire [4-1:0] node17043;
	wire [4-1:0] node17044;
	wire [4-1:0] node17045;
	wire [4-1:0] node17048;
	wire [4-1:0] node17051;
	wire [4-1:0] node17054;
	wire [4-1:0] node17055;
	wire [4-1:0] node17057;
	wire [4-1:0] node17060;
	wire [4-1:0] node17062;
	wire [4-1:0] node17065;
	wire [4-1:0] node17066;
	wire [4-1:0] node17067;
	wire [4-1:0] node17068;
	wire [4-1:0] node17072;
	wire [4-1:0] node17074;
	wire [4-1:0] node17077;
	wire [4-1:0] node17080;
	wire [4-1:0] node17081;
	wire [4-1:0] node17082;
	wire [4-1:0] node17083;
	wire [4-1:0] node17084;
	wire [4-1:0] node17085;
	wire [4-1:0] node17088;
	wire [4-1:0] node17091;
	wire [4-1:0] node17093;
	wire [4-1:0] node17097;
	wire [4-1:0] node17098;
	wire [4-1:0] node17099;
	wire [4-1:0] node17101;
	wire [4-1:0] node17106;
	wire [4-1:0] node17107;
	wire [4-1:0] node17108;
	wire [4-1:0] node17109;
	wire [4-1:0] node17110;
	wire [4-1:0] node17114;
	wire [4-1:0] node17117;
	wire [4-1:0] node17118;
	wire [4-1:0] node17119;
	wire [4-1:0] node17124;
	wire [4-1:0] node17126;
	wire [4-1:0] node17128;
	wire [4-1:0] node17131;
	wire [4-1:0] node17132;
	wire [4-1:0] node17133;
	wire [4-1:0] node17134;
	wire [4-1:0] node17135;
	wire [4-1:0] node17136;
	wire [4-1:0] node17137;
	wire [4-1:0] node17140;
	wire [4-1:0] node17144;
	wire [4-1:0] node17145;
	wire [4-1:0] node17146;
	wire [4-1:0] node17150;
	wire [4-1:0] node17151;
	wire [4-1:0] node17155;
	wire [4-1:0] node17156;
	wire [4-1:0] node17157;
	wire [4-1:0] node17158;
	wire [4-1:0] node17162;
	wire [4-1:0] node17164;
	wire [4-1:0] node17168;
	wire [4-1:0] node17169;
	wire [4-1:0] node17170;
	wire [4-1:0] node17172;
	wire [4-1:0] node17175;
	wire [4-1:0] node17176;
	wire [4-1:0] node17179;
	wire [4-1:0] node17180;
	wire [4-1:0] node17183;
	wire [4-1:0] node17186;
	wire [4-1:0] node17187;
	wire [4-1:0] node17188;
	wire [4-1:0] node17192;
	wire [4-1:0] node17193;
	wire [4-1:0] node17195;
	wire [4-1:0] node17199;
	wire [4-1:0] node17200;
	wire [4-1:0] node17201;
	wire [4-1:0] node17202;
	wire [4-1:0] node17203;
	wire [4-1:0] node17204;
	wire [4-1:0] node17208;
	wire [4-1:0] node17212;
	wire [4-1:0] node17213;
	wire [4-1:0] node17215;
	wire [4-1:0] node17218;
	wire [4-1:0] node17219;
	wire [4-1:0] node17222;
	wire [4-1:0] node17224;
	wire [4-1:0] node17227;
	wire [4-1:0] node17228;
	wire [4-1:0] node17229;
	wire [4-1:0] node17231;
	wire [4-1:0] node17232;
	wire [4-1:0] node17236;
	wire [4-1:0] node17237;
	wire [4-1:0] node17241;
	wire [4-1:0] node17242;
	wire [4-1:0] node17245;
	wire [4-1:0] node17246;
	wire [4-1:0] node17249;
	wire [4-1:0] node17251;
	wire [4-1:0] node17254;
	wire [4-1:0] node17255;
	wire [4-1:0] node17256;
	wire [4-1:0] node17257;
	wire [4-1:0] node17258;
	wire [4-1:0] node17259;
	wire [4-1:0] node17260;
	wire [4-1:0] node17261;
	wire [4-1:0] node17264;
	wire [4-1:0] node17265;
	wire [4-1:0] node17268;
	wire [4-1:0] node17271;
	wire [4-1:0] node17272;
	wire [4-1:0] node17274;
	wire [4-1:0] node17277;
	wire [4-1:0] node17279;
	wire [4-1:0] node17282;
	wire [4-1:0] node17283;
	wire [4-1:0] node17284;
	wire [4-1:0] node17286;
	wire [4-1:0] node17288;
	wire [4-1:0] node17291;
	wire [4-1:0] node17294;
	wire [4-1:0] node17295;
	wire [4-1:0] node17296;
	wire [4-1:0] node17300;
	wire [4-1:0] node17301;
	wire [4-1:0] node17305;
	wire [4-1:0] node17306;
	wire [4-1:0] node17307;
	wire [4-1:0] node17308;
	wire [4-1:0] node17310;
	wire [4-1:0] node17313;
	wire [4-1:0] node17314;
	wire [4-1:0] node17317;
	wire [4-1:0] node17320;
	wire [4-1:0] node17321;
	wire [4-1:0] node17322;
	wire [4-1:0] node17323;
	wire [4-1:0] node17328;
	wire [4-1:0] node17330;
	wire [4-1:0] node17332;
	wire [4-1:0] node17335;
	wire [4-1:0] node17336;
	wire [4-1:0] node17337;
	wire [4-1:0] node17338;
	wire [4-1:0] node17341;
	wire [4-1:0] node17344;
	wire [4-1:0] node17345;
	wire [4-1:0] node17347;
	wire [4-1:0] node17350;
	wire [4-1:0] node17352;
	wire [4-1:0] node17355;
	wire [4-1:0] node17356;
	wire [4-1:0] node17359;
	wire [4-1:0] node17362;
	wire [4-1:0] node17363;
	wire [4-1:0] node17364;
	wire [4-1:0] node17365;
	wire [4-1:0] node17366;
	wire [4-1:0] node17368;
	wire [4-1:0] node17371;
	wire [4-1:0] node17374;
	wire [4-1:0] node17375;
	wire [4-1:0] node17376;
	wire [4-1:0] node17379;
	wire [4-1:0] node17383;
	wire [4-1:0] node17384;
	wire [4-1:0] node17385;
	wire [4-1:0] node17386;
	wire [4-1:0] node17389;
	wire [4-1:0] node17392;
	wire [4-1:0] node17394;
	wire [4-1:0] node17395;
	wire [4-1:0] node17399;
	wire [4-1:0] node17400;
	wire [4-1:0] node17403;
	wire [4-1:0] node17405;
	wire [4-1:0] node17408;
	wire [4-1:0] node17409;
	wire [4-1:0] node17410;
	wire [4-1:0] node17411;
	wire [4-1:0] node17412;
	wire [4-1:0] node17415;
	wire [4-1:0] node17417;
	wire [4-1:0] node17421;
	wire [4-1:0] node17422;
	wire [4-1:0] node17423;
	wire [4-1:0] node17426;
	wire [4-1:0] node17429;
	wire [4-1:0] node17430;
	wire [4-1:0] node17434;
	wire [4-1:0] node17435;
	wire [4-1:0] node17436;
	wire [4-1:0] node17437;
	wire [4-1:0] node17438;
	wire [4-1:0] node17441;
	wire [4-1:0] node17445;
	wire [4-1:0] node17447;
	wire [4-1:0] node17448;
	wire [4-1:0] node17451;
	wire [4-1:0] node17454;
	wire [4-1:0] node17455;
	wire [4-1:0] node17456;
	wire [4-1:0] node17457;
	wire [4-1:0] node17461;
	wire [4-1:0] node17463;
	wire [4-1:0] node17466;
	wire [4-1:0] node17468;
	wire [4-1:0] node17469;
	wire [4-1:0] node17473;
	wire [4-1:0] node17474;
	wire [4-1:0] node17475;
	wire [4-1:0] node17476;
	wire [4-1:0] node17477;
	wire [4-1:0] node17478;
	wire [4-1:0] node17479;
	wire [4-1:0] node17484;
	wire [4-1:0] node17485;
	wire [4-1:0] node17486;
	wire [4-1:0] node17487;
	wire [4-1:0] node17491;
	wire [4-1:0] node17494;
	wire [4-1:0] node17495;
	wire [4-1:0] node17499;
	wire [4-1:0] node17500;
	wire [4-1:0] node17501;
	wire [4-1:0] node17503;
	wire [4-1:0] node17505;
	wire [4-1:0] node17509;
	wire [4-1:0] node17510;
	wire [4-1:0] node17513;
	wire [4-1:0] node17514;
	wire [4-1:0] node17518;
	wire [4-1:0] node17519;
	wire [4-1:0] node17520;
	wire [4-1:0] node17521;
	wire [4-1:0] node17523;
	wire [4-1:0] node17526;
	wire [4-1:0] node17527;
	wire [4-1:0] node17529;
	wire [4-1:0] node17532;
	wire [4-1:0] node17534;
	wire [4-1:0] node17537;
	wire [4-1:0] node17539;
	wire [4-1:0] node17542;
	wire [4-1:0] node17543;
	wire [4-1:0] node17544;
	wire [4-1:0] node17547;
	wire [4-1:0] node17549;
	wire [4-1:0] node17552;
	wire [4-1:0] node17553;
	wire [4-1:0] node17557;
	wire [4-1:0] node17558;
	wire [4-1:0] node17559;
	wire [4-1:0] node17560;
	wire [4-1:0] node17561;
	wire [4-1:0] node17565;
	wire [4-1:0] node17566;
	wire [4-1:0] node17568;
	wire [4-1:0] node17572;
	wire [4-1:0] node17574;
	wire [4-1:0] node17575;
	wire [4-1:0] node17577;
	wire [4-1:0] node17581;
	wire [4-1:0] node17582;
	wire [4-1:0] node17583;
	wire [4-1:0] node17584;
	wire [4-1:0] node17585;
	wire [4-1:0] node17588;
	wire [4-1:0] node17592;
	wire [4-1:0] node17593;
	wire [4-1:0] node17595;
	wire [4-1:0] node17597;
	wire [4-1:0] node17601;
	wire [4-1:0] node17602;
	wire [4-1:0] node17603;
	wire [4-1:0] node17604;
	wire [4-1:0] node17608;
	wire [4-1:0] node17611;
	wire [4-1:0] node17612;
	wire [4-1:0] node17613;
	wire [4-1:0] node17614;
	wire [4-1:0] node17620;
	wire [4-1:0] node17621;
	wire [4-1:0] node17622;
	wire [4-1:0] node17623;
	wire [4-1:0] node17624;
	wire [4-1:0] node17625;
	wire [4-1:0] node17626;
	wire [4-1:0] node17627;
	wire [4-1:0] node17631;
	wire [4-1:0] node17632;
	wire [4-1:0] node17634;
	wire [4-1:0] node17638;
	wire [4-1:0] node17639;
	wire [4-1:0] node17642;
	wire [4-1:0] node17644;
	wire [4-1:0] node17647;
	wire [4-1:0] node17648;
	wire [4-1:0] node17649;
	wire [4-1:0] node17651;
	wire [4-1:0] node17652;
	wire [4-1:0] node17655;
	wire [4-1:0] node17659;
	wire [4-1:0] node17660;
	wire [4-1:0] node17661;
	wire [4-1:0] node17663;
	wire [4-1:0] node17667;
	wire [4-1:0] node17668;
	wire [4-1:0] node17672;
	wire [4-1:0] node17673;
	wire [4-1:0] node17674;
	wire [4-1:0] node17676;
	wire [4-1:0] node17679;
	wire [4-1:0] node17680;
	wire [4-1:0] node17682;
	wire [4-1:0] node17683;
	wire [4-1:0] node17686;
	wire [4-1:0] node17689;
	wire [4-1:0] node17690;
	wire [4-1:0] node17691;
	wire [4-1:0] node17695;
	wire [4-1:0] node17697;
	wire [4-1:0] node17700;
	wire [4-1:0] node17701;
	wire [4-1:0] node17702;
	wire [4-1:0] node17703;
	wire [4-1:0] node17705;
	wire [4-1:0] node17710;
	wire [4-1:0] node17712;
	wire [4-1:0] node17713;
	wire [4-1:0] node17714;
	wire [4-1:0] node17718;
	wire [4-1:0] node17720;
	wire [4-1:0] node17723;
	wire [4-1:0] node17724;
	wire [4-1:0] node17725;
	wire [4-1:0] node17726;
	wire [4-1:0] node17727;
	wire [4-1:0] node17730;
	wire [4-1:0] node17733;
	wire [4-1:0] node17735;
	wire [4-1:0] node17736;
	wire [4-1:0] node17740;
	wire [4-1:0] node17741;
	wire [4-1:0] node17742;
	wire [4-1:0] node17744;
	wire [4-1:0] node17748;
	wire [4-1:0] node17749;
	wire [4-1:0] node17753;
	wire [4-1:0] node17754;
	wire [4-1:0] node17755;
	wire [4-1:0] node17756;
	wire [4-1:0] node17757;
	wire [4-1:0] node17761;
	wire [4-1:0] node17762;
	wire [4-1:0] node17766;
	wire [4-1:0] node17768;
	wire [4-1:0] node17769;
	wire [4-1:0] node17773;
	wire [4-1:0] node17774;
	wire [4-1:0] node17776;
	wire [4-1:0] node17778;
	wire [4-1:0] node17781;
	wire [4-1:0] node17782;
	wire [4-1:0] node17783;
	wire [4-1:0] node17785;
	wire [4-1:0] node17789;
	wire [4-1:0] node17792;
	wire [4-1:0] node17793;
	wire [4-1:0] node17794;
	wire [4-1:0] node17795;
	wire [4-1:0] node17796;
	wire [4-1:0] node17797;
	wire [4-1:0] node17799;
	wire [4-1:0] node17800;
	wire [4-1:0] node17803;
	wire [4-1:0] node17806;
	wire [4-1:0] node17807;
	wire [4-1:0] node17808;
	wire [4-1:0] node17812;
	wire [4-1:0] node17814;
	wire [4-1:0] node17817;
	wire [4-1:0] node17818;
	wire [4-1:0] node17819;
	wire [4-1:0] node17821;
	wire [4-1:0] node17824;
	wire [4-1:0] node17826;
	wire [4-1:0] node17829;
	wire [4-1:0] node17830;
	wire [4-1:0] node17831;
	wire [4-1:0] node17834;
	wire [4-1:0] node17838;
	wire [4-1:0] node17839;
	wire [4-1:0] node17841;
	wire [4-1:0] node17844;
	wire [4-1:0] node17845;
	wire [4-1:0] node17846;
	wire [4-1:0] node17847;
	wire [4-1:0] node17851;
	wire [4-1:0] node17852;
	wire [4-1:0] node17857;
	wire [4-1:0] node17858;
	wire [4-1:0] node17859;
	wire [4-1:0] node17861;
	wire [4-1:0] node17863;
	wire [4-1:0] node17865;
	wire [4-1:0] node17869;
	wire [4-1:0] node17870;
	wire [4-1:0] node17871;
	wire [4-1:0] node17872;
	wire [4-1:0] node17876;
	wire [4-1:0] node17877;
	wire [4-1:0] node17878;
	wire [4-1:0] node17882;
	wire [4-1:0] node17883;
	wire [4-1:0] node17887;
	wire [4-1:0] node17889;
	wire [4-1:0] node17890;
	wire [4-1:0] node17892;
	wire [4-1:0] node17896;
	wire [4-1:0] node17897;
	wire [4-1:0] node17898;
	wire [4-1:0] node17899;
	wire [4-1:0] node17900;
	wire [4-1:0] node17903;
	wire [4-1:0] node17907;
	wire [4-1:0] node17908;
	wire [4-1:0] node17912;
	wire [4-1:0] node17913;
	wire [4-1:0] node17914;
	wire [4-1:0] node17915;
	wire [4-1:0] node17916;
	wire [4-1:0] node17917;
	wire [4-1:0] node17920;
	wire [4-1:0] node17926;
	wire [4-1:0] node17927;
	wire [4-1:0] node17931;
	wire [4-1:0] node17932;
	wire [4-1:0] node17933;
	wire [4-1:0] node17934;
	wire [4-1:0] node17935;
	wire [4-1:0] node17936;
	wire [4-1:0] node17937;
	wire [4-1:0] node17938;
	wire [4-1:0] node17939;
	wire [4-1:0] node17941;
	wire [4-1:0] node17942;
	wire [4-1:0] node17945;
	wire [4-1:0] node17948;
	wire [4-1:0] node17949;
	wire [4-1:0] node17952;
	wire [4-1:0] node17955;
	wire [4-1:0] node17956;
	wire [4-1:0] node17957;
	wire [4-1:0] node17958;
	wire [4-1:0] node17962;
	wire [4-1:0] node17963;
	wire [4-1:0] node17967;
	wire [4-1:0] node17968;
	wire [4-1:0] node17971;
	wire [4-1:0] node17972;
	wire [4-1:0] node17976;
	wire [4-1:0] node17977;
	wire [4-1:0] node17978;
	wire [4-1:0] node17980;
	wire [4-1:0] node17982;
	wire [4-1:0] node17985;
	wire [4-1:0] node17988;
	wire [4-1:0] node17989;
	wire [4-1:0] node17991;
	wire [4-1:0] node17992;
	wire [4-1:0] node17996;
	wire [4-1:0] node17997;
	wire [4-1:0] node17998;
	wire [4-1:0] node18003;
	wire [4-1:0] node18004;
	wire [4-1:0] node18005;
	wire [4-1:0] node18006;
	wire [4-1:0] node18007;
	wire [4-1:0] node18008;
	wire [4-1:0] node18013;
	wire [4-1:0] node18014;
	wire [4-1:0] node18017;
	wire [4-1:0] node18018;
	wire [4-1:0] node18022;
	wire [4-1:0] node18023;
	wire [4-1:0] node18025;
	wire [4-1:0] node18026;
	wire [4-1:0] node18030;
	wire [4-1:0] node18032;
	wire [4-1:0] node18035;
	wire [4-1:0] node18036;
	wire [4-1:0] node18037;
	wire [4-1:0] node18040;
	wire [4-1:0] node18043;
	wire [4-1:0] node18044;
	wire [4-1:0] node18047;
	wire [4-1:0] node18048;
	wire [4-1:0] node18049;
	wire [4-1:0] node18054;
	wire [4-1:0] node18055;
	wire [4-1:0] node18056;
	wire [4-1:0] node18057;
	wire [4-1:0] node18058;
	wire [4-1:0] node18059;
	wire [4-1:0] node18060;
	wire [4-1:0] node18064;
	wire [4-1:0] node18065;
	wire [4-1:0] node18068;
	wire [4-1:0] node18072;
	wire [4-1:0] node18073;
	wire [4-1:0] node18074;
	wire [4-1:0] node18076;
	wire [4-1:0] node18080;
	wire [4-1:0] node18082;
	wire [4-1:0] node18083;
	wire [4-1:0] node18087;
	wire [4-1:0] node18088;
	wire [4-1:0] node18089;
	wire [4-1:0] node18091;
	wire [4-1:0] node18092;
	wire [4-1:0] node18095;
	wire [4-1:0] node18098;
	wire [4-1:0] node18099;
	wire [4-1:0] node18102;
	wire [4-1:0] node18104;
	wire [4-1:0] node18107;
	wire [4-1:0] node18108;
	wire [4-1:0] node18109;
	wire [4-1:0] node18112;
	wire [4-1:0] node18113;
	wire [4-1:0] node18117;
	wire [4-1:0] node18118;
	wire [4-1:0] node18122;
	wire [4-1:0] node18123;
	wire [4-1:0] node18124;
	wire [4-1:0] node18125;
	wire [4-1:0] node18126;
	wire [4-1:0] node18128;
	wire [4-1:0] node18131;
	wire [4-1:0] node18132;
	wire [4-1:0] node18136;
	wire [4-1:0] node18139;
	wire [4-1:0] node18140;
	wire [4-1:0] node18141;
	wire [4-1:0] node18145;
	wire [4-1:0] node18146;
	wire [4-1:0] node18148;
	wire [4-1:0] node18152;
	wire [4-1:0] node18153;
	wire [4-1:0] node18155;
	wire [4-1:0] node18158;
	wire [4-1:0] node18159;
	wire [4-1:0] node18160;
	wire [4-1:0] node18164;
	wire [4-1:0] node18165;
	wire [4-1:0] node18168;
	wire [4-1:0] node18171;
	wire [4-1:0] node18172;
	wire [4-1:0] node18173;
	wire [4-1:0] node18174;
	wire [4-1:0] node18175;
	wire [4-1:0] node18176;
	wire [4-1:0] node18179;
	wire [4-1:0] node18180;
	wire [4-1:0] node18181;
	wire [4-1:0] node18185;
	wire [4-1:0] node18186;
	wire [4-1:0] node18189;
	wire [4-1:0] node18192;
	wire [4-1:0] node18193;
	wire [4-1:0] node18194;
	wire [4-1:0] node18197;
	wire [4-1:0] node18199;
	wire [4-1:0] node18202;
	wire [4-1:0] node18204;
	wire [4-1:0] node18207;
	wire [4-1:0] node18208;
	wire [4-1:0] node18209;
	wire [4-1:0] node18212;
	wire [4-1:0] node18213;
	wire [4-1:0] node18214;
	wire [4-1:0] node18218;
	wire [4-1:0] node18219;
	wire [4-1:0] node18223;
	wire [4-1:0] node18224;
	wire [4-1:0] node18225;
	wire [4-1:0] node18228;
	wire [4-1:0] node18231;
	wire [4-1:0] node18232;
	wire [4-1:0] node18233;
	wire [4-1:0] node18236;
	wire [4-1:0] node18239;
	wire [4-1:0] node18242;
	wire [4-1:0] node18243;
	wire [4-1:0] node18244;
	wire [4-1:0] node18245;
	wire [4-1:0] node18247;
	wire [4-1:0] node18250;
	wire [4-1:0] node18251;
	wire [4-1:0] node18252;
	wire [4-1:0] node18255;
	wire [4-1:0] node18258;
	wire [4-1:0] node18261;
	wire [4-1:0] node18262;
	wire [4-1:0] node18263;
	wire [4-1:0] node18264;
	wire [4-1:0] node18268;
	wire [4-1:0] node18269;
	wire [4-1:0] node18273;
	wire [4-1:0] node18274;
	wire [4-1:0] node18277;
	wire [4-1:0] node18278;
	wire [4-1:0] node18281;
	wire [4-1:0] node18284;
	wire [4-1:0] node18285;
	wire [4-1:0] node18286;
	wire [4-1:0] node18288;
	wire [4-1:0] node18290;
	wire [4-1:0] node18293;
	wire [4-1:0] node18294;
	wire [4-1:0] node18298;
	wire [4-1:0] node18299;
	wire [4-1:0] node18301;
	wire [4-1:0] node18304;
	wire [4-1:0] node18305;
	wire [4-1:0] node18307;
	wire [4-1:0] node18310;
	wire [4-1:0] node18311;
	wire [4-1:0] node18315;
	wire [4-1:0] node18316;
	wire [4-1:0] node18317;
	wire [4-1:0] node18318;
	wire [4-1:0] node18319;
	wire [4-1:0] node18321;
	wire [4-1:0] node18324;
	wire [4-1:0] node18325;
	wire [4-1:0] node18329;
	wire [4-1:0] node18330;
	wire [4-1:0] node18331;
	wire [4-1:0] node18334;
	wire [4-1:0] node18336;
	wire [4-1:0] node18339;
	wire [4-1:0] node18340;
	wire [4-1:0] node18343;
	wire [4-1:0] node18344;
	wire [4-1:0] node18347;
	wire [4-1:0] node18350;
	wire [4-1:0] node18351;
	wire [4-1:0] node18352;
	wire [4-1:0] node18353;
	wire [4-1:0] node18354;
	wire [4-1:0] node18357;
	wire [4-1:0] node18360;
	wire [4-1:0] node18361;
	wire [4-1:0] node18364;
	wire [4-1:0] node18367;
	wire [4-1:0] node18368;
	wire [4-1:0] node18372;
	wire [4-1:0] node18373;
	wire [4-1:0] node18374;
	wire [4-1:0] node18376;
	wire [4-1:0] node18379;
	wire [4-1:0] node18380;
	wire [4-1:0] node18383;
	wire [4-1:0] node18386;
	wire [4-1:0] node18387;
	wire [4-1:0] node18388;
	wire [4-1:0] node18391;
	wire [4-1:0] node18395;
	wire [4-1:0] node18396;
	wire [4-1:0] node18397;
	wire [4-1:0] node18398;
	wire [4-1:0] node18399;
	wire [4-1:0] node18400;
	wire [4-1:0] node18403;
	wire [4-1:0] node18406;
	wire [4-1:0] node18407;
	wire [4-1:0] node18411;
	wire [4-1:0] node18414;
	wire [4-1:0] node18415;
	wire [4-1:0] node18417;
	wire [4-1:0] node18418;
	wire [4-1:0] node18421;
	wire [4-1:0] node18424;
	wire [4-1:0] node18425;
	wire [4-1:0] node18426;
	wire [4-1:0] node18431;
	wire [4-1:0] node18432;
	wire [4-1:0] node18433;
	wire [4-1:0] node18434;
	wire [4-1:0] node18439;
	wire [4-1:0] node18440;
	wire [4-1:0] node18441;
	wire [4-1:0] node18444;
	wire [4-1:0] node18447;
	wire [4-1:0] node18448;
	wire [4-1:0] node18452;
	wire [4-1:0] node18453;
	wire [4-1:0] node18454;
	wire [4-1:0] node18455;
	wire [4-1:0] node18456;
	wire [4-1:0] node18457;
	wire [4-1:0] node18458;
	wire [4-1:0] node18460;
	wire [4-1:0] node18463;
	wire [4-1:0] node18465;
	wire [4-1:0] node18468;
	wire [4-1:0] node18469;
	wire [4-1:0] node18472;
	wire [4-1:0] node18474;
	wire [4-1:0] node18477;
	wire [4-1:0] node18478;
	wire [4-1:0] node18479;
	wire [4-1:0] node18482;
	wire [4-1:0] node18484;
	wire [4-1:0] node18486;
	wire [4-1:0] node18489;
	wire [4-1:0] node18490;
	wire [4-1:0] node18493;
	wire [4-1:0] node18494;
	wire [4-1:0] node18496;
	wire [4-1:0] node18499;
	wire [4-1:0] node18501;
	wire [4-1:0] node18504;
	wire [4-1:0] node18505;
	wire [4-1:0] node18506;
	wire [4-1:0] node18507;
	wire [4-1:0] node18508;
	wire [4-1:0] node18509;
	wire [4-1:0] node18514;
	wire [4-1:0] node18515;
	wire [4-1:0] node18516;
	wire [4-1:0] node18520;
	wire [4-1:0] node18521;
	wire [4-1:0] node18524;
	wire [4-1:0] node18527;
	wire [4-1:0] node18528;
	wire [4-1:0] node18529;
	wire [4-1:0] node18531;
	wire [4-1:0] node18534;
	wire [4-1:0] node18535;
	wire [4-1:0] node18538;
	wire [4-1:0] node18542;
	wire [4-1:0] node18543;
	wire [4-1:0] node18545;
	wire [4-1:0] node18548;
	wire [4-1:0] node18549;
	wire [4-1:0] node18550;
	wire [4-1:0] node18552;
	wire [4-1:0] node18556;
	wire [4-1:0] node18557;
	wire [4-1:0] node18558;
	wire [4-1:0] node18561;
	wire [4-1:0] node18564;
	wire [4-1:0] node18566;
	wire [4-1:0] node18569;
	wire [4-1:0] node18570;
	wire [4-1:0] node18571;
	wire [4-1:0] node18572;
	wire [4-1:0] node18575;
	wire [4-1:0] node18576;
	wire [4-1:0] node18579;
	wire [4-1:0] node18582;
	wire [4-1:0] node18583;
	wire [4-1:0] node18584;
	wire [4-1:0] node18585;
	wire [4-1:0] node18587;
	wire [4-1:0] node18590;
	wire [4-1:0] node18591;
	wire [4-1:0] node18596;
	wire [4-1:0] node18597;
	wire [4-1:0] node18598;
	wire [4-1:0] node18602;
	wire [4-1:0] node18603;
	wire [4-1:0] node18607;
	wire [4-1:0] node18608;
	wire [4-1:0] node18609;
	wire [4-1:0] node18610;
	wire [4-1:0] node18612;
	wire [4-1:0] node18613;
	wire [4-1:0] node18617;
	wire [4-1:0] node18619;
	wire [4-1:0] node18622;
	wire [4-1:0] node18623;
	wire [4-1:0] node18625;
	wire [4-1:0] node18628;
	wire [4-1:0] node18630;
	wire [4-1:0] node18633;
	wire [4-1:0] node18634;
	wire [4-1:0] node18635;
	wire [4-1:0] node18636;
	wire [4-1:0] node18638;
	wire [4-1:0] node18642;
	wire [4-1:0] node18643;
	wire [4-1:0] node18645;
	wire [4-1:0] node18649;
	wire [4-1:0] node18650;
	wire [4-1:0] node18651;
	wire [4-1:0] node18654;
	wire [4-1:0] node18655;
	wire [4-1:0] node18659;
	wire [4-1:0] node18660;
	wire [4-1:0] node18662;
	wire [4-1:0] node18665;
	wire [4-1:0] node18666;
	wire [4-1:0] node18670;
	wire [4-1:0] node18671;
	wire [4-1:0] node18672;
	wire [4-1:0] node18673;
	wire [4-1:0] node18674;
	wire [4-1:0] node18675;
	wire [4-1:0] node18676;
	wire [4-1:0] node18679;
	wire [4-1:0] node18680;
	wire [4-1:0] node18683;
	wire [4-1:0] node18686;
	wire [4-1:0] node18687;
	wire [4-1:0] node18688;
	wire [4-1:0] node18692;
	wire [4-1:0] node18695;
	wire [4-1:0] node18696;
	wire [4-1:0] node18697;
	wire [4-1:0] node18698;
	wire [4-1:0] node18701;
	wire [4-1:0] node18705;
	wire [4-1:0] node18706;
	wire [4-1:0] node18709;
	wire [4-1:0] node18712;
	wire [4-1:0] node18713;
	wire [4-1:0] node18714;
	wire [4-1:0] node18715;
	wire [4-1:0] node18717;
	wire [4-1:0] node18720;
	wire [4-1:0] node18723;
	wire [4-1:0] node18724;
	wire [4-1:0] node18725;
	wire [4-1:0] node18729;
	wire [4-1:0] node18732;
	wire [4-1:0] node18733;
	wire [4-1:0] node18734;
	wire [4-1:0] node18737;
	wire [4-1:0] node18739;
	wire [4-1:0] node18742;
	wire [4-1:0] node18743;
	wire [4-1:0] node18744;
	wire [4-1:0] node18747;
	wire [4-1:0] node18751;
	wire [4-1:0] node18752;
	wire [4-1:0] node18753;
	wire [4-1:0] node18754;
	wire [4-1:0] node18755;
	wire [4-1:0] node18759;
	wire [4-1:0] node18761;
	wire [4-1:0] node18763;
	wire [4-1:0] node18766;
	wire [4-1:0] node18767;
	wire [4-1:0] node18768;
	wire [4-1:0] node18769;
	wire [4-1:0] node18773;
	wire [4-1:0] node18776;
	wire [4-1:0] node18777;
	wire [4-1:0] node18781;
	wire [4-1:0] node18782;
	wire [4-1:0] node18783;
	wire [4-1:0] node18784;
	wire [4-1:0] node18785;
	wire [4-1:0] node18788;
	wire [4-1:0] node18791;
	wire [4-1:0] node18792;
	wire [4-1:0] node18795;
	wire [4-1:0] node18798;
	wire [4-1:0] node18801;
	wire [4-1:0] node18802;
	wire [4-1:0] node18803;
	wire [4-1:0] node18804;
	wire [4-1:0] node18809;
	wire [4-1:0] node18810;
	wire [4-1:0] node18813;
	wire [4-1:0] node18816;
	wire [4-1:0] node18817;
	wire [4-1:0] node18818;
	wire [4-1:0] node18819;
	wire [4-1:0] node18820;
	wire [4-1:0] node18822;
	wire [4-1:0] node18825;
	wire [4-1:0] node18826;
	wire [4-1:0] node18828;
	wire [4-1:0] node18832;
	wire [4-1:0] node18833;
	wire [4-1:0] node18834;
	wire [4-1:0] node18835;
	wire [4-1:0] node18840;
	wire [4-1:0] node18842;
	wire [4-1:0] node18843;
	wire [4-1:0] node18847;
	wire [4-1:0] node18848;
	wire [4-1:0] node18849;
	wire [4-1:0] node18850;
	wire [4-1:0] node18853;
	wire [4-1:0] node18854;
	wire [4-1:0] node18858;
	wire [4-1:0] node18859;
	wire [4-1:0] node18863;
	wire [4-1:0] node18864;
	wire [4-1:0] node18866;
	wire [4-1:0] node18868;
	wire [4-1:0] node18872;
	wire [4-1:0] node18873;
	wire [4-1:0] node18874;
	wire [4-1:0] node18875;
	wire [4-1:0] node18878;
	wire [4-1:0] node18879;
	wire [4-1:0] node18882;
	wire [4-1:0] node18885;
	wire [4-1:0] node18887;
	wire [4-1:0] node18888;
	wire [4-1:0] node18889;
	wire [4-1:0] node18894;
	wire [4-1:0] node18895;
	wire [4-1:0] node18896;
	wire [4-1:0] node18897;
	wire [4-1:0] node18899;
	wire [4-1:0] node18902;
	wire [4-1:0] node18903;
	wire [4-1:0] node18906;
	wire [4-1:0] node18909;
	wire [4-1:0] node18912;
	wire [4-1:0] node18913;
	wire [4-1:0] node18914;
	wire [4-1:0] node18918;
	wire [4-1:0] node18919;
	wire [4-1:0] node18922;
	wire [4-1:0] node18923;
	wire [4-1:0] node18927;
	wire [4-1:0] node18928;
	wire [4-1:0] node18929;
	wire [4-1:0] node18930;
	wire [4-1:0] node18931;
	wire [4-1:0] node18932;
	wire [4-1:0] node18933;
	wire [4-1:0] node18935;
	wire [4-1:0] node18936;
	wire [4-1:0] node18938;
	wire [4-1:0] node18941;
	wire [4-1:0] node18942;
	wire [4-1:0] node18945;
	wire [4-1:0] node18948;
	wire [4-1:0] node18950;
	wire [4-1:0] node18953;
	wire [4-1:0] node18954;
	wire [4-1:0] node18956;
	wire [4-1:0] node18959;
	wire [4-1:0] node18960;
	wire [4-1:0] node18962;
	wire [4-1:0] node18964;
	wire [4-1:0] node18967;
	wire [4-1:0] node18969;
	wire [4-1:0] node18972;
	wire [4-1:0] node18973;
	wire [4-1:0] node18974;
	wire [4-1:0] node18976;
	wire [4-1:0] node18978;
	wire [4-1:0] node18981;
	wire [4-1:0] node18982;
	wire [4-1:0] node18986;
	wire [4-1:0] node18987;
	wire [4-1:0] node18988;
	wire [4-1:0] node18989;
	wire [4-1:0] node18992;
	wire [4-1:0] node18995;
	wire [4-1:0] node18997;
	wire [4-1:0] node18998;
	wire [4-1:0] node19002;
	wire [4-1:0] node19003;
	wire [4-1:0] node19005;
	wire [4-1:0] node19006;
	wire [4-1:0] node19009;
	wire [4-1:0] node19013;
	wire [4-1:0] node19014;
	wire [4-1:0] node19015;
	wire [4-1:0] node19016;
	wire [4-1:0] node19017;
	wire [4-1:0] node19019;
	wire [4-1:0] node19022;
	wire [4-1:0] node19023;
	wire [4-1:0] node19024;
	wire [4-1:0] node19028;
	wire [4-1:0] node19029;
	wire [4-1:0] node19033;
	wire [4-1:0] node19034;
	wire [4-1:0] node19035;
	wire [4-1:0] node19040;
	wire [4-1:0] node19041;
	wire [4-1:0] node19042;
	wire [4-1:0] node19043;
	wire [4-1:0] node19045;
	wire [4-1:0] node19050;
	wire [4-1:0] node19051;
	wire [4-1:0] node19055;
	wire [4-1:0] node19056;
	wire [4-1:0] node19057;
	wire [4-1:0] node19058;
	wire [4-1:0] node19062;
	wire [4-1:0] node19063;
	wire [4-1:0] node19066;
	wire [4-1:0] node19069;
	wire [4-1:0] node19070;
	wire [4-1:0] node19071;
	wire [4-1:0] node19072;
	wire [4-1:0] node19075;
	wire [4-1:0] node19078;
	wire [4-1:0] node19080;
	wire [4-1:0] node19083;
	wire [4-1:0] node19084;
	wire [4-1:0] node19085;
	wire [4-1:0] node19086;
	wire [4-1:0] node19089;
	wire [4-1:0] node19093;
	wire [4-1:0] node19095;
	wire [4-1:0] node19098;
	wire [4-1:0] node19099;
	wire [4-1:0] node19100;
	wire [4-1:0] node19101;
	wire [4-1:0] node19102;
	wire [4-1:0] node19103;
	wire [4-1:0] node19104;
	wire [4-1:0] node19108;
	wire [4-1:0] node19109;
	wire [4-1:0] node19112;
	wire [4-1:0] node19115;
	wire [4-1:0] node19116;
	wire [4-1:0] node19118;
	wire [4-1:0] node19123;
	wire [4-1:0] node19124;
	wire [4-1:0] node19125;
	wire [4-1:0] node19126;
	wire [4-1:0] node19127;
	wire [4-1:0] node19130;
	wire [4-1:0] node19134;
	wire [4-1:0] node19136;
	wire [4-1:0] node19137;
	wire [4-1:0] node19138;
	wire [4-1:0] node19142;
	wire [4-1:0] node19143;
	wire [4-1:0] node19146;
	wire [4-1:0] node19150;
	wire [4-1:0] node19151;
	wire [4-1:0] node19152;
	wire [4-1:0] node19156;
	wire [4-1:0] node19157;
	wire [4-1:0] node19161;
	wire [4-1:0] node19162;
	wire [4-1:0] node19163;
	wire [4-1:0] node19164;
	wire [4-1:0] node19165;
	wire [4-1:0] node19166;
	wire [4-1:0] node19167;
	wire [4-1:0] node19168;
	wire [4-1:0] node19172;
	wire [4-1:0] node19173;
	wire [4-1:0] node19175;
	wire [4-1:0] node19179;
	wire [4-1:0] node19180;
	wire [4-1:0] node19181;
	wire [4-1:0] node19185;
	wire [4-1:0] node19186;
	wire [4-1:0] node19190;
	wire [4-1:0] node19191;
	wire [4-1:0] node19192;
	wire [4-1:0] node19193;
	wire [4-1:0] node19195;
	wire [4-1:0] node19198;
	wire [4-1:0] node19202;
	wire [4-1:0] node19203;
	wire [4-1:0] node19204;
	wire [4-1:0] node19205;
	wire [4-1:0] node19209;
	wire [4-1:0] node19210;
	wire [4-1:0] node19215;
	wire [4-1:0] node19216;
	wire [4-1:0] node19217;
	wire [4-1:0] node19219;
	wire [4-1:0] node19221;
	wire [4-1:0] node19224;
	wire [4-1:0] node19225;
	wire [4-1:0] node19226;
	wire [4-1:0] node19227;
	wire [4-1:0] node19230;
	wire [4-1:0] node19233;
	wire [4-1:0] node19234;
	wire [4-1:0] node19237;
	wire [4-1:0] node19240;
	wire [4-1:0] node19242;
	wire [4-1:0] node19245;
	wire [4-1:0] node19246;
	wire [4-1:0] node19247;
	wire [4-1:0] node19248;
	wire [4-1:0] node19249;
	wire [4-1:0] node19252;
	wire [4-1:0] node19256;
	wire [4-1:0] node19257;
	wire [4-1:0] node19258;
	wire [4-1:0] node19261;
	wire [4-1:0] node19265;
	wire [4-1:0] node19266;
	wire [4-1:0] node19267;
	wire [4-1:0] node19271;
	wire [4-1:0] node19273;
	wire [4-1:0] node19274;
	wire [4-1:0] node19277;
	wire [4-1:0] node19280;
	wire [4-1:0] node19281;
	wire [4-1:0] node19282;
	wire [4-1:0] node19283;
	wire [4-1:0] node19284;
	wire [4-1:0] node19286;
	wire [4-1:0] node19289;
	wire [4-1:0] node19292;
	wire [4-1:0] node19294;
	wire [4-1:0] node19296;
	wire [4-1:0] node19299;
	wire [4-1:0] node19300;
	wire [4-1:0] node19302;
	wire [4-1:0] node19303;
	wire [4-1:0] node19305;
	wire [4-1:0] node19308;
	wire [4-1:0] node19309;
	wire [4-1:0] node19312;
	wire [4-1:0] node19315;
	wire [4-1:0] node19316;
	wire [4-1:0] node19317;
	wire [4-1:0] node19322;
	wire [4-1:0] node19323;
	wire [4-1:0] node19324;
	wire [4-1:0] node19325;
	wire [4-1:0] node19326;
	wire [4-1:0] node19327;
	wire [4-1:0] node19330;
	wire [4-1:0] node19333;
	wire [4-1:0] node19335;
	wire [4-1:0] node19338;
	wire [4-1:0] node19339;
	wire [4-1:0] node19341;
	wire [4-1:0] node19345;
	wire [4-1:0] node19346;
	wire [4-1:0] node19349;
	wire [4-1:0] node19352;
	wire [4-1:0] node19353;
	wire [4-1:0] node19354;
	wire [4-1:0] node19357;
	wire [4-1:0] node19358;
	wire [4-1:0] node19361;
	wire [4-1:0] node19362;
	wire [4-1:0] node19366;
	wire [4-1:0] node19367;
	wire [4-1:0] node19369;
	wire [4-1:0] node19370;
	wire [4-1:0] node19375;
	wire [4-1:0] node19376;
	wire [4-1:0] node19377;
	wire [4-1:0] node19378;
	wire [4-1:0] node19379;
	wire [4-1:0] node19383;
	wire [4-1:0] node19384;
	wire [4-1:0] node19389;
	wire [4-1:0] node19390;
	wire [4-1:0] node19391;
	wire [4-1:0] node19392;
	wire [4-1:0] node19396;
	wire [4-1:0] node19397;
	wire [4-1:0] node19402;
	wire [4-1:0] node19403;
	wire [4-1:0] node19404;
	wire [4-1:0] node19405;
	wire [4-1:0] node19406;
	wire [4-1:0] node19407;
	wire [4-1:0] node19408;
	wire [4-1:0] node19409;
	wire [4-1:0] node19410;
	wire [4-1:0] node19411;
	wire [4-1:0] node19412;
	wire [4-1:0] node19414;
	wire [4-1:0] node19415;
	wire [4-1:0] node19420;
	wire [4-1:0] node19421;
	wire [4-1:0] node19422;
	wire [4-1:0] node19426;
	wire [4-1:0] node19427;
	wire [4-1:0] node19430;
	wire [4-1:0] node19432;
	wire [4-1:0] node19435;
	wire [4-1:0] node19436;
	wire [4-1:0] node19437;
	wire [4-1:0] node19438;
	wire [4-1:0] node19442;
	wire [4-1:0] node19443;
	wire [4-1:0] node19444;
	wire [4-1:0] node19449;
	wire [4-1:0] node19450;
	wire [4-1:0] node19452;
	wire [4-1:0] node19453;
	wire [4-1:0] node19456;
	wire [4-1:0] node19459;
	wire [4-1:0] node19460;
	wire [4-1:0] node19463;
	wire [4-1:0] node19466;
	wire [4-1:0] node19467;
	wire [4-1:0] node19468;
	wire [4-1:0] node19469;
	wire [4-1:0] node19472;
	wire [4-1:0] node19475;
	wire [4-1:0] node19477;
	wire [4-1:0] node19478;
	wire [4-1:0] node19482;
	wire [4-1:0] node19483;
	wire [4-1:0] node19484;
	wire [4-1:0] node19485;
	wire [4-1:0] node19486;
	wire [4-1:0] node19490;
	wire [4-1:0] node19493;
	wire [4-1:0] node19494;
	wire [4-1:0] node19498;
	wire [4-1:0] node19499;
	wire [4-1:0] node19500;
	wire [4-1:0] node19501;
	wire [4-1:0] node19505;
	wire [4-1:0] node19508;
	wire [4-1:0] node19509;
	wire [4-1:0] node19511;
	wire [4-1:0] node19514;
	wire [4-1:0] node19516;
	wire [4-1:0] node19519;
	wire [4-1:0] node19520;
	wire [4-1:0] node19521;
	wire [4-1:0] node19522;
	wire [4-1:0] node19524;
	wire [4-1:0] node19525;
	wire [4-1:0] node19526;
	wire [4-1:0] node19530;
	wire [4-1:0] node19531;
	wire [4-1:0] node19534;
	wire [4-1:0] node19537;
	wire [4-1:0] node19538;
	wire [4-1:0] node19539;
	wire [4-1:0] node19540;
	wire [4-1:0] node19545;
	wire [4-1:0] node19546;
	wire [4-1:0] node19547;
	wire [4-1:0] node19550;
	wire [4-1:0] node19554;
	wire [4-1:0] node19555;
	wire [4-1:0] node19556;
	wire [4-1:0] node19557;
	wire [4-1:0] node19558;
	wire [4-1:0] node19562;
	wire [4-1:0] node19566;
	wire [4-1:0] node19567;
	wire [4-1:0] node19568;
	wire [4-1:0] node19570;
	wire [4-1:0] node19573;
	wire [4-1:0] node19575;
	wire [4-1:0] node19578;
	wire [4-1:0] node19579;
	wire [4-1:0] node19581;
	wire [4-1:0] node19584;
	wire [4-1:0] node19585;
	wire [4-1:0] node19589;
	wire [4-1:0] node19590;
	wire [4-1:0] node19591;
	wire [4-1:0] node19592;
	wire [4-1:0] node19593;
	wire [4-1:0] node19597;
	wire [4-1:0] node19598;
	wire [4-1:0] node19602;
	wire [4-1:0] node19603;
	wire [4-1:0] node19604;
	wire [4-1:0] node19607;
	wire [4-1:0] node19610;
	wire [4-1:0] node19611;
	wire [4-1:0] node19615;
	wire [4-1:0] node19616;
	wire [4-1:0] node19617;
	wire [4-1:0] node19618;
	wire [4-1:0] node19619;
	wire [4-1:0] node19623;
	wire [4-1:0] node19626;
	wire [4-1:0] node19627;
	wire [4-1:0] node19629;
	wire [4-1:0] node19632;
	wire [4-1:0] node19633;
	wire [4-1:0] node19637;
	wire [4-1:0] node19638;
	wire [4-1:0] node19641;
	wire [4-1:0] node19642;
	wire [4-1:0] node19644;
	wire [4-1:0] node19648;
	wire [4-1:0] node19649;
	wire [4-1:0] node19650;
	wire [4-1:0] node19651;
	wire [4-1:0] node19652;
	wire [4-1:0] node19653;
	wire [4-1:0] node19655;
	wire [4-1:0] node19658;
	wire [4-1:0] node19660;
	wire [4-1:0] node19661;
	wire [4-1:0] node19665;
	wire [4-1:0] node19666;
	wire [4-1:0] node19669;
	wire [4-1:0] node19672;
	wire [4-1:0] node19673;
	wire [4-1:0] node19675;
	wire [4-1:0] node19678;
	wire [4-1:0] node19679;
	wire [4-1:0] node19681;
	wire [4-1:0] node19684;
	wire [4-1:0] node19685;
	wire [4-1:0] node19688;
	wire [4-1:0] node19691;
	wire [4-1:0] node19692;
	wire [4-1:0] node19693;
	wire [4-1:0] node19694;
	wire [4-1:0] node19696;
	wire [4-1:0] node19699;
	wire [4-1:0] node19701;
	wire [4-1:0] node19704;
	wire [4-1:0] node19705;
	wire [4-1:0] node19706;
	wire [4-1:0] node19710;
	wire [4-1:0] node19711;
	wire [4-1:0] node19714;
	wire [4-1:0] node19717;
	wire [4-1:0] node19718;
	wire [4-1:0] node19719;
	wire [4-1:0] node19720;
	wire [4-1:0] node19724;
	wire [4-1:0] node19727;
	wire [4-1:0] node19728;
	wire [4-1:0] node19729;
	wire [4-1:0] node19731;
	wire [4-1:0] node19735;
	wire [4-1:0] node19737;
	wire [4-1:0] node19738;
	wire [4-1:0] node19741;
	wire [4-1:0] node19744;
	wire [4-1:0] node19745;
	wire [4-1:0] node19746;
	wire [4-1:0] node19747;
	wire [4-1:0] node19748;
	wire [4-1:0] node19751;
	wire [4-1:0] node19754;
	wire [4-1:0] node19755;
	wire [4-1:0] node19757;
	wire [4-1:0] node19760;
	wire [4-1:0] node19763;
	wire [4-1:0] node19764;
	wire [4-1:0] node19765;
	wire [4-1:0] node19766;
	wire [4-1:0] node19767;
	wire [4-1:0] node19771;
	wire [4-1:0] node19772;
	wire [4-1:0] node19775;
	wire [4-1:0] node19778;
	wire [4-1:0] node19780;
	wire [4-1:0] node19781;
	wire [4-1:0] node19784;
	wire [4-1:0] node19787;
	wire [4-1:0] node19788;
	wire [4-1:0] node19789;
	wire [4-1:0] node19793;
	wire [4-1:0] node19796;
	wire [4-1:0] node19797;
	wire [4-1:0] node19798;
	wire [4-1:0] node19799;
	wire [4-1:0] node19800;
	wire [4-1:0] node19802;
	wire [4-1:0] node19807;
	wire [4-1:0] node19808;
	wire [4-1:0] node19811;
	wire [4-1:0] node19813;
	wire [4-1:0] node19816;
	wire [4-1:0] node19817;
	wire [4-1:0] node19818;
	wire [4-1:0] node19820;
	wire [4-1:0] node19821;
	wire [4-1:0] node19824;
	wire [4-1:0] node19828;
	wire [4-1:0] node19829;
	wire [4-1:0] node19832;
	wire [4-1:0] node19833;
	wire [4-1:0] node19834;
	wire [4-1:0] node19839;
	wire [4-1:0] node19840;
	wire [4-1:0] node19841;
	wire [4-1:0] node19842;
	wire [4-1:0] node19843;
	wire [4-1:0] node19844;
	wire [4-1:0] node19846;
	wire [4-1:0] node19847;
	wire [4-1:0] node19848;
	wire [4-1:0] node19853;
	wire [4-1:0] node19854;
	wire [4-1:0] node19857;
	wire [4-1:0] node19860;
	wire [4-1:0] node19861;
	wire [4-1:0] node19862;
	wire [4-1:0] node19864;
	wire [4-1:0] node19868;
	wire [4-1:0] node19869;
	wire [4-1:0] node19872;
	wire [4-1:0] node19875;
	wire [4-1:0] node19876;
	wire [4-1:0] node19877;
	wire [4-1:0] node19878;
	wire [4-1:0] node19881;
	wire [4-1:0] node19882;
	wire [4-1:0] node19883;
	wire [4-1:0] node19887;
	wire [4-1:0] node19889;
	wire [4-1:0] node19892;
	wire [4-1:0] node19893;
	wire [4-1:0] node19894;
	wire [4-1:0] node19897;
	wire [4-1:0] node19900;
	wire [4-1:0] node19903;
	wire [4-1:0] node19904;
	wire [4-1:0] node19906;
	wire [4-1:0] node19909;
	wire [4-1:0] node19910;
	wire [4-1:0] node19911;
	wire [4-1:0] node19912;
	wire [4-1:0] node19916;
	wire [4-1:0] node19917;
	wire [4-1:0] node19920;
	wire [4-1:0] node19923;
	wire [4-1:0] node19925;
	wire [4-1:0] node19928;
	wire [4-1:0] node19929;
	wire [4-1:0] node19930;
	wire [4-1:0] node19931;
	wire [4-1:0] node19932;
	wire [4-1:0] node19933;
	wire [4-1:0] node19937;
	wire [4-1:0] node19939;
	wire [4-1:0] node19942;
	wire [4-1:0] node19943;
	wire [4-1:0] node19944;
	wire [4-1:0] node19948;
	wire [4-1:0] node19949;
	wire [4-1:0] node19953;
	wire [4-1:0] node19954;
	wire [4-1:0] node19955;
	wire [4-1:0] node19959;
	wire [4-1:0] node19960;
	wire [4-1:0] node19961;
	wire [4-1:0] node19963;
	wire [4-1:0] node19967;
	wire [4-1:0] node19968;
	wire [4-1:0] node19972;
	wire [4-1:0] node19973;
	wire [4-1:0] node19974;
	wire [4-1:0] node19975;
	wire [4-1:0] node19976;
	wire [4-1:0] node19979;
	wire [4-1:0] node19982;
	wire [4-1:0] node19985;
	wire [4-1:0] node19986;
	wire [4-1:0] node19988;
	wire [4-1:0] node19991;
	wire [4-1:0] node19994;
	wire [4-1:0] node19995;
	wire [4-1:0] node19996;
	wire [4-1:0] node19997;
	wire [4-1:0] node20001;
	wire [4-1:0] node20004;
	wire [4-1:0] node20005;
	wire [4-1:0] node20006;
	wire [4-1:0] node20010;
	wire [4-1:0] node20013;
	wire [4-1:0] node20014;
	wire [4-1:0] node20015;
	wire [4-1:0] node20016;
	wire [4-1:0] node20017;
	wire [4-1:0] node20019;
	wire [4-1:0] node20022;
	wire [4-1:0] node20023;
	wire [4-1:0] node20024;
	wire [4-1:0] node20028;
	wire [4-1:0] node20031;
	wire [4-1:0] node20032;
	wire [4-1:0] node20033;
	wire [4-1:0] node20034;
	wire [4-1:0] node20038;
	wire [4-1:0] node20039;
	wire [4-1:0] node20041;
	wire [4-1:0] node20045;
	wire [4-1:0] node20046;
	wire [4-1:0] node20049;
	wire [4-1:0] node20052;
	wire [4-1:0] node20053;
	wire [4-1:0] node20054;
	wire [4-1:0] node20056;
	wire [4-1:0] node20059;
	wire [4-1:0] node20060;
	wire [4-1:0] node20064;
	wire [4-1:0] node20065;
	wire [4-1:0] node20066;
	wire [4-1:0] node20069;
	wire [4-1:0] node20072;
	wire [4-1:0] node20074;
	wire [4-1:0] node20077;
	wire [4-1:0] node20078;
	wire [4-1:0] node20079;
	wire [4-1:0] node20080;
	wire [4-1:0] node20083;
	wire [4-1:0] node20084;
	wire [4-1:0] node20087;
	wire [4-1:0] node20089;
	wire [4-1:0] node20092;
	wire [4-1:0] node20093;
	wire [4-1:0] node20094;
	wire [4-1:0] node20096;
	wire [4-1:0] node20097;
	wire [4-1:0] node20101;
	wire [4-1:0] node20103;
	wire [4-1:0] node20106;
	wire [4-1:0] node20108;
	wire [4-1:0] node20111;
	wire [4-1:0] node20112;
	wire [4-1:0] node20113;
	wire [4-1:0] node20114;
	wire [4-1:0] node20117;
	wire [4-1:0] node20118;
	wire [4-1:0] node20122;
	wire [4-1:0] node20125;
	wire [4-1:0] node20126;
	wire [4-1:0] node20127;
	wire [4-1:0] node20129;
	wire [4-1:0] node20132;
	wire [4-1:0] node20135;
	wire [4-1:0] node20136;
	wire [4-1:0] node20137;
	wire [4-1:0] node20140;
	wire [4-1:0] node20143;
	wire [4-1:0] node20144;
	wire [4-1:0] node20146;
	wire [4-1:0] node20150;
	wire [4-1:0] node20151;
	wire [4-1:0] node20152;
	wire [4-1:0] node20153;
	wire [4-1:0] node20154;
	wire [4-1:0] node20155;
	wire [4-1:0] node20156;
	wire [4-1:0] node20159;
	wire [4-1:0] node20160;
	wire [4-1:0] node20161;
	wire [4-1:0] node20162;
	wire [4-1:0] node20165;
	wire [4-1:0] node20169;
	wire [4-1:0] node20172;
	wire [4-1:0] node20173;
	wire [4-1:0] node20174;
	wire [4-1:0] node20176;
	wire [4-1:0] node20178;
	wire [4-1:0] node20182;
	wire [4-1:0] node20183;
	wire [4-1:0] node20184;
	wire [4-1:0] node20189;
	wire [4-1:0] node20190;
	wire [4-1:0] node20191;
	wire [4-1:0] node20192;
	wire [4-1:0] node20193;
	wire [4-1:0] node20194;
	wire [4-1:0] node20197;
	wire [4-1:0] node20200;
	wire [4-1:0] node20203;
	wire [4-1:0] node20204;
	wire [4-1:0] node20206;
	wire [4-1:0] node20209;
	wire [4-1:0] node20211;
	wire [4-1:0] node20214;
	wire [4-1:0] node20215;
	wire [4-1:0] node20216;
	wire [4-1:0] node20219;
	wire [4-1:0] node20222;
	wire [4-1:0] node20223;
	wire [4-1:0] node20224;
	wire [4-1:0] node20227;
	wire [4-1:0] node20231;
	wire [4-1:0] node20232;
	wire [4-1:0] node20235;
	wire [4-1:0] node20236;
	wire [4-1:0] node20240;
	wire [4-1:0] node20241;
	wire [4-1:0] node20242;
	wire [4-1:0] node20243;
	wire [4-1:0] node20244;
	wire [4-1:0] node20246;
	wire [4-1:0] node20248;
	wire [4-1:0] node20251;
	wire [4-1:0] node20253;
	wire [4-1:0] node20256;
	wire [4-1:0] node20258;
	wire [4-1:0] node20261;
	wire [4-1:0] node20262;
	wire [4-1:0] node20264;
	wire [4-1:0] node20265;
	wire [4-1:0] node20269;
	wire [4-1:0] node20270;
	wire [4-1:0] node20272;
	wire [4-1:0] node20275;
	wire [4-1:0] node20276;
	wire [4-1:0] node20280;
	wire [4-1:0] node20281;
	wire [4-1:0] node20282;
	wire [4-1:0] node20283;
	wire [4-1:0] node20284;
	wire [4-1:0] node20287;
	wire [4-1:0] node20290;
	wire [4-1:0] node20291;
	wire [4-1:0] node20295;
	wire [4-1:0] node20296;
	wire [4-1:0] node20298;
	wire [4-1:0] node20301;
	wire [4-1:0] node20302;
	wire [4-1:0] node20306;
	wire [4-1:0] node20307;
	wire [4-1:0] node20308;
	wire [4-1:0] node20311;
	wire [4-1:0] node20312;
	wire [4-1:0] node20316;
	wire [4-1:0] node20319;
	wire [4-1:0] node20320;
	wire [4-1:0] node20321;
	wire [4-1:0] node20322;
	wire [4-1:0] node20323;
	wire [4-1:0] node20324;
	wire [4-1:0] node20326;
	wire [4-1:0] node20330;
	wire [4-1:0] node20332;
	wire [4-1:0] node20334;
	wire [4-1:0] node20335;
	wire [4-1:0] node20338;
	wire [4-1:0] node20341;
	wire [4-1:0] node20343;
	wire [4-1:0] node20344;
	wire [4-1:0] node20348;
	wire [4-1:0] node20349;
	wire [4-1:0] node20350;
	wire [4-1:0] node20352;
	wire [4-1:0] node20353;
	wire [4-1:0] node20356;
	wire [4-1:0] node20357;
	wire [4-1:0] node20361;
	wire [4-1:0] node20362;
	wire [4-1:0] node20363;
	wire [4-1:0] node20364;
	wire [4-1:0] node20367;
	wire [4-1:0] node20371;
	wire [4-1:0] node20372;
	wire [4-1:0] node20376;
	wire [4-1:0] node20377;
	wire [4-1:0] node20379;
	wire [4-1:0] node20380;
	wire [4-1:0] node20381;
	wire [4-1:0] node20386;
	wire [4-1:0] node20387;
	wire [4-1:0] node20391;
	wire [4-1:0] node20392;
	wire [4-1:0] node20393;
	wire [4-1:0] node20394;
	wire [4-1:0] node20396;
	wire [4-1:0] node20399;
	wire [4-1:0] node20401;
	wire [4-1:0] node20403;
	wire [4-1:0] node20406;
	wire [4-1:0] node20407;
	wire [4-1:0] node20408;
	wire [4-1:0] node20409;
	wire [4-1:0] node20411;
	wire [4-1:0] node20415;
	wire [4-1:0] node20416;
	wire [4-1:0] node20417;
	wire [4-1:0] node20421;
	wire [4-1:0] node20423;
	wire [4-1:0] node20426;
	wire [4-1:0] node20428;
	wire [4-1:0] node20429;
	wire [4-1:0] node20433;
	wire [4-1:0] node20434;
	wire [4-1:0] node20435;
	wire [4-1:0] node20436;
	wire [4-1:0] node20437;
	wire [4-1:0] node20439;
	wire [4-1:0] node20444;
	wire [4-1:0] node20446;
	wire [4-1:0] node20448;
	wire [4-1:0] node20450;
	wire [4-1:0] node20453;
	wire [4-1:0] node20454;
	wire [4-1:0] node20455;
	wire [4-1:0] node20456;
	wire [4-1:0] node20461;
	wire [4-1:0] node20463;
	wire [4-1:0] node20465;
	wire [4-1:0] node20466;
	wire [4-1:0] node20470;
	wire [4-1:0] node20471;
	wire [4-1:0] node20472;
	wire [4-1:0] node20473;
	wire [4-1:0] node20474;
	wire [4-1:0] node20475;
	wire [4-1:0] node20477;
	wire [4-1:0] node20479;
	wire [4-1:0] node20482;
	wire [4-1:0] node20484;
	wire [4-1:0] node20485;
	wire [4-1:0] node20487;
	wire [4-1:0] node20491;
	wire [4-1:0] node20492;
	wire [4-1:0] node20495;
	wire [4-1:0] node20496;
	wire [4-1:0] node20498;
	wire [4-1:0] node20502;
	wire [4-1:0] node20503;
	wire [4-1:0] node20504;
	wire [4-1:0] node20505;
	wire [4-1:0] node20508;
	wire [4-1:0] node20510;
	wire [4-1:0] node20513;
	wire [4-1:0] node20515;
	wire [4-1:0] node20517;
	wire [4-1:0] node20518;
	wire [4-1:0] node20521;
	wire [4-1:0] node20524;
	wire [4-1:0] node20525;
	wire [4-1:0] node20526;
	wire [4-1:0] node20528;
	wire [4-1:0] node20531;
	wire [4-1:0] node20532;
	wire [4-1:0] node20533;
	wire [4-1:0] node20536;
	wire [4-1:0] node20540;
	wire [4-1:0] node20541;
	wire [4-1:0] node20542;
	wire [4-1:0] node20546;
	wire [4-1:0] node20549;
	wire [4-1:0] node20550;
	wire [4-1:0] node20551;
	wire [4-1:0] node20553;
	wire [4-1:0] node20555;
	wire [4-1:0] node20557;
	wire [4-1:0] node20558;
	wire [4-1:0] node20561;
	wire [4-1:0] node20564;
	wire [4-1:0] node20565;
	wire [4-1:0] node20566;
	wire [4-1:0] node20567;
	wire [4-1:0] node20569;
	wire [4-1:0] node20572;
	wire [4-1:0] node20573;
	wire [4-1:0] node20577;
	wire [4-1:0] node20578;
	wire [4-1:0] node20582;
	wire [4-1:0] node20584;
	wire [4-1:0] node20587;
	wire [4-1:0] node20588;
	wire [4-1:0] node20589;
	wire [4-1:0] node20590;
	wire [4-1:0] node20591;
	wire [4-1:0] node20593;
	wire [4-1:0] node20597;
	wire [4-1:0] node20598;
	wire [4-1:0] node20603;
	wire [4-1:0] node20604;
	wire [4-1:0] node20605;
	wire [4-1:0] node20606;
	wire [4-1:0] node20610;
	wire [4-1:0] node20611;
	wire [4-1:0] node20612;
	wire [4-1:0] node20615;
	wire [4-1:0] node20619;
	wire [4-1:0] node20620;
	wire [4-1:0] node20622;
	wire [4-1:0] node20626;
	wire [4-1:0] node20627;
	wire [4-1:0] node20628;
	wire [4-1:0] node20629;
	wire [4-1:0] node20630;
	wire [4-1:0] node20633;
	wire [4-1:0] node20635;
	wire [4-1:0] node20636;
	wire [4-1:0] node20640;
	wire [4-1:0] node20641;
	wire [4-1:0] node20642;
	wire [4-1:0] node20644;
	wire [4-1:0] node20647;
	wire [4-1:0] node20650;
	wire [4-1:0] node20651;
	wire [4-1:0] node20652;
	wire [4-1:0] node20655;
	wire [4-1:0] node20658;
	wire [4-1:0] node20660;
	wire [4-1:0] node20663;
	wire [4-1:0] node20664;
	wire [4-1:0] node20665;
	wire [4-1:0] node20666;
	wire [4-1:0] node20667;
	wire [4-1:0] node20668;
	wire [4-1:0] node20673;
	wire [4-1:0] node20674;
	wire [4-1:0] node20675;
	wire [4-1:0] node20680;
	wire [4-1:0] node20681;
	wire [4-1:0] node20683;
	wire [4-1:0] node20686;
	wire [4-1:0] node20687;
	wire [4-1:0] node20690;
	wire [4-1:0] node20692;
	wire [4-1:0] node20695;
	wire [4-1:0] node20696;
	wire [4-1:0] node20697;
	wire [4-1:0] node20699;
	wire [4-1:0] node20702;
	wire [4-1:0] node20703;
	wire [4-1:0] node20707;
	wire [4-1:0] node20710;
	wire [4-1:0] node20711;
	wire [4-1:0] node20712;
	wire [4-1:0] node20713;
	wire [4-1:0] node20714;
	wire [4-1:0] node20717;
	wire [4-1:0] node20718;
	wire [4-1:0] node20720;
	wire [4-1:0] node20724;
	wire [4-1:0] node20725;
	wire [4-1:0] node20728;
	wire [4-1:0] node20730;
	wire [4-1:0] node20733;
	wire [4-1:0] node20734;
	wire [4-1:0] node20735;
	wire [4-1:0] node20737;
	wire [4-1:0] node20738;
	wire [4-1:0] node20741;
	wire [4-1:0] node20744;
	wire [4-1:0] node20745;
	wire [4-1:0] node20747;
	wire [4-1:0] node20751;
	wire [4-1:0] node20752;
	wire [4-1:0] node20753;
	wire [4-1:0] node20757;
	wire [4-1:0] node20758;
	wire [4-1:0] node20762;
	wire [4-1:0] node20763;
	wire [4-1:0] node20764;
	wire [4-1:0] node20765;
	wire [4-1:0] node20766;
	wire [4-1:0] node20769;
	wire [4-1:0] node20772;
	wire [4-1:0] node20774;
	wire [4-1:0] node20776;
	wire [4-1:0] node20779;
	wire [4-1:0] node20780;
	wire [4-1:0] node20781;
	wire [4-1:0] node20782;
	wire [4-1:0] node20786;
	wire [4-1:0] node20787;
	wire [4-1:0] node20792;
	wire [4-1:0] node20793;
	wire [4-1:0] node20794;
	wire [4-1:0] node20795;
	wire [4-1:0] node20798;
	wire [4-1:0] node20800;
	wire [4-1:0] node20803;
	wire [4-1:0] node20805;
	wire [4-1:0] node20808;
	wire [4-1:0] node20809;
	wire [4-1:0] node20810;
	wire [4-1:0] node20813;
	wire [4-1:0] node20815;
	wire [4-1:0] node20818;
	wire [4-1:0] node20819;
	wire [4-1:0] node20822;
	wire [4-1:0] node20825;
	wire [4-1:0] node20826;
	wire [4-1:0] node20827;
	wire [4-1:0] node20828;
	wire [4-1:0] node20829;
	wire [4-1:0] node20830;
	wire [4-1:0] node20831;
	wire [4-1:0] node20832;
	wire [4-1:0] node20833;
	wire [4-1:0] node20837;
	wire [4-1:0] node20839;
	wire [4-1:0] node20842;
	wire [4-1:0] node20843;
	wire [4-1:0] node20845;
	wire [4-1:0] node20848;
	wire [4-1:0] node20849;
	wire [4-1:0] node20850;
	wire [4-1:0] node20853;
	wire [4-1:0] node20856;
	wire [4-1:0] node20859;
	wire [4-1:0] node20860;
	wire [4-1:0] node20861;
	wire [4-1:0] node20863;
	wire [4-1:0] node20865;
	wire [4-1:0] node20868;
	wire [4-1:0] node20869;
	wire [4-1:0] node20870;
	wire [4-1:0] node20871;
	wire [4-1:0] node20876;
	wire [4-1:0] node20877;
	wire [4-1:0] node20880;
	wire [4-1:0] node20883;
	wire [4-1:0] node20884;
	wire [4-1:0] node20885;
	wire [4-1:0] node20886;
	wire [4-1:0] node20890;
	wire [4-1:0] node20892;
	wire [4-1:0] node20895;
	wire [4-1:0] node20896;
	wire [4-1:0] node20897;
	wire [4-1:0] node20902;
	wire [4-1:0] node20903;
	wire [4-1:0] node20904;
	wire [4-1:0] node20905;
	wire [4-1:0] node20906;
	wire [4-1:0] node20908;
	wire [4-1:0] node20912;
	wire [4-1:0] node20913;
	wire [4-1:0] node20915;
	wire [4-1:0] node20917;
	wire [4-1:0] node20921;
	wire [4-1:0] node20922;
	wire [4-1:0] node20925;
	wire [4-1:0] node20928;
	wire [4-1:0] node20929;
	wire [4-1:0] node20930;
	wire [4-1:0] node20931;
	wire [4-1:0] node20932;
	wire [4-1:0] node20934;
	wire [4-1:0] node20937;
	wire [4-1:0] node20939;
	wire [4-1:0] node20943;
	wire [4-1:0] node20944;
	wire [4-1:0] node20945;
	wire [4-1:0] node20949;
	wire [4-1:0] node20950;
	wire [4-1:0] node20954;
	wire [4-1:0] node20955;
	wire [4-1:0] node20956;
	wire [4-1:0] node20958;
	wire [4-1:0] node20961;
	wire [4-1:0] node20963;
	wire [4-1:0] node20966;
	wire [4-1:0] node20967;
	wire [4-1:0] node20970;
	wire [4-1:0] node20972;
	wire [4-1:0] node20974;
	wire [4-1:0] node20977;
	wire [4-1:0] node20978;
	wire [4-1:0] node20979;
	wire [4-1:0] node20980;
	wire [4-1:0] node20981;
	wire [4-1:0] node20983;
	wire [4-1:0] node20985;
	wire [4-1:0] node20988;
	wire [4-1:0] node20989;
	wire [4-1:0] node20990;
	wire [4-1:0] node20991;
	wire [4-1:0] node20995;
	wire [4-1:0] node20997;
	wire [4-1:0] node21000;
	wire [4-1:0] node21003;
	wire [4-1:0] node21004;
	wire [4-1:0] node21006;
	wire [4-1:0] node21007;
	wire [4-1:0] node21008;
	wire [4-1:0] node21011;
	wire [4-1:0] node21014;
	wire [4-1:0] node21016;
	wire [4-1:0] node21019;
	wire [4-1:0] node21020;
	wire [4-1:0] node21021;
	wire [4-1:0] node21023;
	wire [4-1:0] node21027;
	wire [4-1:0] node21028;
	wire [4-1:0] node21030;
	wire [4-1:0] node21033;
	wire [4-1:0] node21034;
	wire [4-1:0] node21038;
	wire [4-1:0] node21039;
	wire [4-1:0] node21040;
	wire [4-1:0] node21041;
	wire [4-1:0] node21042;
	wire [4-1:0] node21044;
	wire [4-1:0] node21048;
	wire [4-1:0] node21050;
	wire [4-1:0] node21053;
	wire [4-1:0] node21054;
	wire [4-1:0] node21055;
	wire [4-1:0] node21058;
	wire [4-1:0] node21061;
	wire [4-1:0] node21064;
	wire [4-1:0] node21065;
	wire [4-1:0] node21066;
	wire [4-1:0] node21069;
	wire [4-1:0] node21070;
	wire [4-1:0] node21071;
	wire [4-1:0] node21075;
	wire [4-1:0] node21078;
	wire [4-1:0] node21079;
	wire [4-1:0] node21080;
	wire [4-1:0] node21083;
	wire [4-1:0] node21086;
	wire [4-1:0] node21087;
	wire [4-1:0] node21089;
	wire [4-1:0] node21093;
	wire [4-1:0] node21094;
	wire [4-1:0] node21095;
	wire [4-1:0] node21096;
	wire [4-1:0] node21097;
	wire [4-1:0] node21098;
	wire [4-1:0] node21102;
	wire [4-1:0] node21103;
	wire [4-1:0] node21104;
	wire [4-1:0] node21107;
	wire [4-1:0] node21110;
	wire [4-1:0] node21113;
	wire [4-1:0] node21114;
	wire [4-1:0] node21115;
	wire [4-1:0] node21118;
	wire [4-1:0] node21121;
	wire [4-1:0] node21123;
	wire [4-1:0] node21124;
	wire [4-1:0] node21128;
	wire [4-1:0] node21129;
	wire [4-1:0] node21130;
	wire [4-1:0] node21132;
	wire [4-1:0] node21134;
	wire [4-1:0] node21138;
	wire [4-1:0] node21140;
	wire [4-1:0] node21142;
	wire [4-1:0] node21145;
	wire [4-1:0] node21146;
	wire [4-1:0] node21147;
	wire [4-1:0] node21148;
	wire [4-1:0] node21150;
	wire [4-1:0] node21153;
	wire [4-1:0] node21156;
	wire [4-1:0] node21157;
	wire [4-1:0] node21158;
	wire [4-1:0] node21159;
	wire [4-1:0] node21165;
	wire [4-1:0] node21166;
	wire [4-1:0] node21167;
	wire [4-1:0] node21168;
	wire [4-1:0] node21169;
	wire [4-1:0] node21173;
	wire [4-1:0] node21176;
	wire [4-1:0] node21177;
	wire [4-1:0] node21180;
	wire [4-1:0] node21182;
	wire [4-1:0] node21185;
	wire [4-1:0] node21186;
	wire [4-1:0] node21187;
	wire [4-1:0] node21190;
	wire [4-1:0] node21193;
	wire [4-1:0] node21194;
	wire [4-1:0] node21198;
	wire [4-1:0] node21199;
	wire [4-1:0] node21200;
	wire [4-1:0] node21201;
	wire [4-1:0] node21202;
	wire [4-1:0] node21203;
	wire [4-1:0] node21204;
	wire [4-1:0] node21207;
	wire [4-1:0] node21210;
	wire [4-1:0] node21212;
	wire [4-1:0] node21213;
	wire [4-1:0] node21217;
	wire [4-1:0] node21218;
	wire [4-1:0] node21219;
	wire [4-1:0] node21221;
	wire [4-1:0] node21225;
	wire [4-1:0] node21226;
	wire [4-1:0] node21229;
	wire [4-1:0] node21232;
	wire [4-1:0] node21233;
	wire [4-1:0] node21234;
	wire [4-1:0] node21235;
	wire [4-1:0] node21237;
	wire [4-1:0] node21240;
	wire [4-1:0] node21243;
	wire [4-1:0] node21245;
	wire [4-1:0] node21247;
	wire [4-1:0] node21250;
	wire [4-1:0] node21251;
	wire [4-1:0] node21252;
	wire [4-1:0] node21254;
	wire [4-1:0] node21255;
	wire [4-1:0] node21258;
	wire [4-1:0] node21261;
	wire [4-1:0] node21263;
	wire [4-1:0] node21265;
	wire [4-1:0] node21268;
	wire [4-1:0] node21270;
	wire [4-1:0] node21273;
	wire [4-1:0] node21274;
	wire [4-1:0] node21275;
	wire [4-1:0] node21276;
	wire [4-1:0] node21278;
	wire [4-1:0] node21279;
	wire [4-1:0] node21282;
	wire [4-1:0] node21284;
	wire [4-1:0] node21287;
	wire [4-1:0] node21288;
	wire [4-1:0] node21289;
	wire [4-1:0] node21290;
	wire [4-1:0] node21295;
	wire [4-1:0] node21297;
	wire [4-1:0] node21299;
	wire [4-1:0] node21302;
	wire [4-1:0] node21303;
	wire [4-1:0] node21304;
	wire [4-1:0] node21308;
	wire [4-1:0] node21310;
	wire [4-1:0] node21311;
	wire [4-1:0] node21312;
	wire [4-1:0] node21316;
	wire [4-1:0] node21319;
	wire [4-1:0] node21320;
	wire [4-1:0] node21321;
	wire [4-1:0] node21322;
	wire [4-1:0] node21325;
	wire [4-1:0] node21328;
	wire [4-1:0] node21330;
	wire [4-1:0] node21331;
	wire [4-1:0] node21334;
	wire [4-1:0] node21337;
	wire [4-1:0] node21338;
	wire [4-1:0] node21339;
	wire [4-1:0] node21342;
	wire [4-1:0] node21345;
	wire [4-1:0] node21346;
	wire [4-1:0] node21347;
	wire [4-1:0] node21350;
	wire [4-1:0] node21353;
	wire [4-1:0] node21354;
	wire [4-1:0] node21358;
	wire [4-1:0] node21359;
	wire [4-1:0] node21360;
	wire [4-1:0] node21361;
	wire [4-1:0] node21362;
	wire [4-1:0] node21363;
	wire [4-1:0] node21366;
	wire [4-1:0] node21369;
	wire [4-1:0] node21370;
	wire [4-1:0] node21372;
	wire [4-1:0] node21375;
	wire [4-1:0] node21376;
	wire [4-1:0] node21378;
	wire [4-1:0] node21382;
	wire [4-1:0] node21383;
	wire [4-1:0] node21385;
	wire [4-1:0] node21388;
	wire [4-1:0] node21389;
	wire [4-1:0] node21392;
	wire [4-1:0] node21395;
	wire [4-1:0] node21396;
	wire [4-1:0] node21397;
	wire [4-1:0] node21398;
	wire [4-1:0] node21399;
	wire [4-1:0] node21400;
	wire [4-1:0] node21403;
	wire [4-1:0] node21407;
	wire [4-1:0] node21408;
	wire [4-1:0] node21411;
	wire [4-1:0] node21414;
	wire [4-1:0] node21415;
	wire [4-1:0] node21417;
	wire [4-1:0] node21418;
	wire [4-1:0] node21423;
	wire [4-1:0] node21424;
	wire [4-1:0] node21425;
	wire [4-1:0] node21427;
	wire [4-1:0] node21428;
	wire [4-1:0] node21432;
	wire [4-1:0] node21434;
	wire [4-1:0] node21437;
	wire [4-1:0] node21438;
	wire [4-1:0] node21441;
	wire [4-1:0] node21442;
	wire [4-1:0] node21444;
	wire [4-1:0] node21448;
	wire [4-1:0] node21449;
	wire [4-1:0] node21450;
	wire [4-1:0] node21453;
	wire [4-1:0] node21456;
	wire [4-1:0] node21457;
	wire [4-1:0] node21458;
	wire [4-1:0] node21460;
	wire [4-1:0] node21463;
	wire [4-1:0] node21464;
	wire [4-1:0] node21465;
	wire [4-1:0] node21466;
	wire [4-1:0] node21471;
	wire [4-1:0] node21472;
	wire [4-1:0] node21476;
	wire [4-1:0] node21477;
	wire [4-1:0] node21478;
	wire [4-1:0] node21479;
	wire [4-1:0] node21482;
	wire [4-1:0] node21485;
	wire [4-1:0] node21487;
	wire [4-1:0] node21490;
	wire [4-1:0] node21491;
	wire [4-1:0] node21493;
	wire [4-1:0] node21496;
	wire [4-1:0] node21497;
	wire [4-1:0] node21500;
	wire [4-1:0] node21501;
	wire [4-1:0] node21505;
	wire [4-1:0] node21506;
	wire [4-1:0] node21507;
	wire [4-1:0] node21508;
	wire [4-1:0] node21509;
	wire [4-1:0] node21510;
	wire [4-1:0] node21511;
	wire [4-1:0] node21512;
	wire [4-1:0] node21513;
	wire [4-1:0] node21514;
	wire [4-1:0] node21517;
	wire [4-1:0] node21522;
	wire [4-1:0] node21524;
	wire [4-1:0] node21527;
	wire [4-1:0] node21528;
	wire [4-1:0] node21531;
	wire [4-1:0] node21532;
	wire [4-1:0] node21536;
	wire [4-1:0] node21537;
	wire [4-1:0] node21538;
	wire [4-1:0] node21539;
	wire [4-1:0] node21540;
	wire [4-1:0] node21541;
	wire [4-1:0] node21544;
	wire [4-1:0] node21549;
	wire [4-1:0] node21550;
	wire [4-1:0] node21552;
	wire [4-1:0] node21553;
	wire [4-1:0] node21557;
	wire [4-1:0] node21558;
	wire [4-1:0] node21559;
	wire [4-1:0] node21564;
	wire [4-1:0] node21565;
	wire [4-1:0] node21567;
	wire [4-1:0] node21570;
	wire [4-1:0] node21571;
	wire [4-1:0] node21573;
	wire [4-1:0] node21576;
	wire [4-1:0] node21578;
	wire [4-1:0] node21581;
	wire [4-1:0] node21582;
	wire [4-1:0] node21583;
	wire [4-1:0] node21584;
	wire [4-1:0] node21585;
	wire [4-1:0] node21586;
	wire [4-1:0] node21587;
	wire [4-1:0] node21592;
	wire [4-1:0] node21593;
	wire [4-1:0] node21594;
	wire [4-1:0] node21599;
	wire [4-1:0] node21600;
	wire [4-1:0] node21601;
	wire [4-1:0] node21602;
	wire [4-1:0] node21607;
	wire [4-1:0] node21608;
	wire [4-1:0] node21611;
	wire [4-1:0] node21614;
	wire [4-1:0] node21615;
	wire [4-1:0] node21617;
	wire [4-1:0] node21620;
	wire [4-1:0] node21621;
	wire [4-1:0] node21622;
	wire [4-1:0] node21627;
	wire [4-1:0] node21628;
	wire [4-1:0] node21629;
	wire [4-1:0] node21631;
	wire [4-1:0] node21632;
	wire [4-1:0] node21635;
	wire [4-1:0] node21638;
	wire [4-1:0] node21640;
	wire [4-1:0] node21643;
	wire [4-1:0] node21644;
	wire [4-1:0] node21645;
	wire [4-1:0] node21647;
	wire [4-1:0] node21650;
	wire [4-1:0] node21651;
	wire [4-1:0] node21654;
	wire [4-1:0] node21657;
	wire [4-1:0] node21658;
	wire [4-1:0] node21661;
	wire [4-1:0] node21664;
	wire [4-1:0] node21665;
	wire [4-1:0] node21666;
	wire [4-1:0] node21667;
	wire [4-1:0] node21668;
	wire [4-1:0] node21669;
	wire [4-1:0] node21673;
	wire [4-1:0] node21674;
	wire [4-1:0] node21676;
	wire [4-1:0] node21678;
	wire [4-1:0] node21681;
	wire [4-1:0] node21684;
	wire [4-1:0] node21685;
	wire [4-1:0] node21686;
	wire [4-1:0] node21687;
	wire [4-1:0] node21688;
	wire [4-1:0] node21692;
	wire [4-1:0] node21696;
	wire [4-1:0] node21697;
	wire [4-1:0] node21698;
	wire [4-1:0] node21700;
	wire [4-1:0] node21704;
	wire [4-1:0] node21705;
	wire [4-1:0] node21709;
	wire [4-1:0] node21710;
	wire [4-1:0] node21711;
	wire [4-1:0] node21712;
	wire [4-1:0] node21713;
	wire [4-1:0] node21716;
	wire [4-1:0] node21717;
	wire [4-1:0] node21722;
	wire [4-1:0] node21723;
	wire [4-1:0] node21727;
	wire [4-1:0] node21728;
	wire [4-1:0] node21729;
	wire [4-1:0] node21730;
	wire [4-1:0] node21733;
	wire [4-1:0] node21737;
	wire [4-1:0] node21738;
	wire [4-1:0] node21742;
	wire [4-1:0] node21743;
	wire [4-1:0] node21744;
	wire [4-1:0] node21745;
	wire [4-1:0] node21746;
	wire [4-1:0] node21748;
	wire [4-1:0] node21751;
	wire [4-1:0] node21752;
	wire [4-1:0] node21756;
	wire [4-1:0] node21759;
	wire [4-1:0] node21761;
	wire [4-1:0] node21763;
	wire [4-1:0] node21766;
	wire [4-1:0] node21767;
	wire [4-1:0] node21768;
	wire [4-1:0] node21771;
	wire [4-1:0] node21773;
	wire [4-1:0] node21776;
	wire [4-1:0] node21777;
	wire [4-1:0] node21778;
	wire [4-1:0] node21781;
	wire [4-1:0] node21782;
	wire [4-1:0] node21786;
	wire [4-1:0] node21787;
	wire [4-1:0] node21788;
	wire [4-1:0] node21789;
	wire [4-1:0] node21793;
	wire [4-1:0] node21796;
	wire [4-1:0] node21797;
	wire [4-1:0] node21801;
	wire [4-1:0] node21802;
	wire [4-1:0] node21803;
	wire [4-1:0] node21804;
	wire [4-1:0] node21805;
	wire [4-1:0] node21806;
	wire [4-1:0] node21807;
	wire [4-1:0] node21808;
	wire [4-1:0] node21810;
	wire [4-1:0] node21814;
	wire [4-1:0] node21816;
	wire [4-1:0] node21817;
	wire [4-1:0] node21820;
	wire [4-1:0] node21823;
	wire [4-1:0] node21824;
	wire [4-1:0] node21827;
	wire [4-1:0] node21830;
	wire [4-1:0] node21831;
	wire [4-1:0] node21832;
	wire [4-1:0] node21836;
	wire [4-1:0] node21837;
	wire [4-1:0] node21838;
	wire [4-1:0] node21841;
	wire [4-1:0] node21844;
	wire [4-1:0] node21845;
	wire [4-1:0] node21846;
	wire [4-1:0] node21851;
	wire [4-1:0] node21852;
	wire [4-1:0] node21853;
	wire [4-1:0] node21854;
	wire [4-1:0] node21856;
	wire [4-1:0] node21857;
	wire [4-1:0] node21861;
	wire [4-1:0] node21862;
	wire [4-1:0] node21866;
	wire [4-1:0] node21867;
	wire [4-1:0] node21868;
	wire [4-1:0] node21873;
	wire [4-1:0] node21874;
	wire [4-1:0] node21876;
	wire [4-1:0] node21878;
	wire [4-1:0] node21879;
	wire [4-1:0] node21883;
	wire [4-1:0] node21884;
	wire [4-1:0] node21885;
	wire [4-1:0] node21888;
	wire [4-1:0] node21891;
	wire [4-1:0] node21892;
	wire [4-1:0] node21896;
	wire [4-1:0] node21897;
	wire [4-1:0] node21898;
	wire [4-1:0] node21899;
	wire [4-1:0] node21900;
	wire [4-1:0] node21902;
	wire [4-1:0] node21905;
	wire [4-1:0] node21906;
	wire [4-1:0] node21907;
	wire [4-1:0] node21910;
	wire [4-1:0] node21914;
	wire [4-1:0] node21916;
	wire [4-1:0] node21917;
	wire [4-1:0] node21919;
	wire [4-1:0] node21923;
	wire [4-1:0] node21924;
	wire [4-1:0] node21925;
	wire [4-1:0] node21926;
	wire [4-1:0] node21927;
	wire [4-1:0] node21932;
	wire [4-1:0] node21936;
	wire [4-1:0] node21937;
	wire [4-1:0] node21938;
	wire [4-1:0] node21939;
	wire [4-1:0] node21940;
	wire [4-1:0] node21943;
	wire [4-1:0] node21946;
	wire [4-1:0] node21949;
	wire [4-1:0] node21950;
	wire [4-1:0] node21952;
	wire [4-1:0] node21955;
	wire [4-1:0] node21956;
	wire [4-1:0] node21959;
	wire [4-1:0] node21962;
	wire [4-1:0] node21963;
	wire [4-1:0] node21964;
	wire [4-1:0] node21968;
	wire [4-1:0] node21969;
	wire [4-1:0] node21970;
	wire [4-1:0] node21974;
	wire [4-1:0] node21975;
	wire [4-1:0] node21979;
	wire [4-1:0] node21980;
	wire [4-1:0] node21981;
	wire [4-1:0] node21982;
	wire [4-1:0] node21983;
	wire [4-1:0] node21987;
	wire [4-1:0] node21988;
	wire [4-1:0] node21993;
	wire [4-1:0] node21994;
	wire [4-1:0] node21995;
	wire [4-1:0] node21996;
	wire [4-1:0] node22000;
	wire [4-1:0] node22001;
	wire [4-1:0] node22006;
	wire [4-1:0] node22007;
	wire [4-1:0] node22008;
	wire [4-1:0] node22009;
	wire [4-1:0] node22010;
	wire [4-1:0] node22011;
	wire [4-1:0] node22012;
	wire [4-1:0] node22013;
	wire [4-1:0] node22014;
	wire [4-1:0] node22015;
	wire [4-1:0] node22018;
	wire [4-1:0] node22019;
	wire [4-1:0] node22023;
	wire [4-1:0] node22024;
	wire [4-1:0] node22025;
	wire [4-1:0] node22027;
	wire [4-1:0] node22031;
	wire [4-1:0] node22032;
	wire [4-1:0] node22035;
	wire [4-1:0] node22036;
	wire [4-1:0] node22040;
	wire [4-1:0] node22041;
	wire [4-1:0] node22042;
	wire [4-1:0] node22044;
	wire [4-1:0] node22045;
	wire [4-1:0] node22049;
	wire [4-1:0] node22050;
	wire [4-1:0] node22053;
	wire [4-1:0] node22056;
	wire [4-1:0] node22057;
	wire [4-1:0] node22058;
	wire [4-1:0] node22061;
	wire [4-1:0] node22064;
	wire [4-1:0] node22065;
	wire [4-1:0] node22066;
	wire [4-1:0] node22071;
	wire [4-1:0] node22072;
	wire [4-1:0] node22073;
	wire [4-1:0] node22076;
	wire [4-1:0] node22077;
	wire [4-1:0] node22079;
	wire [4-1:0] node22082;
	wire [4-1:0] node22083;
	wire [4-1:0] node22087;
	wire [4-1:0] node22088;
	wire [4-1:0] node22089;
	wire [4-1:0] node22092;
	wire [4-1:0] node22094;
	wire [4-1:0] node22097;
	wire [4-1:0] node22100;
	wire [4-1:0] node22101;
	wire [4-1:0] node22102;
	wire [4-1:0] node22103;
	wire [4-1:0] node22104;
	wire [4-1:0] node22105;
	wire [4-1:0] node22108;
	wire [4-1:0] node22110;
	wire [4-1:0] node22113;
	wire [4-1:0] node22114;
	wire [4-1:0] node22118;
	wire [4-1:0] node22119;
	wire [4-1:0] node22122;
	wire [4-1:0] node22124;
	wire [4-1:0] node22127;
	wire [4-1:0] node22128;
	wire [4-1:0] node22129;
	wire [4-1:0] node22131;
	wire [4-1:0] node22132;
	wire [4-1:0] node22136;
	wire [4-1:0] node22138;
	wire [4-1:0] node22139;
	wire [4-1:0] node22143;
	wire [4-1:0] node22144;
	wire [4-1:0] node22146;
	wire [4-1:0] node22149;
	wire [4-1:0] node22150;
	wire [4-1:0] node22151;
	wire [4-1:0] node22154;
	wire [4-1:0] node22158;
	wire [4-1:0] node22159;
	wire [4-1:0] node22160;
	wire [4-1:0] node22161;
	wire [4-1:0] node22162;
	wire [4-1:0] node22165;
	wire [4-1:0] node22166;
	wire [4-1:0] node22171;
	wire [4-1:0] node22174;
	wire [4-1:0] node22175;
	wire [4-1:0] node22176;
	wire [4-1:0] node22177;
	wire [4-1:0] node22181;
	wire [4-1:0] node22182;
	wire [4-1:0] node22186;
	wire [4-1:0] node22187;
	wire [4-1:0] node22188;
	wire [4-1:0] node22189;
	wire [4-1:0] node22195;
	wire [4-1:0] node22196;
	wire [4-1:0] node22197;
	wire [4-1:0] node22198;
	wire [4-1:0] node22199;
	wire [4-1:0] node22200;
	wire [4-1:0] node22201;
	wire [4-1:0] node22203;
	wire [4-1:0] node22207;
	wire [4-1:0] node22208;
	wire [4-1:0] node22209;
	wire [4-1:0] node22213;
	wire [4-1:0] node22215;
	wire [4-1:0] node22218;
	wire [4-1:0] node22219;
	wire [4-1:0] node22220;
	wire [4-1:0] node22221;
	wire [4-1:0] node22224;
	wire [4-1:0] node22229;
	wire [4-1:0] node22230;
	wire [4-1:0] node22231;
	wire [4-1:0] node22232;
	wire [4-1:0] node22234;
	wire [4-1:0] node22237;
	wire [4-1:0] node22238;
	wire [4-1:0] node22243;
	wire [4-1:0] node22244;
	wire [4-1:0] node22247;
	wire [4-1:0] node22248;
	wire [4-1:0] node22250;
	wire [4-1:0] node22254;
	wire [4-1:0] node22255;
	wire [4-1:0] node22256;
	wire [4-1:0] node22257;
	wire [4-1:0] node22258;
	wire [4-1:0] node22261;
	wire [4-1:0] node22265;
	wire [4-1:0] node22266;
	wire [4-1:0] node22269;
	wire [4-1:0] node22270;
	wire [4-1:0] node22274;
	wire [4-1:0] node22275;
	wire [4-1:0] node22276;
	wire [4-1:0] node22279;
	wire [4-1:0] node22280;
	wire [4-1:0] node22281;
	wire [4-1:0] node22284;
	wire [4-1:0] node22288;
	wire [4-1:0] node22289;
	wire [4-1:0] node22290;
	wire [4-1:0] node22292;
	wire [4-1:0] node22296;
	wire [4-1:0] node22299;
	wire [4-1:0] node22300;
	wire [4-1:0] node22301;
	wire [4-1:0] node22302;
	wire [4-1:0] node22303;
	wire [4-1:0] node22306;
	wire [4-1:0] node22309;
	wire [4-1:0] node22310;
	wire [4-1:0] node22311;
	wire [4-1:0] node22314;
	wire [4-1:0] node22316;
	wire [4-1:0] node22320;
	wire [4-1:0] node22321;
	wire [4-1:0] node22322;
	wire [4-1:0] node22323;
	wire [4-1:0] node22327;
	wire [4-1:0] node22328;
	wire [4-1:0] node22329;
	wire [4-1:0] node22334;
	wire [4-1:0] node22336;
	wire [4-1:0] node22339;
	wire [4-1:0] node22340;
	wire [4-1:0] node22341;
	wire [4-1:0] node22342;
	wire [4-1:0] node22343;
	wire [4-1:0] node22344;
	wire [4-1:0] node22350;
	wire [4-1:0] node22351;
	wire [4-1:0] node22355;
	wire [4-1:0] node22356;
	wire [4-1:0] node22357;
	wire [4-1:0] node22358;
	wire [4-1:0] node22360;
	wire [4-1:0] node22363;
	wire [4-1:0] node22364;
	wire [4-1:0] node22368;
	wire [4-1:0] node22370;
	wire [4-1:0] node22374;
	wire [4-1:0] node22375;
	wire [4-1:0] node22376;
	wire [4-1:0] node22377;
	wire [4-1:0] node22378;
	wire [4-1:0] node22379;
	wire [4-1:0] node22382;
	wire [4-1:0] node22385;
	wire [4-1:0] node22386;
	wire [4-1:0] node22387;
	wire [4-1:0] node22388;
	wire [4-1:0] node22392;
	wire [4-1:0] node22395;
	wire [4-1:0] node22398;
	wire [4-1:0] node22399;
	wire [4-1:0] node22400;
	wire [4-1:0] node22401;
	wire [4-1:0] node22405;
	wire [4-1:0] node22406;
	wire [4-1:0] node22407;
	wire [4-1:0] node22408;
	wire [4-1:0] node22412;
	wire [4-1:0] node22413;
	wire [4-1:0] node22416;
	wire [4-1:0] node22420;
	wire [4-1:0] node22421;
	wire [4-1:0] node22423;
	wire [4-1:0] node22424;
	wire [4-1:0] node22428;
	wire [4-1:0] node22430;
	wire [4-1:0] node22432;
	wire [4-1:0] node22435;
	wire [4-1:0] node22436;
	wire [4-1:0] node22437;
	wire [4-1:0] node22438;
	wire [4-1:0] node22441;
	wire [4-1:0] node22442;
	wire [4-1:0] node22443;
	wire [4-1:0] node22444;
	wire [4-1:0] node22449;
	wire [4-1:0] node22452;
	wire [4-1:0] node22453;
	wire [4-1:0] node22454;
	wire [4-1:0] node22455;
	wire [4-1:0] node22459;
	wire [4-1:0] node22460;
	wire [4-1:0] node22463;
	wire [4-1:0] node22466;
	wire [4-1:0] node22467;
	wire [4-1:0] node22469;
	wire [4-1:0] node22470;
	wire [4-1:0] node22475;
	wire [4-1:0] node22476;
	wire [4-1:0] node22477;
	wire [4-1:0] node22478;
	wire [4-1:0] node22481;
	wire [4-1:0] node22483;
	wire [4-1:0] node22486;
	wire [4-1:0] node22487;
	wire [4-1:0] node22489;
	wire [4-1:0] node22493;
	wire [4-1:0] node22494;
	wire [4-1:0] node22497;
	wire [4-1:0] node22500;
	wire [4-1:0] node22501;
	wire [4-1:0] node22502;
	wire [4-1:0] node22503;
	wire [4-1:0] node22504;
	wire [4-1:0] node22505;
	wire [4-1:0] node22507;
	wire [4-1:0] node22510;
	wire [4-1:0] node22514;
	wire [4-1:0] node22516;
	wire [4-1:0] node22517;
	wire [4-1:0] node22518;
	wire [4-1:0] node22522;
	wire [4-1:0] node22523;
	wire [4-1:0] node22527;
	wire [4-1:0] node22528;
	wire [4-1:0] node22530;
	wire [4-1:0] node22531;
	wire [4-1:0] node22533;
	wire [4-1:0] node22537;
	wire [4-1:0] node22538;
	wire [4-1:0] node22539;
	wire [4-1:0] node22540;
	wire [4-1:0] node22541;
	wire [4-1:0] node22544;
	wire [4-1:0] node22548;
	wire [4-1:0] node22549;
	wire [4-1:0] node22553;
	wire [4-1:0] node22554;
	wire [4-1:0] node22555;
	wire [4-1:0] node22560;
	wire [4-1:0] node22561;
	wire [4-1:0] node22562;
	wire [4-1:0] node22563;
	wire [4-1:0] node22566;
	wire [4-1:0] node22567;
	wire [4-1:0] node22570;
	wire [4-1:0] node22571;
	wire [4-1:0] node22575;
	wire [4-1:0] node22576;
	wire [4-1:0] node22577;
	wire [4-1:0] node22579;
	wire [4-1:0] node22580;
	wire [4-1:0] node22584;
	wire [4-1:0] node22586;
	wire [4-1:0] node22589;
	wire [4-1:0] node22590;
	wire [4-1:0] node22593;
	wire [4-1:0] node22594;
	wire [4-1:0] node22598;
	wire [4-1:0] node22599;
	wire [4-1:0] node22600;
	wire [4-1:0] node22601;
	wire [4-1:0] node22605;
	wire [4-1:0] node22606;
	wire [4-1:0] node22607;
	wire [4-1:0] node22610;
	wire [4-1:0] node22613;
	wire [4-1:0] node22615;
	wire [4-1:0] node22618;
	wire [4-1:0] node22619;
	wire [4-1:0] node22620;
	wire [4-1:0] node22621;
	wire [4-1:0] node22624;
	wire [4-1:0] node22627;
	wire [4-1:0] node22628;
	wire [4-1:0] node22632;
	wire [4-1:0] node22634;
	wire [4-1:0] node22635;
	wire [4-1:0] node22636;
	wire [4-1:0] node22641;
	wire [4-1:0] node22642;
	wire [4-1:0] node22643;
	wire [4-1:0] node22644;
	wire [4-1:0] node22645;
	wire [4-1:0] node22646;
	wire [4-1:0] node22648;
	wire [4-1:0] node22651;
	wire [4-1:0] node22653;
	wire [4-1:0] node22656;
	wire [4-1:0] node22657;
	wire [4-1:0] node22659;
	wire [4-1:0] node22662;
	wire [4-1:0] node22664;
	wire [4-1:0] node22667;
	wire [4-1:0] node22668;
	wire [4-1:0] node22671;
	wire [4-1:0] node22674;
	wire [4-1:0] node22675;
	wire [4-1:0] node22676;
	wire [4-1:0] node22677;
	wire [4-1:0] node22678;
	wire [4-1:0] node22679;
	wire [4-1:0] node22682;
	wire [4-1:0] node22684;
	wire [4-1:0] node22685;
	wire [4-1:0] node22689;
	wire [4-1:0] node22690;
	wire [4-1:0] node22691;
	wire [4-1:0] node22695;
	wire [4-1:0] node22697;
	wire [4-1:0] node22700;
	wire [4-1:0] node22701;
	wire [4-1:0] node22702;
	wire [4-1:0] node22704;
	wire [4-1:0] node22707;
	wire [4-1:0] node22708;
	wire [4-1:0] node22710;
	wire [4-1:0] node22713;
	wire [4-1:0] node22716;
	wire [4-1:0] node22717;
	wire [4-1:0] node22718;
	wire [4-1:0] node22720;
	wire [4-1:0] node22723;
	wire [4-1:0] node22724;
	wire [4-1:0] node22728;
	wire [4-1:0] node22729;
	wire [4-1:0] node22733;
	wire [4-1:0] node22734;
	wire [4-1:0] node22735;
	wire [4-1:0] node22736;
	wire [4-1:0] node22740;
	wire [4-1:0] node22741;
	wire [4-1:0] node22745;
	wire [4-1:0] node22746;
	wire [4-1:0] node22747;
	wire [4-1:0] node22751;
	wire [4-1:0] node22752;
	wire [4-1:0] node22756;
	wire [4-1:0] node22757;
	wire [4-1:0] node22758;
	wire [4-1:0] node22759;
	wire [4-1:0] node22761;
	wire [4-1:0] node22762;
	wire [4-1:0] node22766;
	wire [4-1:0] node22767;
	wire [4-1:0] node22768;
	wire [4-1:0] node22772;
	wire [4-1:0] node22775;
	wire [4-1:0] node22776;
	wire [4-1:0] node22777;
	wire [4-1:0] node22780;
	wire [4-1:0] node22783;
	wire [4-1:0] node22784;
	wire [4-1:0] node22786;
	wire [4-1:0] node22789;
	wire [4-1:0] node22790;
	wire [4-1:0] node22791;
	wire [4-1:0] node22796;
	wire [4-1:0] node22797;
	wire [4-1:0] node22798;
	wire [4-1:0] node22800;
	wire [4-1:0] node22803;
	wire [4-1:0] node22804;
	wire [4-1:0] node22805;
	wire [4-1:0] node22810;
	wire [4-1:0] node22811;
	wire [4-1:0] node22812;
	wire [4-1:0] node22813;
	wire [4-1:0] node22817;
	wire [4-1:0] node22818;
	wire [4-1:0] node22822;
	wire [4-1:0] node22823;
	wire [4-1:0] node22827;
	wire [4-1:0] node22828;
	wire [4-1:0] node22829;
	wire [4-1:0] node22830;
	wire [4-1:0] node22831;
	wire [4-1:0] node22833;
	wire [4-1:0] node22836;
	wire [4-1:0] node22838;
	wire [4-1:0] node22841;
	wire [4-1:0] node22842;
	wire [4-1:0] node22844;
	wire [4-1:0] node22847;
	wire [4-1:0] node22849;
	wire [4-1:0] node22852;
	wire [4-1:0] node22853;
	wire [4-1:0] node22856;
	wire [4-1:0] node22859;
	wire [4-1:0] node22860;
	wire [4-1:0] node22861;
	wire [4-1:0] node22862;
	wire [4-1:0] node22863;
	wire [4-1:0] node22867;
	wire [4-1:0] node22868;
	wire [4-1:0] node22873;
	wire [4-1:0] node22874;
	wire [4-1:0] node22875;
	wire [4-1:0] node22876;
	wire [4-1:0] node22880;
	wire [4-1:0] node22881;
	wire [4-1:0] node22886;
	wire [4-1:0] node22887;
	wire [4-1:0] node22888;
	wire [4-1:0] node22889;
	wire [4-1:0] node22890;
	wire [4-1:0] node22891;
	wire [4-1:0] node22892;
	wire [4-1:0] node22893;
	wire [4-1:0] node22894;
	wire [4-1:0] node22895;
	wire [4-1:0] node22898;
	wire [4-1:0] node22901;
	wire [4-1:0] node22903;
	wire [4-1:0] node22906;
	wire [4-1:0] node22907;
	wire [4-1:0] node22909;
	wire [4-1:0] node22911;
	wire [4-1:0] node22914;
	wire [4-1:0] node22915;
	wire [4-1:0] node22917;
	wire [4-1:0] node22920;
	wire [4-1:0] node22921;
	wire [4-1:0] node22924;
	wire [4-1:0] node22927;
	wire [4-1:0] node22928;
	wire [4-1:0] node22929;
	wire [4-1:0] node22930;
	wire [4-1:0] node22934;
	wire [4-1:0] node22936;
	wire [4-1:0] node22937;
	wire [4-1:0] node22940;
	wire [4-1:0] node22943;
	wire [4-1:0] node22944;
	wire [4-1:0] node22945;
	wire [4-1:0] node22946;
	wire [4-1:0] node22951;
	wire [4-1:0] node22953;
	wire [4-1:0] node22956;
	wire [4-1:0] node22957;
	wire [4-1:0] node22958;
	wire [4-1:0] node22959;
	wire [4-1:0] node22960;
	wire [4-1:0] node22961;
	wire [4-1:0] node22964;
	wire [4-1:0] node22968;
	wire [4-1:0] node22969;
	wire [4-1:0] node22970;
	wire [4-1:0] node22973;
	wire [4-1:0] node22978;
	wire [4-1:0] node22979;
	wire [4-1:0] node22980;
	wire [4-1:0] node22982;
	wire [4-1:0] node22985;
	wire [4-1:0] node22987;
	wire [4-1:0] node22990;
	wire [4-1:0] node22992;
	wire [4-1:0] node22994;
	wire [4-1:0] node22996;
	wire [4-1:0] node22999;
	wire [4-1:0] node23000;
	wire [4-1:0] node23001;
	wire [4-1:0] node23002;
	wire [4-1:0] node23003;
	wire [4-1:0] node23007;
	wire [4-1:0] node23008;
	wire [4-1:0] node23010;
	wire [4-1:0] node23013;
	wire [4-1:0] node23015;
	wire [4-1:0] node23018;
	wire [4-1:0] node23019;
	wire [4-1:0] node23022;
	wire [4-1:0] node23023;
	wire [4-1:0] node23024;
	wire [4-1:0] node23028;
	wire [4-1:0] node23029;
	wire [4-1:0] node23031;
	wire [4-1:0] node23035;
	wire [4-1:0] node23036;
	wire [4-1:0] node23037;
	wire [4-1:0] node23038;
	wire [4-1:0] node23041;
	wire [4-1:0] node23043;
	wire [4-1:0] node23046;
	wire [4-1:0] node23047;
	wire [4-1:0] node23048;
	wire [4-1:0] node23050;
	wire [4-1:0] node23053;
	wire [4-1:0] node23055;
	wire [4-1:0] node23058;
	wire [4-1:0] node23060;
	wire [4-1:0] node23063;
	wire [4-1:0] node23064;
	wire [4-1:0] node23067;
	wire [4-1:0] node23070;
	wire [4-1:0] node23071;
	wire [4-1:0] node23072;
	wire [4-1:0] node23073;
	wire [4-1:0] node23074;
	wire [4-1:0] node23075;
	wire [4-1:0] node23078;
	wire [4-1:0] node23081;
	wire [4-1:0] node23082;
	wire [4-1:0] node23083;
	wire [4-1:0] node23086;
	wire [4-1:0] node23089;
	wire [4-1:0] node23090;
	wire [4-1:0] node23094;
	wire [4-1:0] node23095;
	wire [4-1:0] node23096;
	wire [4-1:0] node23099;
	wire [4-1:0] node23102;
	wire [4-1:0] node23104;
	wire [4-1:0] node23107;
	wire [4-1:0] node23108;
	wire [4-1:0] node23109;
	wire [4-1:0] node23110;
	wire [4-1:0] node23114;
	wire [4-1:0] node23115;
	wire [4-1:0] node23117;
	wire [4-1:0] node23120;
	wire [4-1:0] node23121;
	wire [4-1:0] node23125;
	wire [4-1:0] node23126;
	wire [4-1:0] node23127;
	wire [4-1:0] node23129;
	wire [4-1:0] node23132;
	wire [4-1:0] node23133;
	wire [4-1:0] node23136;
	wire [4-1:0] node23139;
	wire [4-1:0] node23140;
	wire [4-1:0] node23143;
	wire [4-1:0] node23146;
	wire [4-1:0] node23147;
	wire [4-1:0] node23148;
	wire [4-1:0] node23149;
	wire [4-1:0] node23152;
	wire [4-1:0] node23155;
	wire [4-1:0] node23156;
	wire [4-1:0] node23157;
	wire [4-1:0] node23158;
	wire [4-1:0] node23161;
	wire [4-1:0] node23164;
	wire [4-1:0] node23166;
	wire [4-1:0] node23170;
	wire [4-1:0] node23171;
	wire [4-1:0] node23174;
	wire [4-1:0] node23177;
	wire [4-1:0] node23178;
	wire [4-1:0] node23179;
	wire [4-1:0] node23180;
	wire [4-1:0] node23181;
	wire [4-1:0] node23182;
	wire [4-1:0] node23183;
	wire [4-1:0] node23186;
	wire [4-1:0] node23189;
	wire [4-1:0] node23191;
	wire [4-1:0] node23194;
	wire [4-1:0] node23195;
	wire [4-1:0] node23196;
	wire [4-1:0] node23199;
	wire [4-1:0] node23202;
	wire [4-1:0] node23203;
	wire [4-1:0] node23206;
	wire [4-1:0] node23209;
	wire [4-1:0] node23210;
	wire [4-1:0] node23213;
	wire [4-1:0] node23216;
	wire [4-1:0] node23217;
	wire [4-1:0] node23218;
	wire [4-1:0] node23219;
	wire [4-1:0] node23220;
	wire [4-1:0] node23221;
	wire [4-1:0] node23224;
	wire [4-1:0] node23227;
	wire [4-1:0] node23229;
	wire [4-1:0] node23232;
	wire [4-1:0] node23234;
	wire [4-1:0] node23236;
	wire [4-1:0] node23239;
	wire [4-1:0] node23240;
	wire [4-1:0] node23243;
	wire [4-1:0] node23246;
	wire [4-1:0] node23247;
	wire [4-1:0] node23250;
	wire [4-1:0] node23253;
	wire [4-1:0] node23254;
	wire [4-1:0] node23255;
	wire [4-1:0] node23259;
	wire [4-1:0] node23260;
	wire [4-1:0] node23264;
	wire [4-1:0] node23265;
	wire [4-1:0] node23266;
	wire [4-1:0] node23267;
	wire [4-1:0] node23268;
	wire [4-1:0] node23269;
	wire [4-1:0] node23270;
	wire [4-1:0] node23272;
	wire [4-1:0] node23275;
	wire [4-1:0] node23276;
	wire [4-1:0] node23279;
	wire [4-1:0] node23282;
	wire [4-1:0] node23283;
	wire [4-1:0] node23285;
	wire [4-1:0] node23288;
	wire [4-1:0] node23291;
	wire [4-1:0] node23292;
	wire [4-1:0] node23293;
	wire [4-1:0] node23297;
	wire [4-1:0] node23300;
	wire [4-1:0] node23301;
	wire [4-1:0] node23302;
	wire [4-1:0] node23303;
	wire [4-1:0] node23308;
	wire [4-1:0] node23309;
	wire [4-1:0] node23310;
	wire [4-1:0] node23315;
	wire [4-1:0] node23316;
	wire [4-1:0] node23317;
	wire [4-1:0] node23321;
	wire [4-1:0] node23322;
	wire [4-1:0] node23326;
	wire [4-1:0] node23327;
	wire [4-1:0] node23328;
	wire [4-1:0] node23329;
	wire [4-1:0] node23330;
	wire [4-1:0] node23331;
	wire [4-1:0] node23335;
	wire [4-1:0] node23336;
	wire [4-1:0] node23341;
	wire [4-1:0] node23342;
	wire [4-1:0] node23346;
	wire [4-1:0] node23347;
	wire [4-1:0] node23348;
	wire [4-1:0] node23349;
	wire [4-1:0] node23350;
	wire [4-1:0] node23355;
	wire [4-1:0] node23356;
	wire [4-1:0] node23357;

	assign outp = (inp[3]) ? node12656 : node1;
		assign node1 = (inp[6]) ? node7165 : node2;
			assign node2 = (inp[8]) ? node3708 : node3;
				assign node3 = (inp[14]) ? node1905 : node4;
					assign node4 = (inp[15]) ? node988 : node5;
						assign node5 = (inp[5]) ? node469 : node6;
							assign node6 = (inp[11]) ? node232 : node7;
								assign node7 = (inp[2]) ? node117 : node8;
									assign node8 = (inp[13]) ? node70 : node9;
										assign node9 = (inp[12]) ? node39 : node10;
											assign node10 = (inp[7]) ? node26 : node11;
												assign node11 = (inp[0]) ? node17 : node12;
													assign node12 = (inp[9]) ? node14 : 4'b0000;
														assign node14 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node17 = (inp[1]) ? node23 : node18;
														assign node18 = (inp[9]) ? node20 : 4'b0001;
															assign node20 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node23 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node26 = (inp[1]) ? node32 : node27;
													assign node27 = (inp[10]) ? 4'b0011 : node28;
														assign node28 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node32 = (inp[0]) ? node34 : 4'b0010;
														assign node34 = (inp[9]) ? 4'b0011 : node35;
															assign node35 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node39 = (inp[7]) ? node59 : node40;
												assign node40 = (inp[4]) ? node48 : node41;
													assign node41 = (inp[1]) ? 4'b0011 : node42;
														assign node42 = (inp[10]) ? 4'b0011 : node43;
															assign node43 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node48 = (inp[9]) ? node54 : node49;
														assign node49 = (inp[0]) ? node51 : 4'b0111;
															assign node51 = (inp[1]) ? 4'b0110 : 4'b0110;
														assign node54 = (inp[1]) ? 4'b0110 : node55;
															assign node55 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node59 = (inp[9]) ? node67 : node60;
													assign node60 = (inp[10]) ? node62 : 4'b0000;
														assign node62 = (inp[0]) ? 4'b0101 : node63;
															assign node63 = (inp[1]) ? 4'b0001 : 4'b0001;
													assign node67 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node70 = (inp[12]) ? node80 : node71;
											assign node71 = (inp[7]) ? node75 : node72;
												assign node72 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node75 = (inp[10]) ? node77 : 4'b0110;
													assign node77 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node80 = (inp[7]) ? node100 : node81;
												assign node81 = (inp[4]) ? node93 : node82;
													assign node82 = (inp[9]) ? node88 : node83;
														assign node83 = (inp[10]) ? node85 : 4'b0110;
															assign node85 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node88 = (inp[1]) ? 4'b0111 : node89;
															assign node89 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node93 = (inp[9]) ? 4'b0011 : node94;
														assign node94 = (inp[10]) ? node96 : 4'b0010;
															assign node96 = (inp[1]) ? 4'b0010 : 4'b0010;
												assign node100 = (inp[1]) ? node108 : node101;
													assign node101 = (inp[4]) ? 4'b0001 : node102;
														assign node102 = (inp[10]) ? node104 : 4'b0101;
															assign node104 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node108 = (inp[4]) ? node114 : node109;
														assign node109 = (inp[10]) ? 4'b0000 : node110;
															assign node110 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node114 = (inp[9]) ? 4'b0101 : 4'b0100;
									assign node117 = (inp[13]) ? node173 : node118;
										assign node118 = (inp[12]) ? node148 : node119;
											assign node119 = (inp[7]) ? node135 : node120;
												assign node120 = (inp[10]) ? node128 : node121;
													assign node121 = (inp[9]) ? node125 : node122;
														assign node122 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node125 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node128 = (inp[4]) ? node132 : node129;
														assign node129 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node132 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node135 = (inp[10]) ? 4'b0111 : node136;
													assign node136 = (inp[1]) ? node142 : node137;
														assign node137 = (inp[0]) ? 4'b0111 : node138;
															assign node138 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node142 = (inp[9]) ? 4'b0110 : node143;
															assign node143 = (inp[4]) ? 4'b0111 : 4'b0110;
											assign node148 = (inp[7]) ? node158 : node149;
												assign node149 = (inp[4]) ? node153 : node150;
													assign node150 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node153 = (inp[9]) ? node155 : 4'b0011;
														assign node155 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node158 = (inp[4]) ? node170 : node159;
													assign node159 = (inp[1]) ? node167 : node160;
														assign node160 = (inp[10]) ? node164 : node161;
															assign node161 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node164 = (inp[9]) ? 4'b0100 : 4'b0100;
														assign node167 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node170 = (inp[1]) ? 4'b0101 : 4'b0000;
										assign node173 = (inp[4]) ? node207 : node174;
											assign node174 = (inp[0]) ? node190 : node175;
												assign node175 = (inp[10]) ? node181 : node176;
													assign node176 = (inp[1]) ? node178 : 4'b0001;
														assign node178 = (inp[12]) ? 4'b0010 : 4'b0001;
													assign node181 = (inp[1]) ? 4'b0011 : node182;
														assign node182 = (inp[9]) ? node186 : node183;
															assign node183 = (inp[7]) ? 4'b0011 : 4'b0001;
															assign node186 = (inp[12]) ? 4'b0001 : 4'b0010;
												assign node190 = (inp[9]) ? node200 : node191;
													assign node191 = (inp[10]) ? node197 : node192;
														assign node192 = (inp[12]) ? 4'b0001 : node193;
															assign node193 = (inp[1]) ? 4'b0001 : 4'b0011;
														assign node197 = (inp[12]) ? 4'b0011 : 4'b0000;
													assign node200 = (inp[12]) ? 4'b0010 : node201;
														assign node201 = (inp[10]) ? 4'b0001 : node202;
															assign node202 = (inp[7]) ? 4'b0010 : 4'b0000;
											assign node207 = (inp[12]) ? node221 : node208;
												assign node208 = (inp[7]) ? node214 : node209;
													assign node209 = (inp[9]) ? 4'b0000 : node210;
														assign node210 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node214 = (inp[9]) ? 4'b0010 : node215;
														assign node215 = (inp[1]) ? 4'b0011 : node216;
															assign node216 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node221 = (inp[7]) ? node229 : node222;
													assign node222 = (inp[9]) ? node224 : 4'b0110;
														assign node224 = (inp[1]) ? node226 : 4'b0111;
															assign node226 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node229 = (inp[0]) ? 4'b0100 : 4'b0001;
								assign node232 = (inp[10]) ? node352 : node233;
									assign node233 = (inp[7]) ? node289 : node234;
										assign node234 = (inp[12]) ? node252 : node235;
											assign node235 = (inp[2]) ? node247 : node236;
												assign node236 = (inp[13]) ? node242 : node237;
													assign node237 = (inp[1]) ? node239 : 4'b0000;
														assign node239 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node242 = (inp[1]) ? node244 : 4'b0101;
														assign node244 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node247 = (inp[4]) ? node249 : 4'b0101;
													assign node249 = (inp[13]) ? 4'b0000 : 4'b0100;
											assign node252 = (inp[4]) ? node278 : node253;
												assign node253 = (inp[0]) ? node265 : node254;
													assign node254 = (inp[2]) ? node262 : node255;
														assign node255 = (inp[9]) ? node259 : node256;
															assign node256 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node259 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node262 = (inp[13]) ? 4'b0010 : 4'b0111;
													assign node265 = (inp[1]) ? node273 : node266;
														assign node266 = (inp[2]) ? node270 : node267;
															assign node267 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node270 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node273 = (inp[9]) ? node275 : 4'b0110;
															assign node275 = (inp[13]) ? 4'b0011 : 4'b0111;
												assign node278 = (inp[2]) ? node282 : node279;
													assign node279 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node282 = (inp[13]) ? 4'b0111 : node283;
														assign node283 = (inp[0]) ? 4'b0010 : node284;
															assign node284 = (inp[9]) ? 4'b0011 : 4'b0010;
										assign node289 = (inp[12]) ? node327 : node290;
											assign node290 = (inp[1]) ? node310 : node291;
												assign node291 = (inp[13]) ? node301 : node292;
													assign node292 = (inp[2]) ? node298 : node293;
														assign node293 = (inp[0]) ? 4'b0010 : node294;
															assign node294 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node298 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node301 = (inp[2]) ? 4'b0010 : node302;
														assign node302 = (inp[4]) ? node306 : node303;
															assign node303 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node306 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node310 = (inp[2]) ? node320 : node311;
													assign node311 = (inp[13]) ? 4'b0110 : node312;
														assign node312 = (inp[9]) ? node316 : node313;
															assign node313 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node316 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node320 = (inp[13]) ? node322 : 4'b0111;
														assign node322 = (inp[9]) ? 4'b0011 : node323;
															assign node323 = (inp[4]) ? 4'b0010 : 4'b0011;
											assign node327 = (inp[0]) ? node343 : node328;
												assign node328 = (inp[2]) ? node336 : node329;
													assign node329 = (inp[9]) ? node331 : 4'b0000;
														assign node331 = (inp[1]) ? node333 : 4'b0000;
															assign node333 = (inp[4]) ? 4'b0001 : 4'b0001;
													assign node336 = (inp[4]) ? 4'b0100 : node337;
														assign node337 = (inp[9]) ? 4'b0000 : node338;
															assign node338 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node343 = (inp[9]) ? node349 : node344;
													assign node344 = (inp[13]) ? node346 : 4'b0001;
														assign node346 = (inp[1]) ? 4'b0000 : 4'b0101;
													assign node349 = (inp[13]) ? 4'b0001 : 4'b0000;
									assign node352 = (inp[12]) ? node414 : node353;
										assign node353 = (inp[7]) ? node389 : node354;
											assign node354 = (inp[1]) ? node378 : node355;
												assign node355 = (inp[4]) ? node365 : node356;
													assign node356 = (inp[9]) ? node362 : node357;
														assign node357 = (inp[0]) ? 4'b0000 : node358;
															assign node358 = (inp[2]) ? 4'b0000 : 4'b0101;
														assign node362 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node365 = (inp[0]) ? node371 : node366;
														assign node366 = (inp[2]) ? node368 : 4'b0101;
															assign node368 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node371 = (inp[9]) ? node375 : node372;
															assign node372 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node375 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node378 = (inp[13]) ? node384 : node379;
													assign node379 = (inp[2]) ? node381 : 4'b0001;
														assign node381 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node384 = (inp[0]) ? node386 : 4'b0101;
														assign node386 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node389 = (inp[0]) ? node403 : node390;
												assign node390 = (inp[9]) ? node398 : node391;
													assign node391 = (inp[13]) ? node395 : node392;
														assign node392 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node395 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node398 = (inp[4]) ? 4'b0010 : node399;
														assign node399 = (inp[2]) ? 4'b0011 : 4'b0110;
												assign node403 = (inp[9]) ? node407 : node404;
													assign node404 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node407 = (inp[4]) ? 4'b0111 : node408;
														assign node408 = (inp[1]) ? 4'b0011 : node409;
															assign node409 = (inp[2]) ? 4'b0011 : 4'b0011;
										assign node414 = (inp[7]) ? node436 : node415;
											assign node415 = (inp[2]) ? node427 : node416;
												assign node416 = (inp[13]) ? node422 : node417;
													assign node417 = (inp[1]) ? 4'b0011 : node418;
														assign node418 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node422 = (inp[4]) ? 4'b0010 : node423;
														assign node423 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node427 = (inp[1]) ? 4'b0011 : node428;
													assign node428 = (inp[4]) ? 4'b0111 : node429;
														assign node429 = (inp[13]) ? node431 : 4'b0111;
															assign node431 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node436 = (inp[0]) ? node452 : node437;
												assign node437 = (inp[1]) ? node443 : node438;
													assign node438 = (inp[9]) ? 4'b0001 : node439;
														assign node439 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node443 = (inp[9]) ? node449 : node444;
														assign node444 = (inp[2]) ? node446 : 4'b0001;
															assign node446 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node449 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node452 = (inp[9]) ? node464 : node453;
													assign node453 = (inp[13]) ? node459 : node454;
														assign node454 = (inp[2]) ? node456 : 4'b0000;
															assign node456 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node459 = (inp[2]) ? node461 : 4'b0100;
															assign node461 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node464 = (inp[1]) ? 4'b0100 : node465;
														assign node465 = (inp[13]) ? 4'b0101 : 4'b0001;
							assign node469 = (inp[1]) ? node717 : node470;
								assign node470 = (inp[0]) ? node600 : node471;
									assign node471 = (inp[9]) ? node533 : node472;
										assign node472 = (inp[7]) ? node502 : node473;
											assign node473 = (inp[12]) ? node485 : node474;
												assign node474 = (inp[13]) ? node478 : node475;
													assign node475 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node478 = (inp[2]) ? node482 : node479;
														assign node479 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node482 = (inp[4]) ? 4'b0001 : 4'b0000;
												assign node485 = (inp[11]) ? node495 : node486;
													assign node486 = (inp[2]) ? 4'b0111 : node487;
														assign node487 = (inp[4]) ? node491 : node488;
															assign node488 = (inp[13]) ? 4'b0111 : 4'b0010;
															assign node491 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node495 = (inp[4]) ? node497 : 4'b0110;
														assign node497 = (inp[2]) ? 4'b0011 : node498;
															assign node498 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node502 = (inp[12]) ? node516 : node503;
												assign node503 = (inp[4]) ? 4'b0111 : node504;
													assign node504 = (inp[2]) ? node510 : node505;
														assign node505 = (inp[13]) ? node507 : 4'b0011;
															assign node507 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node510 = (inp[11]) ? node512 : 4'b0010;
															assign node512 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node516 = (inp[13]) ? node526 : node517;
													assign node517 = (inp[2]) ? node523 : node518;
														assign node518 = (inp[4]) ? node520 : 4'b0100;
															assign node520 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node523 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node526 = (inp[4]) ? 4'b0100 : node527;
														assign node527 = (inp[2]) ? node529 : 4'b0001;
															assign node529 = (inp[10]) ? 4'b0101 : 4'b0100;
										assign node533 = (inp[7]) ? node569 : node534;
											assign node534 = (inp[12]) ? node550 : node535;
												assign node535 = (inp[10]) ? node545 : node536;
													assign node536 = (inp[4]) ? node540 : node537;
														assign node537 = (inp[2]) ? 4'b0001 : 4'b0101;
														assign node540 = (inp[11]) ? node542 : 4'b0100;
															assign node542 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node545 = (inp[13]) ? 4'b0100 : node546;
														assign node546 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node550 = (inp[13]) ? node560 : node551;
													assign node551 = (inp[10]) ? node557 : node552;
														assign node552 = (inp[11]) ? node554 : 4'b0111;
															assign node554 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node557 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node560 = (inp[4]) ? node566 : node561;
														assign node561 = (inp[2]) ? node563 : 4'b0110;
															assign node563 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node566 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node569 = (inp[12]) ? node591 : node570;
												assign node570 = (inp[10]) ? node582 : node571;
													assign node571 = (inp[11]) ? node577 : node572;
														assign node572 = (inp[2]) ? 4'b0111 : node573;
															assign node573 = (inp[13]) ? 4'b0110 : 4'b0010;
														assign node577 = (inp[13]) ? node579 : 4'b0110;
															assign node579 = (inp[2]) ? 4'b0010 : 4'b0111;
													assign node582 = (inp[4]) ? node588 : node583;
														assign node583 = (inp[2]) ? node585 : 4'b0011;
															assign node585 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node588 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node591 = (inp[11]) ? node597 : node592;
													assign node592 = (inp[10]) ? 4'b0100 : node593;
														assign node593 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node597 = (inp[4]) ? 4'b0001 : 4'b0101;
									assign node600 = (inp[7]) ? node648 : node601;
										assign node601 = (inp[12]) ? node633 : node602;
											assign node602 = (inp[9]) ? node616 : node603;
												assign node603 = (inp[10]) ? node609 : node604;
													assign node604 = (inp[11]) ? 4'b0101 : node605;
														assign node605 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node609 = (inp[2]) ? node613 : node610;
														assign node610 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node613 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node616 = (inp[10]) ? node624 : node617;
													assign node617 = (inp[13]) ? node621 : node618;
														assign node618 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node621 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node624 = (inp[2]) ? node630 : node625;
														assign node625 = (inp[13]) ? node627 : 4'b0001;
															assign node627 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node630 = (inp[4]) ? 4'b0100 : 4'b0101;
											assign node633 = (inp[10]) ? node645 : node634;
												assign node634 = (inp[4]) ? node642 : node635;
													assign node635 = (inp[9]) ? 4'b0011 : node636;
														assign node636 = (inp[13]) ? node638 : 4'b0110;
															assign node638 = (inp[2]) ? 4'b0011 : 4'b0110;
													assign node642 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node645 = (inp[11]) ? 4'b0010 : 4'b0110;
										assign node648 = (inp[12]) ? node686 : node649;
											assign node649 = (inp[9]) ? node667 : node650;
												assign node650 = (inp[10]) ? node660 : node651;
													assign node651 = (inp[11]) ? 4'b0110 : node652;
														assign node652 = (inp[13]) ? node656 : node653;
															assign node653 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node656 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node660 = (inp[11]) ? 4'b0011 : node661;
														assign node661 = (inp[2]) ? node663 : 4'b0110;
															assign node663 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node667 = (inp[4]) ? node675 : node668;
													assign node668 = (inp[2]) ? node672 : node669;
														assign node669 = (inp[13]) ? 4'b0110 : 4'b0010;
														assign node672 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node675 = (inp[2]) ? node681 : node676;
														assign node676 = (inp[13]) ? 4'b0110 : node677;
															assign node677 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node681 = (inp[10]) ? node683 : 4'b0110;
															assign node683 = (inp[13]) ? 4'b0011 : 4'b0111;
											assign node686 = (inp[10]) ? node700 : node687;
												assign node687 = (inp[9]) ? node697 : node688;
													assign node688 = (inp[11]) ? 4'b0100 : node689;
														assign node689 = (inp[4]) ? node693 : node690;
															assign node690 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node693 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node697 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node700 = (inp[11]) ? node712 : node701;
													assign node701 = (inp[9]) ? node705 : node702;
														assign node702 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node705 = (inp[4]) ? node709 : node706;
															assign node706 = (inp[2]) ? 4'b0000 : 4'b0000;
															assign node709 = (inp[2]) ? 4'b0100 : 4'b0001;
													assign node712 = (inp[9]) ? node714 : 4'b0101;
														assign node714 = (inp[4]) ? 4'b0101 : 4'b0001;
								assign node717 = (inp[7]) ? node859 : node718;
									assign node718 = (inp[12]) ? node792 : node719;
										assign node719 = (inp[11]) ? node747 : node720;
											assign node720 = (inp[10]) ? node734 : node721;
												assign node721 = (inp[13]) ? node731 : node722;
													assign node722 = (inp[2]) ? node728 : node723;
														assign node723 = (inp[0]) ? node725 : 4'b0100;
															assign node725 = (inp[4]) ? 4'b0100 : 4'b0100;
														assign node728 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node731 = (inp[2]) ? 4'b0101 : 4'b0001;
												assign node734 = (inp[2]) ? node740 : node735;
													assign node735 = (inp[13]) ? node737 : 4'b0101;
														assign node737 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node740 = (inp[13]) ? node742 : 4'b0000;
														assign node742 = (inp[0]) ? 4'b0100 : node743;
															assign node743 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node747 = (inp[4]) ? node769 : node748;
												assign node748 = (inp[0]) ? node758 : node749;
													assign node749 = (inp[9]) ? 4'b0000 : node750;
														assign node750 = (inp[10]) ? node754 : node751;
															assign node751 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node754 = (inp[2]) ? 4'b0000 : 4'b0000;
													assign node758 = (inp[2]) ? node764 : node759;
														assign node759 = (inp[10]) ? node761 : 4'b0001;
															assign node761 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node764 = (inp[13]) ? 4'b0101 : node765;
															assign node765 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node769 = (inp[13]) ? node781 : node770;
													assign node770 = (inp[2]) ? node778 : node771;
														assign node771 = (inp[0]) ? node775 : node772;
															assign node772 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node775 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node778 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node781 = (inp[2]) ? node787 : node782;
														assign node782 = (inp[10]) ? node784 : 4'b0000;
															assign node784 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node787 = (inp[10]) ? 4'b0101 : node788;
															assign node788 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node792 = (inp[4]) ? node826 : node793;
											assign node793 = (inp[0]) ? node813 : node794;
												assign node794 = (inp[11]) ? node804 : node795;
													assign node795 = (inp[9]) ? node801 : node796;
														assign node796 = (inp[2]) ? 4'b0111 : node797;
															assign node797 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node801 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node804 = (inp[10]) ? node806 : 4'b0010;
														assign node806 = (inp[13]) ? node810 : node807;
															assign node807 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node810 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node813 = (inp[13]) ? node819 : node814;
													assign node814 = (inp[2]) ? 4'b0011 : node815;
														assign node815 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node819 = (inp[2]) ? node821 : 4'b0010;
														assign node821 = (inp[11]) ? node823 : 4'b0110;
															assign node823 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node826 = (inp[0]) ? node844 : node827;
												assign node827 = (inp[10]) ? node835 : node828;
													assign node828 = (inp[11]) ? node830 : 4'b0010;
														assign node830 = (inp[13]) ? node832 : 4'b0010;
															assign node832 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node835 = (inp[2]) ? node839 : node836;
														assign node836 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node839 = (inp[13]) ? 4'b0011 : node840;
															assign node840 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node844 = (inp[11]) ? node854 : node845;
													assign node845 = (inp[13]) ? node849 : node846;
														assign node846 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node849 = (inp[2]) ? node851 : 4'b0111;
															assign node851 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node854 = (inp[2]) ? 4'b0011 : node855;
														assign node855 = (inp[13]) ? 4'b0111 : 4'b0011;
									assign node859 = (inp[12]) ? node915 : node860;
										assign node860 = (inp[2]) ? node888 : node861;
											assign node861 = (inp[13]) ? node875 : node862;
												assign node862 = (inp[9]) ? node864 : 4'b0110;
													assign node864 = (inp[10]) ? node870 : node865;
														assign node865 = (inp[11]) ? node867 : 4'b0110;
															assign node867 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node870 = (inp[4]) ? node872 : 4'b0111;
															assign node872 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node875 = (inp[10]) ? node881 : node876;
													assign node876 = (inp[4]) ? node878 : 4'b0011;
														assign node878 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node881 = (inp[11]) ? 4'b0011 : node882;
														assign node882 = (inp[4]) ? 4'b0011 : node883;
															assign node883 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node888 = (inp[13]) ? node906 : node889;
												assign node889 = (inp[11]) ? node891 : 4'b0010;
													assign node891 = (inp[9]) ? node899 : node892;
														assign node892 = (inp[0]) ? node896 : node893;
															assign node893 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node896 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node899 = (inp[10]) ? node903 : node900;
															assign node900 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node903 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node906 = (inp[10]) ? 4'b0110 : node907;
													assign node907 = (inp[9]) ? node911 : node908;
														assign node908 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node911 = (inp[4]) ? 4'b0110 : 4'b0111;
										assign node915 = (inp[13]) ? node947 : node916;
											assign node916 = (inp[2]) ? node934 : node917;
												assign node917 = (inp[4]) ? node925 : node918;
													assign node918 = (inp[0]) ? 4'b0101 : node919;
														assign node919 = (inp[10]) ? node921 : 4'b0101;
															assign node921 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node925 = (inp[0]) ? node931 : node926;
														assign node926 = (inp[11]) ? node928 : 4'b0001;
															assign node928 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node931 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node934 = (inp[4]) ? node944 : node935;
													assign node935 = (inp[11]) ? node941 : node936;
														assign node936 = (inp[0]) ? node938 : 4'b0000;
															assign node938 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node941 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node944 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node947 = (inp[11]) ? node971 : node948;
												assign node948 = (inp[9]) ? node962 : node949;
													assign node949 = (inp[4]) ? node957 : node950;
														assign node950 = (inp[10]) ? node954 : node951;
															assign node951 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node954 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node957 = (inp[10]) ? 4'b0101 : node958;
															assign node958 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node962 = (inp[10]) ? node968 : node963;
														assign node963 = (inp[4]) ? node965 : 4'b0100;
															assign node965 = (inp[0]) ? 4'b0000 : 4'b0100;
														assign node968 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node971 = (inp[0]) ? node979 : node972;
													assign node972 = (inp[10]) ? 4'b0000 : node973;
														assign node973 = (inp[2]) ? node975 : 4'b0100;
															assign node975 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node979 = (inp[4]) ? node985 : node980;
														assign node980 = (inp[2]) ? node982 : 4'b0000;
															assign node982 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node985 = (inp[10]) ? 4'b0001 : 4'b0000;
						assign node988 = (inp[13]) ? node1440 : node989;
							assign node989 = (inp[2]) ? node1227 : node990;
								assign node990 = (inp[12]) ? node1116 : node991;
									assign node991 = (inp[5]) ? node1053 : node992;
										assign node992 = (inp[7]) ? node1032 : node993;
											assign node993 = (inp[4]) ? node1007 : node994;
												assign node994 = (inp[9]) ? node1000 : node995;
													assign node995 = (inp[1]) ? 4'b0000 : node996;
														assign node996 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node1000 = (inp[10]) ? 4'b0001 : node1001;
														assign node1001 = (inp[11]) ? node1003 : 4'b0001;
															assign node1003 = (inp[1]) ? 4'b0000 : 4'b0000;
												assign node1007 = (inp[1]) ? node1021 : node1008;
													assign node1008 = (inp[9]) ? node1014 : node1009;
														assign node1009 = (inp[11]) ? 4'b0010 : node1010;
															assign node1010 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node1014 = (inp[0]) ? node1018 : node1015;
															assign node1015 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node1018 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node1021 = (inp[0]) ? node1027 : node1022;
														assign node1022 = (inp[10]) ? node1024 : 4'b0111;
															assign node1024 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node1027 = (inp[10]) ? 4'b0110 : node1028;
															assign node1028 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node1032 = (inp[4]) ? node1048 : node1033;
												assign node1033 = (inp[11]) ? node1041 : node1034;
													assign node1034 = (inp[0]) ? 4'b0110 : node1035;
														assign node1035 = (inp[1]) ? node1037 : 4'b0110;
															assign node1037 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node1041 = (inp[1]) ? node1043 : 4'b0111;
														assign node1043 = (inp[10]) ? node1045 : 4'b0110;
															assign node1045 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node1048 = (inp[9]) ? node1050 : 4'b0000;
													assign node1050 = (inp[10]) ? 4'b0001 : 4'b0000;
										assign node1053 = (inp[4]) ? node1093 : node1054;
											assign node1054 = (inp[7]) ? node1068 : node1055;
												assign node1055 = (inp[1]) ? node1061 : node1056;
													assign node1056 = (inp[0]) ? node1058 : 4'b0000;
														assign node1058 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node1061 = (inp[9]) ? 4'b0100 : node1062;
														assign node1062 = (inp[0]) ? 4'b0101 : node1063;
															assign node1063 = (inp[10]) ? 4'b0100 : 4'b0100;
												assign node1068 = (inp[1]) ? node1080 : node1069;
													assign node1069 = (inp[9]) ? node1077 : node1070;
														assign node1070 = (inp[11]) ? node1074 : node1071;
															assign node1071 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node1074 = (inp[0]) ? 4'b0110 : 4'b0110;
														assign node1077 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node1080 = (inp[11]) ? node1088 : node1081;
														assign node1081 = (inp[10]) ? node1085 : node1082;
															assign node1082 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node1085 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node1088 = (inp[0]) ? 4'b0010 : node1089;
															assign node1089 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node1093 = (inp[7]) ? node1105 : node1094;
												assign node1094 = (inp[9]) ? node1100 : node1095;
													assign node1095 = (inp[11]) ? node1097 : 4'b0110;
														assign node1097 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node1100 = (inp[11]) ? node1102 : 4'b0111;
														assign node1102 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node1105 = (inp[1]) ? node1107 : 4'b0000;
													assign node1107 = (inp[9]) ? node1111 : node1108;
														assign node1108 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node1111 = (inp[11]) ? node1113 : 4'b0101;
															assign node1113 = (inp[0]) ? 4'b0101 : 4'b0100;
									assign node1116 = (inp[4]) ? node1164 : node1117;
										assign node1117 = (inp[7]) ? node1145 : node1118;
											assign node1118 = (inp[5]) ? node1136 : node1119;
												assign node1119 = (inp[0]) ? node1129 : node1120;
													assign node1120 = (inp[11]) ? node1122 : 4'b0010;
														assign node1122 = (inp[9]) ? node1126 : node1123;
															assign node1123 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node1126 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node1129 = (inp[10]) ? 4'b0011 : node1130;
														assign node1130 = (inp[1]) ? node1132 : 4'b0011;
															assign node1132 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node1136 = (inp[1]) ? node1140 : node1137;
													assign node1137 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node1140 = (inp[11]) ? 4'b0111 : node1141;
														assign node1141 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node1145 = (inp[5]) ? node1153 : node1146;
												assign node1146 = (inp[1]) ? node1148 : 4'b0100;
													assign node1148 = (inp[0]) ? 4'b0000 : node1149;
														assign node1149 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node1153 = (inp[9]) ? node1159 : node1154;
													assign node1154 = (inp[10]) ? 4'b0001 : node1155;
														assign node1155 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node1159 = (inp[11]) ? node1161 : 4'b0000;
														assign node1161 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node1164 = (inp[7]) ? node1196 : node1165;
											assign node1165 = (inp[1]) ? node1183 : node1166;
												assign node1166 = (inp[0]) ? node1174 : node1167;
													assign node1167 = (inp[5]) ? 4'b0000 : node1168;
														assign node1168 = (inp[11]) ? node1170 : 4'b0000;
															assign node1170 = (inp[9]) ? 4'b0000 : 4'b0000;
													assign node1174 = (inp[5]) ? node1176 : 4'b0001;
														assign node1176 = (inp[9]) ? node1180 : node1177;
															assign node1177 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node1180 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node1183 = (inp[5]) ? node1191 : node1184;
													assign node1184 = (inp[10]) ? node1188 : node1185;
														assign node1185 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node1188 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node1191 = (inp[0]) ? 4'b0101 : node1192;
														assign node1192 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node1196 = (inp[1]) ? node1212 : node1197;
												assign node1197 = (inp[0]) ? node1207 : node1198;
													assign node1198 = (inp[10]) ? node1200 : 4'b0111;
														assign node1200 = (inp[5]) ? node1204 : node1201;
															assign node1201 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node1204 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node1207 = (inp[5]) ? node1209 : 4'b0110;
														assign node1209 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node1212 = (inp[5]) ? node1218 : node1213;
													assign node1213 = (inp[0]) ? node1215 : 4'b0111;
														assign node1215 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node1218 = (inp[10]) ? 4'b0011 : node1219;
														assign node1219 = (inp[0]) ? node1223 : node1220;
															assign node1220 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node1223 = (inp[9]) ? 4'b0010 : 4'b0011;
								assign node1227 = (inp[4]) ? node1337 : node1228;
									assign node1228 = (inp[12]) ? node1278 : node1229;
										assign node1229 = (inp[7]) ? node1253 : node1230;
											assign node1230 = (inp[1]) ? node1238 : node1231;
												assign node1231 = (inp[10]) ? 4'b0100 : node1232;
													assign node1232 = (inp[11]) ? node1234 : 4'b0100;
														assign node1234 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node1238 = (inp[5]) ? node1244 : node1239;
													assign node1239 = (inp[9]) ? 4'b0101 : node1240;
														assign node1240 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node1244 = (inp[10]) ? 4'b0000 : node1245;
														assign node1245 = (inp[0]) ? node1249 : node1246;
															assign node1246 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node1249 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node1253 = (inp[5]) ? node1269 : node1254;
												assign node1254 = (inp[1]) ? node1262 : node1255;
													assign node1255 = (inp[11]) ? 4'b0010 : node1256;
														assign node1256 = (inp[9]) ? 4'b0010 : node1257;
															assign node1257 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node1262 = (inp[9]) ? node1266 : node1263;
														assign node1263 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node1266 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node1269 = (inp[1]) ? node1271 : 4'b0011;
													assign node1271 = (inp[10]) ? 4'b0110 : node1272;
														assign node1272 = (inp[11]) ? node1274 : 4'b0111;
															assign node1274 = (inp[9]) ? 4'b0110 : 4'b0110;
										assign node1278 = (inp[7]) ? node1306 : node1279;
											assign node1279 = (inp[5]) ? node1295 : node1280;
												assign node1280 = (inp[9]) ? node1286 : node1281;
													assign node1281 = (inp[10]) ? node1283 : 4'b0110;
														assign node1283 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node1286 = (inp[0]) ? 4'b0110 : node1287;
														assign node1287 = (inp[1]) ? node1291 : node1288;
															assign node1288 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node1291 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node1295 = (inp[1]) ? node1299 : node1296;
													assign node1296 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node1299 = (inp[10]) ? 4'b0011 : node1300;
														assign node1300 = (inp[9]) ? node1302 : 4'b0010;
															assign node1302 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node1306 = (inp[0]) ? node1320 : node1307;
												assign node1307 = (inp[5]) ? node1309 : 4'b0101;
													assign node1309 = (inp[11]) ? node1315 : node1310;
														assign node1310 = (inp[9]) ? node1312 : 4'b0101;
															assign node1312 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node1315 = (inp[1]) ? node1317 : 4'b0100;
															assign node1317 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node1320 = (inp[1]) ? node1328 : node1321;
													assign node1321 = (inp[5]) ? node1325 : node1322;
														assign node1322 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node1325 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node1328 = (inp[9]) ? 4'b0100 : node1329;
														assign node1329 = (inp[5]) ? node1333 : node1330;
															assign node1330 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node1333 = (inp[10]) ? 4'b0101 : 4'b0100;
									assign node1337 = (inp[5]) ? node1389 : node1338;
										assign node1338 = (inp[7]) ? node1360 : node1339;
											assign node1339 = (inp[12]) ? node1347 : node1340;
												assign node1340 = (inp[1]) ? node1342 : 4'b0110;
													assign node1342 = (inp[11]) ? 4'b0011 : node1343;
														assign node1343 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node1347 = (inp[11]) ? node1351 : node1348;
													assign node1348 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node1351 = (inp[0]) ? node1353 : 4'b0100;
														assign node1353 = (inp[10]) ? node1357 : node1354;
															assign node1354 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node1357 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node1360 = (inp[12]) ? node1374 : node1361;
												assign node1361 = (inp[11]) ? node1369 : node1362;
													assign node1362 = (inp[1]) ? 4'b0100 : node1363;
														assign node1363 = (inp[9]) ? 4'b0100 : node1364;
															assign node1364 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node1369 = (inp[10]) ? node1371 : 4'b0101;
														assign node1371 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node1374 = (inp[10]) ? node1384 : node1375;
													assign node1375 = (inp[9]) ? node1379 : node1376;
														assign node1376 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node1379 = (inp[1]) ? node1381 : 4'b0010;
															assign node1381 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node1384 = (inp[11]) ? 4'b0010 : node1385;
														assign node1385 = (inp[9]) ? 4'b0010 : 4'b0011;
										assign node1389 = (inp[7]) ? node1415 : node1390;
											assign node1390 = (inp[12]) ? node1404 : node1391;
												assign node1391 = (inp[1]) ? node1397 : node1392;
													assign node1392 = (inp[10]) ? 4'b0010 : node1393;
														assign node1393 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node1397 = (inp[9]) ? node1399 : 4'b0011;
														assign node1399 = (inp[10]) ? node1401 : 4'b0010;
															assign node1401 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node1404 = (inp[1]) ? node1408 : node1405;
													assign node1405 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node1408 = (inp[10]) ? node1410 : 4'b0001;
														assign node1410 = (inp[11]) ? 4'b0001 : node1411;
															assign node1411 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node1415 = (inp[12]) ? node1425 : node1416;
												assign node1416 = (inp[1]) ? node1420 : node1417;
													assign node1417 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node1420 = (inp[11]) ? 4'b0001 : node1421;
														assign node1421 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node1425 = (inp[1]) ? node1433 : node1426;
													assign node1426 = (inp[0]) ? node1428 : 4'b0011;
														assign node1428 = (inp[10]) ? 4'b0010 : node1429;
															assign node1429 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node1433 = (inp[10]) ? node1435 : 4'b0111;
														assign node1435 = (inp[0]) ? 4'b0110 : node1436;
															assign node1436 = (inp[9]) ? 4'b0110 : 4'b0111;
							assign node1440 = (inp[2]) ? node1698 : node1441;
								assign node1441 = (inp[4]) ? node1567 : node1442;
									assign node1442 = (inp[12]) ? node1494 : node1443;
										assign node1443 = (inp[7]) ? node1475 : node1444;
											assign node1444 = (inp[5]) ? node1462 : node1445;
												assign node1445 = (inp[0]) ? node1453 : node1446;
													assign node1446 = (inp[9]) ? node1448 : 4'b0100;
														assign node1448 = (inp[1]) ? node1450 : 4'b0101;
															assign node1450 = (inp[11]) ? 4'b0100 : 4'b0100;
													assign node1453 = (inp[9]) ? 4'b0101 : node1454;
														assign node1454 = (inp[10]) ? node1458 : node1455;
															assign node1455 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node1458 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node1462 = (inp[1]) ? node1470 : node1463;
													assign node1463 = (inp[11]) ? 4'b0100 : node1464;
														assign node1464 = (inp[10]) ? 4'b0101 : node1465;
															assign node1465 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node1470 = (inp[9]) ? node1472 : 4'b0000;
														assign node1472 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node1475 = (inp[5]) ? node1485 : node1476;
												assign node1476 = (inp[9]) ? 4'b0010 : node1477;
													assign node1477 = (inp[10]) ? 4'b0011 : node1478;
														assign node1478 = (inp[1]) ? node1480 : 4'b0010;
															assign node1480 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node1485 = (inp[1]) ? node1491 : node1486;
													assign node1486 = (inp[9]) ? node1488 : 4'b0011;
														assign node1488 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node1491 = (inp[0]) ? 4'b0111 : 4'b0110;
										assign node1494 = (inp[7]) ? node1524 : node1495;
											assign node1495 = (inp[5]) ? node1511 : node1496;
												assign node1496 = (inp[1]) ? node1506 : node1497;
													assign node1497 = (inp[0]) ? 4'b0110 : node1498;
														assign node1498 = (inp[10]) ? node1502 : node1499;
															assign node1499 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node1502 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node1506 = (inp[10]) ? node1508 : 4'b0111;
														assign node1508 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node1511 = (inp[1]) ? node1519 : node1512;
													assign node1512 = (inp[9]) ? node1516 : node1513;
														assign node1513 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node1516 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node1519 = (inp[0]) ? 4'b0010 : node1520;
														assign node1520 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node1524 = (inp[1]) ? node1542 : node1525;
												assign node1525 = (inp[5]) ? node1533 : node1526;
													assign node1526 = (inp[9]) ? node1528 : 4'b0000;
														assign node1528 = (inp[11]) ? 4'b0001 : node1529;
															assign node1529 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node1533 = (inp[10]) ? node1539 : node1534;
														assign node1534 = (inp[0]) ? node1536 : 4'b0100;
															assign node1536 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node1539 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node1542 = (inp[0]) ? node1552 : node1543;
													assign node1543 = (inp[11]) ? node1545 : 4'b0100;
														assign node1545 = (inp[10]) ? node1549 : node1546;
															assign node1546 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node1549 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node1552 = (inp[10]) ? node1560 : node1553;
														assign node1553 = (inp[5]) ? node1557 : node1554;
															assign node1554 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node1557 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node1560 = (inp[5]) ? node1564 : node1561;
															assign node1561 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node1564 = (inp[9]) ? 4'b0101 : 4'b0100;
									assign node1567 = (inp[5]) ? node1629 : node1568;
										assign node1568 = (inp[7]) ? node1598 : node1569;
											assign node1569 = (inp[12]) ? node1581 : node1570;
												assign node1570 = (inp[1]) ? node1578 : node1571;
													assign node1571 = (inp[0]) ? 4'b0111 : node1572;
														assign node1572 = (inp[10]) ? 4'b0110 : node1573;
															assign node1573 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node1578 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node1581 = (inp[1]) ? node1589 : node1582;
													assign node1582 = (inp[10]) ? node1586 : node1583;
														assign node1583 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node1586 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node1589 = (inp[11]) ? 4'b0101 : node1590;
														assign node1590 = (inp[9]) ? node1594 : node1591;
															assign node1591 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node1594 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node1598 = (inp[12]) ? node1614 : node1599;
												assign node1599 = (inp[0]) ? node1607 : node1600;
													assign node1600 = (inp[9]) ? 4'b0101 : node1601;
														assign node1601 = (inp[10]) ? node1603 : 4'b0100;
															assign node1603 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node1607 = (inp[1]) ? node1609 : 4'b0100;
														assign node1609 = (inp[10]) ? 4'b0101 : node1610;
															assign node1610 = (inp[11]) ? 4'b0100 : 4'b0100;
												assign node1614 = (inp[0]) ? node1620 : node1615;
													assign node1615 = (inp[9]) ? 4'b0010 : node1616;
														assign node1616 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node1620 = (inp[1]) ? node1622 : 4'b0011;
														assign node1622 = (inp[11]) ? node1626 : node1623;
															assign node1623 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node1626 = (inp[9]) ? 4'b0010 : 4'b0010;
										assign node1629 = (inp[0]) ? node1655 : node1630;
											assign node1630 = (inp[1]) ? node1636 : node1631;
												assign node1631 = (inp[9]) ? 4'b0010 : node1632;
													assign node1632 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node1636 = (inp[12]) ? node1644 : node1637;
													assign node1637 = (inp[7]) ? node1639 : 4'b0010;
														assign node1639 = (inp[9]) ? node1641 : 4'b0000;
															assign node1641 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node1644 = (inp[7]) ? node1650 : node1645;
														assign node1645 = (inp[11]) ? 4'b0001 : node1646;
															assign node1646 = (inp[10]) ? 4'b0000 : 4'b0000;
														assign node1650 = (inp[10]) ? node1652 : 4'b0110;
															assign node1652 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node1655 = (inp[1]) ? node1679 : node1656;
												assign node1656 = (inp[10]) ? node1664 : node1657;
													assign node1657 = (inp[7]) ? node1659 : 4'b0101;
														assign node1659 = (inp[11]) ? node1661 : 4'b0100;
															assign node1661 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node1664 = (inp[9]) ? node1672 : node1665;
														assign node1665 = (inp[12]) ? node1669 : node1666;
															assign node1666 = (inp[7]) ? 4'b0100 : 4'b0011;
															assign node1669 = (inp[7]) ? 4'b0011 : 4'b0101;
														assign node1672 = (inp[12]) ? node1676 : node1673;
															assign node1673 = (inp[7]) ? 4'b0101 : 4'b0011;
															assign node1676 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node1679 = (inp[12]) ? node1689 : node1680;
													assign node1680 = (inp[7]) ? node1686 : node1681;
														assign node1681 = (inp[11]) ? 4'b0011 : node1682;
															assign node1682 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node1686 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node1689 = (inp[7]) ? node1695 : node1690;
														assign node1690 = (inp[11]) ? node1692 : 4'b0000;
															assign node1692 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node1695 = (inp[11]) ? 4'b0110 : 4'b0111;
								assign node1698 = (inp[1]) ? node1802 : node1699;
									assign node1699 = (inp[7]) ? node1757 : node1700;
										assign node1700 = (inp[4]) ? node1728 : node1701;
											assign node1701 = (inp[12]) ? node1719 : node1702;
												assign node1702 = (inp[5]) ? node1708 : node1703;
													assign node1703 = (inp[10]) ? 4'b0001 : node1704;
														assign node1704 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node1708 = (inp[10]) ? node1714 : node1709;
														assign node1709 = (inp[0]) ? node1711 : 4'b0001;
															assign node1711 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node1714 = (inp[0]) ? 4'b0000 : node1715;
															assign node1715 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node1719 = (inp[9]) ? 4'b0010 : node1720;
													assign node1720 = (inp[11]) ? 4'b0011 : node1721;
														assign node1721 = (inp[5]) ? node1723 : 4'b0011;
															assign node1723 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node1728 = (inp[12]) ? node1744 : node1729;
												assign node1729 = (inp[5]) ? node1741 : node1730;
													assign node1730 = (inp[0]) ? node1736 : node1731;
														assign node1731 = (inp[11]) ? 4'b0010 : node1732;
															assign node1732 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node1736 = (inp[9]) ? 4'b0011 : node1737;
															assign node1737 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node1741 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node1744 = (inp[5]) ? node1752 : node1745;
													assign node1745 = (inp[11]) ? node1747 : 4'b0001;
														assign node1747 = (inp[10]) ? node1749 : 4'b0000;
															assign node1749 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node1752 = (inp[10]) ? 4'b0000 : node1753;
														assign node1753 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node1757 = (inp[12]) ? node1779 : node1758;
											assign node1758 = (inp[4]) ? node1766 : node1759;
												assign node1759 = (inp[0]) ? 4'b0110 : node1760;
													assign node1760 = (inp[5]) ? 4'b0111 : node1761;
														assign node1761 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node1766 = (inp[9]) ? node1768 : 4'b0001;
													assign node1768 = (inp[10]) ? node1774 : node1769;
														assign node1769 = (inp[11]) ? node1771 : 4'b0000;
															assign node1771 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node1774 = (inp[11]) ? 4'b0001 : node1775;
															assign node1775 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node1779 = (inp[4]) ? node1785 : node1780;
												assign node1780 = (inp[5]) ? node1782 : 4'b0100;
													assign node1782 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node1785 = (inp[11]) ? node1791 : node1786;
													assign node1786 = (inp[10]) ? node1788 : 4'b0111;
														assign node1788 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node1791 = (inp[5]) ? node1797 : node1792;
														assign node1792 = (inp[10]) ? node1794 : 4'b0110;
															assign node1794 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node1797 = (inp[0]) ? node1799 : 4'b0111;
															assign node1799 = (inp[9]) ? 4'b0111 : 4'b0110;
									assign node1802 = (inp[4]) ? node1858 : node1803;
										assign node1803 = (inp[12]) ? node1825 : node1804;
											assign node1804 = (inp[7]) ? node1812 : node1805;
												assign node1805 = (inp[0]) ? node1809 : node1806;
													assign node1806 = (inp[5]) ? 4'b0100 : 4'b0000;
													assign node1809 = (inp[5]) ? 4'b0101 : 4'b0001;
												assign node1812 = (inp[5]) ? node1820 : node1813;
													assign node1813 = (inp[9]) ? 4'b0110 : node1814;
														assign node1814 = (inp[10]) ? node1816 : 4'b0110;
															assign node1816 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node1820 = (inp[0]) ? 4'b0010 : node1821;
														assign node1821 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node1825 = (inp[7]) ? node1845 : node1826;
												assign node1826 = (inp[5]) ? node1838 : node1827;
													assign node1827 = (inp[11]) ? node1833 : node1828;
														assign node1828 = (inp[9]) ? 4'b0010 : node1829;
															assign node1829 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node1833 = (inp[9]) ? 4'b0011 : node1834;
															assign node1834 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node1838 = (inp[0]) ? 4'b0110 : node1839;
														assign node1839 = (inp[10]) ? 4'b0111 : node1840;
															assign node1840 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node1845 = (inp[9]) ? node1853 : node1846;
													assign node1846 = (inp[0]) ? 4'b0000 : node1847;
														assign node1847 = (inp[5]) ? node1849 : 4'b0001;
															assign node1849 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node1853 = (inp[0]) ? node1855 : 4'b0000;
														assign node1855 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node1858 = (inp[0]) ? node1888 : node1859;
											assign node1859 = (inp[5]) ? node1873 : node1860;
												assign node1860 = (inp[9]) ? node1864 : node1861;
													assign node1861 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node1864 = (inp[11]) ? node1866 : 4'b0111;
														assign node1866 = (inp[10]) ? node1870 : node1867;
															assign node1867 = (inp[7]) ? 4'b0001 : 4'b0110;
															assign node1870 = (inp[7]) ? 4'b0111 : 4'b0001;
												assign node1873 = (inp[12]) ? node1883 : node1874;
													assign node1874 = (inp[7]) ? node1876 : 4'b0111;
														assign node1876 = (inp[9]) ? node1880 : node1877;
															assign node1877 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node1880 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node1883 = (inp[7]) ? node1885 : 4'b0100;
														assign node1885 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node1888 = (inp[12]) ? node1898 : node1889;
												assign node1889 = (inp[7]) ? 4'b0000 : node1890;
													assign node1890 = (inp[11]) ? 4'b0111 : node1891;
														assign node1891 = (inp[5]) ? 4'b0110 : node1892;
															assign node1892 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node1898 = (inp[7]) ? node1902 : node1899;
													assign node1899 = (inp[5]) ? 4'b0100 : 4'b0000;
													assign node1902 = (inp[9]) ? 4'b0010 : 4'b0110;
					assign node1905 = (inp[13]) ? node2849 : node1906;
						assign node1906 = (inp[2]) ? node2376 : node1907;
							assign node1907 = (inp[1]) ? node2131 : node1908;
								assign node1908 = (inp[5]) ? node2012 : node1909;
									assign node1909 = (inp[15]) ? node1959 : node1910;
										assign node1910 = (inp[12]) ? node1938 : node1911;
											assign node1911 = (inp[7]) ? node1925 : node1912;
												assign node1912 = (inp[11]) ? node1920 : node1913;
													assign node1913 = (inp[9]) ? node1917 : node1914;
														assign node1914 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node1917 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node1920 = (inp[4]) ? node1922 : 4'b1000;
														assign node1922 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node1925 = (inp[10]) ? node1931 : node1926;
													assign node1926 = (inp[11]) ? node1928 : 4'b1010;
														assign node1928 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node1931 = (inp[9]) ? node1933 : 4'b1011;
														assign node1933 = (inp[0]) ? 4'b1010 : node1934;
															assign node1934 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node1938 = (inp[7]) ? node1950 : node1939;
												assign node1939 = (inp[4]) ? node1943 : node1940;
													assign node1940 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node1943 = (inp[11]) ? node1945 : 4'b1110;
														assign node1945 = (inp[10]) ? 4'b1111 : node1946;
															assign node1946 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node1950 = (inp[4]) ? node1956 : node1951;
													assign node1951 = (inp[11]) ? node1953 : 4'b1101;
														assign node1953 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node1956 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node1959 = (inp[7]) ? node1987 : node1960;
											assign node1960 = (inp[9]) ? node1978 : node1961;
												assign node1961 = (inp[11]) ? node1965 : node1962;
													assign node1962 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node1965 = (inp[0]) ? node1973 : node1966;
														assign node1966 = (inp[4]) ? node1970 : node1967;
															assign node1967 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node1970 = (inp[12]) ? 4'b1011 : 4'b1100;
														assign node1973 = (inp[12]) ? 4'b1011 : node1974;
															assign node1974 = (inp[4]) ? 4'b1101 : 4'b1011;
												assign node1978 = (inp[10]) ? node1982 : node1979;
													assign node1979 = (inp[0]) ? 4'b1101 : 4'b1011;
													assign node1982 = (inp[12]) ? 4'b1100 : node1983;
														assign node1983 = (inp[4]) ? 4'b1100 : 4'b1010;
											assign node1987 = (inp[12]) ? node2001 : node1988;
												assign node1988 = (inp[4]) ? node1998 : node1989;
													assign node1989 = (inp[11]) ? node1993 : node1990;
														assign node1990 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node1993 = (inp[0]) ? node1995 : 4'b1101;
															assign node1995 = (inp[10]) ? 4'b1100 : 4'b1100;
													assign node1998 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node2001 = (inp[4]) ? node2009 : node2002;
													assign node2002 = (inp[10]) ? 4'b1011 : node2003;
														assign node2003 = (inp[0]) ? 4'b1010 : node2004;
															assign node2004 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node2009 = (inp[10]) ? 4'b1001 : 4'b1000;
									assign node2012 = (inp[7]) ? node2072 : node2013;
										assign node2013 = (inp[12]) ? node2043 : node2014;
											assign node2014 = (inp[4]) ? node2032 : node2015;
												assign node2015 = (inp[15]) ? node2023 : node2016;
													assign node2016 = (inp[10]) ? 4'b1100 : node2017;
														assign node2017 = (inp[9]) ? node2019 : 4'b1100;
															assign node2019 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node2023 = (inp[10]) ? node2027 : node2024;
														assign node2024 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node2027 = (inp[9]) ? 4'b1110 : node2028;
															assign node2028 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node2032 = (inp[15]) ? node2036 : node2033;
													assign node2033 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node2036 = (inp[0]) ? node2038 : 4'b1000;
														assign node2038 = (inp[10]) ? node2040 : 4'b1001;
															assign node2040 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node2043 = (inp[4]) ? node2059 : node2044;
												assign node2044 = (inp[15]) ? node2056 : node2045;
													assign node2045 = (inp[10]) ? node2049 : node2046;
														assign node2046 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node2049 = (inp[11]) ? node2053 : node2050;
															assign node2050 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node2053 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node2056 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node2059 = (inp[15]) ? node2065 : node2060;
													assign node2060 = (inp[11]) ? node2062 : 4'b1110;
														assign node2062 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node2065 = (inp[9]) ? 4'b1010 : node2066;
														assign node2066 = (inp[10]) ? node2068 : 4'b1011;
															assign node2068 = (inp[11]) ? 4'b1010 : 4'b1011;
										assign node2072 = (inp[12]) ? node2096 : node2073;
											assign node2073 = (inp[15]) ? node2087 : node2074;
												assign node2074 = (inp[10]) ? node2082 : node2075;
													assign node2075 = (inp[9]) ? node2077 : 4'b1111;
														assign node2077 = (inp[4]) ? 4'b1111 : node2078;
															assign node2078 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node2082 = (inp[4]) ? 4'b1110 : node2083;
														assign node2083 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node2087 = (inp[4]) ? node2093 : node2088;
													assign node2088 = (inp[11]) ? 4'b1100 : node2089;
														assign node2089 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node2093 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node2096 = (inp[4]) ? node2110 : node2097;
												assign node2097 = (inp[15]) ? node2105 : node2098;
													assign node2098 = (inp[11]) ? 4'b1001 : node2099;
														assign node2099 = (inp[10]) ? node2101 : 4'b1000;
															assign node2101 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node2105 = (inp[0]) ? 4'b1111 : node2106;
														assign node2106 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node2110 = (inp[11]) ? node2124 : node2111;
													assign node2111 = (inp[15]) ? node2119 : node2112;
														assign node2112 = (inp[0]) ? node2116 : node2113;
															assign node2113 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node2116 = (inp[9]) ? 4'b1100 : 4'b1100;
														assign node2119 = (inp[0]) ? 4'b1101 : node2120;
															assign node2120 = (inp[10]) ? 4'b1100 : 4'b1100;
													assign node2124 = (inp[0]) ? 4'b1100 : node2125;
														assign node2125 = (inp[15]) ? 4'b1101 : node2126;
															assign node2126 = (inp[10]) ? 4'b1100 : 4'b1100;
								assign node2131 = (inp[12]) ? node2249 : node2132;
									assign node2132 = (inp[7]) ? node2196 : node2133;
										assign node2133 = (inp[15]) ? node2167 : node2134;
											assign node2134 = (inp[4]) ? node2150 : node2135;
												assign node2135 = (inp[10]) ? node2143 : node2136;
													assign node2136 = (inp[5]) ? node2138 : 4'b1001;
														assign node2138 = (inp[0]) ? node2140 : 4'b1000;
															assign node2140 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node2143 = (inp[9]) ? node2145 : 4'b1001;
														assign node2145 = (inp[5]) ? 4'b1001 : node2146;
															assign node2146 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node2150 = (inp[9]) ? node2162 : node2151;
													assign node2151 = (inp[10]) ? node2157 : node2152;
														assign node2152 = (inp[11]) ? 4'b1000 : node2153;
															assign node2153 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node2157 = (inp[0]) ? 4'b1001 : node2158;
															assign node2158 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node2162 = (inp[5]) ? 4'b1000 : node2163;
														assign node2163 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node2167 = (inp[4]) ? node2183 : node2168;
												assign node2168 = (inp[11]) ? 4'b1010 : node2169;
													assign node2169 = (inp[5]) ? node2175 : node2170;
														assign node2170 = (inp[9]) ? 4'b1011 : node2171;
															assign node2171 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node2175 = (inp[10]) ? node2179 : node2176;
															assign node2176 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node2179 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node2183 = (inp[5]) ? node2191 : node2184;
													assign node2184 = (inp[11]) ? 4'b1100 : node2185;
														assign node2185 = (inp[9]) ? node2187 : 4'b1101;
															assign node2187 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node2191 = (inp[9]) ? node2193 : 4'b1100;
														assign node2193 = (inp[10]) ? 4'b1101 : 4'b1100;
										assign node2196 = (inp[4]) ? node2222 : node2197;
											assign node2197 = (inp[15]) ? node2209 : node2198;
												assign node2198 = (inp[9]) ? 4'b1010 : node2199;
													assign node2199 = (inp[11]) ? node2205 : node2200;
														assign node2200 = (inp[10]) ? node2202 : 4'b1010;
															assign node2202 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node2205 = (inp[5]) ? 4'b1010 : 4'b1011;
												assign node2209 = (inp[5]) ? node2213 : node2210;
													assign node2210 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node2213 = (inp[11]) ? node2217 : node2214;
														assign node2214 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node2217 = (inp[9]) ? node2219 : 4'b1101;
															assign node2219 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node2222 = (inp[11]) ? node2238 : node2223;
												assign node2223 = (inp[15]) ? node2231 : node2224;
													assign node2224 = (inp[5]) ? 4'b1011 : node2225;
														assign node2225 = (inp[9]) ? 4'b1010 : node2226;
															assign node2226 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node2231 = (inp[5]) ? 4'b1010 : node2232;
														assign node2232 = (inp[10]) ? 4'b1011 : node2233;
															assign node2233 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node2238 = (inp[0]) ? node2240 : 4'b1011;
													assign node2240 = (inp[9]) ? node2246 : node2241;
														assign node2241 = (inp[15]) ? 4'b1011 : node2242;
															assign node2242 = (inp[5]) ? 4'b1011 : 4'b1010;
														assign node2246 = (inp[5]) ? 4'b1010 : 4'b1011;
									assign node2249 = (inp[7]) ? node2319 : node2250;
										assign node2250 = (inp[4]) ? node2284 : node2251;
											assign node2251 = (inp[15]) ? node2263 : node2252;
												assign node2252 = (inp[5]) ? node2260 : node2253;
													assign node2253 = (inp[0]) ? 4'b1110 : node2254;
														assign node2254 = (inp[10]) ? node2256 : 4'b1110;
															assign node2256 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node2260 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node2263 = (inp[5]) ? node2275 : node2264;
													assign node2264 = (inp[10]) ? node2270 : node2265;
														assign node2265 = (inp[11]) ? 4'b1101 : node2266;
															assign node2266 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node2270 = (inp[11]) ? 4'b1100 : node2271;
															assign node2271 = (inp[0]) ? 4'b1100 : 4'b1100;
													assign node2275 = (inp[0]) ? 4'b1100 : node2276;
														assign node2276 = (inp[9]) ? node2280 : node2277;
															assign node2277 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node2280 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node2284 = (inp[11]) ? node2298 : node2285;
												assign node2285 = (inp[15]) ? node2289 : node2286;
													assign node2286 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node2289 = (inp[5]) ? 4'b1011 : node2290;
														assign node2290 = (inp[10]) ? node2294 : node2291;
															assign node2291 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node2294 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node2298 = (inp[15]) ? node2310 : node2299;
													assign node2299 = (inp[5]) ? node2305 : node2300;
														assign node2300 = (inp[10]) ? 4'b1010 : node2301;
															assign node2301 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node2305 = (inp[9]) ? node2307 : 4'b1110;
															assign node2307 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node2310 = (inp[5]) ? node2314 : node2311;
														assign node2311 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node2314 = (inp[0]) ? node2316 : 4'b1011;
															assign node2316 = (inp[10]) ? 4'b1010 : 4'b1010;
										assign node2319 = (inp[4]) ? node2347 : node2320;
											assign node2320 = (inp[15]) ? node2336 : node2321;
												assign node2321 = (inp[11]) ? node2325 : node2322;
													assign node2322 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node2325 = (inp[9]) ? node2331 : node2326;
														assign node2326 = (inp[10]) ? 4'b1101 : node2327;
															assign node2327 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node2331 = (inp[0]) ? 4'b1100 : node2332;
															assign node2332 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node2336 = (inp[11]) ? node2342 : node2337;
													assign node2337 = (inp[5]) ? node2339 : 4'b1011;
														assign node2339 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node2342 = (inp[10]) ? node2344 : 4'b1011;
														assign node2344 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node2347 = (inp[5]) ? node2361 : node2348;
												assign node2348 = (inp[0]) ? node2354 : node2349;
													assign node2349 = (inp[10]) ? node2351 : 4'b1001;
														assign node2351 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node2354 = (inp[9]) ? 4'b1001 : node2355;
														assign node2355 = (inp[11]) ? node2357 : 4'b1000;
															assign node2357 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node2361 = (inp[9]) ? node2371 : node2362;
													assign node2362 = (inp[11]) ? node2368 : node2363;
														assign node2363 = (inp[0]) ? 4'b1001 : node2364;
															assign node2364 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node2368 = (inp[15]) ? 4'b1001 : 4'b1000;
													assign node2371 = (inp[10]) ? 4'b1000 : node2372;
														assign node2372 = (inp[15]) ? 4'b1000 : 4'b1001;
							assign node2376 = (inp[1]) ? node2618 : node2377;
								assign node2377 = (inp[5]) ? node2489 : node2378;
									assign node2378 = (inp[4]) ? node2446 : node2379;
										assign node2379 = (inp[7]) ? node2407 : node2380;
											assign node2380 = (inp[0]) ? node2390 : node2381;
												assign node2381 = (inp[15]) ? 4'b1110 : node2382;
													assign node2382 = (inp[12]) ? 4'b1110 : node2383;
														assign node2383 = (inp[11]) ? node2385 : 4'b1100;
															assign node2385 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node2390 = (inp[15]) ? node2400 : node2391;
													assign node2391 = (inp[12]) ? node2397 : node2392;
														assign node2392 = (inp[9]) ? node2394 : 4'b1101;
															assign node2394 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node2397 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node2400 = (inp[12]) ? node2402 : 4'b1111;
														assign node2402 = (inp[9]) ? 4'b1001 : node2403;
															assign node2403 = (inp[10]) ? 4'b1000 : 4'b1001;
											assign node2407 = (inp[9]) ? node2425 : node2408;
												assign node2408 = (inp[12]) ? node2418 : node2409;
													assign node2409 = (inp[15]) ? node2413 : node2410;
														assign node2410 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node2413 = (inp[11]) ? node2415 : 4'b1001;
															assign node2415 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node2418 = (inp[0]) ? node2420 : 4'b1110;
														assign node2420 = (inp[11]) ? node2422 : 4'b1111;
															assign node2422 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node2425 = (inp[10]) ? node2435 : node2426;
													assign node2426 = (inp[0]) ? node2428 : 4'b1000;
														assign node2428 = (inp[12]) ? node2432 : node2429;
															assign node2429 = (inp[15]) ? 4'b1000 : 4'b1110;
															assign node2432 = (inp[15]) ? 4'b1110 : 4'b1000;
													assign node2435 = (inp[11]) ? node2441 : node2436;
														assign node2436 = (inp[15]) ? 4'b1001 : node2437;
															assign node2437 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node2441 = (inp[0]) ? 4'b1001 : node2442;
															assign node2442 = (inp[15]) ? 4'b1000 : 4'b1001;
										assign node2446 = (inp[7]) ? node2466 : node2447;
											assign node2447 = (inp[12]) ? node2457 : node2448;
												assign node2448 = (inp[15]) ? 4'b1001 : node2449;
													assign node2449 = (inp[11]) ? node2451 : 4'b1101;
														assign node2451 = (inp[10]) ? node2453 : 4'b1100;
															assign node2453 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node2457 = (inp[15]) ? node2461 : node2458;
													assign node2458 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node2461 = (inp[0]) ? 4'b1110 : node2462;
														assign node2462 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node2466 = (inp[12]) ? node2484 : node2467;
												assign node2467 = (inp[15]) ? node2473 : node2468;
													assign node2468 = (inp[11]) ? 4'b1110 : node2469;
														assign node2469 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node2473 = (inp[0]) ? node2479 : node2474;
														assign node2474 = (inp[9]) ? node2476 : 4'b1111;
															assign node2476 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node2479 = (inp[9]) ? node2481 : 4'b1110;
															assign node2481 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node2484 = (inp[0]) ? node2486 : 4'b1100;
													assign node2486 = (inp[9]) ? 4'b1101 : 4'b1100;
									assign node2489 = (inp[7]) ? node2553 : node2490;
										assign node2490 = (inp[12]) ? node2522 : node2491;
											assign node2491 = (inp[4]) ? node2511 : node2492;
												assign node2492 = (inp[15]) ? node2500 : node2493;
													assign node2493 = (inp[11]) ? node2495 : 4'b1000;
														assign node2495 = (inp[10]) ? 4'b1001 : node2496;
															assign node2496 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node2500 = (inp[11]) ? node2506 : node2501;
														assign node2501 = (inp[0]) ? node2503 : 4'b1011;
															assign node2503 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node2506 = (inp[10]) ? node2508 : 4'b1010;
															assign node2508 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node2511 = (inp[15]) ? node2515 : node2512;
													assign node2512 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node2515 = (inp[0]) ? 4'b1101 : node2516;
														assign node2516 = (inp[11]) ? node2518 : 4'b1101;
															assign node2518 = (inp[10]) ? 4'b1100 : 4'b1100;
											assign node2522 = (inp[15]) ? node2534 : node2523;
												assign node2523 = (inp[4]) ? node2531 : node2524;
													assign node2524 = (inp[10]) ? node2526 : 4'b1111;
														assign node2526 = (inp[11]) ? 4'b1111 : node2527;
															assign node2527 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node2531 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node2534 = (inp[4]) ? node2542 : node2535;
													assign node2535 = (inp[10]) ? node2539 : node2536;
														assign node2536 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node2539 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node2542 = (inp[9]) ? node2548 : node2543;
														assign node2543 = (inp[0]) ? 4'b1111 : node2544;
															assign node2544 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node2548 = (inp[10]) ? node2550 : 4'b1110;
															assign node2550 = (inp[11]) ? 4'b1110 : 4'b1111;
										assign node2553 = (inp[12]) ? node2581 : node2554;
											assign node2554 = (inp[15]) ? node2574 : node2555;
												assign node2555 = (inp[4]) ? node2563 : node2556;
													assign node2556 = (inp[10]) ? 4'b1011 : node2557;
														assign node2557 = (inp[9]) ? node2559 : 4'b1010;
															assign node2559 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node2563 = (inp[0]) ? node2569 : node2564;
														assign node2564 = (inp[9]) ? node2566 : 4'b1011;
															assign node2566 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node2569 = (inp[10]) ? 4'b1010 : node2570;
															assign node2570 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node2574 = (inp[4]) ? node2578 : node2575;
													assign node2575 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node2578 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node2581 = (inp[4]) ? node2599 : node2582;
												assign node2582 = (inp[15]) ? node2588 : node2583;
													assign node2583 = (inp[9]) ? 4'b1101 : node2584;
														assign node2584 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node2588 = (inp[9]) ? node2594 : node2589;
														assign node2589 = (inp[11]) ? 4'b1011 : node2590;
															assign node2590 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node2594 = (inp[0]) ? 4'b1010 : node2595;
															assign node2595 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node2599 = (inp[15]) ? node2607 : node2600;
													assign node2600 = (inp[11]) ? node2602 : 4'b1000;
														assign node2602 = (inp[10]) ? node2604 : 4'b1000;
															assign node2604 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node2607 = (inp[11]) ? node2613 : node2608;
														assign node2608 = (inp[9]) ? node2610 : 4'b1001;
															assign node2610 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node2613 = (inp[0]) ? node2615 : 4'b1000;
															assign node2615 = (inp[10]) ? 4'b1000 : 4'b1001;
								assign node2618 = (inp[7]) ? node2736 : node2619;
									assign node2619 = (inp[12]) ? node2677 : node2620;
										assign node2620 = (inp[15]) ? node2652 : node2621;
											assign node2621 = (inp[10]) ? node2633 : node2622;
												assign node2622 = (inp[0]) ? 4'b1101 : node2623;
													assign node2623 = (inp[5]) ? 4'b1101 : node2624;
														assign node2624 = (inp[4]) ? node2628 : node2625;
															assign node2625 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node2628 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node2633 = (inp[5]) ? node2643 : node2634;
													assign node2634 = (inp[0]) ? node2640 : node2635;
														assign node2635 = (inp[11]) ? node2637 : 4'b1101;
															assign node2637 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node2640 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node2643 = (inp[4]) ? node2645 : 4'b1100;
														assign node2645 = (inp[9]) ? node2649 : node2646;
															assign node2646 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node2649 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node2652 = (inp[4]) ? node2664 : node2653;
												assign node2653 = (inp[11]) ? 4'b1110 : node2654;
													assign node2654 = (inp[5]) ? node2658 : node2655;
														assign node2655 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node2658 = (inp[9]) ? node2660 : 4'b1110;
															assign node2660 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node2664 = (inp[5]) ? node2666 : 4'b1001;
													assign node2666 = (inp[9]) ? node2672 : node2667;
														assign node2667 = (inp[10]) ? 4'b1000 : node2668;
															assign node2668 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node2672 = (inp[10]) ? 4'b1001 : node2673;
															assign node2673 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node2677 = (inp[4]) ? node2705 : node2678;
											assign node2678 = (inp[15]) ? node2692 : node2679;
												assign node2679 = (inp[5]) ? node2685 : node2680;
													assign node2680 = (inp[11]) ? 4'b1011 : node2681;
														assign node2681 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node2685 = (inp[9]) ? node2689 : node2686;
														assign node2686 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node2689 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node2692 = (inp[10]) ? node2700 : node2693;
													assign node2693 = (inp[11]) ? node2695 : 4'b1001;
														assign node2695 = (inp[9]) ? node2697 : 4'b1000;
															assign node2697 = (inp[5]) ? 4'b1000 : 4'b1001;
													assign node2700 = (inp[9]) ? 4'b1000 : node2701;
														assign node2701 = (inp[5]) ? 4'b1000 : 4'b1001;
											assign node2705 = (inp[0]) ? node2717 : node2706;
												assign node2706 = (inp[11]) ? node2712 : node2707;
													assign node2707 = (inp[10]) ? 4'b1111 : node2708;
														assign node2708 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node2712 = (inp[9]) ? node2714 : 4'b1010;
														assign node2714 = (inp[5]) ? 4'b1111 : 4'b1011;
												assign node2717 = (inp[11]) ? node2725 : node2718;
													assign node2718 = (inp[15]) ? node2722 : node2719;
														assign node2719 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node2722 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node2725 = (inp[15]) ? node2731 : node2726;
														assign node2726 = (inp[10]) ? node2728 : 4'b1011;
															assign node2728 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node2731 = (inp[5]) ? node2733 : 4'b1011;
															assign node2733 = (inp[10]) ? 4'b1110 : 4'b1110;
									assign node2736 = (inp[12]) ? node2796 : node2737;
										assign node2737 = (inp[15]) ? node2775 : node2738;
											assign node2738 = (inp[4]) ? node2760 : node2739;
												assign node2739 = (inp[10]) ? node2751 : node2740;
													assign node2740 = (inp[9]) ? node2746 : node2741;
														assign node2741 = (inp[5]) ? node2743 : 4'b1110;
															assign node2743 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node2746 = (inp[11]) ? node2748 : 4'b1111;
															assign node2748 = (inp[5]) ? 4'b1110 : 4'b1111;
													assign node2751 = (inp[9]) ? 4'b1110 : node2752;
														assign node2752 = (inp[0]) ? node2756 : node2753;
															assign node2753 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node2756 = (inp[5]) ? 4'b1111 : 4'b1110;
												assign node2760 = (inp[0]) ? node2768 : node2761;
													assign node2761 = (inp[5]) ? node2763 : 4'b1111;
														assign node2763 = (inp[9]) ? 4'b1110 : node2764;
															assign node2764 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node2768 = (inp[5]) ? node2770 : 4'b1110;
														assign node2770 = (inp[9]) ? 4'b1110 : node2771;
															assign node2771 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node2775 = (inp[4]) ? node2785 : node2776;
												assign node2776 = (inp[5]) ? node2780 : node2777;
													assign node2777 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node2780 = (inp[10]) ? node2782 : 4'b1000;
														assign node2782 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node2785 = (inp[5]) ? 4'b1110 : node2786;
													assign node2786 = (inp[0]) ? 4'b1111 : node2787;
														assign node2787 = (inp[11]) ? node2791 : node2788;
															assign node2788 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node2791 = (inp[10]) ? 4'b1110 : 4'b1111;
										assign node2796 = (inp[4]) ? node2814 : node2797;
											assign node2797 = (inp[15]) ? node2807 : node2798;
												assign node2798 = (inp[9]) ? node2804 : node2799;
													assign node2799 = (inp[0]) ? 4'b1001 : node2800;
														assign node2800 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node2804 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node2807 = (inp[10]) ? node2809 : 4'b1111;
													assign node2809 = (inp[5]) ? node2811 : 4'b1111;
														assign node2811 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node2814 = (inp[0]) ? node2828 : node2815;
												assign node2815 = (inp[10]) ? node2821 : node2816;
													assign node2816 = (inp[15]) ? 4'b1101 : node2817;
														assign node2817 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node2821 = (inp[11]) ? 4'b1101 : node2822;
														assign node2822 = (inp[15]) ? 4'b1100 : node2823;
															assign node2823 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node2828 = (inp[15]) ? node2836 : node2829;
													assign node2829 = (inp[9]) ? node2831 : 4'b1100;
														assign node2831 = (inp[11]) ? 4'b1101 : node2832;
															assign node2832 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node2836 = (inp[11]) ? node2844 : node2837;
														assign node2837 = (inp[5]) ? node2841 : node2838;
															assign node2838 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node2841 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node2844 = (inp[9]) ? 4'b1100 : node2845;
															assign node2845 = (inp[10]) ? 4'b1101 : 4'b1100;
						assign node2849 = (inp[2]) ? node3291 : node2850;
							assign node2850 = (inp[5]) ? node3070 : node2851;
								assign node2851 = (inp[7]) ? node2961 : node2852;
									assign node2852 = (inp[12]) ? node2902 : node2853;
										assign node2853 = (inp[4]) ? node2883 : node2854;
											assign node2854 = (inp[15]) ? node2870 : node2855;
												assign node2855 = (inp[0]) ? node2861 : node2856;
													assign node2856 = (inp[10]) ? node2858 : 4'b1101;
														assign node2858 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node2861 = (inp[11]) ? node2865 : node2862;
														assign node2862 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node2865 = (inp[10]) ? node2867 : 4'b1100;
															assign node2867 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node2870 = (inp[1]) ? node2878 : node2871;
													assign node2871 = (inp[11]) ? node2873 : 4'b1111;
														assign node2873 = (inp[10]) ? node2875 : 4'b1110;
															assign node2875 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node2878 = (inp[10]) ? 4'b1110 : node2879;
														assign node2879 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node2883 = (inp[15]) ? node2893 : node2884;
												assign node2884 = (inp[9]) ? 4'b1100 : node2885;
													assign node2885 = (inp[10]) ? 4'b1101 : node2886;
														assign node2886 = (inp[11]) ? node2888 : 4'b1100;
															assign node2888 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node2893 = (inp[9]) ? node2899 : node2894;
													assign node2894 = (inp[11]) ? 4'b1000 : node2895;
														assign node2895 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node2899 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node2902 = (inp[1]) ? node2930 : node2903;
											assign node2903 = (inp[11]) ? node2919 : node2904;
												assign node2904 = (inp[9]) ? node2910 : node2905;
													assign node2905 = (inp[15]) ? 4'b1000 : node2906;
														assign node2906 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node2910 = (inp[15]) ? node2914 : node2911;
														assign node2911 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node2914 = (inp[10]) ? 4'b1111 : node2915;
															assign node2915 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node2919 = (inp[15]) ? node2927 : node2920;
													assign node2920 = (inp[4]) ? node2922 : 4'b1110;
														assign node2922 = (inp[9]) ? node2924 : 4'b1010;
															assign node2924 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node2927 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node2930 = (inp[4]) ? node2942 : node2931;
												assign node2931 = (inp[15]) ? node2935 : node2932;
													assign node2932 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node2935 = (inp[11]) ? 4'b1001 : node2936;
														assign node2936 = (inp[0]) ? 4'b1000 : node2937;
															assign node2937 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node2942 = (inp[15]) ? node2950 : node2943;
													assign node2943 = (inp[10]) ? node2945 : 4'b1110;
														assign node2945 = (inp[0]) ? 4'b1111 : node2946;
															assign node2946 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node2950 = (inp[9]) ? node2956 : node2951;
														assign node2951 = (inp[0]) ? 4'b1011 : node2952;
															assign node2952 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node2956 = (inp[10]) ? 4'b1010 : node2957;
															assign node2957 = (inp[0]) ? 4'b1010 : 4'b1010;
									assign node2961 = (inp[12]) ? node3021 : node2962;
										assign node2962 = (inp[15]) ? node2998 : node2963;
											assign node2963 = (inp[4]) ? node2983 : node2964;
												assign node2964 = (inp[0]) ? node2974 : node2965;
													assign node2965 = (inp[9]) ? node2967 : 4'b1111;
														assign node2967 = (inp[10]) ? node2971 : node2968;
															assign node2968 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node2971 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node2974 = (inp[1]) ? node2976 : 4'b1110;
														assign node2976 = (inp[11]) ? node2980 : node2977;
															assign node2977 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node2980 = (inp[9]) ? 4'b1110 : 4'b1110;
												assign node2983 = (inp[10]) ? node2991 : node2984;
													assign node2984 = (inp[1]) ? node2986 : 4'b1111;
														assign node2986 = (inp[11]) ? node2988 : 4'b1111;
															assign node2988 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node2991 = (inp[0]) ? 4'b1110 : node2992;
														assign node2992 = (inp[1]) ? 4'b1111 : node2993;
															assign node2993 = (inp[9]) ? 4'b1110 : 4'b1110;
											assign node2998 = (inp[4]) ? node3010 : node2999;
												assign node2999 = (inp[1]) ? node3003 : node3000;
													assign node3000 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node3003 = (inp[10]) ? node3007 : node3004;
														assign node3004 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node3007 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node3010 = (inp[0]) ? node3012 : 4'b1110;
													assign node3012 = (inp[11]) ? 4'b1111 : node3013;
														assign node3013 = (inp[10]) ? node3017 : node3014;
															assign node3014 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node3017 = (inp[9]) ? 4'b1110 : 4'b1111;
										assign node3021 = (inp[15]) ? node3047 : node3022;
											assign node3022 = (inp[4]) ? node3032 : node3023;
												assign node3023 = (inp[1]) ? node3025 : 4'b1000;
													assign node3025 = (inp[10]) ? 4'b1001 : node3026;
														assign node3026 = (inp[9]) ? node3028 : 4'b1000;
															assign node3028 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node3032 = (inp[11]) ? node3034 : 4'b1100;
													assign node3034 = (inp[9]) ? node3042 : node3035;
														assign node3035 = (inp[0]) ? node3039 : node3036;
															assign node3036 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node3039 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node3042 = (inp[10]) ? node3044 : 4'b1101;
															assign node3044 = (inp[1]) ? 4'b1100 : 4'b1101;
											assign node3047 = (inp[4]) ? node3061 : node3048;
												assign node3048 = (inp[0]) ? node3056 : node3049;
													assign node3049 = (inp[9]) ? 4'b1111 : node3050;
														assign node3050 = (inp[10]) ? node3052 : 4'b1111;
															assign node3052 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node3056 = (inp[9]) ? 4'b1110 : node3057;
														assign node3057 = (inp[1]) ? 4'b1110 : 4'b1111;
												assign node3061 = (inp[0]) ? node3063 : 4'b1100;
													assign node3063 = (inp[10]) ? node3065 : 4'b1101;
														assign node3065 = (inp[1]) ? 4'b1100 : node3066;
															assign node3066 = (inp[9]) ? 4'b1100 : 4'b1100;
								assign node3070 = (inp[1]) ? node3186 : node3071;
									assign node3071 = (inp[7]) ? node3129 : node3072;
										assign node3072 = (inp[12]) ? node3106 : node3073;
											assign node3073 = (inp[4]) ? node3089 : node3074;
												assign node3074 = (inp[15]) ? node3082 : node3075;
													assign node3075 = (inp[9]) ? node3077 : 4'b1000;
														assign node3077 = (inp[0]) ? node3079 : 4'b1001;
															assign node3079 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node3082 = (inp[9]) ? node3086 : node3083;
														assign node3083 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node3086 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node3089 = (inp[15]) ? node3097 : node3090;
													assign node3090 = (inp[9]) ? 4'b1001 : node3091;
														assign node3091 = (inp[10]) ? 4'b1000 : node3092;
															assign node3092 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node3097 = (inp[10]) ? node3103 : node3098;
														assign node3098 = (inp[9]) ? 4'b1101 : node3099;
															assign node3099 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node3103 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node3106 = (inp[4]) ? node3118 : node3107;
												assign node3107 = (inp[15]) ? 4'b1101 : node3108;
													assign node3108 = (inp[10]) ? node3112 : node3109;
														assign node3109 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node3112 = (inp[9]) ? node3114 : 4'b1111;
															assign node3114 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node3118 = (inp[15]) ? node3126 : node3119;
													assign node3119 = (inp[9]) ? node3121 : 4'b1011;
														assign node3121 = (inp[11]) ? 4'b1010 : node3122;
															assign node3122 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node3126 = (inp[9]) ? 4'b1110 : 4'b1111;
										assign node3129 = (inp[12]) ? node3157 : node3130;
											assign node3130 = (inp[4]) ? node3146 : node3131;
												assign node3131 = (inp[15]) ? node3139 : node3132;
													assign node3132 = (inp[0]) ? 4'b1010 : node3133;
														assign node3133 = (inp[11]) ? node3135 : 4'b1011;
															assign node3135 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node3139 = (inp[9]) ? node3143 : node3140;
														assign node3140 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node3143 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node3146 = (inp[15]) ? node3154 : node3147;
													assign node3147 = (inp[10]) ? node3149 : 4'b1010;
														assign node3149 = (inp[0]) ? 4'b1010 : node3150;
															assign node3150 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node3154 = (inp[10]) ? 4'b1010 : 4'b1011;
											assign node3157 = (inp[4]) ? node3167 : node3158;
												assign node3158 = (inp[15]) ? node3164 : node3159;
													assign node3159 = (inp[10]) ? 4'b1101 : node3160;
														assign node3160 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node3164 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node3167 = (inp[0]) ? node3179 : node3168;
													assign node3168 = (inp[11]) ? node3174 : node3169;
														assign node3169 = (inp[10]) ? node3171 : 4'b1000;
															assign node3171 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node3174 = (inp[10]) ? node3176 : 4'b1001;
															assign node3176 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node3179 = (inp[15]) ? node3181 : 4'b1001;
														assign node3181 = (inp[9]) ? 4'b1000 : node3182;
															assign node3182 = (inp[11]) ? 4'b1000 : 4'b1001;
									assign node3186 = (inp[9]) ? node3230 : node3187;
										assign node3187 = (inp[15]) ? node3211 : node3188;
											assign node3188 = (inp[12]) ? node3198 : node3189;
												assign node3189 = (inp[7]) ? node3195 : node3190;
													assign node3190 = (inp[10]) ? 4'b1101 : node3191;
														assign node3191 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node3195 = (inp[4]) ? 4'b1111 : 4'b1110;
												assign node3198 = (inp[7]) ? node3200 : 4'b1111;
													assign node3200 = (inp[4]) ? node3208 : node3201;
														assign node3201 = (inp[10]) ? node3205 : node3202;
															assign node3202 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node3205 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node3208 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node3211 = (inp[4]) ? node3223 : node3212;
												assign node3212 = (inp[10]) ? node3218 : node3213;
													assign node3213 = (inp[11]) ? 4'b1001 : node3214;
														assign node3214 = (inp[12]) ? 4'b1111 : 4'b1110;
													assign node3218 = (inp[7]) ? 4'b1110 : node3219;
														assign node3219 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node3223 = (inp[10]) ? node3225 : 4'b1110;
													assign node3225 = (inp[11]) ? node3227 : 4'b1000;
														assign node3227 = (inp[0]) ? 4'b1000 : 4'b1110;
										assign node3230 = (inp[15]) ? node3268 : node3231;
											assign node3231 = (inp[12]) ? node3253 : node3232;
												assign node3232 = (inp[7]) ? node3242 : node3233;
													assign node3233 = (inp[4]) ? node3237 : node3234;
														assign node3234 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node3237 = (inp[10]) ? 4'b1101 : node3238;
															assign node3238 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node3242 = (inp[10]) ? node3248 : node3243;
														assign node3243 = (inp[11]) ? 4'b1110 : node3244;
															assign node3244 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node3248 = (inp[0]) ? node3250 : 4'b1111;
															assign node3250 = (inp[4]) ? 4'b1110 : 4'b1111;
												assign node3253 = (inp[7]) ? node3259 : node3254;
													assign node3254 = (inp[4]) ? node3256 : 4'b1111;
														assign node3256 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node3259 = (inp[4]) ? node3263 : node3260;
														assign node3260 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node3263 = (inp[10]) ? 4'b1100 : node3264;
															assign node3264 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node3268 = (inp[12]) ? node3282 : node3269;
												assign node3269 = (inp[7]) ? node3279 : node3270;
													assign node3270 = (inp[4]) ? node3274 : node3271;
														assign node3271 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node3274 = (inp[0]) ? 4'b1001 : node3275;
															assign node3275 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node3279 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node3282 = (inp[11]) ? node3284 : 4'b1001;
													assign node3284 = (inp[0]) ? 4'b1100 : node3285;
														assign node3285 = (inp[7]) ? node3287 : 4'b1111;
															assign node3287 = (inp[4]) ? 4'b1100 : 4'b1111;
							assign node3291 = (inp[1]) ? node3483 : node3292;
								assign node3292 = (inp[5]) ? node3386 : node3293;
									assign node3293 = (inp[15]) ? node3325 : node3294;
										assign node3294 = (inp[12]) ? node3310 : node3295;
											assign node3295 = (inp[7]) ? node3301 : node3296;
												assign node3296 = (inp[10]) ? node3298 : 4'b1001;
													assign node3298 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node3301 = (inp[11]) ? node3303 : 4'b1011;
													assign node3303 = (inp[10]) ? node3305 : 4'b1011;
														assign node3305 = (inp[9]) ? 4'b1010 : node3306;
															assign node3306 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node3310 = (inp[7]) ? node3318 : node3311;
												assign node3311 = (inp[4]) ? 4'b1111 : node3312;
													assign node3312 = (inp[10]) ? node3314 : 4'b1011;
														assign node3314 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node3318 = (inp[4]) ? node3322 : node3319;
													assign node3319 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node3322 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node3325 = (inp[7]) ? node3361 : node3326;
											assign node3326 = (inp[9]) ? node3342 : node3327;
												assign node3327 = (inp[11]) ? node3335 : node3328;
													assign node3328 = (inp[0]) ? node3330 : 4'b1101;
														assign node3330 = (inp[10]) ? node3332 : 4'b1010;
															assign node3332 = (inp[4]) ? 4'b1011 : 4'b1101;
													assign node3335 = (inp[4]) ? node3339 : node3336;
														assign node3336 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node3339 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node3342 = (inp[0]) ? node3350 : node3343;
													assign node3343 = (inp[12]) ? node3347 : node3344;
														assign node3344 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node3347 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node3350 = (inp[10]) ? node3356 : node3351;
														assign node3351 = (inp[4]) ? node3353 : 4'b1101;
															assign node3353 = (inp[12]) ? 4'b1010 : 4'b1100;
														assign node3356 = (inp[11]) ? node3358 : 4'b1010;
															assign node3358 = (inp[12]) ? 4'b1100 : 4'b1101;
											assign node3361 = (inp[12]) ? node3371 : node3362;
												assign node3362 = (inp[4]) ? node3368 : node3363;
													assign node3363 = (inp[0]) ? 4'b1100 : node3364;
														assign node3364 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node3368 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node3371 = (inp[4]) ? node3383 : node3372;
													assign node3372 = (inp[9]) ? node3378 : node3373;
														assign node3373 = (inp[11]) ? node3375 : 4'b1010;
															assign node3375 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node3378 = (inp[0]) ? 4'b1011 : node3379;
															assign node3379 = (inp[10]) ? 4'b1010 : 4'b1010;
													assign node3383 = (inp[9]) ? 4'b1001 : 4'b1000;
									assign node3386 = (inp[12]) ? node3438 : node3387;
										assign node3387 = (inp[7]) ? node3413 : node3388;
											assign node3388 = (inp[4]) ? node3396 : node3389;
												assign node3389 = (inp[15]) ? node3391 : 4'b1101;
													assign node3391 = (inp[10]) ? 4'b1111 : node3392;
														assign node3392 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node3396 = (inp[15]) ? node3406 : node3397;
													assign node3397 = (inp[11]) ? node3403 : node3398;
														assign node3398 = (inp[0]) ? 4'b1101 : node3399;
															assign node3399 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node3403 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node3406 = (inp[10]) ? node3408 : 4'b1001;
														assign node3408 = (inp[0]) ? 4'b1000 : node3409;
															assign node3409 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node3413 = (inp[15]) ? node3429 : node3414;
												assign node3414 = (inp[4]) ? node3424 : node3415;
													assign node3415 = (inp[0]) ? node3417 : 4'b1111;
														assign node3417 = (inp[11]) ? node3421 : node3418;
															assign node3418 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node3421 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node3424 = (inp[10]) ? 4'b1110 : node3425;
														assign node3425 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node3429 = (inp[4]) ? node3435 : node3430;
													assign node3430 = (inp[0]) ? node3432 : 4'b1100;
														assign node3432 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node3435 = (inp[0]) ? 4'b1111 : 4'b1110;
										assign node3438 = (inp[7]) ? node3460 : node3439;
											assign node3439 = (inp[4]) ? node3453 : node3440;
												assign node3440 = (inp[15]) ? node3446 : node3441;
													assign node3441 = (inp[10]) ? 4'b1011 : node3442;
														assign node3442 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node3446 = (inp[0]) ? node3448 : 4'b1000;
														assign node3448 = (inp[9]) ? 4'b1001 : node3449;
															assign node3449 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node3453 = (inp[15]) ? node3457 : node3454;
													assign node3454 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node3457 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node3460 = (inp[4]) ? node3470 : node3461;
												assign node3461 = (inp[15]) ? 4'b1111 : node3462;
													assign node3462 = (inp[11]) ? 4'b1001 : node3463;
														assign node3463 = (inp[9]) ? 4'b1000 : node3464;
															assign node3464 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node3470 = (inp[10]) ? node3478 : node3471;
													assign node3471 = (inp[9]) ? 4'b1101 : node3472;
														assign node3472 = (inp[0]) ? 4'b1101 : node3473;
															assign node3473 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node3478 = (inp[9]) ? 4'b1100 : node3479;
														assign node3479 = (inp[11]) ? 4'b1101 : 4'b1100;
								assign node3483 = (inp[7]) ? node3623 : node3484;
									assign node3484 = (inp[12]) ? node3536 : node3485;
										assign node3485 = (inp[4]) ? node3511 : node3486;
											assign node3486 = (inp[15]) ? node3496 : node3487;
												assign node3487 = (inp[11]) ? 4'b1001 : node3488;
													assign node3488 = (inp[9]) ? node3490 : 4'b1000;
														assign node3490 = (inp[10]) ? 4'b1001 : node3491;
															assign node3491 = (inp[5]) ? 4'b1000 : 4'b1000;
												assign node3496 = (inp[5]) ? node3502 : node3497;
													assign node3497 = (inp[0]) ? node3499 : 4'b1010;
														assign node3499 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node3502 = (inp[11]) ? node3508 : node3503;
														assign node3503 = (inp[10]) ? node3505 : 4'b1011;
															assign node3505 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node3508 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node3511 = (inp[15]) ? node3523 : node3512;
												assign node3512 = (inp[5]) ? node3518 : node3513;
													assign node3513 = (inp[10]) ? node3515 : 4'b1001;
														assign node3515 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node3518 = (inp[11]) ? 4'b1000 : node3519;
														assign node3519 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node3523 = (inp[9]) ? node3531 : node3524;
													assign node3524 = (inp[10]) ? 4'b1100 : node3525;
														assign node3525 = (inp[11]) ? 4'b1101 : node3526;
															assign node3526 = (inp[5]) ? 4'b1100 : 4'b1100;
													assign node3531 = (inp[0]) ? 4'b1101 : node3532;
														assign node3532 = (inp[10]) ? 4'b1101 : 4'b1100;
										assign node3536 = (inp[4]) ? node3570 : node3537;
											assign node3537 = (inp[15]) ? node3553 : node3538;
												assign node3538 = (inp[5]) ? node3544 : node3539;
													assign node3539 = (inp[11]) ? node3541 : 4'b1111;
														assign node3541 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node3544 = (inp[11]) ? node3546 : 4'b1011;
														assign node3546 = (inp[0]) ? node3550 : node3547;
															assign node3547 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node3550 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node3553 = (inp[5]) ? node3559 : node3554;
													assign node3554 = (inp[0]) ? node3556 : 4'b1101;
														assign node3556 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node3559 = (inp[11]) ? node3565 : node3560;
														assign node3560 = (inp[9]) ? 4'b1101 : node3561;
															assign node3561 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node3565 = (inp[9]) ? 4'b1100 : node3566;
															assign node3566 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node3570 = (inp[11]) ? node3598 : node3571;
												assign node3571 = (inp[15]) ? node3583 : node3572;
													assign node3572 = (inp[5]) ? node3578 : node3573;
														assign node3573 = (inp[10]) ? 4'b1011 : node3574;
															assign node3574 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node3578 = (inp[9]) ? node3580 : 4'b1111;
															assign node3580 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node3583 = (inp[5]) ? node3591 : node3584;
														assign node3584 = (inp[0]) ? node3588 : node3585;
															assign node3585 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node3588 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node3591 = (inp[9]) ? node3595 : node3592;
															assign node3592 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node3595 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node3598 = (inp[10]) ? node3610 : node3599;
													assign node3599 = (inp[5]) ? node3605 : node3600;
														assign node3600 = (inp[15]) ? 4'b1110 : node3601;
															assign node3601 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node3605 = (inp[15]) ? 4'b1010 : node3606;
															assign node3606 = (inp[0]) ? 4'b1110 : 4'b1110;
													assign node3610 = (inp[0]) ? node3616 : node3611;
														assign node3611 = (inp[5]) ? node3613 : 4'b1111;
															assign node3613 = (inp[15]) ? 4'b1010 : 4'b1110;
														assign node3616 = (inp[15]) ? node3620 : node3617;
															assign node3617 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node3620 = (inp[9]) ? 4'b1010 : 4'b1011;
									assign node3623 = (inp[12]) ? node3667 : node3624;
										assign node3624 = (inp[15]) ? node3652 : node3625;
											assign node3625 = (inp[4]) ? node3639 : node3626;
												assign node3626 = (inp[10]) ? node3634 : node3627;
													assign node3627 = (inp[9]) ? 4'b1011 : node3628;
														assign node3628 = (inp[11]) ? node3630 : 4'b1011;
															assign node3630 = (inp[5]) ? 4'b1010 : 4'b1011;
													assign node3634 = (inp[5]) ? node3636 : 4'b1010;
														assign node3636 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node3639 = (inp[9]) ? node3643 : node3640;
													assign node3640 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node3643 = (inp[0]) ? node3649 : node3644;
														assign node3644 = (inp[11]) ? node3646 : 4'b1010;
															assign node3646 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node3649 = (inp[10]) ? 4'b1010 : 4'b1011;
											assign node3652 = (inp[4]) ? node3660 : node3653;
												assign node3653 = (inp[10]) ? 4'b1100 : node3654;
													assign node3654 = (inp[9]) ? 4'b1000 : node3655;
														assign node3655 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node3660 = (inp[0]) ? 4'b1011 : node3661;
													assign node3661 = (inp[9]) ? 4'b1010 : node3662;
														assign node3662 = (inp[10]) ? 4'b1011 : 4'b1010;
										assign node3667 = (inp[4]) ? node3693 : node3668;
											assign node3668 = (inp[15]) ? node3676 : node3669;
												assign node3669 = (inp[10]) ? 4'b1100 : node3670;
													assign node3670 = (inp[9]) ? 4'b1101 : node3671;
														assign node3671 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node3676 = (inp[10]) ? node3686 : node3677;
													assign node3677 = (inp[11]) ? 4'b1011 : node3678;
														assign node3678 = (inp[5]) ? node3682 : node3679;
															assign node3679 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node3682 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node3686 = (inp[5]) ? 4'b1010 : node3687;
														assign node3687 = (inp[0]) ? 4'b1011 : node3688;
															assign node3688 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node3693 = (inp[10]) ? node3703 : node3694;
												assign node3694 = (inp[9]) ? node3698 : node3695;
													assign node3695 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node3698 = (inp[0]) ? 4'b1001 : node3699;
														assign node3699 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node3703 = (inp[0]) ? node3705 : 4'b1001;
													assign node3705 = (inp[9]) ? 4'b1000 : 4'b1001;
				assign node3708 = (inp[7]) ? node5458 : node3709;
					assign node3709 = (inp[10]) ? node4555 : node3710;
						assign node3710 = (inp[0]) ? node4148 : node3711;
							assign node3711 = (inp[13]) ? node3921 : node3712;
								assign node3712 = (inp[14]) ? node3800 : node3713;
									assign node3713 = (inp[15]) ? node3749 : node3714;
										assign node3714 = (inp[12]) ? node3734 : node3715;
											assign node3715 = (inp[4]) ? node3727 : node3716;
												assign node3716 = (inp[11]) ? node3722 : node3717;
													assign node3717 = (inp[1]) ? node3719 : 4'b1000;
														assign node3719 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node3722 = (inp[1]) ? 4'b1001 : node3723;
														assign node3723 = (inp[2]) ? 4'b1100 : 4'b1000;
												assign node3727 = (inp[9]) ? 4'b1010 : node3728;
													assign node3728 = (inp[1]) ? node3730 : 4'b1111;
														assign node3730 = (inp[2]) ? 4'b1010 : 4'b1110;
											assign node3734 = (inp[4]) ? node3740 : node3735;
												assign node3735 = (inp[11]) ? 4'b1010 : node3736;
													assign node3736 = (inp[1]) ? 4'b1011 : 4'b1110;
												assign node3740 = (inp[5]) ? 4'b1001 : node3741;
													assign node3741 = (inp[1]) ? node3743 : 4'b1100;
														assign node3743 = (inp[2]) ? 4'b1100 : node3744;
															assign node3744 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node3749 = (inp[2]) ? node3781 : node3750;
											assign node3750 = (inp[1]) ? node3762 : node3751;
												assign node3751 = (inp[4]) ? node3755 : node3752;
													assign node3752 = (inp[12]) ? 4'b1010 : 4'b1000;
													assign node3755 = (inp[12]) ? 4'b1001 : node3756;
														assign node3756 = (inp[11]) ? 4'b1111 : node3757;
															assign node3757 = (inp[5]) ? 4'b1110 : 4'b1010;
												assign node3762 = (inp[5]) ? node3772 : node3763;
													assign node3763 = (inp[9]) ? node3767 : node3764;
														assign node3764 = (inp[4]) ? 4'b1111 : 4'b1101;
														assign node3767 = (inp[11]) ? 4'b1110 : node3768;
															assign node3768 = (inp[4]) ? 4'b1110 : 4'b1111;
													assign node3772 = (inp[4]) ? node3776 : node3773;
														assign node3773 = (inp[11]) ? 4'b1110 : 4'b1100;
														assign node3776 = (inp[12]) ? node3778 : 4'b1011;
															assign node3778 = (inp[9]) ? 4'b1101 : 4'b1100;
											assign node3781 = (inp[1]) ? node3793 : node3782;
												assign node3782 = (inp[5]) ? node3788 : node3783;
													assign node3783 = (inp[11]) ? 4'b1100 : node3784;
														assign node3784 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node3788 = (inp[12]) ? node3790 : 4'b1010;
														assign node3790 = (inp[4]) ? 4'b1100 : 4'b1110;
												assign node3793 = (inp[4]) ? node3797 : node3794;
													assign node3794 = (inp[9]) ? 4'b1001 : 4'b1010;
													assign node3797 = (inp[12]) ? 4'b1000 : 4'b1010;
									assign node3800 = (inp[1]) ? node3864 : node3801;
										assign node3801 = (inp[15]) ? node3837 : node3802;
											assign node3802 = (inp[5]) ? node3822 : node3803;
												assign node3803 = (inp[2]) ? node3813 : node3804;
													assign node3804 = (inp[11]) ? node3810 : node3805;
														assign node3805 = (inp[4]) ? node3807 : 4'b1000;
															assign node3807 = (inp[12]) ? 4'b1000 : 4'b1010;
														assign node3810 = (inp[4]) ? 4'b1011 : 4'b1001;
													assign node3813 = (inp[4]) ? node3817 : node3814;
														assign node3814 = (inp[12]) ? 4'b1110 : 4'b1100;
														assign node3817 = (inp[12]) ? node3819 : 4'b1111;
															assign node3819 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node3822 = (inp[2]) ? node3830 : node3823;
													assign node3823 = (inp[11]) ? node3825 : 4'b1100;
														assign node3825 = (inp[4]) ? node3827 : 4'b1010;
															assign node3827 = (inp[12]) ? 4'b1100 : 4'b1110;
													assign node3830 = (inp[4]) ? node3834 : node3831;
														assign node3831 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node3834 = (inp[12]) ? 4'b1000 : 4'b1010;
											assign node3837 = (inp[9]) ? node3851 : node3838;
												assign node3838 = (inp[5]) ? node3848 : node3839;
													assign node3839 = (inp[2]) ? node3843 : node3840;
														assign node3840 = (inp[11]) ? 4'b1111 : 4'b1100;
														assign node3843 = (inp[11]) ? 4'b1011 : node3844;
															assign node3844 = (inp[12]) ? 4'b1011 : 4'b1010;
													assign node3848 = (inp[12]) ? 4'b1110 : 4'b1010;
												assign node3851 = (inp[4]) ? node3859 : node3852;
													assign node3852 = (inp[12]) ? 4'b1111 : node3853;
														assign node3853 = (inp[5]) ? node3855 : 4'b1001;
															assign node3855 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node3859 = (inp[12]) ? node3861 : 4'b1011;
														assign node3861 = (inp[5]) ? 4'b1001 : 4'b1000;
										assign node3864 = (inp[2]) ? node3888 : node3865;
											assign node3865 = (inp[4]) ? node3877 : node3866;
												assign node3866 = (inp[12]) ? node3872 : node3867;
													assign node3867 = (inp[11]) ? 4'b1100 : node3868;
														assign node3868 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node3872 = (inp[15]) ? node3874 : 4'b1111;
														assign node3874 = (inp[5]) ? 4'b1110 : 4'b1010;
												assign node3877 = (inp[12]) ? node3885 : node3878;
													assign node3878 = (inp[15]) ? node3882 : node3879;
														assign node3879 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node3882 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node3885 = (inp[5]) ? 4'b1000 : 4'b1101;
											assign node3888 = (inp[4]) ? node3908 : node3889;
												assign node3889 = (inp[12]) ? node3899 : node3890;
													assign node3890 = (inp[15]) ? node3894 : node3891;
														assign node3891 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node3894 = (inp[11]) ? 4'b1001 : node3895;
															assign node3895 = (inp[5]) ? 4'b1000 : 4'b1001;
													assign node3899 = (inp[9]) ? node3901 : 4'b1010;
														assign node3901 = (inp[11]) ? node3905 : node3902;
															assign node3902 = (inp[5]) ? 4'b1011 : 4'b1110;
															assign node3905 = (inp[5]) ? 4'b1010 : 4'b1011;
												assign node3908 = (inp[12]) ? node3914 : node3909;
													assign node3909 = (inp[15]) ? 4'b1110 : node3910;
														assign node3910 = (inp[9]) ? 4'b1110 : 4'b1011;
													assign node3914 = (inp[15]) ? node3918 : node3915;
														assign node3915 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node3918 = (inp[9]) ? 4'b1000 : 4'b1100;
								assign node3921 = (inp[4]) ? node4015 : node3922;
									assign node3922 = (inp[12]) ? node3972 : node3923;
										assign node3923 = (inp[2]) ? node3949 : node3924;
											assign node3924 = (inp[1]) ? node3940 : node3925;
												assign node3925 = (inp[15]) ? node3931 : node3926;
													assign node3926 = (inp[14]) ? 4'b1000 : node3927;
														assign node3927 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node3931 = (inp[9]) ? 4'b1001 : node3932;
														assign node3932 = (inp[11]) ? node3936 : node3933;
															assign node3933 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node3936 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node3940 = (inp[11]) ? node3942 : 4'b1100;
													assign node3942 = (inp[9]) ? 4'b1101 : node3943;
														assign node3943 = (inp[14]) ? 4'b1000 : node3944;
															assign node3944 = (inp[15]) ? 4'b1100 : 4'b1101;
											assign node3949 = (inp[1]) ? node3959 : node3950;
												assign node3950 = (inp[14]) ? node3952 : 4'b1101;
													assign node3952 = (inp[15]) ? node3954 : 4'b1001;
														assign node3954 = (inp[11]) ? node3956 : 4'b1100;
															assign node3956 = (inp[5]) ? 4'b1100 : 4'b1101;
												assign node3959 = (inp[15]) ? node3965 : node3960;
													assign node3960 = (inp[14]) ? node3962 : 4'b1001;
														assign node3962 = (inp[5]) ? 4'b1101 : 4'b1001;
													assign node3965 = (inp[14]) ? node3969 : node3966;
														assign node3966 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node3969 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node3972 = (inp[1]) ? node3992 : node3973;
											assign node3973 = (inp[2]) ? node3989 : node3974;
												assign node3974 = (inp[15]) ? node3980 : node3975;
													assign node3975 = (inp[11]) ? node3977 : 4'b1010;
														assign node3977 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node3980 = (inp[9]) ? node3986 : node3981;
														assign node3981 = (inp[5]) ? 4'b1011 : node3982;
															assign node3982 = (inp[14]) ? 4'b1111 : 4'b1011;
														assign node3986 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node3989 = (inp[15]) ? 4'b1010 : 4'b1111;
											assign node3992 = (inp[2]) ? node4004 : node3993;
												assign node3993 = (inp[15]) ? 4'b1111 : node3994;
													assign node3994 = (inp[11]) ? node4000 : node3995;
														assign node3995 = (inp[14]) ? node3997 : 4'b1111;
															assign node3997 = (inp[5]) ? 4'b1110 : 4'b1111;
														assign node4000 = (inp[14]) ? 4'b1111 : 4'b1110;
												assign node4004 = (inp[15]) ? node4010 : node4005;
													assign node4005 = (inp[9]) ? node4007 : 4'b1010;
														assign node4007 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node4010 = (inp[14]) ? node4012 : 4'b1011;
														assign node4012 = (inp[11]) ? 4'b1111 : 4'b1110;
									assign node4015 = (inp[12]) ? node4077 : node4016;
										assign node4016 = (inp[15]) ? node4042 : node4017;
											assign node4017 = (inp[9]) ? node4027 : node4018;
												assign node4018 = (inp[14]) ? node4024 : node4019;
													assign node4019 = (inp[5]) ? node4021 : 4'b1110;
														assign node4021 = (inp[1]) ? 4'b1111 : 4'b1110;
													assign node4024 = (inp[1]) ? 4'b1010 : 4'b1111;
												assign node4027 = (inp[11]) ? node4037 : node4028;
													assign node4028 = (inp[5]) ? node4034 : node4029;
														assign node4029 = (inp[1]) ? node4031 : 4'b1010;
															assign node4031 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node4034 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node4037 = (inp[2]) ? 4'b1110 : node4038;
														assign node4038 = (inp[5]) ? 4'b1110 : 4'b1010;
											assign node4042 = (inp[14]) ? node4060 : node4043;
												assign node4043 = (inp[11]) ? node4053 : node4044;
													assign node4044 = (inp[9]) ? node4050 : node4045;
														assign node4045 = (inp[2]) ? 4'b1011 : node4046;
															assign node4046 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node4050 = (inp[1]) ? 4'b1110 : 4'b1011;
													assign node4053 = (inp[9]) ? node4055 : 4'b1110;
														assign node4055 = (inp[5]) ? 4'b1011 : node4056;
															assign node4056 = (inp[1]) ? 4'b1010 : 4'b1010;
												assign node4060 = (inp[1]) ? node4070 : node4061;
													assign node4061 = (inp[11]) ? node4065 : node4062;
														assign node4062 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node4065 = (inp[5]) ? 4'b1111 : node4066;
															assign node4066 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node4070 = (inp[2]) ? node4072 : 4'b1010;
														assign node4072 = (inp[5]) ? node4074 : 4'b1111;
															assign node4074 = (inp[11]) ? 4'b1010 : 4'b1011;
										assign node4077 = (inp[11]) ? node4111 : node4078;
											assign node4078 = (inp[9]) ? node4088 : node4079;
												assign node4079 = (inp[5]) ? 4'b1001 : node4080;
													assign node4080 = (inp[1]) ? node4082 : 4'b1100;
														assign node4082 = (inp[2]) ? node4084 : 4'b1000;
															assign node4084 = (inp[14]) ? 4'b1101 : 4'b1001;
												assign node4088 = (inp[15]) ? node4098 : node4089;
													assign node4089 = (inp[2]) ? node4091 : 4'b1001;
														assign node4091 = (inp[14]) ? node4095 : node4092;
															assign node4092 = (inp[5]) ? 4'b1000 : 4'b1000;
															assign node4095 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node4098 = (inp[2]) ? node4104 : node4099;
														assign node4099 = (inp[5]) ? node4101 : 4'b1000;
															assign node4101 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node4104 = (inp[14]) ? node4108 : node4105;
															assign node4105 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node4108 = (inp[5]) ? 4'b1100 : 4'b1000;
											assign node4111 = (inp[5]) ? node4127 : node4112;
												assign node4112 = (inp[2]) ? node4122 : node4113;
													assign node4113 = (inp[1]) ? node4119 : node4114;
														assign node4114 = (inp[15]) ? 4'b1000 : node4115;
															assign node4115 = (inp[14]) ? 4'b1000 : 4'b1101;
														assign node4119 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node4122 = (inp[1]) ? 4'b1001 : node4123;
														assign node4123 = (inp[15]) ? 4'b1101 : 4'b1100;
												assign node4127 = (inp[9]) ? node4141 : node4128;
													assign node4128 = (inp[1]) ? node4136 : node4129;
														assign node4129 = (inp[2]) ? node4133 : node4130;
															assign node4130 = (inp[14]) ? 4'b1000 : 4'b1000;
															assign node4133 = (inp[15]) ? 4'b1100 : 4'b1101;
														assign node4136 = (inp[2]) ? 4'b1000 : node4137;
															assign node4137 = (inp[14]) ? 4'b1000 : 4'b1100;
													assign node4141 = (inp[2]) ? 4'b1100 : node4142;
														assign node4142 = (inp[1]) ? node4144 : 4'b1101;
															assign node4144 = (inp[14]) ? 4'b1000 : 4'b1101;
							assign node4148 = (inp[5]) ? node4342 : node4149;
								assign node4149 = (inp[1]) ? node4247 : node4150;
									assign node4150 = (inp[2]) ? node4196 : node4151;
										assign node4151 = (inp[14]) ? node4169 : node4152;
											assign node4152 = (inp[15]) ? node4156 : node4153;
												assign node4153 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node4156 = (inp[4]) ? node4160 : node4157;
													assign node4157 = (inp[12]) ? 4'b1011 : 4'b1001;
													assign node4160 = (inp[12]) ? node4164 : node4161;
														assign node4161 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node4164 = (inp[13]) ? 4'b1001 : node4165;
															assign node4165 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node4169 = (inp[15]) ? node4183 : node4170;
												assign node4170 = (inp[4]) ? node4174 : node4171;
													assign node4171 = (inp[12]) ? 4'b1011 : 4'b1001;
													assign node4174 = (inp[12]) ? node4180 : node4175;
														assign node4175 = (inp[11]) ? node4177 : 4'b1011;
															assign node4177 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node4180 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node4183 = (inp[12]) ? node4189 : node4184;
													assign node4184 = (inp[4]) ? node4186 : 4'b1000;
														assign node4186 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node4189 = (inp[4]) ? node4191 : 4'b1111;
														assign node4191 = (inp[9]) ? 4'b1100 : node4192;
															assign node4192 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node4196 = (inp[15]) ? node4222 : node4197;
											assign node4197 = (inp[14]) ? node4205 : node4198;
												assign node4198 = (inp[13]) ? node4200 : 4'b1111;
													assign node4200 = (inp[9]) ? 4'b1110 : node4201;
														assign node4201 = (inp[12]) ? 4'b1110 : 4'b1101;
												assign node4205 = (inp[4]) ? node4213 : node4206;
													assign node4206 = (inp[12]) ? 4'b1111 : node4207;
														assign node4207 = (inp[13]) ? node4209 : 4'b1101;
															assign node4209 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node4213 = (inp[12]) ? node4217 : node4214;
														assign node4214 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node4217 = (inp[13]) ? 4'b1101 : node4218;
															assign node4218 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node4222 = (inp[14]) ? node4240 : node4223;
												assign node4223 = (inp[11]) ? node4231 : node4224;
													assign node4224 = (inp[4]) ? node4226 : 4'b1100;
														assign node4226 = (inp[12]) ? 4'b1100 : node4227;
															assign node4227 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node4231 = (inp[13]) ? node4237 : node4232;
														assign node4232 = (inp[12]) ? node4234 : 4'b1101;
															assign node4234 = (inp[4]) ? 4'b1101 : 4'b1111;
														assign node4237 = (inp[12]) ? 4'b1111 : 4'b1110;
												assign node4240 = (inp[4]) ? node4244 : node4241;
													assign node4241 = (inp[12]) ? 4'b1011 : 4'b1101;
													assign node4244 = (inp[12]) ? 4'b1001 : 4'b1011;
									assign node4247 = (inp[2]) ? node4287 : node4248;
										assign node4248 = (inp[12]) ? node4260 : node4249;
											assign node4249 = (inp[4]) ? node4251 : 4'b1101;
												assign node4251 = (inp[14]) ? node4253 : 4'b1111;
													assign node4253 = (inp[15]) ? node4255 : 4'b1111;
														assign node4255 = (inp[9]) ? node4257 : 4'b1011;
															assign node4257 = (inp[13]) ? 4'b1011 : 4'b1010;
											assign node4260 = (inp[4]) ? node4270 : node4261;
												assign node4261 = (inp[15]) ? node4263 : 4'b1110;
													assign node4263 = (inp[13]) ? node4267 : node4264;
														assign node4264 = (inp[14]) ? 4'b1011 : 4'b1111;
														assign node4267 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node4270 = (inp[15]) ? node4280 : node4271;
													assign node4271 = (inp[14]) ? node4277 : node4272;
														assign node4272 = (inp[13]) ? 4'b1001 : node4273;
															assign node4273 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node4277 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node4280 = (inp[14]) ? 4'b1001 : node4281;
														assign node4281 = (inp[13]) ? node4283 : 4'b1101;
															assign node4283 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node4287 = (inp[11]) ? node4317 : node4288;
											assign node4288 = (inp[15]) ? node4306 : node4289;
												assign node4289 = (inp[14]) ? node4299 : node4290;
													assign node4290 = (inp[4]) ? node4294 : node4291;
														assign node4291 = (inp[12]) ? 4'b1011 : 4'b1001;
														assign node4294 = (inp[12]) ? 4'b1100 : node4295;
															assign node4295 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node4299 = (inp[4]) ? node4301 : 4'b1000;
														assign node4301 = (inp[12]) ? node4303 : 4'b1011;
															assign node4303 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node4306 = (inp[14]) ? 4'b1000 : node4307;
													assign node4307 = (inp[12]) ? node4313 : node4308;
														assign node4308 = (inp[4]) ? node4310 : 4'b1001;
															assign node4310 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node4313 = (inp[4]) ? 4'b1000 : 4'b1010;
											assign node4317 = (inp[14]) ? node4327 : node4318;
												assign node4318 = (inp[9]) ? 4'b1011 : node4319;
													assign node4319 = (inp[4]) ? node4323 : node4320;
														assign node4320 = (inp[12]) ? 4'b1011 : 4'b1000;
														assign node4323 = (inp[12]) ? 4'b1001 : 4'b1011;
												assign node4327 = (inp[4]) ? node4337 : node4328;
													assign node4328 = (inp[12]) ? node4332 : node4329;
														assign node4329 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node4332 = (inp[15]) ? 4'b1111 : node4333;
															assign node4333 = (inp[13]) ? 4'b1011 : 4'b1010;
													assign node4337 = (inp[9]) ? 4'b1000 : node4338;
														assign node4338 = (inp[12]) ? 4'b1100 : 4'b1110;
								assign node4342 = (inp[11]) ? node4450 : node4343;
									assign node4343 = (inp[4]) ? node4387 : node4344;
										assign node4344 = (inp[12]) ? node4358 : node4345;
											assign node4345 = (inp[2]) ? 4'b1000 : node4346;
												assign node4346 = (inp[9]) ? node4348 : 4'b1000;
													assign node4348 = (inp[13]) ? node4354 : node4349;
														assign node4349 = (inp[15]) ? 4'b1001 : node4350;
															assign node4350 = (inp[14]) ? 4'b1001 : 4'b1101;
														assign node4354 = (inp[1]) ? 4'b1000 : 4'b1101;
											assign node4358 = (inp[2]) ? node4374 : node4359;
												assign node4359 = (inp[1]) ? node4367 : node4360;
													assign node4360 = (inp[9]) ? 4'b1011 : node4361;
														assign node4361 = (inp[15]) ? node4363 : 4'b1011;
															assign node4363 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node4367 = (inp[14]) ? node4369 : 4'b1110;
														assign node4369 = (inp[13]) ? node4371 : 4'b1111;
															assign node4371 = (inp[15]) ? 4'b1110 : 4'b1111;
												assign node4374 = (inp[1]) ? node4380 : node4375;
													assign node4375 = (inp[14]) ? 4'b1110 : node4376;
														assign node4376 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node4380 = (inp[9]) ? 4'b1010 : node4381;
														assign node4381 = (inp[14]) ? 4'b1011 : node4382;
															assign node4382 = (inp[15]) ? 4'b1011 : 4'b1010;
										assign node4387 = (inp[12]) ? node4423 : node4388;
											assign node4388 = (inp[13]) ? node4406 : node4389;
												assign node4389 = (inp[15]) ? node4397 : node4390;
													assign node4390 = (inp[14]) ? 4'b1111 : node4391;
														assign node4391 = (inp[2]) ? 4'b1011 : node4392;
															assign node4392 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node4397 = (inp[1]) ? node4399 : 4'b1111;
														assign node4399 = (inp[2]) ? node4403 : node4400;
															assign node4400 = (inp[14]) ? 4'b1110 : 4'b1010;
															assign node4403 = (inp[14]) ? 4'b1010 : 4'b1111;
												assign node4406 = (inp[9]) ? node4416 : node4407;
													assign node4407 = (inp[15]) ? node4413 : node4408;
														assign node4408 = (inp[14]) ? 4'b1110 : node4409;
															assign node4409 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node4413 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node4416 = (inp[14]) ? 4'b1010 : node4417;
														assign node4417 = (inp[2]) ? node4419 : 4'b1111;
															assign node4419 = (inp[15]) ? 4'b1010 : 4'b1011;
											assign node4423 = (inp[13]) ? node4439 : node4424;
												assign node4424 = (inp[14]) ? node4430 : node4425;
													assign node4425 = (inp[1]) ? node4427 : 4'b1000;
														assign node4427 = (inp[2]) ? 4'b1000 : 4'b1101;
													assign node4430 = (inp[15]) ? node4432 : 4'b1101;
														assign node4432 = (inp[2]) ? node4436 : node4433;
															assign node4433 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node4436 = (inp[1]) ? 4'b1000 : 4'b1100;
												assign node4439 = (inp[9]) ? 4'b1101 : node4440;
													assign node4440 = (inp[2]) ? node4442 : 4'b1101;
														assign node4442 = (inp[15]) ? node4446 : node4443;
															assign node4443 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node4446 = (inp[1]) ? 4'b1000 : 4'b1101;
									assign node4450 = (inp[15]) ? node4502 : node4451;
										assign node4451 = (inp[4]) ? node4475 : node4452;
											assign node4452 = (inp[12]) ? node4468 : node4453;
												assign node4453 = (inp[2]) ? node4459 : node4454;
													assign node4454 = (inp[14]) ? node4456 : 4'b1000;
														assign node4456 = (inp[1]) ? 4'b1001 : 4'b1101;
													assign node4459 = (inp[13]) ? node4463 : node4460;
														assign node4460 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node4463 = (inp[9]) ? node4465 : 4'b1000;
															assign node4465 = (inp[14]) ? 4'b1000 : 4'b1000;
												assign node4468 = (inp[1]) ? node4472 : node4469;
													assign node4469 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node4472 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node4475 = (inp[12]) ? node4487 : node4476;
												assign node4476 = (inp[9]) ? node4484 : node4477;
													assign node4477 = (inp[2]) ? node4479 : 4'b1010;
														assign node4479 = (inp[1]) ? node4481 : 4'b1011;
															assign node4481 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node4484 = (inp[1]) ? 4'b1011 : 4'b1111;
												assign node4487 = (inp[9]) ? node4497 : node4488;
													assign node4488 = (inp[13]) ? 4'b1001 : node4489;
														assign node4489 = (inp[1]) ? node4493 : node4490;
															assign node4490 = (inp[2]) ? 4'b1101 : 4'b1000;
															assign node4493 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node4497 = (inp[2]) ? 4'b1100 : node4498;
														assign node4498 = (inp[13]) ? 4'b1001 : 4'b1000;
										assign node4502 = (inp[1]) ? node4522 : node4503;
											assign node4503 = (inp[2]) ? node4519 : node4504;
												assign node4504 = (inp[12]) ? node4516 : node4505;
													assign node4505 = (inp[4]) ? node4511 : node4506;
														assign node4506 = (inp[14]) ? node4508 : 4'b1001;
															assign node4508 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node4511 = (inp[14]) ? 4'b1011 : node4512;
															assign node4512 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node4516 = (inp[4]) ? 4'b1000 : 4'b1011;
												assign node4519 = (inp[9]) ? 4'b1111 : 4'b1101;
											assign node4522 = (inp[2]) ? node4544 : node4523;
												assign node4523 = (inp[12]) ? node4537 : node4524;
													assign node4524 = (inp[4]) ? node4530 : node4525;
														assign node4525 = (inp[9]) ? 4'b1101 : node4526;
															assign node4526 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node4530 = (inp[14]) ? node4534 : node4531;
															assign node4531 = (inp[13]) ? 4'b1010 : 4'b1011;
															assign node4534 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node4537 = (inp[4]) ? node4539 : 4'b1110;
														assign node4539 = (inp[9]) ? node4541 : 4'b1100;
															assign node4541 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node4544 = (inp[12]) ? node4552 : node4545;
													assign node4545 = (inp[9]) ? node4547 : 4'b1000;
														assign node4547 = (inp[13]) ? 4'b1111 : node4548;
															assign node4548 = (inp[14]) ? 4'b1010 : 4'b1110;
													assign node4552 = (inp[4]) ? 4'b1001 : 4'b1011;
						assign node4555 = (inp[0]) ? node5003 : node4556;
							assign node4556 = (inp[13]) ? node4762 : node4557;
								assign node4557 = (inp[14]) ? node4643 : node4558;
									assign node4558 = (inp[1]) ? node4594 : node4559;
										assign node4559 = (inp[2]) ? node4573 : node4560;
											assign node4560 = (inp[4]) ? node4564 : node4561;
												assign node4561 = (inp[12]) ? 4'b1011 : 4'b1001;
												assign node4564 = (inp[12]) ? node4570 : node4565;
													assign node4565 = (inp[15]) ? node4567 : 4'b1011;
														assign node4567 = (inp[11]) ? 4'b1011 : 4'b1111;
													assign node4570 = (inp[11]) ? 4'b1101 : 4'b1000;
											assign node4573 = (inp[9]) ? node4583 : node4574;
												assign node4574 = (inp[11]) ? node4580 : node4575;
													assign node4575 = (inp[12]) ? node4577 : 4'b1101;
														assign node4577 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node4580 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node4583 = (inp[15]) ? node4589 : node4584;
													assign node4584 = (inp[4]) ? 4'b1110 : node4585;
														assign node4585 = (inp[12]) ? 4'b1111 : 4'b1101;
													assign node4589 = (inp[12]) ? 4'b1101 : node4590;
														assign node4590 = (inp[4]) ? 4'b1011 : 4'b1101;
										assign node4594 = (inp[2]) ? node4620 : node4595;
											assign node4595 = (inp[11]) ? node4605 : node4596;
												assign node4596 = (inp[12]) ? node4598 : 4'b1101;
													assign node4598 = (inp[4]) ? node4600 : 4'b1110;
														assign node4600 = (inp[15]) ? 4'b1101 : node4601;
															assign node4601 = (inp[9]) ? 4'b1101 : 4'b1000;
												assign node4605 = (inp[15]) ? node4615 : node4606;
													assign node4606 = (inp[9]) ? node4612 : node4607;
														assign node4607 = (inp[12]) ? 4'b1110 : node4608;
															assign node4608 = (inp[4]) ? 4'b1110 : 4'b1101;
														assign node4612 = (inp[5]) ? 4'b1101 : 4'b1001;
													assign node4615 = (inp[4]) ? node4617 : 4'b1111;
														assign node4617 = (inp[5]) ? 4'b1011 : 4'b1110;
											assign node4620 = (inp[5]) ? node4632 : node4621;
												assign node4621 = (inp[11]) ? 4'b1011 : node4622;
													assign node4622 = (inp[4]) ? node4626 : node4623;
														assign node4623 = (inp[12]) ? 4'b1011 : 4'b1001;
														assign node4626 = (inp[12]) ? 4'b1000 : node4627;
															assign node4627 = (inp[15]) ? 4'b1011 : 4'b1010;
												assign node4632 = (inp[12]) ? node4636 : node4633;
													assign node4633 = (inp[4]) ? 4'b1011 : 4'b1000;
													assign node4636 = (inp[4]) ? 4'b1001 : node4637;
														assign node4637 = (inp[11]) ? 4'b1011 : node4638;
															assign node4638 = (inp[15]) ? 4'b1011 : 4'b1010;
									assign node4643 = (inp[4]) ? node4705 : node4644;
										assign node4644 = (inp[12]) ? node4676 : node4645;
											assign node4645 = (inp[15]) ? node4665 : node4646;
												assign node4646 = (inp[1]) ? node4656 : node4647;
													assign node4647 = (inp[9]) ? 4'b1100 : node4648;
														assign node4648 = (inp[11]) ? node4652 : node4649;
															assign node4649 = (inp[5]) ? 4'b1000 : 4'b1001;
															assign node4652 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node4656 = (inp[9]) ? 4'b1001 : node4657;
														assign node4657 = (inp[5]) ? node4661 : node4658;
															assign node4658 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node4661 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node4665 = (inp[1]) ? node4673 : node4666;
													assign node4666 = (inp[2]) ? node4668 : 4'b1001;
														assign node4668 = (inp[5]) ? node4670 : 4'b1101;
															assign node4670 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node4673 = (inp[5]) ? 4'b1100 : 4'b1000;
											assign node4676 = (inp[11]) ? node4688 : node4677;
												assign node4677 = (inp[1]) ? node4681 : node4678;
													assign node4678 = (inp[2]) ? 4'b1110 : 4'b1011;
													assign node4681 = (inp[2]) ? node4685 : node4682;
														assign node4682 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node4685 = (inp[15]) ? 4'b1010 : 4'b1011;
												assign node4688 = (inp[1]) ? node4696 : node4689;
													assign node4689 = (inp[15]) ? node4691 : 4'b1111;
														assign node4691 = (inp[9]) ? node4693 : 4'b1011;
															assign node4693 = (inp[2]) ? 4'b1111 : 4'b1011;
													assign node4696 = (inp[2]) ? node4700 : node4697;
														assign node4697 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node4700 = (inp[5]) ? 4'b1011 : node4701;
															assign node4701 = (inp[15]) ? 4'b1111 : 4'b1010;
										assign node4705 = (inp[12]) ? node4739 : node4706;
											assign node4706 = (inp[2]) ? node4722 : node4707;
												assign node4707 = (inp[9]) ? node4719 : node4708;
													assign node4708 = (inp[11]) ? node4714 : node4709;
														assign node4709 = (inp[1]) ? node4711 : 4'b1111;
															assign node4711 = (inp[15]) ? 4'b1010 : 4'b1010;
														assign node4714 = (inp[5]) ? 4'b1111 : node4715;
															assign node4715 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node4719 = (inp[1]) ? 4'b1110 : 4'b1010;
												assign node4722 = (inp[9]) ? node4734 : node4723;
													assign node4723 = (inp[1]) ? node4729 : node4724;
														assign node4724 = (inp[5]) ? node4726 : 4'b1110;
															assign node4726 = (inp[11]) ? 4'b1111 : 4'b1011;
														assign node4729 = (inp[11]) ? 4'b1010 : node4730;
															assign node4730 = (inp[15]) ? 4'b1010 : 4'b1011;
													assign node4734 = (inp[5]) ? node4736 : 4'b1011;
														assign node4736 = (inp[1]) ? 4'b1010 : 4'b1011;
											assign node4739 = (inp[11]) ? node4749 : node4740;
												assign node4740 = (inp[9]) ? node4742 : 4'b1100;
													assign node4742 = (inp[15]) ? 4'b1101 : node4743;
														assign node4743 = (inp[2]) ? node4745 : 4'b1100;
															assign node4745 = (inp[1]) ? 4'b1101 : 4'b1000;
												assign node4749 = (inp[5]) ? node4755 : node4750;
													assign node4750 = (inp[9]) ? 4'b1100 : node4751;
														assign node4751 = (inp[2]) ? 4'b1100 : 4'b1001;
													assign node4755 = (inp[9]) ? node4759 : node4756;
														assign node4756 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node4759 = (inp[1]) ? 4'b1001 : 4'b1101;
								assign node4762 = (inp[9]) ? node4890 : node4763;
									assign node4763 = (inp[15]) ? node4823 : node4764;
										assign node4764 = (inp[4]) ? node4794 : node4765;
											assign node4765 = (inp[12]) ? node4783 : node4766;
												assign node4766 = (inp[14]) ? node4772 : node4767;
													assign node4767 = (inp[2]) ? node4769 : 4'b1000;
														assign node4769 = (inp[11]) ? 4'b1100 : 4'b1000;
													assign node4772 = (inp[5]) ? node4778 : node4773;
														assign node4773 = (inp[11]) ? node4775 : 4'b1001;
															assign node4775 = (inp[1]) ? 4'b1000 : 4'b1101;
														assign node4778 = (inp[1]) ? node4780 : 4'b1000;
															assign node4780 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node4783 = (inp[14]) ? 4'b1110 : node4784;
													assign node4784 = (inp[5]) ? node4790 : node4785;
														assign node4785 = (inp[2]) ? 4'b1011 : node4786;
															assign node4786 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node4790 = (inp[1]) ? 4'b1111 : 4'b1110;
											assign node4794 = (inp[12]) ? node4812 : node4795;
												assign node4795 = (inp[14]) ? node4803 : node4796;
													assign node4796 = (inp[2]) ? node4800 : node4797;
														assign node4797 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node4800 = (inp[5]) ? 4'b1111 : 4'b1110;
													assign node4803 = (inp[2]) ? 4'b1011 : node4804;
														assign node4804 = (inp[5]) ? node4808 : node4805;
															assign node4805 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node4808 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node4812 = (inp[14]) ? node4816 : node4813;
													assign node4813 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node4816 = (inp[5]) ? 4'b1000 : node4817;
														assign node4817 = (inp[1]) ? 4'b1001 : node4818;
															assign node4818 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node4823 = (inp[1]) ? node4861 : node4824;
											assign node4824 = (inp[2]) ? node4842 : node4825;
												assign node4825 = (inp[11]) ? node4837 : node4826;
													assign node4826 = (inp[14]) ? node4834 : node4827;
														assign node4827 = (inp[4]) ? node4831 : node4828;
															assign node4828 = (inp[12]) ? 4'b1010 : 4'b1000;
															assign node4831 = (inp[12]) ? 4'b1001 : 4'b1010;
														assign node4834 = (inp[4]) ? 4'b1011 : 4'b1001;
													assign node4837 = (inp[14]) ? 4'b1100 : node4838;
														assign node4838 = (inp[5]) ? 4'b1000 : 4'b1001;
												assign node4842 = (inp[4]) ? node4850 : node4843;
													assign node4843 = (inp[12]) ? node4845 : 4'b1101;
														assign node4845 = (inp[5]) ? 4'b1111 : node4846;
															assign node4846 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node4850 = (inp[12]) ? node4856 : node4851;
														assign node4851 = (inp[14]) ? node4853 : 4'b1010;
															assign node4853 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node4856 = (inp[14]) ? node4858 : 4'b1100;
															assign node4858 = (inp[5]) ? 4'b1101 : 4'b1001;
											assign node4861 = (inp[2]) ? node4877 : node4862;
												assign node4862 = (inp[12]) ? node4866 : node4863;
													assign node4863 = (inp[5]) ? 4'b1010 : 4'b1101;
													assign node4866 = (inp[4]) ? node4872 : node4867;
														assign node4867 = (inp[14]) ? node4869 : 4'b1110;
															assign node4869 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node4872 = (inp[11]) ? 4'b1000 : node4873;
															assign node4873 = (inp[5]) ? 4'b1101 : 4'b1100;
												assign node4877 = (inp[14]) ? node4883 : node4878;
													assign node4878 = (inp[11]) ? node4880 : 4'b1000;
														assign node4880 = (inp[4]) ? 4'b1011 : 4'b1000;
													assign node4883 = (inp[5]) ? node4887 : node4884;
														assign node4884 = (inp[12]) ? 4'b1100 : 4'b1110;
														assign node4887 = (inp[12]) ? 4'b1001 : 4'b1000;
									assign node4890 = (inp[1]) ? node4958 : node4891;
										assign node4891 = (inp[2]) ? node4923 : node4892;
											assign node4892 = (inp[14]) ? node4908 : node4893;
												assign node4893 = (inp[5]) ? 4'b1001 : node4894;
													assign node4894 = (inp[15]) ? node4900 : node4895;
														assign node4895 = (inp[11]) ? 4'b1010 : node4896;
															assign node4896 = (inp[4]) ? 4'b1001 : 4'b1011;
														assign node4900 = (inp[12]) ? node4904 : node4901;
															assign node4901 = (inp[11]) ? 4'b1001 : 4'b1010;
															assign node4904 = (inp[4]) ? 4'b1001 : 4'b1011;
												assign node4908 = (inp[11]) ? node4918 : node4909;
													assign node4909 = (inp[12]) ? node4913 : node4910;
														assign node4910 = (inp[5]) ? 4'b1101 : 4'b1110;
														assign node4913 = (inp[15]) ? 4'b1101 : node4914;
															assign node4914 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node4918 = (inp[4]) ? 4'b1011 : node4919;
														assign node4919 = (inp[15]) ? 4'b1000 : 4'b1001;
											assign node4923 = (inp[11]) ? node4931 : node4924;
												assign node4924 = (inp[5]) ? 4'b1101 : node4925;
													assign node4925 = (inp[15]) ? node4927 : 4'b1100;
														assign node4927 = (inp[4]) ? 4'b1111 : 4'b1101;
												assign node4931 = (inp[15]) ? node4947 : node4932;
													assign node4932 = (inp[5]) ? node4940 : node4933;
														assign node4933 = (inp[12]) ? node4937 : node4934;
															assign node4934 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node4937 = (inp[14]) ? 4'b1101 : 4'b1110;
														assign node4940 = (inp[12]) ? node4944 : node4941;
															assign node4941 = (inp[4]) ? 4'b1111 : 4'b1100;
															assign node4944 = (inp[4]) ? 4'b1000 : 4'b1110;
													assign node4947 = (inp[14]) ? node4953 : node4948;
														assign node4948 = (inp[5]) ? node4950 : 4'b1101;
															assign node4950 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node4953 = (inp[5]) ? 4'b1101 : node4954;
															assign node4954 = (inp[12]) ? 4'b1000 : 4'b1010;
										assign node4958 = (inp[2]) ? node4978 : node4959;
											assign node4959 = (inp[4]) ? node4969 : node4960;
												assign node4960 = (inp[12]) ? node4966 : node4961;
													assign node4961 = (inp[15]) ? 4'b1101 : node4962;
														assign node4962 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node4966 = (inp[5]) ? 4'b1111 : 4'b1110;
												assign node4969 = (inp[12]) ? node4975 : node4970;
													assign node4970 = (inp[15]) ? node4972 : 4'b1111;
														assign node4972 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node4975 = (inp[11]) ? 4'b1101 : 4'b1001;
											assign node4978 = (inp[12]) ? node4992 : node4979;
												assign node4979 = (inp[4]) ? node4985 : node4980;
													assign node4980 = (inp[14]) ? node4982 : 4'b1000;
														assign node4982 = (inp[5]) ? 4'b1100 : 4'b1000;
													assign node4985 = (inp[11]) ? node4989 : node4986;
														assign node4986 = (inp[15]) ? 4'b1010 : 4'b1011;
														assign node4989 = (inp[15]) ? 4'b1011 : 4'b1111;
												assign node4992 = (inp[4]) ? node5000 : node4993;
													assign node4993 = (inp[11]) ? 4'b1011 : node4994;
														assign node4994 = (inp[14]) ? node4996 : 4'b1010;
															assign node4996 = (inp[15]) ? 4'b1011 : 4'b1010;
													assign node5000 = (inp[14]) ? 4'b1001 : 4'b1000;
							assign node5003 = (inp[13]) ? node5223 : node5004;
								assign node5004 = (inp[14]) ? node5104 : node5005;
									assign node5005 = (inp[11]) ? node5055 : node5006;
										assign node5006 = (inp[1]) ? node5026 : node5007;
											assign node5007 = (inp[2]) ? node5017 : node5008;
												assign node5008 = (inp[4]) ? node5012 : node5009;
													assign node5009 = (inp[12]) ? 4'b1010 : 4'b1000;
													assign node5012 = (inp[12]) ? node5014 : 4'b1010;
														assign node5014 = (inp[5]) ? 4'b1001 : 4'b1100;
												assign node5017 = (inp[4]) ? node5021 : node5018;
													assign node5018 = (inp[12]) ? 4'b1110 : 4'b1100;
													assign node5021 = (inp[15]) ? node5023 : 4'b1111;
														assign node5023 = (inp[5]) ? 4'b1010 : 4'b1111;
											assign node5026 = (inp[2]) ? node5038 : node5027;
												assign node5027 = (inp[15]) ? node5033 : node5028;
													assign node5028 = (inp[12]) ? 4'b1111 : node5029;
														assign node5029 = (inp[4]) ? 4'b1110 : 4'b1100;
													assign node5033 = (inp[12]) ? 4'b1100 : node5034;
														assign node5034 = (inp[4]) ? 4'b1011 : 4'b1100;
												assign node5038 = (inp[4]) ? node5044 : node5039;
													assign node5039 = (inp[12]) ? 4'b1011 : node5040;
														assign node5040 = (inp[15]) ? 4'b1001 : 4'b1000;
													assign node5044 = (inp[12]) ? node5052 : node5045;
														assign node5045 = (inp[15]) ? node5049 : node5046;
															assign node5046 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node5049 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node5052 = (inp[15]) ? 4'b1000 : 4'b1001;
										assign node5055 = (inp[9]) ? node5081 : node5056;
											assign node5056 = (inp[2]) ? node5076 : node5057;
												assign node5057 = (inp[1]) ? node5069 : node5058;
													assign node5058 = (inp[4]) ? node5062 : node5059;
														assign node5059 = (inp[12]) ? 4'b1010 : 4'b1000;
														assign node5062 = (inp[12]) ? node5066 : node5063;
															assign node5063 = (inp[5]) ? 4'b1011 : 4'b1010;
															assign node5066 = (inp[15]) ? 4'b1001 : 4'b1100;
													assign node5069 = (inp[4]) ? 4'b1000 : node5070;
														assign node5070 = (inp[12]) ? 4'b1111 : node5071;
															assign node5071 = (inp[15]) ? 4'b1101 : 4'b1100;
												assign node5076 = (inp[1]) ? node5078 : 4'b1100;
													assign node5078 = (inp[4]) ? 4'b1010 : 4'b1001;
											assign node5081 = (inp[2]) ? node5093 : node5082;
												assign node5082 = (inp[1]) ? node5088 : node5083;
													assign node5083 = (inp[4]) ? 4'b1100 : node5084;
														assign node5084 = (inp[12]) ? 4'b1010 : 4'b1000;
													assign node5088 = (inp[15]) ? node5090 : 4'b1100;
														assign node5090 = (inp[4]) ? 4'b1100 : 4'b1110;
												assign node5093 = (inp[1]) ? node5099 : node5094;
													assign node5094 = (inp[4]) ? node5096 : 4'b1100;
														assign node5096 = (inp[5]) ? 4'b1010 : 4'b1111;
													assign node5099 = (inp[15]) ? 4'b1010 : node5100;
														assign node5100 = (inp[12]) ? 4'b1000 : 4'b1010;
									assign node5104 = (inp[1]) ? node5156 : node5105;
										assign node5105 = (inp[2]) ? node5133 : node5106;
											assign node5106 = (inp[11]) ? node5114 : node5107;
												assign node5107 = (inp[4]) ? 4'b1110 : node5108;
													assign node5108 = (inp[15]) ? 4'b1000 : node5109;
														assign node5109 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node5114 = (inp[12]) ? node5124 : node5115;
													assign node5115 = (inp[4]) ? node5119 : node5116;
														assign node5116 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node5119 = (inp[5]) ? 4'b1110 : node5120;
															assign node5120 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node5124 = (inp[4]) ? node5126 : 4'b1010;
														assign node5126 = (inp[9]) ? node5130 : node5127;
															assign node5127 = (inp[5]) ? 4'b1001 : 4'b1000;
															assign node5130 = (inp[5]) ? 4'b1000 : 4'b1100;
											assign node5133 = (inp[4]) ? node5145 : node5134;
												assign node5134 = (inp[12]) ? node5136 : 4'b1100;
													assign node5136 = (inp[11]) ? node5140 : node5137;
														assign node5137 = (inp[5]) ? 4'b1111 : 4'b1110;
														assign node5140 = (inp[5]) ? 4'b1110 : node5141;
															assign node5141 = (inp[15]) ? 4'b1010 : 4'b1110;
												assign node5145 = (inp[12]) ? node5151 : node5146;
													assign node5146 = (inp[5]) ? 4'b1010 : node5147;
														assign node5147 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node5151 = (inp[5]) ? 4'b1101 : node5152;
														assign node5152 = (inp[15]) ? 4'b1000 : 4'b1100;
										assign node5156 = (inp[2]) ? node5202 : node5157;
											assign node5157 = (inp[15]) ? node5181 : node5158;
												assign node5158 = (inp[5]) ? node5172 : node5159;
													assign node5159 = (inp[9]) ? node5165 : node5160;
														assign node5160 = (inp[11]) ? node5162 : 4'b1110;
															assign node5162 = (inp[4]) ? 4'b1101 : 4'b1110;
														assign node5165 = (inp[4]) ? node5169 : node5166;
															assign node5166 = (inp[12]) ? 4'b1110 : 4'b1101;
															assign node5169 = (inp[12]) ? 4'b1101 : 4'b1110;
													assign node5172 = (inp[9]) ? node5176 : node5173;
														assign node5173 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node5176 = (inp[4]) ? 4'b1000 : node5177;
															assign node5177 = (inp[12]) ? 4'b1111 : 4'b1000;
												assign node5181 = (inp[5]) ? node5193 : node5182;
													assign node5182 = (inp[9]) ? node5190 : node5183;
														assign node5183 = (inp[11]) ? node5187 : node5184;
															assign node5184 = (inp[12]) ? 4'b1010 : 4'b1011;
															assign node5187 = (inp[4]) ? 4'b1010 : 4'b1011;
														assign node5190 = (inp[12]) ? 4'b1000 : 4'b1010;
													assign node5193 = (inp[4]) ? 4'b1111 : node5194;
														assign node5194 = (inp[12]) ? node5198 : node5195;
															assign node5195 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node5198 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node5202 = (inp[5]) ? node5216 : node5203;
												assign node5203 = (inp[15]) ? node5209 : node5204;
													assign node5204 = (inp[12]) ? node5206 : 4'b1000;
														assign node5206 = (inp[9]) ? 4'b1001 : 4'b1011;
													assign node5209 = (inp[4]) ? node5211 : 4'b1110;
														assign node5211 = (inp[12]) ? node5213 : 4'b1110;
															assign node5213 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node5216 = (inp[11]) ? node5218 : 4'b1011;
													assign node5218 = (inp[12]) ? node5220 : 4'b1011;
														assign node5220 = (inp[9]) ? 4'b1010 : 4'b1000;
								assign node5223 = (inp[14]) ? node5355 : node5224;
									assign node5224 = (inp[9]) ? node5290 : node5225;
										assign node5225 = (inp[12]) ? node5255 : node5226;
											assign node5226 = (inp[4]) ? node5240 : node5227;
												assign node5227 = (inp[2]) ? node5233 : node5228;
													assign node5228 = (inp[1]) ? 4'b1100 : node5229;
														assign node5229 = (inp[15]) ? 4'b1001 : 4'b1000;
													assign node5233 = (inp[1]) ? 4'b1001 : node5234;
														assign node5234 = (inp[11]) ? 4'b1100 : node5235;
															assign node5235 = (inp[15]) ? 4'b1101 : 4'b1100;
												assign node5240 = (inp[5]) ? node5246 : node5241;
													assign node5241 = (inp[1]) ? node5243 : 4'b1111;
														assign node5243 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node5246 = (inp[11]) ? node5250 : node5247;
														assign node5247 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node5250 = (inp[1]) ? node5252 : 4'b1011;
															assign node5252 = (inp[2]) ? 4'b1011 : 4'b1111;
											assign node5255 = (inp[4]) ? node5277 : node5256;
												assign node5256 = (inp[11]) ? node5264 : node5257;
													assign node5257 = (inp[15]) ? node5259 : 4'b1010;
														assign node5259 = (inp[5]) ? node5261 : 4'b1111;
															assign node5261 = (inp[1]) ? 4'b1011 : 4'b1011;
													assign node5264 = (inp[1]) ? node5272 : node5265;
														assign node5265 = (inp[15]) ? node5269 : node5266;
															assign node5266 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node5269 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node5272 = (inp[2]) ? 4'b1010 : node5273;
															assign node5273 = (inp[15]) ? 4'b1111 : 4'b1110;
												assign node5277 = (inp[11]) ? node5279 : 4'b1100;
													assign node5279 = (inp[2]) ? node5283 : node5280;
														assign node5280 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node5283 = (inp[5]) ? node5287 : node5284;
															assign node5284 = (inp[1]) ? 4'b1101 : 4'b1000;
															assign node5287 = (inp[15]) ? 4'b1100 : 4'b1000;
										assign node5290 = (inp[1]) ? node5330 : node5291;
											assign node5291 = (inp[2]) ? node5309 : node5292;
												assign node5292 = (inp[11]) ? node5304 : node5293;
													assign node5293 = (inp[5]) ? node5297 : node5294;
														assign node5294 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node5297 = (inp[4]) ? node5301 : node5298;
															assign node5298 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node5301 = (inp[12]) ? 4'b1001 : 4'b1011;
													assign node5304 = (inp[12]) ? node5306 : 4'b1110;
														assign node5306 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node5309 = (inp[5]) ? node5323 : node5310;
													assign node5310 = (inp[11]) ? node5316 : node5311;
														assign node5311 = (inp[15]) ? node5313 : 4'b1111;
															assign node5313 = (inp[12]) ? 4'b1111 : 4'b1101;
														assign node5316 = (inp[4]) ? node5320 : node5317;
															assign node5317 = (inp[12]) ? 4'b1110 : 4'b1100;
															assign node5320 = (inp[12]) ? 4'b1101 : 4'b1111;
													assign node5323 = (inp[4]) ? 4'b1100 : node5324;
														assign node5324 = (inp[12]) ? 4'b1111 : node5325;
															assign node5325 = (inp[15]) ? 4'b1101 : 4'b1100;
											assign node5330 = (inp[2]) ? node5342 : node5331;
												assign node5331 = (inp[4]) ? node5335 : node5332;
													assign node5332 = (inp[12]) ? 4'b1111 : 4'b1100;
													assign node5335 = (inp[12]) ? node5339 : node5336;
														assign node5336 = (inp[15]) ? 4'b1011 : 4'b1111;
														assign node5339 = (inp[5]) ? 4'b1100 : 4'b1101;
												assign node5342 = (inp[4]) ? node5348 : node5343;
													assign node5343 = (inp[12]) ? 4'b1011 : node5344;
														assign node5344 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node5348 = (inp[12]) ? node5352 : node5349;
														assign node5349 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node5352 = (inp[15]) ? 4'b1001 : 4'b1101;
									assign node5355 = (inp[4]) ? node5405 : node5356;
										assign node5356 = (inp[12]) ? node5376 : node5357;
											assign node5357 = (inp[9]) ? node5367 : node5358;
												assign node5358 = (inp[2]) ? 4'b1001 : node5359;
													assign node5359 = (inp[11]) ? node5361 : 4'b1000;
														assign node5361 = (inp[1]) ? 4'b1100 : node5362;
															assign node5362 = (inp[15]) ? 4'b1001 : 4'b1100;
												assign node5367 = (inp[11]) ? node5369 : 4'b1100;
													assign node5369 = (inp[1]) ? 4'b1000 : node5370;
														assign node5370 = (inp[15]) ? node5372 : 4'b1100;
															assign node5372 = (inp[2]) ? 4'b1101 : 4'b1001;
											assign node5376 = (inp[9]) ? node5384 : node5377;
												assign node5377 = (inp[2]) ? 4'b1111 : node5378;
													assign node5378 = (inp[15]) ? node5380 : 4'b1010;
														assign node5380 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node5384 = (inp[11]) ? node5394 : node5385;
													assign node5385 = (inp[15]) ? node5391 : node5386;
														assign node5386 = (inp[1]) ? node5388 : 4'b1111;
															assign node5388 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node5391 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node5394 = (inp[1]) ? node5400 : node5395;
														assign node5395 = (inp[5]) ? node5397 : 4'b1010;
															assign node5397 = (inp[2]) ? 4'b1111 : 4'b1010;
														assign node5400 = (inp[5]) ? 4'b1111 : node5401;
															assign node5401 = (inp[2]) ? 4'b1111 : 4'b1011;
										assign node5405 = (inp[12]) ? node5435 : node5406;
											assign node5406 = (inp[11]) ? node5420 : node5407;
												assign node5407 = (inp[5]) ? 4'b1111 : node5408;
													assign node5408 = (inp[1]) ? node5414 : node5409;
														assign node5409 = (inp[15]) ? node5411 : 4'b1010;
															assign node5411 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node5414 = (inp[9]) ? 4'b1010 : node5415;
															assign node5415 = (inp[2]) ? 4'b1010 : 4'b1110;
												assign node5420 = (inp[2]) ? node5430 : node5421;
													assign node5421 = (inp[9]) ? 4'b1010 : node5422;
														assign node5422 = (inp[5]) ? node5426 : node5423;
															assign node5423 = (inp[15]) ? 4'b1111 : 4'b1010;
															assign node5426 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node5430 = (inp[15]) ? node5432 : 4'b1010;
														assign node5432 = (inp[5]) ? 4'b1010 : 4'b1011;
											assign node5435 = (inp[9]) ? node5447 : node5436;
												assign node5436 = (inp[5]) ? node5442 : node5437;
													assign node5437 = (inp[1]) ? node5439 : 4'b1000;
														assign node5439 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node5442 = (inp[2]) ? 4'b1000 : node5443;
														assign node5443 = (inp[15]) ? 4'b1100 : 4'b1101;
												assign node5447 = (inp[2]) ? node5451 : node5448;
													assign node5448 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node5451 = (inp[1]) ? node5453 : 4'b1100;
														assign node5453 = (inp[5]) ? node5455 : 4'b1101;
															assign node5455 = (inp[15]) ? 4'b1000 : 4'b1100;
					assign node5458 = (inp[13]) ? node6374 : node5459;
						assign node5459 = (inp[1]) ? node5895 : node5460;
							assign node5460 = (inp[2]) ? node5658 : node5461;
								assign node5461 = (inp[14]) ? node5575 : node5462;
									assign node5462 = (inp[12]) ? node5524 : node5463;
										assign node5463 = (inp[4]) ? node5493 : node5464;
											assign node5464 = (inp[11]) ? node5478 : node5465;
												assign node5465 = (inp[10]) ? node5471 : node5466;
													assign node5466 = (inp[15]) ? node5468 : 4'b1001;
														assign node5468 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node5471 = (inp[5]) ? node5475 : node5472;
														assign node5472 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node5475 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node5478 = (inp[5]) ? node5486 : node5479;
													assign node5479 = (inp[15]) ? 4'b1101 : node5480;
														assign node5480 = (inp[10]) ? node5482 : 4'b1000;
															assign node5482 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node5486 = (inp[15]) ? 4'b1000 : node5487;
														assign node5487 = (inp[9]) ? 4'b1101 : node5488;
															assign node5488 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node5493 = (inp[15]) ? node5511 : node5494;
												assign node5494 = (inp[5]) ? node5500 : node5495;
													assign node5495 = (inp[10]) ? node5497 : 4'b1011;
														assign node5497 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node5500 = (inp[0]) ? node5504 : node5501;
														assign node5501 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node5504 = (inp[9]) ? node5508 : node5505;
															assign node5505 = (inp[11]) ? 4'b1110 : 4'b1110;
															assign node5508 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node5511 = (inp[10]) ? node5519 : node5512;
													assign node5512 = (inp[0]) ? node5514 : 4'b1010;
														assign node5514 = (inp[11]) ? node5516 : 4'b1011;
															assign node5516 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node5519 = (inp[0]) ? 4'b1010 : node5520;
														assign node5520 = (inp[5]) ? 4'b1011 : 4'b1010;
										assign node5524 = (inp[4]) ? node5548 : node5525;
											assign node5525 = (inp[9]) ? node5539 : node5526;
												assign node5526 = (inp[10]) ? node5534 : node5527;
													assign node5527 = (inp[11]) ? node5529 : 4'b1110;
														assign node5529 = (inp[0]) ? 4'b1010 : node5530;
															assign node5530 = (inp[5]) ? 4'b1010 : 4'b1011;
													assign node5534 = (inp[15]) ? node5536 : 4'b1011;
														assign node5536 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node5539 = (inp[15]) ? node5545 : node5540;
													assign node5540 = (inp[10]) ? 4'b1111 : node5541;
														assign node5541 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node5545 = (inp[5]) ? 4'b1010 : 4'b1111;
											assign node5548 = (inp[15]) ? node5562 : node5549;
												assign node5549 = (inp[10]) ? node5551 : 4'b1000;
													assign node5551 = (inp[0]) ? node5557 : node5552;
														assign node5552 = (inp[11]) ? 4'b1000 : node5553;
															assign node5553 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node5557 = (inp[5]) ? node5559 : 4'b1001;
															assign node5559 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node5562 = (inp[5]) ? node5570 : node5563;
													assign node5563 = (inp[9]) ? 4'b1101 : node5564;
														assign node5564 = (inp[11]) ? node5566 : 4'b1100;
															assign node5566 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node5570 = (inp[10]) ? 4'b1001 : node5571;
														assign node5571 = (inp[0]) ? 4'b1000 : 4'b1001;
									assign node5575 = (inp[4]) ? node5623 : node5576;
										assign node5576 = (inp[12]) ? node5604 : node5577;
											assign node5577 = (inp[9]) ? node5591 : node5578;
												assign node5578 = (inp[0]) ? node5586 : node5579;
													assign node5579 = (inp[5]) ? 4'b1000 : node5580;
														assign node5580 = (inp[15]) ? 4'b1001 : node5581;
															assign node5581 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node5586 = (inp[5]) ? node5588 : 4'b1000;
														assign node5588 = (inp[15]) ? 4'b1100 : 4'b1000;
												assign node5591 = (inp[11]) ? node5595 : node5592;
													assign node5592 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node5595 = (inp[15]) ? node5601 : node5596;
														assign node5596 = (inp[5]) ? node5598 : 4'b1001;
															assign node5598 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node5601 = (inp[5]) ? 4'b1101 : 4'b1001;
											assign node5604 = (inp[15]) ? node5614 : node5605;
												assign node5605 = (inp[5]) ? node5611 : node5606;
													assign node5606 = (inp[0]) ? 4'b1111 : node5607;
														assign node5607 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node5611 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node5614 = (inp[0]) ? 4'b1011 : node5615;
													assign node5615 = (inp[11]) ? 4'b1010 : node5616;
														assign node5616 = (inp[5]) ? 4'b1010 : node5617;
															assign node5617 = (inp[10]) ? 4'b1010 : 4'b1011;
										assign node5623 = (inp[12]) ? node5643 : node5624;
											assign node5624 = (inp[11]) ? node5630 : node5625;
												assign node5625 = (inp[5]) ? 4'b1011 : node5626;
													assign node5626 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node5630 = (inp[15]) ? node5636 : node5631;
													assign node5631 = (inp[5]) ? node5633 : 4'b1010;
														assign node5633 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node5636 = (inp[5]) ? node5638 : 4'b1011;
														assign node5638 = (inp[10]) ? 4'b1010 : node5639;
															assign node5639 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node5643 = (inp[15]) ? node5651 : node5644;
												assign node5644 = (inp[0]) ? 4'b1001 : node5645;
													assign node5645 = (inp[5]) ? node5647 : 4'b1000;
														assign node5647 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node5651 = (inp[10]) ? node5655 : node5652;
													assign node5652 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node5655 = (inp[0]) ? 4'b1001 : 4'b1000;
								assign node5658 = (inp[4]) ? node5772 : node5659;
									assign node5659 = (inp[12]) ? node5717 : node5660;
										assign node5660 = (inp[15]) ? node5690 : node5661;
											assign node5661 = (inp[14]) ? node5677 : node5662;
												assign node5662 = (inp[5]) ? node5670 : node5663;
													assign node5663 = (inp[9]) ? node5665 : 4'b1100;
														assign node5665 = (inp[10]) ? node5667 : 4'b1101;
															assign node5667 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node5670 = (inp[10]) ? 4'b1000 : node5671;
														assign node5671 = (inp[11]) ? 4'b1001 : node5672;
															assign node5672 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node5677 = (inp[10]) ? 4'b1100 : node5678;
													assign node5678 = (inp[9]) ? node5684 : node5679;
														assign node5679 = (inp[0]) ? node5681 : 4'b1101;
															assign node5681 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node5684 = (inp[5]) ? 4'b1100 : node5685;
															assign node5685 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node5690 = (inp[11]) ? node5708 : node5691;
												assign node5691 = (inp[9]) ? node5701 : node5692;
													assign node5692 = (inp[10]) ? 4'b1001 : node5693;
														assign node5693 = (inp[5]) ? node5697 : node5694;
															assign node5694 = (inp[14]) ? 4'b1101 : 4'b1000;
															assign node5697 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node5701 = (inp[0]) ? node5703 : 4'b1000;
														assign node5703 = (inp[5]) ? 4'b1101 : node5704;
															assign node5704 = (inp[14]) ? 4'b1100 : 4'b1000;
												assign node5708 = (inp[14]) ? node5714 : node5709;
													assign node5709 = (inp[9]) ? 4'b1001 : node5710;
														assign node5710 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node5714 = (inp[5]) ? 4'b1001 : 4'b1100;
										assign node5717 = (inp[5]) ? node5739 : node5718;
											assign node5718 = (inp[14]) ? node5732 : node5719;
												assign node5719 = (inp[15]) ? node5727 : node5720;
													assign node5720 = (inp[9]) ? 4'b1110 : node5721;
														assign node5721 = (inp[0]) ? 4'b1111 : node5722;
															assign node5722 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node5727 = (inp[0]) ? node5729 : 4'b1011;
														assign node5729 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node5732 = (inp[15]) ? 4'b1110 : node5733;
													assign node5733 = (inp[0]) ? node5735 : 4'b1010;
														assign node5735 = (inp[10]) ? 4'b1011 : 4'b1010;
											assign node5739 = (inp[15]) ? node5753 : node5740;
												assign node5740 = (inp[14]) ? node5744 : node5741;
													assign node5741 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node5744 = (inp[9]) ? node5746 : 4'b1111;
														assign node5746 = (inp[0]) ? node5750 : node5747;
															assign node5747 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node5750 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node5753 = (inp[0]) ? node5759 : node5754;
													assign node5754 = (inp[10]) ? node5756 : 4'b1110;
														assign node5756 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node5759 = (inp[9]) ? node5767 : node5760;
														assign node5760 = (inp[10]) ? node5764 : node5761;
															assign node5761 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node5764 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node5767 = (inp[10]) ? 4'b1110 : node5768;
															assign node5768 = (inp[14]) ? 4'b1110 : 4'b1111;
									assign node5772 = (inp[12]) ? node5840 : node5773;
										assign node5773 = (inp[9]) ? node5809 : node5774;
											assign node5774 = (inp[14]) ? node5788 : node5775;
												assign node5775 = (inp[5]) ? node5781 : node5776;
													assign node5776 = (inp[15]) ? node5778 : 4'b1110;
														assign node5778 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node5781 = (inp[15]) ? 4'b1110 : node5782;
														assign node5782 = (inp[10]) ? 4'b1011 : node5783;
															assign node5783 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node5788 = (inp[15]) ? node5798 : node5789;
													assign node5789 = (inp[5]) ? 4'b1110 : node5790;
														assign node5790 = (inp[0]) ? node5794 : node5791;
															assign node5791 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node5794 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node5798 = (inp[10]) ? node5804 : node5799;
														assign node5799 = (inp[0]) ? node5801 : 4'b1111;
															assign node5801 = (inp[5]) ? 4'b1110 : 4'b1111;
														assign node5804 = (inp[11]) ? node5806 : 4'b1110;
															assign node5806 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node5809 = (inp[5]) ? node5825 : node5810;
												assign node5810 = (inp[14]) ? node5818 : node5811;
													assign node5811 = (inp[11]) ? 4'b1111 : node5812;
														assign node5812 = (inp[15]) ? node5814 : 4'b1110;
															assign node5814 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node5818 = (inp[15]) ? node5820 : 4'b1110;
														assign node5820 = (inp[10]) ? node5822 : 4'b1110;
															assign node5822 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node5825 = (inp[11]) ? node5831 : node5826;
													assign node5826 = (inp[14]) ? 4'b1111 : node5827;
														assign node5827 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node5831 = (inp[15]) ? node5837 : node5832;
														assign node5832 = (inp[10]) ? 4'b1111 : node5833;
															assign node5833 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node5837 = (inp[0]) ? 4'b1111 : 4'b1110;
										assign node5840 = (inp[15]) ? node5866 : node5841;
											assign node5841 = (inp[9]) ? node5857 : node5842;
												assign node5842 = (inp[5]) ? node5848 : node5843;
													assign node5843 = (inp[10]) ? node5845 : 4'b1100;
														assign node5845 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node5848 = (inp[11]) ? node5854 : node5849;
														assign node5849 = (inp[0]) ? node5851 : 4'b1101;
															assign node5851 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node5854 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node5857 = (inp[0]) ? node5863 : node5858;
													assign node5858 = (inp[10]) ? 4'b1101 : node5859;
														assign node5859 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node5863 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node5866 = (inp[9]) ? node5878 : node5867;
												assign node5867 = (inp[5]) ? 4'b1101 : node5868;
													assign node5868 = (inp[14]) ? node5874 : node5869;
														assign node5869 = (inp[0]) ? node5871 : 4'b1000;
															assign node5871 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node5874 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node5878 = (inp[10]) ? node5884 : node5879;
													assign node5879 = (inp[14]) ? 4'b1100 : node5880;
														assign node5880 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node5884 = (inp[0]) ? node5890 : node5885;
														assign node5885 = (inp[11]) ? 4'b1101 : node5886;
															assign node5886 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node5890 = (inp[11]) ? 4'b1100 : node5891;
															assign node5891 = (inp[5]) ? 4'b1100 : 4'b1101;
							assign node5895 = (inp[2]) ? node6125 : node5896;
								assign node5896 = (inp[4]) ? node6014 : node5897;
									assign node5897 = (inp[12]) ? node5949 : node5898;
										assign node5898 = (inp[15]) ? node5924 : node5899;
											assign node5899 = (inp[14]) ? node5913 : node5900;
												assign node5900 = (inp[5]) ? node5906 : node5901;
													assign node5901 = (inp[0]) ? 4'b1101 : node5902;
														assign node5902 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node5906 = (inp[10]) ? 4'b1000 : node5907;
														assign node5907 = (inp[9]) ? 4'b1001 : node5908;
															assign node5908 = (inp[11]) ? 4'b1000 : 4'b1000;
												assign node5913 = (inp[9]) ? node5919 : node5914;
													assign node5914 = (inp[5]) ? 4'b1101 : node5915;
														assign node5915 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node5919 = (inp[0]) ? node5921 : 4'b1100;
														assign node5921 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node5924 = (inp[9]) ? node5938 : node5925;
												assign node5925 = (inp[0]) ? node5935 : node5926;
													assign node5926 = (inp[10]) ? node5930 : node5927;
														assign node5927 = (inp[14]) ? 4'b1000 : 4'b1100;
														assign node5930 = (inp[5]) ? 4'b1101 : node5931;
															assign node5931 = (inp[14]) ? 4'b1101 : 4'b1000;
													assign node5935 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node5938 = (inp[5]) ? node5942 : node5939;
													assign node5939 = (inp[14]) ? 4'b1100 : 4'b1000;
													assign node5942 = (inp[14]) ? node5944 : 4'b1100;
														assign node5944 = (inp[11]) ? node5946 : 4'b1000;
															assign node5946 = (inp[10]) ? 4'b1000 : 4'b1000;
										assign node5949 = (inp[15]) ? node5987 : node5950;
											assign node5950 = (inp[0]) ? node5972 : node5951;
												assign node5951 = (inp[10]) ? node5963 : node5952;
													assign node5952 = (inp[5]) ? node5960 : node5953;
														assign node5953 = (inp[14]) ? node5957 : node5954;
															assign node5954 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node5957 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node5960 = (inp[11]) ? 4'b1011 : 4'b1111;
													assign node5963 = (inp[5]) ? node5969 : node5964;
														assign node5964 = (inp[14]) ? 4'b1011 : node5965;
															assign node5965 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node5969 = (inp[14]) ? 4'b1110 : 4'b1010;
												assign node5972 = (inp[10]) ? node5982 : node5973;
													assign node5973 = (inp[5]) ? node5979 : node5974;
														assign node5974 = (inp[14]) ? node5976 : 4'b1111;
															assign node5976 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node5979 = (inp[14]) ? 4'b1110 : 4'b1010;
													assign node5982 = (inp[5]) ? node5984 : 4'b1010;
														assign node5984 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node5987 = (inp[5]) ? node5997 : node5988;
												assign node5988 = (inp[14]) ? 4'b1110 : node5989;
													assign node5989 = (inp[10]) ? 4'b1010 : node5990;
														assign node5990 = (inp[11]) ? 4'b1011 : node5991;
															assign node5991 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node5997 = (inp[0]) ? node6003 : node5998;
													assign node5998 = (inp[14]) ? 4'b1111 : node5999;
														assign node5999 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node6003 = (inp[10]) ? node6009 : node6004;
														assign node6004 = (inp[14]) ? 4'b1110 : node6005;
															assign node6005 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node6009 = (inp[11]) ? node6011 : 4'b1111;
															assign node6011 = (inp[14]) ? 4'b1111 : 4'b1110;
									assign node6014 = (inp[12]) ? node6068 : node6015;
										assign node6015 = (inp[5]) ? node6049 : node6016;
											assign node6016 = (inp[10]) ? node6032 : node6017;
												assign node6017 = (inp[11]) ? node6025 : node6018;
													assign node6018 = (inp[0]) ? node6022 : node6019;
														assign node6019 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node6022 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node6025 = (inp[15]) ? 4'b1110 : node6026;
														assign node6026 = (inp[14]) ? node6028 : 4'b1110;
															assign node6028 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node6032 = (inp[14]) ? node6038 : node6033;
													assign node6033 = (inp[11]) ? node6035 : 4'b1111;
														assign node6035 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node6038 = (inp[15]) ? node6046 : node6039;
														assign node6039 = (inp[11]) ? node6043 : node6040;
															assign node6040 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node6043 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node6046 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node6049 = (inp[15]) ? node6057 : node6050;
												assign node6050 = (inp[14]) ? 4'b1110 : node6051;
													assign node6051 = (inp[10]) ? 4'b1010 : node6052;
														assign node6052 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node6057 = (inp[9]) ? node6061 : node6058;
													assign node6058 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node6061 = (inp[14]) ? 4'b1110 : node6062;
														assign node6062 = (inp[10]) ? node6064 : 4'b1110;
															assign node6064 = (inp[0]) ? 4'b1110 : 4'b1110;
										assign node6068 = (inp[5]) ? node6096 : node6069;
											assign node6069 = (inp[14]) ? node6089 : node6070;
												assign node6070 = (inp[15]) ? node6076 : node6071;
													assign node6071 = (inp[0]) ? 4'b1100 : node6072;
														assign node6072 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node6076 = (inp[11]) ? node6082 : node6077;
														assign node6077 = (inp[10]) ? 4'b1001 : node6078;
															assign node6078 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node6082 = (inp[10]) ? node6086 : node6083;
															assign node6083 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node6086 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node6089 = (inp[15]) ? 4'b1100 : node6090;
													assign node6090 = (inp[9]) ? 4'b1100 : node6091;
														assign node6091 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node6096 = (inp[10]) ? node6110 : node6097;
												assign node6097 = (inp[14]) ? node6103 : node6098;
													assign node6098 = (inp[11]) ? 4'b1101 : node6099;
														assign node6099 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node6103 = (inp[0]) ? node6105 : 4'b1100;
														assign node6105 = (inp[15]) ? 4'b1100 : node6106;
															assign node6106 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node6110 = (inp[14]) ? 4'b1101 : node6111;
													assign node6111 = (inp[0]) ? node6119 : node6112;
														assign node6112 = (inp[9]) ? node6116 : node6113;
															assign node6113 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node6116 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node6119 = (inp[15]) ? node6121 : 4'b1100;
															assign node6121 = (inp[11]) ? 4'b1101 : 4'b1100;
								assign node6125 = (inp[4]) ? node6261 : node6126;
									assign node6126 = (inp[12]) ? node6196 : node6127;
										assign node6127 = (inp[15]) ? node6163 : node6128;
											assign node6128 = (inp[14]) ? node6140 : node6129;
												assign node6129 = (inp[5]) ? node6133 : node6130;
													assign node6130 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node6133 = (inp[10]) ? node6135 : 4'b1100;
														assign node6135 = (inp[0]) ? 4'b1100 : node6136;
															assign node6136 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node6140 = (inp[9]) ? node6152 : node6141;
													assign node6141 = (inp[11]) ? node6147 : node6142;
														assign node6142 = (inp[0]) ? node6144 : 4'b1000;
															assign node6144 = (inp[5]) ? 4'b1000 : 4'b1001;
														assign node6147 = (inp[0]) ? 4'b1000 : node6148;
															assign node6148 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node6152 = (inp[11]) ? node6160 : node6153;
														assign node6153 = (inp[10]) ? node6157 : node6154;
															assign node6154 = (inp[5]) ? 4'b1000 : 4'b1001;
															assign node6157 = (inp[0]) ? 4'b1000 : 4'b1000;
														assign node6160 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node6163 = (inp[0]) ? node6179 : node6164;
												assign node6164 = (inp[9]) ? node6168 : node6165;
													assign node6165 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node6168 = (inp[11]) ? node6174 : node6169;
														assign node6169 = (inp[14]) ? node6171 : 4'b1000;
															assign node6171 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node6174 = (inp[5]) ? 4'b1101 : node6175;
															assign node6175 = (inp[14]) ? 4'b1001 : 4'b1101;
												assign node6179 = (inp[10]) ? node6185 : node6180;
													assign node6180 = (inp[9]) ? 4'b1100 : node6181;
														assign node6181 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node6185 = (inp[14]) ? node6191 : node6186;
														assign node6186 = (inp[5]) ? node6188 : 4'b1101;
															assign node6188 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node6191 = (inp[5]) ? node6193 : 4'b1000;
															assign node6193 = (inp[9]) ? 4'b1100 : 4'b1101;
										assign node6196 = (inp[5]) ? node6232 : node6197;
											assign node6197 = (inp[9]) ? node6217 : node6198;
												assign node6198 = (inp[0]) ? node6208 : node6199;
													assign node6199 = (inp[15]) ? node6203 : node6200;
														assign node6200 = (inp[11]) ? 4'b1010 : 4'b1110;
														assign node6203 = (inp[14]) ? 4'b1010 : node6204;
															assign node6204 = (inp[11]) ? 4'b1110 : 4'b1110;
													assign node6208 = (inp[10]) ? node6212 : node6209;
														assign node6209 = (inp[15]) ? 4'b1111 : 4'b1011;
														assign node6212 = (inp[15]) ? node6214 : 4'b1110;
															assign node6214 = (inp[14]) ? 4'b1011 : 4'b1110;
												assign node6217 = (inp[10]) ? node6227 : node6218;
													assign node6218 = (inp[11]) ? node6220 : 4'b1111;
														assign node6220 = (inp[14]) ? node6224 : node6221;
															assign node6221 = (inp[15]) ? 4'b1110 : 4'b1011;
															assign node6224 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node6227 = (inp[14]) ? node6229 : 4'b1011;
														assign node6229 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node6232 = (inp[15]) ? node6244 : node6233;
												assign node6233 = (inp[14]) ? node6237 : node6234;
													assign node6234 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node6237 = (inp[10]) ? 4'b1011 : node6238;
														assign node6238 = (inp[9]) ? 4'b1010 : node6239;
															assign node6239 = (inp[11]) ? 4'b1010 : 4'b1010;
												assign node6244 = (inp[14]) ? node6254 : node6245;
													assign node6245 = (inp[11]) ? node6249 : node6246;
														assign node6246 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node6249 = (inp[9]) ? node6251 : 4'b1011;
															assign node6251 = (inp[0]) ? 4'b1010 : 4'b1010;
													assign node6254 = (inp[10]) ? node6256 : 4'b1010;
														assign node6256 = (inp[0]) ? 4'b1010 : node6257;
															assign node6257 = (inp[11]) ? 4'b1011 : 4'b1010;
									assign node6261 = (inp[12]) ? node6317 : node6262;
										assign node6262 = (inp[5]) ? node6296 : node6263;
											assign node6263 = (inp[9]) ? node6279 : node6264;
												assign node6264 = (inp[10]) ? node6272 : node6265;
													assign node6265 = (inp[0]) ? node6267 : 4'b1010;
														assign node6267 = (inp[15]) ? 4'b1011 : node6268;
															assign node6268 = (inp[14]) ? 4'b1011 : 4'b1010;
													assign node6272 = (inp[14]) ? 4'b1011 : node6273;
														assign node6273 = (inp[11]) ? 4'b1011 : node6274;
															assign node6274 = (inp[15]) ? 4'b1010 : 4'b1010;
												assign node6279 = (inp[0]) ? node6283 : node6280;
													assign node6280 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node6283 = (inp[15]) ? node6289 : node6284;
														assign node6284 = (inp[10]) ? 4'b1010 : node6285;
															assign node6285 = (inp[14]) ? 4'b1010 : 4'b1010;
														assign node6289 = (inp[11]) ? node6293 : node6290;
															assign node6290 = (inp[14]) ? 4'b1010 : 4'b1010;
															assign node6293 = (inp[10]) ? 4'b1011 : 4'b1010;
											assign node6296 = (inp[14]) ? node6304 : node6297;
												assign node6297 = (inp[15]) ? node6299 : 4'b1110;
													assign node6299 = (inp[9]) ? node6301 : 4'b1011;
														assign node6301 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node6304 = (inp[10]) ? node6312 : node6305;
													assign node6305 = (inp[11]) ? node6307 : 4'b1011;
														assign node6307 = (inp[9]) ? 4'b1011 : node6308;
															assign node6308 = (inp[0]) ? 4'b1010 : 4'b1010;
													assign node6312 = (inp[11]) ? 4'b1010 : node6313;
														assign node6313 = (inp[15]) ? 4'b1010 : 4'b1011;
										assign node6317 = (inp[15]) ? node6349 : node6318;
											assign node6318 = (inp[10]) ? node6332 : node6319;
												assign node6319 = (inp[11]) ? node6325 : node6320;
													assign node6320 = (inp[9]) ? node6322 : 4'b1000;
														assign node6322 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node6325 = (inp[0]) ? node6329 : node6326;
														assign node6326 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node6329 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node6332 = (inp[9]) ? node6344 : node6333;
													assign node6333 = (inp[11]) ? node6339 : node6334;
														assign node6334 = (inp[5]) ? 4'b1000 : node6335;
															assign node6335 = (inp[14]) ? 4'b1000 : 4'b1000;
														assign node6339 = (inp[0]) ? 4'b1001 : node6340;
															assign node6340 = (inp[5]) ? 4'b1000 : 4'b1000;
													assign node6344 = (inp[11]) ? 4'b1000 : node6345;
														assign node6345 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node6349 = (inp[5]) ? node6359 : node6350;
												assign node6350 = (inp[14]) ? node6356 : node6351;
													assign node6351 = (inp[0]) ? 4'b1101 : node6352;
														assign node6352 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node6356 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node6359 = (inp[0]) ? node6369 : node6360;
													assign node6360 = (inp[11]) ? node6366 : node6361;
														assign node6361 = (inp[10]) ? node6363 : 4'b1001;
															assign node6363 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node6366 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node6369 = (inp[10]) ? node6371 : 4'b1001;
														assign node6371 = (inp[14]) ? 4'b1001 : 4'b1000;
						assign node6374 = (inp[1]) ? node6784 : node6375;
							assign node6375 = (inp[2]) ? node6587 : node6376;
								assign node6376 = (inp[14]) ? node6490 : node6377;
									assign node6377 = (inp[4]) ? node6437 : node6378;
										assign node6378 = (inp[12]) ? node6404 : node6379;
											assign node6379 = (inp[0]) ? node6389 : node6380;
												assign node6380 = (inp[5]) ? node6384 : node6381;
													assign node6381 = (inp[15]) ? 4'b1101 : 4'b1001;
													assign node6384 = (inp[15]) ? node6386 : 4'b1101;
														assign node6386 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node6389 = (inp[15]) ? node6399 : node6390;
													assign node6390 = (inp[5]) ? node6392 : 4'b1000;
														assign node6392 = (inp[9]) ? node6396 : node6393;
															assign node6393 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node6396 = (inp[10]) ? 4'b1100 : 4'b1100;
													assign node6399 = (inp[5]) ? node6401 : 4'b1101;
														assign node6401 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node6404 = (inp[9]) ? node6414 : node6405;
												assign node6405 = (inp[5]) ? node6411 : node6406;
													assign node6406 = (inp[0]) ? node6408 : 4'b1111;
														assign node6408 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node6411 = (inp[15]) ? 4'b1010 : 4'b1110;
												assign node6414 = (inp[5]) ? node6426 : node6415;
													assign node6415 = (inp[15]) ? node6421 : node6416;
														assign node6416 = (inp[10]) ? 4'b1010 : node6417;
															assign node6417 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node6421 = (inp[0]) ? node6423 : 4'b1110;
															assign node6423 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node6426 = (inp[15]) ? node6432 : node6427;
														assign node6427 = (inp[11]) ? 4'b1111 : node6428;
															assign node6428 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node6432 = (inp[10]) ? 4'b1011 : node6433;
															assign node6433 = (inp[0]) ? 4'b1011 : 4'b1010;
										assign node6437 = (inp[12]) ? node6461 : node6438;
											assign node6438 = (inp[15]) ? node6450 : node6439;
												assign node6439 = (inp[5]) ? node6443 : node6440;
													assign node6440 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node6443 = (inp[0]) ? node6447 : node6444;
														assign node6444 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node6447 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node6450 = (inp[10]) ? 4'b1011 : node6451;
													assign node6451 = (inp[5]) ? node6455 : node6452;
														assign node6452 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node6455 = (inp[9]) ? 4'b1010 : node6456;
															assign node6456 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node6461 = (inp[15]) ? node6481 : node6462;
												assign node6462 = (inp[10]) ? node6470 : node6463;
													assign node6463 = (inp[9]) ? node6465 : 4'b1000;
														assign node6465 = (inp[11]) ? node6467 : 4'b1000;
															assign node6467 = (inp[5]) ? 4'b1000 : 4'b1001;
													assign node6470 = (inp[11]) ? node6474 : node6471;
														assign node6471 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node6474 = (inp[9]) ? node6478 : node6475;
															assign node6475 = (inp[5]) ? 4'b1001 : 4'b1000;
															assign node6478 = (inp[5]) ? 4'b1000 : 4'b1000;
												assign node6481 = (inp[5]) ? node6487 : node6482;
													assign node6482 = (inp[9]) ? 4'b1100 : node6483;
														assign node6483 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node6487 = (inp[10]) ? 4'b1001 : 4'b1000;
									assign node6490 = (inp[4]) ? node6550 : node6491;
										assign node6491 = (inp[12]) ? node6521 : node6492;
											assign node6492 = (inp[5]) ? node6504 : node6493;
												assign node6493 = (inp[0]) ? node6499 : node6494;
													assign node6494 = (inp[11]) ? node6496 : 4'b1000;
														assign node6496 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node6499 = (inp[15]) ? 4'b1001 : node6500;
														assign node6500 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node6504 = (inp[15]) ? node6510 : node6505;
													assign node6505 = (inp[0]) ? node6507 : 4'b1000;
														assign node6507 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node6510 = (inp[0]) ? node6516 : node6511;
														assign node6511 = (inp[10]) ? 4'b1100 : node6512;
															assign node6512 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node6516 = (inp[11]) ? 4'b1101 : node6517;
															assign node6517 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node6521 = (inp[15]) ? node6537 : node6522;
												assign node6522 = (inp[5]) ? node6530 : node6523;
													assign node6523 = (inp[11]) ? 4'b1111 : node6524;
														assign node6524 = (inp[9]) ? node6526 : 4'b1110;
															assign node6526 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node6530 = (inp[11]) ? node6532 : 4'b1011;
														assign node6532 = (inp[9]) ? 4'b1011 : node6533;
															assign node6533 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node6537 = (inp[11]) ? node6545 : node6538;
													assign node6538 = (inp[0]) ? node6542 : node6539;
														assign node6539 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node6542 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node6545 = (inp[0]) ? 4'b1010 : node6546;
														assign node6546 = (inp[5]) ? 4'b1011 : 4'b1010;
										assign node6550 = (inp[12]) ? node6568 : node6551;
											assign node6551 = (inp[15]) ? node6559 : node6552;
												assign node6552 = (inp[0]) ? node6556 : node6553;
													assign node6553 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node6556 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node6559 = (inp[0]) ? 4'b1010 : node6560;
													assign node6560 = (inp[9]) ? node6562 : 4'b1011;
														assign node6562 = (inp[11]) ? 4'b1010 : node6563;
															assign node6563 = (inp[10]) ? 4'b1011 : 4'b1010;
											assign node6568 = (inp[11]) ? node6576 : node6569;
												assign node6569 = (inp[0]) ? node6573 : node6570;
													assign node6570 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node6573 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node6576 = (inp[0]) ? node6582 : node6577;
													assign node6577 = (inp[10]) ? 4'b1000 : node6578;
														assign node6578 = (inp[15]) ? 4'b1000 : 4'b1001;
													assign node6582 = (inp[10]) ? node6584 : 4'b1001;
														assign node6584 = (inp[15]) ? 4'b1000 : 4'b1001;
								assign node6587 = (inp[4]) ? node6705 : node6588;
									assign node6588 = (inp[12]) ? node6652 : node6589;
										assign node6589 = (inp[9]) ? node6621 : node6590;
											assign node6590 = (inp[0]) ? node6608 : node6591;
												assign node6591 = (inp[5]) ? node6599 : node6592;
													assign node6592 = (inp[10]) ? node6594 : 4'b1100;
														assign node6594 = (inp[14]) ? 4'b1101 : node6595;
															assign node6595 = (inp[11]) ? 4'b1001 : 4'b1101;
													assign node6599 = (inp[10]) ? node6603 : node6600;
														assign node6600 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node6603 = (inp[11]) ? node6605 : 4'b1001;
															assign node6605 = (inp[14]) ? 4'b1101 : 4'b1001;
												assign node6608 = (inp[15]) ? node6614 : node6609;
													assign node6609 = (inp[10]) ? node6611 : 4'b1101;
														assign node6611 = (inp[5]) ? 4'b1100 : 4'b1101;
													assign node6614 = (inp[14]) ? node6618 : node6615;
														assign node6615 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node6618 = (inp[10]) ? 4'b1100 : 4'b1001;
											assign node6621 = (inp[15]) ? node6635 : node6622;
												assign node6622 = (inp[14]) ? node6630 : node6623;
													assign node6623 = (inp[5]) ? 4'b1000 : node6624;
														assign node6624 = (inp[10]) ? node6626 : 4'b1100;
															assign node6626 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node6630 = (inp[10]) ? node6632 : 4'b1101;
														assign node6632 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node6635 = (inp[0]) ? node6645 : node6636;
													assign node6636 = (inp[10]) ? node6640 : node6637;
														assign node6637 = (inp[5]) ? 4'b1000 : 4'b1100;
														assign node6640 = (inp[5]) ? node6642 : 4'b1001;
															assign node6642 = (inp[14]) ? 4'b1000 : 4'b1100;
													assign node6645 = (inp[10]) ? node6649 : node6646;
														assign node6646 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node6649 = (inp[14]) ? 4'b1100 : 4'b1000;
										assign node6652 = (inp[14]) ? node6678 : node6653;
											assign node6653 = (inp[9]) ? node6665 : node6654;
												assign node6654 = (inp[10]) ? node6656 : 4'b1010;
													assign node6656 = (inp[15]) ? node6662 : node6657;
														assign node6657 = (inp[5]) ? node6659 : 4'b1111;
															assign node6659 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node6662 = (inp[5]) ? 4'b1110 : 4'b1010;
												assign node6665 = (inp[15]) ? node6675 : node6666;
													assign node6666 = (inp[5]) ? node6670 : node6667;
														assign node6667 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node6670 = (inp[11]) ? node6672 : 4'b1011;
															assign node6672 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node6675 = (inp[5]) ? 4'b1111 : 4'b1011;
											assign node6678 = (inp[15]) ? node6692 : node6679;
												assign node6679 = (inp[5]) ? node6685 : node6680;
													assign node6680 = (inp[11]) ? node6682 : 4'b1011;
														assign node6682 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node6685 = (inp[9]) ? node6687 : 4'b1111;
														assign node6687 = (inp[0]) ? node6689 : 4'b1111;
															assign node6689 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node6692 = (inp[10]) ? node6698 : node6693;
													assign node6693 = (inp[0]) ? node6695 : 4'b1110;
														assign node6695 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node6698 = (inp[0]) ? 4'b1110 : node6699;
														assign node6699 = (inp[5]) ? 4'b1111 : node6700;
															assign node6700 = (inp[11]) ? 4'b1111 : 4'b1110;
									assign node6705 = (inp[12]) ? node6741 : node6706;
										assign node6706 = (inp[5]) ? node6724 : node6707;
											assign node6707 = (inp[0]) ? node6715 : node6708;
												assign node6708 = (inp[10]) ? node6712 : node6709;
													assign node6709 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node6712 = (inp[15]) ? 4'b1110 : 4'b1111;
												assign node6715 = (inp[10]) ? 4'b1111 : node6716;
													assign node6716 = (inp[9]) ? node6718 : 4'b1111;
														assign node6718 = (inp[11]) ? node6720 : 4'b1110;
															assign node6720 = (inp[14]) ? 4'b1110 : 4'b1111;
											assign node6724 = (inp[15]) ? node6736 : node6725;
												assign node6725 = (inp[14]) ? node6733 : node6726;
													assign node6726 = (inp[11]) ? 4'b1010 : node6727;
														assign node6727 = (inp[10]) ? 4'b1011 : node6728;
															assign node6728 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node6733 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node6736 = (inp[0]) ? 4'b1110 : node6737;
													assign node6737 = (inp[9]) ? 4'b1110 : 4'b1111;
										assign node6741 = (inp[10]) ? node6765 : node6742;
											assign node6742 = (inp[0]) ? node6750 : node6743;
												assign node6743 = (inp[11]) ? node6745 : 4'b1101;
													assign node6745 = (inp[5]) ? 4'b1100 : node6746;
														assign node6746 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node6750 = (inp[11]) ? node6758 : node6751;
													assign node6751 = (inp[15]) ? node6755 : node6752;
														assign node6752 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node6755 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node6758 = (inp[14]) ? 4'b1101 : node6759;
														assign node6759 = (inp[15]) ? 4'b1001 : node6760;
															assign node6760 = (inp[5]) ? 4'b1101 : 4'b1100;
											assign node6765 = (inp[0]) ? node6779 : node6766;
												assign node6766 = (inp[11]) ? node6774 : node6767;
													assign node6767 = (inp[15]) ? node6771 : node6768;
														assign node6768 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node6771 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node6774 = (inp[9]) ? node6776 : 4'b1101;
														assign node6776 = (inp[5]) ? 4'b1101 : 4'b1001;
												assign node6779 = (inp[5]) ? 4'b1100 : node6780;
													assign node6780 = (inp[14]) ? 4'b1100 : 4'b1101;
							assign node6784 = (inp[2]) ? node6974 : node6785;
								assign node6785 = (inp[4]) ? node6887 : node6786;
									assign node6786 = (inp[12]) ? node6832 : node6787;
										assign node6787 = (inp[11]) ? node6805 : node6788;
											assign node6788 = (inp[14]) ? node6796 : node6789;
												assign node6789 = (inp[5]) ? node6793 : node6790;
													assign node6790 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node6793 = (inp[15]) ? 4'b1100 : 4'b1000;
												assign node6796 = (inp[0]) ? node6802 : node6797;
													assign node6797 = (inp[10]) ? 4'b1101 : node6798;
														assign node6798 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node6802 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node6805 = (inp[14]) ? node6819 : node6806;
												assign node6806 = (inp[9]) ? node6814 : node6807;
													assign node6807 = (inp[5]) ? node6811 : node6808;
														assign node6808 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node6811 = (inp[15]) ? 4'b1101 : 4'b1001;
													assign node6814 = (inp[0]) ? 4'b1000 : node6815;
														assign node6815 = (inp[5]) ? 4'b1101 : 4'b1000;
												assign node6819 = (inp[15]) ? node6827 : node6820;
													assign node6820 = (inp[0]) ? node6822 : 4'b1101;
														assign node6822 = (inp[5]) ? 4'b1100 : node6823;
															assign node6823 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node6827 = (inp[5]) ? 4'b1000 : node6828;
														assign node6828 = (inp[10]) ? 4'b1101 : 4'b1100;
										assign node6832 = (inp[15]) ? node6868 : node6833;
											assign node6833 = (inp[10]) ? node6855 : node6834;
												assign node6834 = (inp[11]) ? node6846 : node6835;
													assign node6835 = (inp[14]) ? node6839 : node6836;
														assign node6836 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node6839 = (inp[5]) ? node6843 : node6840;
															assign node6840 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node6843 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node6846 = (inp[0]) ? node6852 : node6847;
														assign node6847 = (inp[5]) ? 4'b1111 : node6848;
															assign node6848 = (inp[14]) ? 4'b1010 : 4'b1110;
														assign node6852 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node6855 = (inp[9]) ? node6865 : node6856;
													assign node6856 = (inp[14]) ? node6860 : node6857;
														assign node6857 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node6860 = (inp[5]) ? node6862 : 4'b1010;
															assign node6862 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node6865 = (inp[11]) ? 4'b1010 : 4'b1110;
											assign node6868 = (inp[10]) ? node6876 : node6869;
												assign node6869 = (inp[0]) ? 4'b1110 : node6870;
													assign node6870 = (inp[5]) ? 4'b1111 : node6871;
														assign node6871 = (inp[14]) ? 4'b1110 : 4'b1010;
												assign node6876 = (inp[11]) ? 4'b1111 : node6877;
													assign node6877 = (inp[5]) ? node6883 : node6878;
														assign node6878 = (inp[14]) ? node6880 : 4'b1011;
															assign node6880 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node6883 = (inp[0]) ? 4'b1111 : 4'b1110;
									assign node6887 = (inp[12]) ? node6927 : node6888;
										assign node6888 = (inp[10]) ? node6912 : node6889;
											assign node6889 = (inp[0]) ? node6903 : node6890;
												assign node6890 = (inp[15]) ? node6896 : node6891;
													assign node6891 = (inp[5]) ? node6893 : 4'b1110;
														assign node6893 = (inp[11]) ? 4'b1110 : 4'b1010;
													assign node6896 = (inp[5]) ? 4'b1110 : node6897;
														assign node6897 = (inp[9]) ? 4'b1110 : node6898;
															assign node6898 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node6903 = (inp[14]) ? 4'b1111 : node6904;
													assign node6904 = (inp[15]) ? node6908 : node6905;
														assign node6905 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node6908 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node6912 = (inp[0]) ? node6920 : node6913;
												assign node6913 = (inp[14]) ? 4'b1111 : node6914;
													assign node6914 = (inp[11]) ? node6916 : 4'b1111;
														assign node6916 = (inp[5]) ? 4'b1111 : 4'b1110;
												assign node6920 = (inp[14]) ? 4'b1110 : node6921;
													assign node6921 = (inp[11]) ? node6923 : 4'b1110;
														assign node6923 = (inp[5]) ? 4'b1110 : 4'b1111;
										assign node6927 = (inp[14]) ? node6949 : node6928;
											assign node6928 = (inp[5]) ? node6938 : node6929;
												assign node6929 = (inp[15]) ? node6933 : node6930;
													assign node6930 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node6933 = (inp[9]) ? node6935 : 4'b1001;
														assign node6935 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node6938 = (inp[15]) ? node6940 : 4'b1100;
													assign node6940 = (inp[9]) ? node6946 : node6941;
														assign node6941 = (inp[0]) ? 4'b1100 : node6942;
															assign node6942 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node6946 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node6949 = (inp[9]) ? node6963 : node6950;
												assign node6950 = (inp[5]) ? node6958 : node6951;
													assign node6951 = (inp[0]) ? node6955 : node6952;
														assign node6952 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node6955 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node6958 = (inp[10]) ? 4'b1101 : node6959;
														assign node6959 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node6963 = (inp[11]) ? node6967 : node6964;
													assign node6964 = (inp[5]) ? 4'b1100 : 4'b1101;
													assign node6967 = (inp[5]) ? node6969 : 4'b1100;
														assign node6969 = (inp[15]) ? node6971 : 4'b1101;
															assign node6971 = (inp[0]) ? 4'b1100 : 4'b1100;
								assign node6974 = (inp[4]) ? node7088 : node6975;
									assign node6975 = (inp[12]) ? node7017 : node6976;
										assign node6976 = (inp[14]) ? node7002 : node6977;
											assign node6977 = (inp[9]) ? node6987 : node6978;
												assign node6978 = (inp[0]) ? node6982 : node6979;
													assign node6979 = (inp[15]) ? 4'b1001 : 4'b1100;
													assign node6982 = (inp[15]) ? node6984 : 4'b1000;
														assign node6984 = (inp[5]) ? 4'b1000 : 4'b1100;
												assign node6987 = (inp[11]) ? node6997 : node6988;
													assign node6988 = (inp[15]) ? node6992 : node6989;
														assign node6989 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node6992 = (inp[10]) ? 4'b1100 : node6993;
															assign node6993 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node6997 = (inp[15]) ? node6999 : 4'b1100;
														assign node6999 = (inp[0]) ? 4'b1000 : 4'b1100;
											assign node7002 = (inp[5]) ? node7010 : node7003;
												assign node7003 = (inp[0]) ? node7007 : node7004;
													assign node7004 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node7007 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node7010 = (inp[15]) ? node7012 : 4'b1000;
													assign node7012 = (inp[0]) ? node7014 : 4'b1100;
														assign node7014 = (inp[10]) ? 4'b1100 : 4'b1101;
										assign node7017 = (inp[15]) ? node7057 : node7018;
											assign node7018 = (inp[5]) ? node7042 : node7019;
												assign node7019 = (inp[14]) ? node7031 : node7020;
													assign node7020 = (inp[9]) ? node7026 : node7021;
														assign node7021 = (inp[0]) ? node7023 : 4'b1011;
															assign node7023 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node7026 = (inp[10]) ? node7028 : 4'b1010;
															assign node7028 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node7031 = (inp[9]) ? node7037 : node7032;
														assign node7032 = (inp[0]) ? node7034 : 4'b1110;
															assign node7034 = (inp[10]) ? 4'b1110 : 4'b1110;
														assign node7037 = (inp[0]) ? node7039 : 4'b1111;
															assign node7039 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node7042 = (inp[14]) ? node7054 : node7043;
													assign node7043 = (inp[11]) ? node7049 : node7044;
														assign node7044 = (inp[9]) ? node7046 : 4'b1111;
															assign node7046 = (inp[0]) ? 4'b1110 : 4'b1110;
														assign node7049 = (inp[9]) ? node7051 : 4'b1110;
															assign node7051 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node7054 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node7057 = (inp[14]) ? node7075 : node7058;
												assign node7058 = (inp[5]) ? node7072 : node7059;
													assign node7059 = (inp[9]) ? node7065 : node7060;
														assign node7060 = (inp[10]) ? node7062 : 4'b1110;
															assign node7062 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node7065 = (inp[10]) ? node7069 : node7066;
															assign node7066 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node7069 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node7072 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node7075 = (inp[10]) ? node7079 : node7076;
													assign node7076 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node7079 = (inp[0]) ? node7083 : node7080;
														assign node7080 = (inp[5]) ? 4'b1011 : 4'b1010;
														assign node7083 = (inp[5]) ? 4'b1010 : node7084;
															assign node7084 = (inp[11]) ? 4'b1010 : 4'b1011;
									assign node7088 = (inp[12]) ? node7122 : node7089;
										assign node7089 = (inp[14]) ? node7115 : node7090;
											assign node7090 = (inp[15]) ? node7102 : node7091;
												assign node7091 = (inp[5]) ? node7097 : node7092;
													assign node7092 = (inp[0]) ? node7094 : 4'b1010;
														assign node7094 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node7097 = (inp[9]) ? 4'b1111 : node7098;
														assign node7098 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node7102 = (inp[11]) ? node7110 : node7103;
													assign node7103 = (inp[0]) ? node7105 : 4'b1010;
														assign node7105 = (inp[5]) ? 4'b1011 : node7106;
															assign node7106 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node7110 = (inp[0]) ? node7112 : 4'b1011;
														assign node7112 = (inp[10]) ? 4'b1010 : 4'b1011;
											assign node7115 = (inp[10]) ? node7119 : node7116;
												assign node7116 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node7119 = (inp[0]) ? 4'b1010 : 4'b1011;
										assign node7122 = (inp[15]) ? node7138 : node7123;
											assign node7123 = (inp[0]) ? node7131 : node7124;
												assign node7124 = (inp[10]) ? 4'b1001 : node7125;
													assign node7125 = (inp[5]) ? node7127 : 4'b1000;
														assign node7127 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node7131 = (inp[10]) ? node7133 : 4'b1001;
													assign node7133 = (inp[11]) ? 4'b1000 : node7134;
														assign node7134 = (inp[5]) ? 4'b1001 : 4'b1000;
											assign node7138 = (inp[5]) ? node7156 : node7139;
												assign node7139 = (inp[14]) ? node7149 : node7140;
													assign node7140 = (inp[9]) ? node7142 : 4'b1101;
														assign node7142 = (inp[11]) ? node7146 : node7143;
															assign node7143 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node7146 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node7149 = (inp[11]) ? 4'b1001 : node7150;
														assign node7150 = (inp[0]) ? node7152 : 4'b1000;
															assign node7152 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node7156 = (inp[0]) ? 4'b1000 : node7157;
													assign node7157 = (inp[14]) ? 4'b1000 : node7158;
														assign node7158 = (inp[9]) ? node7160 : 4'b1001;
															assign node7160 = (inp[10]) ? 4'b1000 : 4'b1000;
			assign node7165 = (inp[14]) ? node10463 : node7166;
				assign node7166 = (inp[8]) ? node8866 : node7167;
					assign node7167 = (inp[7]) ? node8059 : node7168;
						assign node7168 = (inp[15]) ? node7634 : node7169;
							assign node7169 = (inp[10]) ? node7429 : node7170;
								assign node7170 = (inp[1]) ? node7294 : node7171;
									assign node7171 = (inp[2]) ? node7237 : node7172;
										assign node7172 = (inp[0]) ? node7200 : node7173;
											assign node7173 = (inp[13]) ? node7185 : node7174;
												assign node7174 = (inp[5]) ? node7180 : node7175;
													assign node7175 = (inp[9]) ? node7177 : 4'b1000;
														assign node7177 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node7180 = (inp[11]) ? 4'b1101 : node7181;
														assign node7181 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node7185 = (inp[12]) ? node7193 : node7186;
													assign node7186 = (inp[9]) ? node7188 : 4'b1001;
														assign node7188 = (inp[4]) ? node7190 : 4'b1001;
															assign node7190 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node7193 = (inp[9]) ? 4'b1100 : node7194;
														assign node7194 = (inp[11]) ? node7196 : 4'b1101;
															assign node7196 = (inp[4]) ? 4'b1000 : 4'b1001;
											assign node7200 = (inp[4]) ? node7222 : node7201;
												assign node7201 = (inp[9]) ? node7209 : node7202;
													assign node7202 = (inp[12]) ? 4'b1000 : node7203;
														assign node7203 = (inp[11]) ? 4'b1101 : node7204;
															assign node7204 = (inp[5]) ? 4'b1100 : 4'b1000;
													assign node7209 = (inp[12]) ? node7217 : node7210;
														assign node7210 = (inp[11]) ? node7214 : node7211;
															assign node7211 = (inp[5]) ? 4'b1000 : 4'b1001;
															assign node7214 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node7217 = (inp[11]) ? node7219 : 4'b1101;
															assign node7219 = (inp[13]) ? 4'b1000 : 4'b1100;
												assign node7222 = (inp[11]) ? node7228 : node7223;
													assign node7223 = (inp[9]) ? node7225 : 4'b1101;
														assign node7225 = (inp[12]) ? 4'b1100 : 4'b1101;
													assign node7228 = (inp[12]) ? node7230 : 4'b1100;
														assign node7230 = (inp[5]) ? node7234 : node7231;
															assign node7231 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node7234 = (inp[13]) ? 4'b1101 : 4'b1001;
										assign node7237 = (inp[5]) ? node7261 : node7238;
											assign node7238 = (inp[13]) ? node7256 : node7239;
												assign node7239 = (inp[12]) ? node7251 : node7240;
													assign node7240 = (inp[0]) ? node7246 : node7241;
														assign node7241 = (inp[9]) ? node7243 : 4'b1001;
															assign node7243 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node7246 = (inp[11]) ? node7248 : 4'b1001;
															assign node7248 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node7251 = (inp[4]) ? 4'b1100 : node7252;
														assign node7252 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node7256 = (inp[12]) ? 4'b1001 : node7257;
													assign node7257 = (inp[4]) ? 4'b1100 : 4'b1101;
											assign node7261 = (inp[13]) ? node7283 : node7262;
												assign node7262 = (inp[4]) ? node7276 : node7263;
													assign node7263 = (inp[9]) ? node7271 : node7264;
														assign node7264 = (inp[0]) ? node7268 : node7265;
															assign node7265 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node7268 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node7271 = (inp[11]) ? 4'b1101 : node7272;
															assign node7272 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node7276 = (inp[12]) ? node7278 : 4'b1101;
														assign node7278 = (inp[11]) ? node7280 : 4'b1000;
															assign node7280 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node7283 = (inp[11]) ? node7291 : node7284;
													assign node7284 = (inp[12]) ? node7286 : 4'b1001;
														assign node7286 = (inp[4]) ? node7288 : 4'b1001;
															assign node7288 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node7291 = (inp[9]) ? 4'b1001 : 4'b1000;
									assign node7294 = (inp[4]) ? node7368 : node7295;
										assign node7295 = (inp[13]) ? node7333 : node7296;
											assign node7296 = (inp[0]) ? node7320 : node7297;
												assign node7297 = (inp[9]) ? node7311 : node7298;
													assign node7298 = (inp[2]) ? node7306 : node7299;
														assign node7299 = (inp[12]) ? node7303 : node7300;
															assign node7300 = (inp[5]) ? 4'b1100 : 4'b1000;
															assign node7303 = (inp[11]) ? 4'b1000 : 4'b1101;
														assign node7306 = (inp[11]) ? node7308 : 4'b1100;
															assign node7308 = (inp[12]) ? 4'b1100 : 4'b1101;
													assign node7311 = (inp[11]) ? node7315 : node7312;
														assign node7312 = (inp[12]) ? 4'b1100 : 4'b1001;
														assign node7315 = (inp[12]) ? 4'b1000 : node7316;
															assign node7316 = (inp[5]) ? 4'b1100 : 4'b1000;
												assign node7320 = (inp[12]) ? node7328 : node7321;
													assign node7321 = (inp[9]) ? 4'b1001 : node7322;
														assign node7322 = (inp[2]) ? node7324 : 4'b1001;
															assign node7324 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node7328 = (inp[5]) ? node7330 : 4'b1100;
														assign node7330 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node7333 = (inp[5]) ? node7349 : node7334;
												assign node7334 = (inp[12]) ? node7344 : node7335;
													assign node7335 = (inp[9]) ? node7341 : node7336;
														assign node7336 = (inp[11]) ? node7338 : 4'b1100;
															assign node7338 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node7341 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node7344 = (inp[9]) ? node7346 : 4'b1000;
														assign node7346 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node7349 = (inp[12]) ? node7357 : node7350;
													assign node7350 = (inp[2]) ? node7352 : 4'b1001;
														assign node7352 = (inp[0]) ? node7354 : 4'b1001;
															assign node7354 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node7357 = (inp[9]) ? node7363 : node7358;
														assign node7358 = (inp[11]) ? 4'b1101 : node7359;
															assign node7359 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node7363 = (inp[0]) ? 4'b1100 : node7364;
															assign node7364 = (inp[2]) ? 4'b1100 : 4'b1101;
										assign node7368 = (inp[9]) ? node7404 : node7369;
											assign node7369 = (inp[11]) ? node7387 : node7370;
												assign node7370 = (inp[0]) ? node7380 : node7371;
													assign node7371 = (inp[5]) ? node7377 : node7372;
														assign node7372 = (inp[13]) ? 4'b1101 : node7373;
															assign node7373 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node7377 = (inp[13]) ? 4'b1000 : 4'b1100;
													assign node7380 = (inp[12]) ? node7384 : node7381;
														assign node7381 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node7384 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node7387 = (inp[12]) ? node7397 : node7388;
													assign node7388 = (inp[13]) ? node7392 : node7389;
														assign node7389 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node7392 = (inp[5]) ? node7394 : 4'b1101;
															assign node7394 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node7397 = (inp[5]) ? node7401 : node7398;
														assign node7398 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node7401 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node7404 = (inp[13]) ? node7420 : node7405;
												assign node7405 = (inp[5]) ? node7413 : node7406;
													assign node7406 = (inp[11]) ? node7410 : node7407;
														assign node7407 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node7410 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node7413 = (inp[12]) ? 4'b1101 : node7414;
														assign node7414 = (inp[0]) ? node7416 : 4'b1100;
															assign node7416 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node7420 = (inp[5]) ? node7422 : 4'b1100;
													assign node7422 = (inp[11]) ? node7424 : 4'b1000;
														assign node7424 = (inp[12]) ? node7426 : 4'b1001;
															assign node7426 = (inp[0]) ? 4'b1001 : 4'b1000;
								assign node7429 = (inp[9]) ? node7521 : node7430;
									assign node7430 = (inp[11]) ? node7476 : node7431;
										assign node7431 = (inp[12]) ? node7443 : node7432;
											assign node7432 = (inp[5]) ? node7436 : node7433;
												assign node7433 = (inp[13]) ? 4'b1100 : 4'b1000;
												assign node7436 = (inp[13]) ? 4'b1001 : node7437;
													assign node7437 = (inp[2]) ? 4'b1101 : node7438;
														assign node7438 = (inp[4]) ? 4'b1101 : 4'b1100;
											assign node7443 = (inp[0]) ? node7463 : node7444;
												assign node7444 = (inp[13]) ? node7450 : node7445;
													assign node7445 = (inp[2]) ? 4'b1101 : node7446;
														assign node7446 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node7450 = (inp[4]) ? node7456 : node7451;
														assign node7451 = (inp[1]) ? node7453 : 4'b1001;
															assign node7453 = (inp[5]) ? 4'b1100 : 4'b1001;
														assign node7456 = (inp[5]) ? node7460 : node7457;
															assign node7457 = (inp[1]) ? 4'b1101 : 4'b1000;
															assign node7460 = (inp[1]) ? 4'b1000 : 4'b1100;
												assign node7463 = (inp[13]) ? node7469 : node7464;
													assign node7464 = (inp[1]) ? node7466 : 4'b1100;
														assign node7466 = (inp[5]) ? 4'b1100 : 4'b1001;
													assign node7469 = (inp[1]) ? node7471 : 4'b1001;
														assign node7471 = (inp[4]) ? 4'b1101 : node7472;
															assign node7472 = (inp[2]) ? 4'b1000 : 4'b1100;
										assign node7476 = (inp[5]) ? node7498 : node7477;
											assign node7477 = (inp[13]) ? node7489 : node7478;
												assign node7478 = (inp[1]) ? node7484 : node7479;
													assign node7479 = (inp[2]) ? node7481 : 4'b1001;
														assign node7481 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node7484 = (inp[0]) ? 4'b1001 : node7485;
														assign node7485 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node7489 = (inp[0]) ? 4'b1101 : node7490;
													assign node7490 = (inp[12]) ? node7492 : 4'b1101;
														assign node7492 = (inp[4]) ? 4'b1001 : node7493;
															assign node7493 = (inp[1]) ? 4'b1001 : 4'b1101;
											assign node7498 = (inp[13]) ? node7512 : node7499;
												assign node7499 = (inp[0]) ? node7501 : 4'b1101;
													assign node7501 = (inp[2]) ? node7509 : node7502;
														assign node7502 = (inp[4]) ? node7506 : node7503;
															assign node7503 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node7506 = (inp[12]) ? 4'b1101 : 4'b1100;
														assign node7509 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node7512 = (inp[1]) ? node7514 : 4'b1100;
													assign node7514 = (inp[12]) ? node7518 : node7515;
														assign node7515 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node7518 = (inp[4]) ? 4'b1001 : 4'b1101;
									assign node7521 = (inp[11]) ? node7587 : node7522;
										assign node7522 = (inp[2]) ? node7556 : node7523;
											assign node7523 = (inp[5]) ? node7539 : node7524;
												assign node7524 = (inp[12]) ? node7528 : node7525;
													assign node7525 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node7528 = (inp[0]) ? node7532 : node7529;
														assign node7529 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node7532 = (inp[13]) ? node7536 : node7533;
															assign node7533 = (inp[4]) ? 4'b1101 : 4'b1100;
															assign node7536 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node7539 = (inp[13]) ? node7549 : node7540;
													assign node7540 = (inp[1]) ? node7546 : node7541;
														assign node7541 = (inp[4]) ? node7543 : 4'b1101;
															assign node7543 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node7546 = (inp[4]) ? 4'b1101 : 4'b1000;
													assign node7549 = (inp[1]) ? node7551 : 4'b1000;
														assign node7551 = (inp[12]) ? node7553 : 4'b1000;
															assign node7553 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node7556 = (inp[0]) ? node7572 : node7557;
												assign node7557 = (inp[4]) ? node7561 : node7558;
													assign node7558 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node7561 = (inp[13]) ? node7567 : node7562;
														assign node7562 = (inp[5]) ? 4'b1100 : node7563;
															assign node7563 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node7567 = (inp[12]) ? node7569 : 4'b1100;
															assign node7569 = (inp[5]) ? 4'b1101 : 4'b1001;
												assign node7572 = (inp[5]) ? node7582 : node7573;
													assign node7573 = (inp[1]) ? node7579 : node7574;
														assign node7574 = (inp[4]) ? node7576 : 4'b1100;
															assign node7576 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node7579 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node7582 = (inp[1]) ? node7584 : 4'b1000;
														assign node7584 = (inp[12]) ? 4'b1101 : 4'b1000;
										assign node7587 = (inp[5]) ? node7599 : node7588;
											assign node7588 = (inp[13]) ? node7594 : node7589;
												assign node7589 = (inp[12]) ? node7591 : 4'b1000;
													assign node7591 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node7594 = (inp[4]) ? node7596 : 4'b1100;
													assign node7596 = (inp[1]) ? 4'b1100 : 4'b1001;
											assign node7599 = (inp[13]) ? node7617 : node7600;
												assign node7600 = (inp[12]) ? node7604 : node7601;
													assign node7601 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node7604 = (inp[0]) ? node7610 : node7605;
														assign node7605 = (inp[1]) ? node7607 : 4'b1000;
															assign node7607 = (inp[4]) ? 4'b1101 : 4'b1000;
														assign node7610 = (inp[1]) ? node7614 : node7611;
															assign node7611 = (inp[4]) ? 4'b1001 : 4'b1100;
															assign node7614 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node7617 = (inp[12]) ? node7625 : node7618;
													assign node7618 = (inp[2]) ? node7620 : 4'b1001;
														assign node7620 = (inp[4]) ? node7622 : 4'b1001;
															assign node7622 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node7625 = (inp[1]) ? node7629 : node7626;
														assign node7626 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node7629 = (inp[4]) ? 4'b1000 : node7630;
															assign node7630 = (inp[2]) ? 4'b1100 : 4'b1101;
							assign node7634 = (inp[5]) ? node7862 : node7635;
								assign node7635 = (inp[13]) ? node7763 : node7636;
									assign node7636 = (inp[1]) ? node7690 : node7637;
										assign node7637 = (inp[10]) ? node7657 : node7638;
											assign node7638 = (inp[4]) ? node7644 : node7639;
												assign node7639 = (inp[9]) ? 4'b1011 : node7640;
													assign node7640 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node7644 = (inp[0]) ? node7646 : 4'b1010;
													assign node7646 = (inp[12]) ? node7652 : node7647;
														assign node7647 = (inp[11]) ? node7649 : 4'b1011;
															assign node7649 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node7652 = (inp[2]) ? node7654 : 4'b1010;
															assign node7654 = (inp[9]) ? 4'b1010 : 4'b1010;
											assign node7657 = (inp[12]) ? node7675 : node7658;
												assign node7658 = (inp[11]) ? node7664 : node7659;
													assign node7659 = (inp[9]) ? 4'b1011 : node7660;
														assign node7660 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node7664 = (inp[9]) ? node7670 : node7665;
														assign node7665 = (inp[2]) ? node7667 : 4'b1011;
															assign node7667 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node7670 = (inp[4]) ? 4'b1010 : node7671;
															assign node7671 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node7675 = (inp[4]) ? node7685 : node7676;
													assign node7676 = (inp[2]) ? node7678 : 4'b1010;
														assign node7678 = (inp[9]) ? node7682 : node7679;
															assign node7679 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node7682 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node7685 = (inp[9]) ? 4'b1011 : node7686;
														assign node7686 = (inp[11]) ? 4'b1011 : 4'b1010;
										assign node7690 = (inp[11]) ? node7720 : node7691;
											assign node7691 = (inp[9]) ? node7709 : node7692;
												assign node7692 = (inp[2]) ? node7702 : node7693;
													assign node7693 = (inp[12]) ? node7699 : node7694;
														assign node7694 = (inp[0]) ? 4'b1111 : node7695;
															assign node7695 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node7699 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node7702 = (inp[10]) ? 4'b1110 : node7703;
														assign node7703 = (inp[12]) ? 4'b1110 : node7704;
															assign node7704 = (inp[4]) ? 4'b1110 : 4'b1011;
												assign node7709 = (inp[4]) ? node7717 : node7710;
													assign node7710 = (inp[12]) ? node7714 : node7711;
														assign node7711 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node7714 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node7717 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node7720 = (inp[10]) ? node7742 : node7721;
												assign node7721 = (inp[9]) ? node7733 : node7722;
													assign node7722 = (inp[4]) ? node7728 : node7723;
														assign node7723 = (inp[12]) ? node7725 : 4'b1010;
															assign node7725 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node7728 = (inp[0]) ? node7730 : 4'b1111;
															assign node7730 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node7733 = (inp[4]) ? node7739 : node7734;
														assign node7734 = (inp[12]) ? node7736 : 4'b1010;
															assign node7736 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node7739 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node7742 = (inp[0]) ? node7754 : node7743;
													assign node7743 = (inp[9]) ? node7747 : node7744;
														assign node7744 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node7747 = (inp[4]) ? node7751 : node7748;
															assign node7748 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node7751 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node7754 = (inp[4]) ? node7758 : node7755;
														assign node7755 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node7758 = (inp[12]) ? node7760 : 4'b1110;
															assign node7760 = (inp[9]) ? 4'b1010 : 4'b1011;
									assign node7763 = (inp[1]) ? node7807 : node7764;
										assign node7764 = (inp[12]) ? node7780 : node7765;
											assign node7765 = (inp[11]) ? node7775 : node7766;
												assign node7766 = (inp[9]) ? node7770 : node7767;
													assign node7767 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node7770 = (inp[0]) ? 4'b1110 : node7771;
														assign node7771 = (inp[4]) ? 4'b1111 : 4'b1110;
												assign node7775 = (inp[9]) ? node7777 : 4'b1110;
													assign node7777 = (inp[10]) ? 4'b1110 : 4'b1111;
											assign node7780 = (inp[2]) ? node7798 : node7781;
												assign node7781 = (inp[10]) ? node7791 : node7782;
													assign node7782 = (inp[4]) ? node7788 : node7783;
														assign node7783 = (inp[0]) ? node7785 : 4'b1110;
															assign node7785 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node7788 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node7791 = (inp[0]) ? node7793 : 4'b1110;
														assign node7793 = (inp[4]) ? node7795 : 4'b1111;
															assign node7795 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node7798 = (inp[4]) ? 4'b1111 : node7799;
													assign node7799 = (inp[10]) ? 4'b1111 : node7800;
														assign node7800 = (inp[11]) ? node7802 : 4'b1111;
															assign node7802 = (inp[9]) ? 4'b1110 : 4'b1110;
										assign node7807 = (inp[12]) ? node7833 : node7808;
											assign node7808 = (inp[4]) ? node7822 : node7809;
												assign node7809 = (inp[2]) ? node7817 : node7810;
													assign node7810 = (inp[10]) ? node7814 : node7811;
														assign node7811 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node7814 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node7817 = (inp[10]) ? node7819 : 4'b1111;
														assign node7819 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node7822 = (inp[11]) ? node7828 : node7823;
													assign node7823 = (inp[9]) ? node7825 : 4'b1010;
														assign node7825 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node7828 = (inp[9]) ? node7830 : 4'b1011;
														assign node7830 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node7833 = (inp[4]) ? node7845 : node7834;
												assign node7834 = (inp[2]) ? node7840 : node7835;
													assign node7835 = (inp[11]) ? 4'b1010 : node7836;
														assign node7836 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node7840 = (inp[9]) ? node7842 : 4'b1011;
														assign node7842 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node7845 = (inp[11]) ? node7853 : node7846;
													assign node7846 = (inp[10]) ? 4'b1111 : node7847;
														assign node7847 = (inp[2]) ? 4'b1110 : node7848;
															assign node7848 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node7853 = (inp[9]) ? node7859 : node7854;
														assign node7854 = (inp[0]) ? 4'b1110 : node7855;
															assign node7855 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node7859 = (inp[2]) ? 4'b1110 : 4'b1111;
								assign node7862 = (inp[13]) ? node7960 : node7863;
									assign node7863 = (inp[1]) ? node7919 : node7864;
										assign node7864 = (inp[12]) ? node7894 : node7865;
											assign node7865 = (inp[9]) ? node7885 : node7866;
												assign node7866 = (inp[11]) ? node7876 : node7867;
													assign node7867 = (inp[0]) ? node7869 : 4'b1110;
														assign node7869 = (inp[4]) ? node7873 : node7870;
															assign node7870 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node7873 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node7876 = (inp[0]) ? node7878 : 4'b1111;
														assign node7878 = (inp[2]) ? node7882 : node7879;
															assign node7879 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node7882 = (inp[4]) ? 4'b1111 : 4'b1110;
												assign node7885 = (inp[11]) ? node7887 : 4'b1111;
													assign node7887 = (inp[0]) ? node7889 : 4'b1110;
														assign node7889 = (inp[10]) ? 4'b1111 : node7890;
															assign node7890 = (inp[4]) ? 4'b1110 : 4'b1110;
											assign node7894 = (inp[2]) ? node7904 : node7895;
												assign node7895 = (inp[9]) ? 4'b1110 : node7896;
													assign node7896 = (inp[10]) ? node7900 : node7897;
														assign node7897 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node7900 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node7904 = (inp[11]) ? node7914 : node7905;
													assign node7905 = (inp[10]) ? node7909 : node7906;
														assign node7906 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node7909 = (inp[9]) ? 4'b1110 : node7910;
															assign node7910 = (inp[4]) ? 4'b1110 : 4'b1111;
													assign node7914 = (inp[0]) ? 4'b1111 : node7915;
														assign node7915 = (inp[9]) ? 4'b1110 : 4'b1111;
										assign node7919 = (inp[0]) ? node7941 : node7920;
											assign node7920 = (inp[10]) ? node7936 : node7921;
												assign node7921 = (inp[12]) ? node7927 : node7922;
													assign node7922 = (inp[4]) ? 4'b1011 : node7923;
														assign node7923 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node7927 = (inp[4]) ? node7933 : node7928;
														assign node7928 = (inp[2]) ? node7930 : 4'b1011;
															assign node7930 = (inp[11]) ? 4'b1010 : 4'b1010;
														assign node7933 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node7936 = (inp[4]) ? 4'b1111 : node7937;
													assign node7937 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node7941 = (inp[11]) ? node7949 : node7942;
												assign node7942 = (inp[9]) ? 4'b1011 : node7943;
													assign node7943 = (inp[2]) ? node7945 : 4'b1111;
														assign node7945 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node7949 = (inp[4]) ? node7955 : node7950;
													assign node7950 = (inp[12]) ? 4'b1011 : node7951;
														assign node7951 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node7955 = (inp[9]) ? node7957 : 4'b1011;
														assign node7957 = (inp[2]) ? 4'b1110 : 4'b1010;
									assign node7960 = (inp[1]) ? node7992 : node7961;
										assign node7961 = (inp[9]) ? node7979 : node7962;
											assign node7962 = (inp[11]) ? node7970 : node7963;
												assign node7963 = (inp[2]) ? 4'b1010 : node7964;
													assign node7964 = (inp[0]) ? 4'b1010 : node7965;
														assign node7965 = (inp[4]) ? 4'b1010 : 4'b1011;
												assign node7970 = (inp[0]) ? node7974 : node7971;
													assign node7971 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node7974 = (inp[4]) ? node7976 : 4'b1011;
														assign node7976 = (inp[12]) ? 4'b1010 : 4'b1011;
											assign node7979 = (inp[11]) ? node7981 : 4'b1011;
												assign node7981 = (inp[2]) ? node7987 : node7982;
													assign node7982 = (inp[0]) ? node7984 : 4'b1011;
														assign node7984 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node7987 = (inp[12]) ? 4'b1010 : node7988;
														assign node7988 = (inp[0]) ? 4'b1010 : 4'b1011;
										assign node7992 = (inp[10]) ? node8020 : node7993;
											assign node7993 = (inp[9]) ? node8009 : node7994;
												assign node7994 = (inp[11]) ? node8002 : node7995;
													assign node7995 = (inp[2]) ? 4'b1110 : node7996;
														assign node7996 = (inp[12]) ? node7998 : 4'b1010;
															assign node7998 = (inp[4]) ? 4'b1010 : 4'b1111;
													assign node8002 = (inp[12]) ? 4'b1110 : node8003;
														assign node8003 = (inp[0]) ? node8005 : 4'b1111;
															assign node8005 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node8009 = (inp[12]) ? node8013 : node8010;
													assign node8010 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node8013 = (inp[4]) ? node8017 : node8014;
														assign node8014 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node8017 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node8020 = (inp[11]) ? node8038 : node8021;
												assign node8021 = (inp[4]) ? node8031 : node8022;
													assign node8022 = (inp[12]) ? node8026 : node8023;
														assign node8023 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node8026 = (inp[2]) ? node8028 : 4'b1111;
															assign node8028 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node8031 = (inp[12]) ? 4'b1011 : node8032;
														assign node8032 = (inp[9]) ? node8034 : 4'b1111;
															assign node8034 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node8038 = (inp[0]) ? node8048 : node8039;
													assign node8039 = (inp[2]) ? node8041 : 4'b1111;
														assign node8041 = (inp[12]) ? node8045 : node8042;
															assign node8042 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node8045 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node8048 = (inp[9]) ? node8056 : node8049;
														assign node8049 = (inp[12]) ? node8053 : node8050;
															assign node8050 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node8053 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node8056 = (inp[2]) ? 4'b1110 : 4'b1010;
						assign node8059 = (inp[15]) ? node8487 : node8060;
							assign node8060 = (inp[4]) ? node8256 : node8061;
								assign node8061 = (inp[12]) ? node8151 : node8062;
									assign node8062 = (inp[11]) ? node8100 : node8063;
										assign node8063 = (inp[9]) ? node8081 : node8064;
											assign node8064 = (inp[5]) ? node8072 : node8065;
												assign node8065 = (inp[13]) ? 4'b1110 : node8066;
													assign node8066 = (inp[10]) ? node8068 : 4'b1010;
														assign node8068 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node8072 = (inp[13]) ? node8078 : node8073;
													assign node8073 = (inp[10]) ? node8075 : 4'b1111;
														assign node8075 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node8078 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node8081 = (inp[5]) ? node8091 : node8082;
												assign node8082 = (inp[13]) ? 4'b1111 : node8083;
													assign node8083 = (inp[1]) ? node8085 : 4'b1011;
														assign node8085 = (inp[0]) ? node8087 : 4'b1011;
															assign node8087 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node8091 = (inp[13]) ? node8097 : node8092;
													assign node8092 = (inp[0]) ? node8094 : 4'b1110;
														assign node8094 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node8097 = (inp[0]) ? 4'b1011 : 4'b1010;
										assign node8100 = (inp[9]) ? node8130 : node8101;
											assign node8101 = (inp[10]) ? node8115 : node8102;
												assign node8102 = (inp[5]) ? node8110 : node8103;
													assign node8103 = (inp[13]) ? 4'b1111 : node8104;
														assign node8104 = (inp[2]) ? node8106 : 4'b1011;
															assign node8106 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node8110 = (inp[2]) ? node8112 : 4'b1110;
														assign node8112 = (inp[13]) ? 4'b1011 : 4'b1111;
												assign node8115 = (inp[13]) ? node8121 : node8116;
													assign node8116 = (inp[2]) ? node8118 : 4'b1110;
														assign node8118 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node8121 = (inp[5]) ? node8125 : node8122;
														assign node8122 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node8125 = (inp[2]) ? 4'b1011 : node8126;
															assign node8126 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node8130 = (inp[13]) ? node8140 : node8131;
												assign node8131 = (inp[5]) ? node8135 : node8132;
													assign node8132 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node8135 = (inp[0]) ? node8137 : 4'b1111;
														assign node8137 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node8140 = (inp[5]) ? node8146 : node8141;
													assign node8141 = (inp[2]) ? node8143 : 4'b1110;
														assign node8143 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node8146 = (inp[0]) ? 4'b1010 : node8147;
														assign node8147 = (inp[2]) ? 4'b1010 : 4'b1011;
									assign node8151 = (inp[11]) ? node8203 : node8152;
										assign node8152 = (inp[2]) ? node8174 : node8153;
											assign node8153 = (inp[9]) ? node8169 : node8154;
												assign node8154 = (inp[1]) ? node8164 : node8155;
													assign node8155 = (inp[5]) ? node8161 : node8156;
														assign node8156 = (inp[0]) ? node8158 : 4'b1110;
															assign node8158 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node8161 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node8164 = (inp[5]) ? 4'b1111 : node8165;
														assign node8165 = (inp[13]) ? 4'b1010 : 4'b1110;
												assign node8169 = (inp[0]) ? node8171 : 4'b1110;
													assign node8171 = (inp[13]) ? 4'b1110 : 4'b1010;
											assign node8174 = (inp[1]) ? node8192 : node8175;
												assign node8175 = (inp[0]) ? node8185 : node8176;
													assign node8176 = (inp[10]) ? node8178 : 4'b1011;
														assign node8178 = (inp[9]) ? node8182 : node8179;
															assign node8179 = (inp[5]) ? 4'b1010 : 4'b1111;
															assign node8182 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node8185 = (inp[9]) ? node8187 : 4'b1110;
														assign node8187 = (inp[13]) ? node8189 : 4'b1010;
															assign node8189 = (inp[5]) ? 4'b1010 : 4'b1110;
												assign node8192 = (inp[5]) ? node8196 : node8193;
													assign node8193 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node8196 = (inp[13]) ? node8198 : 4'b1010;
														assign node8198 = (inp[0]) ? node8200 : 4'b1111;
															assign node8200 = (inp[9]) ? 4'b1111 : 4'b1110;
										assign node8203 = (inp[13]) ? node8235 : node8204;
											assign node8204 = (inp[0]) ? node8220 : node8205;
												assign node8205 = (inp[10]) ? node8211 : node8206;
													assign node8206 = (inp[1]) ? 4'b1110 : node8207;
														assign node8207 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node8211 = (inp[9]) ? 4'b1110 : node8212;
														assign node8212 = (inp[2]) ? node8216 : node8213;
															assign node8213 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node8216 = (inp[1]) ? 4'b1111 : 4'b1010;
												assign node8220 = (inp[5]) ? node8226 : node8221;
													assign node8221 = (inp[1]) ? 4'b1110 : node8222;
														assign node8222 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node8226 = (inp[1]) ? node8228 : 4'b1111;
														assign node8228 = (inp[10]) ? node8232 : node8229;
															assign node8229 = (inp[9]) ? 4'b1010 : 4'b1010;
															assign node8232 = (inp[2]) ? 4'b1010 : 4'b1010;
											assign node8235 = (inp[1]) ? node8245 : node8236;
												assign node8236 = (inp[5]) ? node8240 : node8237;
													assign node8237 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node8240 = (inp[10]) ? 4'b1011 : node8241;
														assign node8241 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node8245 = (inp[5]) ? node8253 : node8246;
													assign node8246 = (inp[9]) ? node8248 : 4'b1011;
														assign node8248 = (inp[0]) ? node8250 : 4'b1010;
															assign node8250 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node8253 = (inp[10]) ? 4'b1111 : 4'b1110;
								assign node8256 = (inp[0]) ? node8376 : node8257;
									assign node8257 = (inp[10]) ? node8325 : node8258;
										assign node8258 = (inp[9]) ? node8294 : node8259;
											assign node8259 = (inp[12]) ? node8271 : node8260;
												assign node8260 = (inp[13]) ? node8264 : node8261;
													assign node8261 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node8264 = (inp[5]) ? node8268 : node8265;
														assign node8265 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node8268 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node8271 = (inp[13]) ? node8283 : node8272;
													assign node8272 = (inp[1]) ? node8280 : node8273;
														assign node8273 = (inp[11]) ? node8277 : node8274;
															assign node8274 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node8277 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node8280 = (inp[5]) ? 4'b1110 : 4'b1010;
													assign node8283 = (inp[5]) ? node8289 : node8284;
														assign node8284 = (inp[1]) ? 4'b1111 : node8285;
															assign node8285 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node8289 = (inp[11]) ? node8291 : 4'b1010;
															assign node8291 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node8294 = (inp[11]) ? node8314 : node8295;
												assign node8295 = (inp[12]) ? node8301 : node8296;
													assign node8296 = (inp[5]) ? node8298 : 4'b1111;
														assign node8298 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node8301 = (inp[1]) ? node8309 : node8302;
														assign node8302 = (inp[13]) ? node8306 : node8303;
															assign node8303 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node8306 = (inp[5]) ? 4'b1111 : 4'b1010;
														assign node8309 = (inp[13]) ? 4'b1011 : node8310;
															assign node8310 = (inp[2]) ? 4'b1010 : 4'b1110;
												assign node8314 = (inp[13]) ? node8320 : node8315;
													assign node8315 = (inp[5]) ? 4'b1111 : node8316;
														assign node8316 = (inp[1]) ? 4'b1011 : 4'b1110;
													assign node8320 = (inp[12]) ? 4'b1110 : node8321;
														assign node8321 = (inp[5]) ? 4'b1010 : 4'b1110;
										assign node8325 = (inp[9]) ? node8347 : node8326;
											assign node8326 = (inp[13]) ? node8338 : node8327;
												assign node8327 = (inp[12]) ? node8331 : node8328;
													assign node8328 = (inp[11]) ? 4'b1011 : 4'b1111;
													assign node8331 = (inp[11]) ? 4'b1110 : node8332;
														assign node8332 = (inp[1]) ? 4'b1011 : node8333;
															assign node8333 = (inp[5]) ? 4'b1010 : 4'b1110;
												assign node8338 = (inp[5]) ? node8340 : 4'b1110;
													assign node8340 = (inp[12]) ? 4'b1011 : node8341;
														assign node8341 = (inp[1]) ? 4'b1010 : node8342;
															assign node8342 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node8347 = (inp[12]) ? node8365 : node8348;
												assign node8348 = (inp[11]) ? node8356 : node8349;
													assign node8349 = (inp[2]) ? node8351 : 4'b1011;
														assign node8351 = (inp[13]) ? 4'b1010 : node8352;
															assign node8352 = (inp[5]) ? 4'b1110 : 4'b1010;
													assign node8356 = (inp[13]) ? node8362 : node8357;
														assign node8357 = (inp[5]) ? 4'b1111 : node8358;
															assign node8358 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node8362 = (inp[5]) ? 4'b1010 : 4'b1110;
												assign node8365 = (inp[1]) ? node8369 : node8366;
													assign node8366 = (inp[13]) ? 4'b1111 : 4'b1011;
													assign node8369 = (inp[2]) ? node8373 : node8370;
														assign node8370 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node8373 = (inp[11]) ? 4'b1011 : 4'b1010;
									assign node8376 = (inp[5]) ? node8430 : node8377;
										assign node8377 = (inp[13]) ? node8407 : node8378;
											assign node8378 = (inp[1]) ? node8392 : node8379;
												assign node8379 = (inp[12]) ? node8385 : node8380;
													assign node8380 = (inp[9]) ? 4'b1010 : node8381;
														assign node8381 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node8385 = (inp[10]) ? node8387 : 4'b1110;
														assign node8387 = (inp[11]) ? 4'b1111 : node8388;
															assign node8388 = (inp[2]) ? 4'b1110 : 4'b1110;
												assign node8392 = (inp[12]) ? node8400 : node8393;
													assign node8393 = (inp[10]) ? node8395 : 4'b1011;
														assign node8395 = (inp[2]) ? node8397 : 4'b1010;
															assign node8397 = (inp[9]) ? 4'b1010 : 4'b1010;
													assign node8400 = (inp[2]) ? node8402 : 4'b1011;
														assign node8402 = (inp[11]) ? node8404 : 4'b1011;
															assign node8404 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node8407 = (inp[1]) ? node8417 : node8408;
												assign node8408 = (inp[12]) ? node8414 : node8409;
													assign node8409 = (inp[11]) ? node8411 : 4'b1111;
														assign node8411 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node8414 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node8417 = (inp[2]) ? node8419 : 4'b1111;
													assign node8419 = (inp[12]) ? node8425 : node8420;
														assign node8420 = (inp[11]) ? node8422 : 4'b1111;
															assign node8422 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node8425 = (inp[11]) ? 4'b1111 : node8426;
															assign node8426 = (inp[9]) ? 4'b1111 : 4'b1110;
										assign node8430 = (inp[13]) ? node8464 : node8431;
											assign node8431 = (inp[1]) ? node8445 : node8432;
												assign node8432 = (inp[12]) ? node8440 : node8433;
													assign node8433 = (inp[11]) ? 4'b1110 : node8434;
														assign node8434 = (inp[9]) ? node8436 : 4'b1111;
															assign node8436 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node8440 = (inp[11]) ? 4'b1011 : node8441;
														assign node8441 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node8445 = (inp[9]) ? node8457 : node8446;
													assign node8446 = (inp[10]) ? node8452 : node8447;
														assign node8447 = (inp[2]) ? node8449 : 4'b1110;
															assign node8449 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node8452 = (inp[12]) ? node8454 : 4'b1110;
															assign node8454 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node8457 = (inp[2]) ? node8461 : node8458;
														assign node8458 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node8461 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node8464 = (inp[1]) ? node8482 : node8465;
												assign node8465 = (inp[12]) ? node8471 : node8466;
													assign node8466 = (inp[2]) ? node8468 : 4'b1011;
														assign node8468 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node8471 = (inp[11]) ? node8477 : node8472;
														assign node8472 = (inp[2]) ? node8474 : 4'b1110;
															assign node8474 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node8477 = (inp[2]) ? node8479 : 4'b1111;
															assign node8479 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node8482 = (inp[11]) ? node8484 : 4'b1011;
													assign node8484 = (inp[9]) ? 4'b1010 : 4'b1011;
							assign node8487 = (inp[5]) ? node8655 : node8488;
								assign node8488 = (inp[13]) ? node8572 : node8489;
									assign node8489 = (inp[1]) ? node8535 : node8490;
										assign node8490 = (inp[4]) ? node8520 : node8491;
											assign node8491 = (inp[12]) ? node8503 : node8492;
												assign node8492 = (inp[11]) ? node8498 : node8493;
													assign node8493 = (inp[9]) ? 4'b1101 : node8494;
														assign node8494 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node8498 = (inp[9]) ? 4'b1100 : node8499;
														assign node8499 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node8503 = (inp[0]) ? node8509 : node8504;
													assign node8504 = (inp[11]) ? 4'b1001 : node8505;
														assign node8505 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node8509 = (inp[9]) ? node8515 : node8510;
														assign node8510 = (inp[10]) ? 4'b1001 : node8511;
															assign node8511 = (inp[11]) ? 4'b1000 : 4'b1000;
														assign node8515 = (inp[10]) ? 4'b1000 : node8516;
															assign node8516 = (inp[11]) ? 4'b1000 : 4'b1000;
											assign node8520 = (inp[12]) ? node8526 : node8521;
												assign node8521 = (inp[11]) ? node8523 : 4'b1001;
													assign node8523 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node8526 = (inp[10]) ? node8528 : 4'b1101;
													assign node8528 = (inp[2]) ? node8530 : 4'b1100;
														assign node8530 = (inp[0]) ? 4'b1101 : node8531;
															assign node8531 = (inp[9]) ? 4'b1101 : 4'b1100;
										assign node8535 = (inp[0]) ? node8555 : node8536;
											assign node8536 = (inp[2]) ? node8546 : node8537;
												assign node8537 = (inp[11]) ? node8543 : node8538;
													assign node8538 = (inp[10]) ? 4'b1000 : node8539;
														assign node8539 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node8543 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node8546 = (inp[11]) ? node8548 : 4'b1000;
													assign node8548 = (inp[4]) ? node8552 : node8549;
														assign node8549 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node8552 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node8555 = (inp[2]) ? node8563 : node8556;
												assign node8556 = (inp[11]) ? node8560 : node8557;
													assign node8557 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node8560 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node8563 = (inp[10]) ? node8567 : node8564;
													assign node8564 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node8567 = (inp[9]) ? node8569 : 4'b1001;
														assign node8569 = (inp[11]) ? 4'b1001 : 4'b1000;
									assign node8572 = (inp[1]) ? node8610 : node8573;
										assign node8573 = (inp[11]) ? node8597 : node8574;
											assign node8574 = (inp[9]) ? node8586 : node8575;
												assign node8575 = (inp[4]) ? node8579 : node8576;
													assign node8576 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node8579 = (inp[12]) ? 4'b1001 : node8580;
														assign node8580 = (inp[0]) ? node8582 : 4'b1101;
															assign node8582 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node8586 = (inp[12]) ? node8592 : node8587;
													assign node8587 = (inp[4]) ? 4'b1100 : node8588;
														assign node8588 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node8592 = (inp[4]) ? 4'b1001 : node8593;
														assign node8593 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node8597 = (inp[0]) ? node8605 : node8598;
												assign node8598 = (inp[9]) ? node8600 : 4'b1101;
													assign node8600 = (inp[2]) ? 4'b1000 : node8601;
														assign node8601 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node8605 = (inp[9]) ? 4'b1000 : node8606;
													assign node8606 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node8610 = (inp[11]) ? node8632 : node8611;
											assign node8611 = (inp[9]) ? node8623 : node8612;
												assign node8612 = (inp[2]) ? node8614 : 4'b1100;
													assign node8614 = (inp[10]) ? node8616 : 4'b1101;
														assign node8616 = (inp[0]) ? node8620 : node8617;
															assign node8617 = (inp[4]) ? 4'b1101 : 4'b1100;
															assign node8620 = (inp[4]) ? 4'b1100 : 4'b1101;
												assign node8623 = (inp[2]) ? node8625 : 4'b1101;
													assign node8625 = (inp[0]) ? node8629 : node8626;
														assign node8626 = (inp[4]) ? 4'b1100 : 4'b1101;
														assign node8629 = (inp[4]) ? 4'b1101 : 4'b1100;
											assign node8632 = (inp[9]) ? node8644 : node8633;
												assign node8633 = (inp[2]) ? node8635 : 4'b1101;
													assign node8635 = (inp[10]) ? node8641 : node8636;
														assign node8636 = (inp[12]) ? 4'b1101 : node8637;
															assign node8637 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node8641 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node8644 = (inp[12]) ? node8646 : 4'b1101;
													assign node8646 = (inp[0]) ? 4'b1100 : node8647;
														assign node8647 = (inp[2]) ? node8651 : node8648;
															assign node8648 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node8651 = (inp[4]) ? 4'b1101 : 4'b1100;
								assign node8655 = (inp[13]) ? node8749 : node8656;
									assign node8656 = (inp[1]) ? node8712 : node8657;
										assign node8657 = (inp[12]) ? node8687 : node8658;
											assign node8658 = (inp[4]) ? node8678 : node8659;
												assign node8659 = (inp[10]) ? node8669 : node8660;
													assign node8660 = (inp[9]) ? node8666 : node8661;
														assign node8661 = (inp[11]) ? 4'b1001 : node8662;
															assign node8662 = (inp[2]) ? 4'b1000 : 4'b1000;
														assign node8666 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node8669 = (inp[11]) ? node8673 : node8670;
														assign node8670 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node8673 = (inp[9]) ? node8675 : 4'b1001;
															assign node8675 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node8678 = (inp[11]) ? 4'b1101 : node8679;
													assign node8679 = (inp[10]) ? 4'b1100 : node8680;
														assign node8680 = (inp[2]) ? node8682 : 4'b1100;
															assign node8682 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node8687 = (inp[4]) ? node8703 : node8688;
												assign node8688 = (inp[0]) ? node8694 : node8689;
													assign node8689 = (inp[11]) ? node8691 : 4'b1101;
														assign node8691 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node8694 = (inp[2]) ? node8696 : 4'b1100;
														assign node8696 = (inp[10]) ? node8700 : node8697;
															assign node8697 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node8700 = (inp[11]) ? 4'b1100 : 4'b1100;
												assign node8703 = (inp[2]) ? node8705 : 4'b1000;
													assign node8705 = (inp[11]) ? 4'b1001 : node8706;
														assign node8706 = (inp[0]) ? 4'b1000 : node8707;
															assign node8707 = (inp[9]) ? 4'b1001 : 4'b1000;
										assign node8712 = (inp[9]) ? node8730 : node8713;
											assign node8713 = (inp[11]) ? node8719 : node8714;
												assign node8714 = (inp[2]) ? 4'b1100 : node8715;
													assign node8715 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node8719 = (inp[0]) ? node8721 : 4'b1101;
													assign node8721 = (inp[12]) ? 4'b1101 : node8722;
														assign node8722 = (inp[4]) ? node8726 : node8723;
															assign node8723 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node8726 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node8730 = (inp[11]) ? node8742 : node8731;
												assign node8731 = (inp[2]) ? 4'b1101 : node8732;
													assign node8732 = (inp[10]) ? node8734 : 4'b1101;
														assign node8734 = (inp[12]) ? node8738 : node8735;
															assign node8735 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node8738 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node8742 = (inp[10]) ? node8744 : 4'b1100;
													assign node8744 = (inp[0]) ? 4'b1100 : node8745;
														assign node8745 = (inp[2]) ? 4'b1100 : 4'b1101;
									assign node8749 = (inp[1]) ? node8823 : node8750;
										assign node8750 = (inp[0]) ? node8786 : node8751;
											assign node8751 = (inp[2]) ? node8765 : node8752;
												assign node8752 = (inp[9]) ? node8760 : node8753;
													assign node8753 = (inp[11]) ? 4'b1000 : node8754;
														assign node8754 = (inp[4]) ? 4'b1001 : node8755;
															assign node8755 = (inp[12]) ? 4'b1001 : 4'b1100;
													assign node8760 = (inp[12]) ? node8762 : 4'b1001;
														assign node8762 = (inp[4]) ? 4'b1100 : 4'b1001;
												assign node8765 = (inp[10]) ? node8777 : node8766;
													assign node8766 = (inp[9]) ? node8772 : node8767;
														assign node8767 = (inp[4]) ? node8769 : 4'b1000;
															assign node8769 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node8772 = (inp[12]) ? node8774 : 4'b1100;
															assign node8774 = (inp[4]) ? 4'b1100 : 4'b1001;
													assign node8777 = (inp[11]) ? node8781 : node8778;
														assign node8778 = (inp[4]) ? 4'b1100 : 4'b1001;
														assign node8781 = (inp[12]) ? 4'b1000 : node8782;
															assign node8782 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node8786 = (inp[12]) ? node8806 : node8787;
												assign node8787 = (inp[4]) ? node8797 : node8788;
													assign node8788 = (inp[2]) ? node8794 : node8789;
														assign node8789 = (inp[11]) ? node8791 : 4'b1100;
															assign node8791 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node8794 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node8797 = (inp[2]) ? node8799 : 4'b1001;
														assign node8799 = (inp[11]) ? node8803 : node8800;
															assign node8800 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node8803 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node8806 = (inp[4]) ? node8814 : node8807;
													assign node8807 = (inp[10]) ? node8809 : 4'b1000;
														assign node8809 = (inp[11]) ? 4'b1001 : node8810;
															assign node8810 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node8814 = (inp[2]) ? node8816 : 4'b1100;
														assign node8816 = (inp[11]) ? node8820 : node8817;
															assign node8817 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node8820 = (inp[9]) ? 4'b1100 : 4'b1101;
										assign node8823 = (inp[9]) ? node8847 : node8824;
											assign node8824 = (inp[0]) ? node8840 : node8825;
												assign node8825 = (inp[2]) ? node8835 : node8826;
													assign node8826 = (inp[12]) ? 4'b1000 : node8827;
														assign node8827 = (inp[11]) ? node8831 : node8828;
															assign node8828 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node8831 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node8835 = (inp[11]) ? node8837 : 4'b1001;
														assign node8837 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node8840 = (inp[11]) ? node8842 : 4'b1000;
													assign node8842 = (inp[12]) ? node8844 : 4'b1001;
														assign node8844 = (inp[4]) ? 4'b1001 : 4'b1000;
											assign node8847 = (inp[11]) ? node8859 : node8848;
												assign node8848 = (inp[0]) ? 4'b1001 : node8849;
													assign node8849 = (inp[2]) ? node8853 : node8850;
														assign node8850 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node8853 = (inp[12]) ? 4'b1000 : node8854;
															assign node8854 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node8859 = (inp[12]) ? node8861 : 4'b1000;
													assign node8861 = (inp[10]) ? 4'b1001 : node8862;
														assign node8862 = (inp[2]) ? 4'b1000 : 4'b1001;
					assign node8866 = (inp[0]) ? node9748 : node8867;
						assign node8867 = (inp[11]) ? node9307 : node8868;
							assign node8868 = (inp[9]) ? node9084 : node8869;
								assign node8869 = (inp[4]) ? node8973 : node8870;
									assign node8870 = (inp[15]) ? node8922 : node8871;
										assign node8871 = (inp[13]) ? node8891 : node8872;
											assign node8872 = (inp[1]) ? node8880 : node8873;
												assign node8873 = (inp[5]) ? node8875 : 4'b0000;
													assign node8875 = (inp[12]) ? node8877 : 4'b0101;
														assign node8877 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node8880 = (inp[2]) ? node8882 : 4'b0101;
													assign node8882 = (inp[10]) ? node8886 : node8883;
														assign node8883 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node8886 = (inp[12]) ? 4'b0000 : node8887;
															assign node8887 = (inp[5]) ? 4'b0000 : 4'b0100;
											assign node8891 = (inp[2]) ? node8913 : node8892;
												assign node8892 = (inp[5]) ? node8902 : node8893;
													assign node8893 = (inp[10]) ? node8897 : node8894;
														assign node8894 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node8897 = (inp[1]) ? node8899 : 4'b0000;
															assign node8899 = (inp[7]) ? 4'b0000 : 4'b0101;
													assign node8902 = (inp[1]) ? node8908 : node8903;
														assign node8903 = (inp[7]) ? node8905 : 4'b0100;
															assign node8905 = (inp[12]) ? 4'b0000 : 4'b0101;
														assign node8908 = (inp[10]) ? node8910 : 4'b0000;
															assign node8910 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node8913 = (inp[1]) ? node8917 : node8914;
													assign node8914 = (inp[5]) ? 4'b0101 : 4'b0001;
													assign node8917 = (inp[12]) ? 4'b0000 : node8918;
														assign node8918 = (inp[5]) ? 4'b0001 : 4'b0101;
										assign node8922 = (inp[5]) ? node8946 : node8923;
											assign node8923 = (inp[1]) ? node8935 : node8924;
												assign node8924 = (inp[12]) ? node8928 : node8925;
													assign node8925 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node8928 = (inp[13]) ? node8930 : 4'b0011;
														assign node8930 = (inp[7]) ? 4'b0010 : node8931;
															assign node8931 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node8935 = (inp[13]) ? node8939 : node8936;
													assign node8936 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node8939 = (inp[2]) ? 4'b0011 : node8940;
														assign node8940 = (inp[7]) ? node8942 : 4'b0110;
															assign node8942 = (inp[12]) ? 4'b0110 : 4'b0010;
											assign node8946 = (inp[2]) ? node8962 : node8947;
												assign node8947 = (inp[13]) ? node8957 : node8948;
													assign node8948 = (inp[12]) ? node8954 : node8949;
														assign node8949 = (inp[1]) ? 4'b0110 : node8950;
															assign node8950 = (inp[7]) ? 4'b0011 : 4'b0110;
														assign node8954 = (inp[1]) ? 4'b0010 : 4'b0110;
													assign node8957 = (inp[12]) ? 4'b0011 : node8958;
														assign node8958 = (inp[7]) ? 4'b0011 : 4'b0111;
												assign node8962 = (inp[12]) ? node8970 : node8963;
													assign node8963 = (inp[13]) ? node8965 : 4'b0110;
														assign node8965 = (inp[1]) ? node8967 : 4'b0011;
															assign node8967 = (inp[7]) ? 4'b0110 : 4'b0011;
													assign node8970 = (inp[1]) ? 4'b0010 : 4'b0110;
									assign node8973 = (inp[15]) ? node9031 : node8974;
										assign node8974 = (inp[2]) ? node9004 : node8975;
											assign node8975 = (inp[5]) ? node8991 : node8976;
												assign node8976 = (inp[1]) ? node8984 : node8977;
													assign node8977 = (inp[7]) ? node8981 : node8978;
														assign node8978 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node8981 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node8984 = (inp[7]) ? 4'b0110 : node8985;
														assign node8985 = (inp[12]) ? node8987 : 4'b0110;
															assign node8987 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node8991 = (inp[7]) ? node8997 : node8992;
													assign node8992 = (inp[1]) ? node8994 : 4'b0011;
														assign node8994 = (inp[12]) ? 4'b0110 : 4'b0011;
													assign node8997 = (inp[1]) ? 4'b0010 : node8998;
														assign node8998 = (inp[10]) ? node9000 : 4'b0110;
															assign node9000 = (inp[12]) ? 4'b0110 : 4'b0111;
											assign node9004 = (inp[13]) ? node9016 : node9005;
												assign node9005 = (inp[10]) ? node9007 : 4'b0111;
													assign node9007 = (inp[7]) ? node9011 : node9008;
														assign node9008 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node9011 = (inp[12]) ? 4'b0011 : node9012;
															assign node9012 = (inp[5]) ? 4'b0111 : 4'b0011;
												assign node9016 = (inp[1]) ? node9022 : node9017;
													assign node9017 = (inp[7]) ? node9019 : 4'b0110;
														assign node9019 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node9022 = (inp[5]) ? node9028 : node9023;
														assign node9023 = (inp[12]) ? node9025 : 4'b0110;
															assign node9025 = (inp[10]) ? 4'b0110 : 4'b0011;
														assign node9028 = (inp[7]) ? 4'b0010 : 4'b0011;
										assign node9031 = (inp[7]) ? node9063 : node9032;
											assign node9032 = (inp[5]) ? node9050 : node9033;
												assign node9033 = (inp[13]) ? node9039 : node9034;
													assign node9034 = (inp[2]) ? node9036 : 4'b0100;
														assign node9036 = (inp[10]) ? 4'b0101 : 4'b0000;
													assign node9039 = (inp[2]) ? node9045 : node9040;
														assign node9040 = (inp[12]) ? node9042 : 4'b0000;
															assign node9042 = (inp[1]) ? 4'b0101 : 4'b0000;
														assign node9045 = (inp[12]) ? node9047 : 4'b0101;
															assign node9047 = (inp[1]) ? 4'b0101 : 4'b0001;
												assign node9050 = (inp[2]) ? node9054 : node9051;
													assign node9051 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node9054 = (inp[13]) ? node9056 : 4'b0100;
														assign node9056 = (inp[12]) ? node9060 : node9057;
															assign node9057 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node9060 = (inp[1]) ? 4'b0000 : 4'b0100;
											assign node9063 = (inp[13]) ? node9075 : node9064;
												assign node9064 = (inp[10]) ? 4'b0101 : node9065;
													assign node9065 = (inp[12]) ? 4'b0001 : node9066;
														assign node9066 = (inp[2]) ? node9070 : node9067;
															assign node9067 = (inp[5]) ? 4'b0001 : 4'b0101;
															assign node9070 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node9075 = (inp[1]) ? node9081 : node9076;
													assign node9076 = (inp[5]) ? node9078 : 4'b0000;
														assign node9078 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node9081 = (inp[5]) ? 4'b0000 : 4'b0100;
								assign node9084 = (inp[10]) ? node9198 : node9085;
									assign node9085 = (inp[15]) ? node9135 : node9086;
										assign node9086 = (inp[4]) ? node9114 : node9087;
											assign node9087 = (inp[2]) ? node9099 : node9088;
												assign node9088 = (inp[5]) ? node9096 : node9089;
													assign node9089 = (inp[13]) ? node9091 : 4'b0100;
														assign node9091 = (inp[12]) ? 4'b0000 : node9092;
															assign node9092 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node9096 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node9099 = (inp[12]) ? node9103 : node9100;
													assign node9100 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node9103 = (inp[5]) ? node9107 : node9104;
														assign node9104 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node9107 = (inp[1]) ? node9111 : node9108;
															assign node9108 = (inp[13]) ? 4'b0101 : 4'b0000;
															assign node9111 = (inp[7]) ? 4'b0100 : 4'b0000;
											assign node9114 = (inp[5]) ? node9122 : node9115;
												assign node9115 = (inp[1]) ? 4'b0110 : node9116;
													assign node9116 = (inp[12]) ? node9118 : 4'b0010;
														assign node9118 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node9122 = (inp[7]) ? node9130 : node9123;
													assign node9123 = (inp[2]) ? node9125 : 4'b0011;
														assign node9125 = (inp[13]) ? node9127 : 4'b0010;
															assign node9127 = (inp[1]) ? 4'b0010 : 4'b0110;
													assign node9130 = (inp[12]) ? 4'b0110 : node9131;
														assign node9131 = (inp[2]) ? 4'b0111 : 4'b0110;
										assign node9135 = (inp[4]) ? node9159 : node9136;
											assign node9136 = (inp[13]) ? node9144 : node9137;
												assign node9137 = (inp[1]) ? node9141 : node9138;
													assign node9138 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node9141 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node9144 = (inp[2]) ? node9152 : node9145;
													assign node9145 = (inp[5]) ? node9149 : node9146;
														assign node9146 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node9149 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node9152 = (inp[7]) ? 4'b0110 : node9153;
														assign node9153 = (inp[1]) ? 4'b0011 : node9154;
															assign node9154 = (inp[5]) ? 4'b0110 : 4'b0010;
											assign node9159 = (inp[7]) ? node9183 : node9160;
												assign node9160 = (inp[12]) ? node9172 : node9161;
													assign node9161 = (inp[2]) ? node9167 : node9162;
														assign node9162 = (inp[13]) ? 4'b0101 : node9163;
															assign node9163 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node9167 = (inp[1]) ? node9169 : 4'b0101;
															assign node9169 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node9172 = (inp[13]) ? node9178 : node9173;
														assign node9173 = (inp[5]) ? node9175 : 4'b0100;
															assign node9175 = (inp[1]) ? 4'b0001 : 4'b0100;
														assign node9178 = (inp[5]) ? 4'b0000 : node9179;
															assign node9179 = (inp[1]) ? 4'b0101 : 4'b0000;
												assign node9183 = (inp[12]) ? node9189 : node9184;
													assign node9184 = (inp[5]) ? 4'b0001 : node9185;
														assign node9185 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node9189 = (inp[2]) ? node9193 : node9190;
														assign node9190 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node9193 = (inp[13]) ? 4'b0000 : node9194;
															assign node9194 = (inp[1]) ? 4'b0000 : 4'b0100;
									assign node9198 = (inp[4]) ? node9258 : node9199;
										assign node9199 = (inp[15]) ? node9225 : node9200;
											assign node9200 = (inp[2]) ? node9214 : node9201;
												assign node9201 = (inp[12]) ? node9205 : node9202;
													assign node9202 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node9205 = (inp[13]) ? 4'b0000 : node9206;
														assign node9206 = (inp[7]) ? node9210 : node9207;
															assign node9207 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node9210 = (inp[5]) ? 4'b0000 : 4'b0100;
												assign node9214 = (inp[7]) ? node9216 : 4'b0101;
													assign node9216 = (inp[12]) ? node9222 : node9217;
														assign node9217 = (inp[13]) ? node9219 : 4'b0101;
															assign node9219 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node9222 = (inp[5]) ? 4'b0101 : 4'b0000;
											assign node9225 = (inp[13]) ? node9239 : node9226;
												assign node9226 = (inp[12]) ? node9228 : 4'b0110;
													assign node9228 = (inp[5]) ? node9236 : node9229;
														assign node9229 = (inp[1]) ? node9233 : node9230;
															assign node9230 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node9233 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node9236 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node9239 = (inp[2]) ? node9247 : node9240;
													assign node9240 = (inp[7]) ? 4'b0111 : node9241;
														assign node9241 = (inp[1]) ? node9243 : 4'b0111;
															assign node9243 = (inp[5]) ? 4'b0011 : 4'b0111;
													assign node9247 = (inp[1]) ? node9253 : node9248;
														assign node9248 = (inp[12]) ? 4'b0110 : node9249;
															assign node9249 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node9253 = (inp[12]) ? node9255 : 4'b0110;
															assign node9255 = (inp[7]) ? 4'b0110 : 4'b0111;
										assign node9258 = (inp[15]) ? node9280 : node9259;
											assign node9259 = (inp[2]) ? node9265 : node9260;
												assign node9260 = (inp[5]) ? 4'b0010 : node9261;
													assign node9261 = (inp[1]) ? 4'b0110 : 4'b0010;
												assign node9265 = (inp[7]) ? node9273 : node9266;
													assign node9266 = (inp[12]) ? 4'b0011 : node9267;
														assign node9267 = (inp[5]) ? node9269 : 4'b0110;
															assign node9269 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node9273 = (inp[1]) ? 4'b0111 : node9274;
														assign node9274 = (inp[5]) ? node9276 : 4'b0010;
															assign node9276 = (inp[12]) ? 4'b0110 : 4'b0111;
											assign node9280 = (inp[2]) ? node9296 : node9281;
												assign node9281 = (inp[5]) ? node9293 : node9282;
													assign node9282 = (inp[13]) ? node9290 : node9283;
														assign node9283 = (inp[1]) ? node9287 : node9284;
															assign node9284 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node9287 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node9290 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node9293 = (inp[7]) ? 4'b0100 : 4'b0000;
												assign node9296 = (inp[12]) ? node9302 : node9297;
													assign node9297 = (inp[7]) ? 4'b0100 : node9298;
														assign node9298 = (inp[5]) ? 4'b0100 : 4'b0000;
													assign node9302 = (inp[5]) ? node9304 : 4'b0000;
														assign node9304 = (inp[13]) ? 4'b0000 : 4'b0100;
							assign node9307 = (inp[9]) ? node9525 : node9308;
								assign node9308 = (inp[15]) ? node9416 : node9309;
									assign node9309 = (inp[4]) ? node9365 : node9310;
										assign node9310 = (inp[13]) ? node9332 : node9311;
											assign node9311 = (inp[5]) ? node9321 : node9312;
												assign node9312 = (inp[12]) ? node9316 : node9313;
													assign node9313 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node9316 = (inp[10]) ? node9318 : 4'b0100;
														assign node9318 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node9321 = (inp[1]) ? node9327 : node9322;
													assign node9322 = (inp[12]) ? node9324 : 4'b0100;
														assign node9324 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node9327 = (inp[7]) ? node9329 : 4'b0000;
														assign node9329 = (inp[12]) ? 4'b0100 : 4'b0000;
											assign node9332 = (inp[2]) ? node9344 : node9333;
												assign node9333 = (inp[1]) ? node9339 : node9334;
													assign node9334 = (inp[7]) ? node9336 : 4'b0101;
														assign node9336 = (inp[12]) ? 4'b0001 : 4'b0100;
													assign node9339 = (inp[12]) ? 4'b0100 : node9340;
														assign node9340 = (inp[5]) ? 4'b0000 : 4'b0101;
												assign node9344 = (inp[5]) ? node9356 : node9345;
													assign node9345 = (inp[7]) ? node9349 : node9346;
														assign node9346 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node9349 = (inp[10]) ? node9353 : node9350;
															assign node9350 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node9353 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node9356 = (inp[1]) ? node9360 : node9357;
														assign node9357 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node9360 = (inp[7]) ? node9362 : 4'b0000;
															assign node9362 = (inp[12]) ? 4'b0101 : 4'b0001;
										assign node9365 = (inp[13]) ? node9391 : node9366;
											assign node9366 = (inp[5]) ? node9380 : node9367;
												assign node9367 = (inp[2]) ? node9373 : node9368;
													assign node9368 = (inp[12]) ? 4'b0010 : node9369;
														assign node9369 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node9373 = (inp[10]) ? node9375 : 4'b0110;
														assign node9375 = (inp[12]) ? node9377 : 4'b0010;
															assign node9377 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node9380 = (inp[1]) ? node9386 : node9381;
													assign node9381 = (inp[12]) ? 4'b0111 : node9382;
														assign node9382 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node9386 = (inp[7]) ? node9388 : 4'b0011;
														assign node9388 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node9391 = (inp[1]) ? node9409 : node9392;
												assign node9392 = (inp[5]) ? node9398 : node9393;
													assign node9393 = (inp[7]) ? node9395 : 4'b0111;
														assign node9395 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node9398 = (inp[7]) ? node9402 : node9399;
														assign node9399 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node9402 = (inp[2]) ? node9406 : node9403;
															assign node9403 = (inp[12]) ? 4'b0110 : 4'b0111;
															assign node9406 = (inp[12]) ? 4'b0111 : 4'b0110;
												assign node9409 = (inp[5]) ? node9411 : 4'b0111;
													assign node9411 = (inp[7]) ? 4'b0011 : node9412;
														assign node9412 = (inp[12]) ? 4'b0111 : 4'b0010;
									assign node9416 = (inp[4]) ? node9470 : node9417;
										assign node9417 = (inp[13]) ? node9439 : node9418;
											assign node9418 = (inp[1]) ? node9430 : node9419;
												assign node9419 = (inp[7]) ? node9423 : node9420;
													assign node9420 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node9423 = (inp[12]) ? 4'b0010 : node9424;
														assign node9424 = (inp[5]) ? node9426 : 4'b0111;
															assign node9426 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node9430 = (inp[5]) ? node9436 : node9431;
													assign node9431 = (inp[7]) ? node9433 : 4'b0111;
														assign node9433 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node9436 = (inp[12]) ? 4'b0011 : 4'b0010;
											assign node9439 = (inp[1]) ? node9451 : node9440;
												assign node9440 = (inp[5]) ? node9446 : node9441;
													assign node9441 = (inp[2]) ? node9443 : 4'b0010;
														assign node9443 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node9446 = (inp[12]) ? node9448 : 4'b0010;
														assign node9448 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node9451 = (inp[5]) ? node9463 : node9452;
													assign node9452 = (inp[10]) ? node9458 : node9453;
														assign node9453 = (inp[2]) ? node9455 : 4'b0111;
															assign node9455 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node9458 = (inp[2]) ? 4'b0111 : node9459;
															assign node9459 = (inp[7]) ? 4'b0011 : 4'b0111;
													assign node9463 = (inp[2]) ? node9467 : node9464;
														assign node9464 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node9467 = (inp[10]) ? 4'b0111 : 4'b0011;
										assign node9470 = (inp[13]) ? node9498 : node9471;
											assign node9471 = (inp[7]) ? node9487 : node9472;
												assign node9472 = (inp[2]) ? node9476 : node9473;
													assign node9473 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node9476 = (inp[5]) ? node9484 : node9477;
														assign node9477 = (inp[1]) ? node9481 : node9478;
															assign node9478 = (inp[10]) ? 4'b0001 : 4'b0100;
															assign node9481 = (inp[12]) ? 4'b0100 : 4'b0001;
														assign node9484 = (inp[1]) ? 4'b0001 : 4'b0101;
												assign node9487 = (inp[12]) ? node9493 : node9488;
													assign node9488 = (inp[1]) ? 4'b0000 : node9489;
														assign node9489 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node9493 = (inp[5]) ? node9495 : 4'b0000;
														assign node9495 = (inp[1]) ? 4'b0000 : 4'b0100;
											assign node9498 = (inp[7]) ? node9516 : node9499;
												assign node9499 = (inp[1]) ? node9509 : node9500;
													assign node9500 = (inp[5]) ? node9506 : node9501;
														assign node9501 = (inp[12]) ? node9503 : 4'b0100;
															assign node9503 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node9506 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node9509 = (inp[2]) ? node9511 : 4'b0100;
														assign node9511 = (inp[12]) ? 4'b0100 : node9512;
															assign node9512 = (inp[5]) ? 4'b0101 : 4'b0001;
												assign node9516 = (inp[1]) ? node9522 : node9517;
													assign node9517 = (inp[5]) ? node9519 : 4'b0001;
														assign node9519 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node9522 = (inp[5]) ? 4'b0001 : 4'b0101;
								assign node9525 = (inp[13]) ? node9661 : node9526;
									assign node9526 = (inp[1]) ? node9584 : node9527;
										assign node9527 = (inp[5]) ? node9559 : node9528;
											assign node9528 = (inp[12]) ? node9540 : node9529;
												assign node9529 = (inp[15]) ? node9535 : node9530;
													assign node9530 = (inp[4]) ? node9532 : 4'b0001;
														assign node9532 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node9535 = (inp[4]) ? 4'b0001 : node9536;
														assign node9536 = (inp[7]) ? 4'b0111 : 4'b0011;
												assign node9540 = (inp[15]) ? node9554 : node9541;
													assign node9541 = (inp[4]) ? node9547 : node9542;
														assign node9542 = (inp[2]) ? 4'b0100 : node9543;
															assign node9543 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node9547 = (inp[7]) ? node9551 : node9548;
															assign node9548 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node9551 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node9554 = (inp[7]) ? node9556 : 4'b0011;
														assign node9556 = (inp[4]) ? 4'b0000 : 4'b0010;
											assign node9559 = (inp[12]) ? node9571 : node9560;
												assign node9560 = (inp[7]) ? node9564 : node9561;
													assign node9561 = (inp[10]) ? 4'b0101 : 4'b0111;
													assign node9564 = (inp[4]) ? node9568 : node9565;
														assign node9565 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node9568 = (inp[15]) ? 4'b0101 : 4'b0110;
												assign node9571 = (inp[10]) ? node9577 : node9572;
													assign node9572 = (inp[4]) ? node9574 : 4'b0101;
														assign node9574 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node9577 = (inp[15]) ? 4'b0111 : node9578;
														assign node9578 = (inp[4]) ? 4'b0011 : node9579;
															assign node9579 = (inp[2]) ? 4'b0101 : 4'b0001;
										assign node9584 = (inp[5]) ? node9628 : node9585;
											assign node9585 = (inp[10]) ? node9605 : node9586;
												assign node9586 = (inp[12]) ? node9592 : node9587;
													assign node9587 = (inp[4]) ? node9589 : 4'b0101;
														assign node9589 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node9592 = (inp[15]) ? node9598 : node9593;
														assign node9593 = (inp[7]) ? node9595 : 4'b0010;
															assign node9595 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node9598 = (inp[4]) ? node9602 : node9599;
															assign node9599 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node9602 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node9605 = (inp[4]) ? node9617 : node9606;
													assign node9606 = (inp[15]) ? node9610 : node9607;
														assign node9607 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node9610 = (inp[7]) ? node9614 : node9611;
															assign node9611 = (inp[12]) ? 4'b0110 : 4'b0110;
															assign node9614 = (inp[12]) ? 4'b0111 : 4'b0010;
													assign node9617 = (inp[15]) ? node9623 : node9618;
														assign node9618 = (inp[7]) ? 4'b0110 : node9619;
															assign node9619 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node9623 = (inp[2]) ? 4'b0101 : node9624;
															assign node9624 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node9628 = (inp[12]) ? node9644 : node9629;
												assign node9629 = (inp[15]) ? node9637 : node9630;
													assign node9630 = (inp[4]) ? node9632 : 4'b0000;
														assign node9632 = (inp[10]) ? node9634 : 4'b0010;
															assign node9634 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node9637 = (inp[4]) ? node9641 : node9638;
														assign node9638 = (inp[7]) ? 4'b0111 : 4'b0010;
														assign node9641 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node9644 = (inp[2]) ? node9654 : node9645;
													assign node9645 = (inp[7]) ? node9649 : node9646;
														assign node9646 = (inp[15]) ? 4'b0011 : 4'b0111;
														assign node9649 = (inp[10]) ? node9651 : 4'b0100;
															assign node9651 = (inp[15]) ? 4'b0000 : 4'b0011;
													assign node9654 = (inp[7]) ? node9656 : 4'b0001;
														assign node9656 = (inp[10]) ? 4'b0010 : node9657;
															assign node9657 = (inp[4]) ? 4'b0001 : 4'b0011;
									assign node9661 = (inp[7]) ? node9705 : node9662;
										assign node9662 = (inp[5]) ? node9686 : node9663;
											assign node9663 = (inp[1]) ? node9677 : node9664;
												assign node9664 = (inp[4]) ? node9670 : node9665;
													assign node9665 = (inp[15]) ? node9667 : 4'b0000;
														assign node9667 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node9670 = (inp[15]) ? node9672 : 4'b0111;
														assign node9672 = (inp[12]) ? node9674 : 4'b0100;
															assign node9674 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node9677 = (inp[15]) ? node9681 : node9678;
													assign node9678 = (inp[4]) ? 4'b0011 : 4'b0101;
													assign node9681 = (inp[4]) ? 4'b0100 : node9682;
														assign node9682 = (inp[12]) ? 4'b0110 : 4'b0111;
											assign node9686 = (inp[1]) ? node9694 : node9687;
												assign node9687 = (inp[2]) ? node9689 : 4'b0101;
													assign node9689 = (inp[15]) ? node9691 : 4'b0100;
														assign node9691 = (inp[4]) ? 4'b0101 : 4'b0111;
												assign node9694 = (inp[4]) ? node9698 : node9695;
													assign node9695 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node9698 = (inp[10]) ? 4'b0010 : node9699;
														assign node9699 = (inp[12]) ? 4'b0111 : node9700;
															assign node9700 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node9705 = (inp[15]) ? node9727 : node9706;
											assign node9706 = (inp[4]) ? node9716 : node9707;
												assign node9707 = (inp[10]) ? 4'b0001 : node9708;
													assign node9708 = (inp[2]) ? node9712 : node9709;
														assign node9709 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node9712 = (inp[1]) ? 4'b0001 : 4'b0101;
												assign node9716 = (inp[1]) ? node9724 : node9717;
													assign node9717 = (inp[5]) ? node9721 : node9718;
														assign node9718 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node9721 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node9724 = (inp[5]) ? 4'b0011 : 4'b0111;
											assign node9727 = (inp[4]) ? node9735 : node9728;
												assign node9728 = (inp[12]) ? node9732 : node9729;
													assign node9729 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node9732 = (inp[2]) ? 4'b0111 : 4'b0011;
												assign node9735 = (inp[1]) ? node9745 : node9736;
													assign node9736 = (inp[5]) ? 4'b0101 : node9737;
														assign node9737 = (inp[12]) ? node9741 : node9738;
															assign node9738 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node9741 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node9745 = (inp[5]) ? 4'b0001 : 4'b0101;
						assign node9748 = (inp[11]) ? node10104 : node9749;
							assign node9749 = (inp[4]) ? node9951 : node9750;
								assign node9750 = (inp[15]) ? node9862 : node9751;
									assign node9751 = (inp[9]) ? node9815 : node9752;
										assign node9752 = (inp[12]) ? node9788 : node9753;
											assign node9753 = (inp[2]) ? node9767 : node9754;
												assign node9754 = (inp[7]) ? node9762 : node9755;
													assign node9755 = (inp[5]) ? node9759 : node9756;
														assign node9756 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node9759 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node9762 = (inp[13]) ? node9764 : 4'b0001;
														assign node9764 = (inp[5]) ? 4'b0001 : 4'b0101;
												assign node9767 = (inp[7]) ? node9777 : node9768;
													assign node9768 = (inp[10]) ? node9774 : node9769;
														assign node9769 = (inp[1]) ? 4'b0000 : node9770;
															assign node9770 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node9774 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node9777 = (inp[10]) ? node9783 : node9778;
														assign node9778 = (inp[13]) ? node9780 : 4'b0001;
															assign node9780 = (inp[5]) ? 4'b0001 : 4'b0100;
														assign node9783 = (inp[5]) ? 4'b0100 : node9784;
															assign node9784 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node9788 = (inp[1]) ? node9798 : node9789;
												assign node9789 = (inp[10]) ? node9793 : node9790;
													assign node9790 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node9793 = (inp[13]) ? node9795 : 4'b0001;
														assign node9795 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node9798 = (inp[2]) ? node9806 : node9799;
													assign node9799 = (inp[7]) ? node9803 : node9800;
														assign node9800 = (inp[5]) ? 4'b0000 : 4'b0100;
														assign node9803 = (inp[5]) ? 4'b0100 : 4'b0001;
													assign node9806 = (inp[7]) ? node9810 : node9807;
														assign node9807 = (inp[5]) ? 4'b0001 : 4'b0101;
														assign node9810 = (inp[5]) ? node9812 : 4'b0001;
															assign node9812 = (inp[13]) ? 4'b0101 : 4'b0100;
										assign node9815 = (inp[2]) ? node9839 : node9816;
											assign node9816 = (inp[5]) ? node9828 : node9817;
												assign node9817 = (inp[1]) ? node9823 : node9818;
													assign node9818 = (inp[13]) ? 4'b0001 : node9819;
														assign node9819 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node9823 = (inp[7]) ? node9825 : 4'b0100;
														assign node9825 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node9828 = (inp[1]) ? node9832 : node9829;
													assign node9829 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node9832 = (inp[10]) ? 4'b0001 : node9833;
														assign node9833 = (inp[12]) ? 4'b0100 : node9834;
															assign node9834 = (inp[13]) ? 4'b0000 : 4'b0000;
											assign node9839 = (inp[13]) ? node9853 : node9840;
												assign node9840 = (inp[12]) ? node9850 : node9841;
													assign node9841 = (inp[5]) ? node9845 : node9842;
														assign node9842 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node9845 = (inp[10]) ? node9847 : 4'b0000;
															assign node9847 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node9850 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node9853 = (inp[5]) ? node9859 : node9854;
													assign node9854 = (inp[1]) ? node9856 : 4'b0000;
														assign node9856 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node9859 = (inp[7]) ? 4'b0101 : 4'b0100;
									assign node9862 = (inp[12]) ? node9918 : node9863;
										assign node9863 = (inp[10]) ? node9889 : node9864;
											assign node9864 = (inp[1]) ? node9876 : node9865;
												assign node9865 = (inp[9]) ? node9871 : node9866;
													assign node9866 = (inp[2]) ? 4'b0010 : node9867;
														assign node9867 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node9871 = (inp[7]) ? 4'b0010 : node9872;
														assign node9872 = (inp[5]) ? 4'b0110 : 4'b0010;
												assign node9876 = (inp[13]) ? node9878 : 4'b0010;
													assign node9878 = (inp[9]) ? node9882 : node9879;
														assign node9879 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node9882 = (inp[5]) ? node9886 : node9883;
															assign node9883 = (inp[7]) ? 4'b0010 : 4'b0111;
															assign node9886 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node9889 = (inp[13]) ? node9901 : node9890;
												assign node9890 = (inp[1]) ? node9898 : node9891;
													assign node9891 = (inp[9]) ? node9893 : 4'b0111;
														assign node9893 = (inp[5]) ? node9895 : 4'b0011;
															assign node9895 = (inp[7]) ? 4'b0011 : 4'b0111;
													assign node9898 = (inp[2]) ? 4'b0010 : 4'b0111;
												assign node9901 = (inp[2]) ? node9907 : node9902;
													assign node9902 = (inp[7]) ? 4'b0010 : node9903;
														assign node9903 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node9907 = (inp[1]) ? node9911 : node9908;
														assign node9908 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node9911 = (inp[5]) ? node9915 : node9912;
															assign node9912 = (inp[7]) ? 4'b0010 : 4'b0111;
															assign node9915 = (inp[7]) ? 4'b0111 : 4'b0010;
										assign node9918 = (inp[5]) ? node9940 : node9919;
											assign node9919 = (inp[1]) ? node9931 : node9920;
												assign node9920 = (inp[13]) ? node9924 : node9921;
													assign node9921 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node9924 = (inp[10]) ? node9928 : node9925;
														assign node9925 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node9928 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node9931 = (inp[7]) ? node9937 : node9932;
													assign node9932 = (inp[13]) ? 4'b0110 : node9933;
														assign node9933 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node9937 = (inp[13]) ? 4'b0111 : 4'b0110;
											assign node9940 = (inp[1]) ? node9946 : node9941;
												assign node9941 = (inp[13]) ? node9943 : 4'b0111;
													assign node9943 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node9946 = (inp[13]) ? node9948 : 4'b0011;
													assign node9948 = (inp[2]) ? 4'b0011 : 4'b0010;
								assign node9951 = (inp[15]) ? node10033 : node9952;
									assign node9952 = (inp[13]) ? node10000 : node9953;
										assign node9953 = (inp[12]) ? node9975 : node9954;
											assign node9954 = (inp[9]) ? node9962 : node9955;
												assign node9955 = (inp[5]) ? node9959 : node9956;
													assign node9956 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node9959 = (inp[7]) ? 4'b0110 : 4'b0010;
												assign node9962 = (inp[10]) ? node9968 : node9963;
													assign node9963 = (inp[1]) ? node9965 : 4'b0011;
														assign node9965 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node9968 = (inp[5]) ? node9970 : 4'b0010;
														assign node9970 = (inp[2]) ? 4'b0011 : node9971;
															assign node9971 = (inp[7]) ? 4'b0011 : 4'b0010;
											assign node9975 = (inp[2]) ? node9983 : node9976;
												assign node9976 = (inp[9]) ? 4'b0111 : node9977;
													assign node9977 = (inp[5]) ? 4'b0111 : node9978;
														assign node9978 = (inp[7]) ? 4'b0111 : 4'b0010;
												assign node9983 = (inp[1]) ? node9993 : node9984;
													assign node9984 = (inp[9]) ? 4'b0111 : node9985;
														assign node9985 = (inp[10]) ? node9989 : node9986;
															assign node9986 = (inp[5]) ? 4'b0011 : 4'b0011;
															assign node9989 = (inp[7]) ? 4'b0011 : 4'b0110;
													assign node9993 = (inp[10]) ? node9995 : 4'b0010;
														assign node9995 = (inp[7]) ? node9997 : 4'b0110;
															assign node9997 = (inp[5]) ? 4'b0010 : 4'b0110;
										assign node10000 = (inp[1]) ? node10020 : node10001;
											assign node10001 = (inp[5]) ? node10009 : node10002;
												assign node10002 = (inp[7]) ? node10006 : node10003;
													assign node10003 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node10006 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node10009 = (inp[12]) ? node10017 : node10010;
													assign node10010 = (inp[10]) ? 4'b0111 : node10011;
														assign node10011 = (inp[9]) ? node10013 : 4'b0110;
															assign node10013 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node10017 = (inp[7]) ? 4'b0110 : 4'b0010;
											assign node10020 = (inp[5]) ? node10028 : node10021;
												assign node10021 = (inp[7]) ? 4'b0111 : node10022;
													assign node10022 = (inp[12]) ? node10024 : 4'b0111;
														assign node10024 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node10028 = (inp[7]) ? 4'b0011 : node10029;
													assign node10029 = (inp[12]) ? 4'b0111 : 4'b0010;
									assign node10033 = (inp[7]) ? node10075 : node10034;
										assign node10034 = (inp[13]) ? node10054 : node10035;
											assign node10035 = (inp[2]) ? node10041 : node10036;
												assign node10036 = (inp[1]) ? 4'b0000 : node10037;
													assign node10037 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node10041 = (inp[1]) ? node10049 : node10042;
													assign node10042 = (inp[5]) ? node10046 : node10043;
														assign node10043 = (inp[12]) ? 4'b0001 : 4'b0100;
														assign node10046 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node10049 = (inp[12]) ? node10051 : 4'b0100;
														assign node10051 = (inp[5]) ? 4'b0001 : 4'b0100;
											assign node10054 = (inp[5]) ? node10064 : node10055;
												assign node10055 = (inp[2]) ? node10061 : node10056;
													assign node10056 = (inp[10]) ? node10058 : 4'b0001;
														assign node10058 = (inp[1]) ? 4'b0001 : 4'b0100;
													assign node10061 = (inp[12]) ? 4'b0100 : 4'b0001;
												assign node10064 = (inp[10]) ? node10070 : node10065;
													assign node10065 = (inp[1]) ? node10067 : 4'b0001;
														assign node10067 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node10070 = (inp[12]) ? node10072 : 4'b0101;
														assign node10072 = (inp[2]) ? 4'b0001 : 4'b0101;
										assign node10075 = (inp[1]) ? node10097 : node10076;
											assign node10076 = (inp[5]) ? node10090 : node10077;
												assign node10077 = (inp[9]) ? node10083 : node10078;
													assign node10078 = (inp[12]) ? 4'b0000 : node10079;
														assign node10079 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node10083 = (inp[13]) ? node10085 : 4'b0001;
														assign node10085 = (inp[12]) ? node10087 : 4'b0000;
															assign node10087 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node10090 = (inp[12]) ? 4'b0101 : node10091;
													assign node10091 = (inp[13]) ? 4'b0100 : node10092;
														assign node10092 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node10097 = (inp[5]) ? 4'b0001 : node10098;
												assign node10098 = (inp[2]) ? 4'b0101 : node10099;
													assign node10099 = (inp[13]) ? 4'b0101 : 4'b0100;
							assign node10104 = (inp[13]) ? node10278 : node10105;
								assign node10105 = (inp[4]) ? node10177 : node10106;
									assign node10106 = (inp[15]) ? node10138 : node10107;
										assign node10107 = (inp[5]) ? node10125 : node10108;
											assign node10108 = (inp[2]) ? node10118 : node10109;
												assign node10109 = (inp[1]) ? node10115 : node10110;
													assign node10110 = (inp[7]) ? node10112 : 4'b0000;
														assign node10112 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node10115 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node10118 = (inp[12]) ? node10122 : node10119;
													assign node10119 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node10122 = (inp[1]) ? 4'b0000 : 4'b0101;
											assign node10125 = (inp[1]) ? node10129 : node10126;
												assign node10126 = (inp[7]) ? 4'b0000 : 4'b0100;
												assign node10129 = (inp[7]) ? node10135 : node10130;
													assign node10130 = (inp[2]) ? node10132 : 4'b0001;
														assign node10132 = (inp[12]) ? 4'b0000 : 4'b0001;
													assign node10135 = (inp[12]) ? 4'b0101 : 4'b0001;
										assign node10138 = (inp[7]) ? node10150 : node10139;
											assign node10139 = (inp[1]) ? node10143 : node10140;
												assign node10140 = (inp[5]) ? 4'b0110 : 4'b0010;
												assign node10143 = (inp[5]) ? node10147 : node10144;
													assign node10144 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node10147 = (inp[12]) ? 4'b0010 : 4'b0011;
											assign node10150 = (inp[9]) ? node10170 : node10151;
												assign node10151 = (inp[12]) ? node10165 : node10152;
													assign node10152 = (inp[2]) ? node10160 : node10153;
														assign node10153 = (inp[1]) ? node10157 : node10154;
															assign node10154 = (inp[5]) ? 4'b0011 : 4'b0110;
															assign node10157 = (inp[10]) ? 4'b0110 : 4'b0011;
														assign node10160 = (inp[5]) ? node10162 : 4'b0110;
															assign node10162 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node10165 = (inp[5]) ? 4'b0010 : node10166;
														assign node10166 = (inp[1]) ? 4'b0111 : 4'b0011;
												assign node10170 = (inp[5]) ? node10172 : 4'b0011;
													assign node10172 = (inp[2]) ? 4'b0010 : node10173;
														assign node10173 = (inp[1]) ? 4'b0010 : 4'b0011;
									assign node10177 = (inp[15]) ? node10227 : node10178;
										assign node10178 = (inp[2]) ? node10200 : node10179;
											assign node10179 = (inp[5]) ? node10189 : node10180;
												assign node10180 = (inp[12]) ? node10184 : node10181;
													assign node10181 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node10184 = (inp[1]) ? 4'b0011 : node10185;
														assign node10185 = (inp[7]) ? 4'b0011 : 4'b0110;
												assign node10189 = (inp[1]) ? node10195 : node10190;
													assign node10190 = (inp[7]) ? node10192 : 4'b0011;
														assign node10192 = (inp[12]) ? 4'b0110 : 4'b0111;
													assign node10195 = (inp[7]) ? 4'b0010 : node10196;
														assign node10196 = (inp[12]) ? 4'b0110 : 4'b0011;
											assign node10200 = (inp[5]) ? node10214 : node10201;
												assign node10201 = (inp[7]) ? node10209 : node10202;
													assign node10202 = (inp[10]) ? 4'b0111 : node10203;
														assign node10203 = (inp[1]) ? 4'b0011 : node10204;
															assign node10204 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node10209 = (inp[1]) ? 4'b0111 : node10210;
														assign node10210 = (inp[12]) ? 4'b0010 : 4'b0011;
												assign node10214 = (inp[1]) ? node10222 : node10215;
													assign node10215 = (inp[7]) ? node10219 : node10216;
														assign node10216 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node10219 = (inp[12]) ? 4'b0110 : 4'b0111;
													assign node10222 = (inp[12]) ? 4'b0111 : node10223;
														assign node10223 = (inp[10]) ? 4'b0011 : 4'b0010;
										assign node10227 = (inp[2]) ? node10251 : node10228;
											assign node10228 = (inp[1]) ? node10240 : node10229;
												assign node10229 = (inp[12]) ? node10237 : node10230;
													assign node10230 = (inp[7]) ? node10234 : node10231;
														assign node10231 = (inp[10]) ? 4'b0001 : 4'b0100;
														assign node10234 = (inp[5]) ? 4'b0100 : 4'b0000;
													assign node10237 = (inp[5]) ? 4'b0101 : 4'b0001;
												assign node10240 = (inp[10]) ? node10246 : node10241;
													assign node10241 = (inp[5]) ? node10243 : 4'b0101;
														assign node10243 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node10246 = (inp[9]) ? node10248 : 4'b0001;
														assign node10248 = (inp[7]) ? 4'b0001 : 4'b0100;
											assign node10251 = (inp[7]) ? node10269 : node10252;
												assign node10252 = (inp[10]) ? node10262 : node10253;
													assign node10253 = (inp[9]) ? node10257 : node10254;
														assign node10254 = (inp[5]) ? 4'b0101 : 4'b0000;
														assign node10257 = (inp[12]) ? node10259 : 4'b0000;
															assign node10259 = (inp[1]) ? 4'b0000 : 4'b0100;
													assign node10262 = (inp[1]) ? 4'b0101 : node10263;
														assign node10263 = (inp[12]) ? node10265 : 4'b0101;
															assign node10265 = (inp[5]) ? 4'b0100 : 4'b0000;
												assign node10269 = (inp[1]) ? node10275 : node10270;
													assign node10270 = (inp[5]) ? node10272 : 4'b0000;
														assign node10272 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node10275 = (inp[5]) ? 4'b0000 : 4'b0100;
								assign node10278 = (inp[4]) ? node10382 : node10279;
									assign node10279 = (inp[15]) ? node10329 : node10280;
										assign node10280 = (inp[2]) ? node10304 : node10281;
											assign node10281 = (inp[12]) ? node10291 : node10282;
												assign node10282 = (inp[1]) ? node10288 : node10283;
													assign node10283 = (inp[7]) ? 4'b0101 : node10284;
														assign node10284 = (inp[5]) ? 4'b0100 : 4'b0000;
													assign node10288 = (inp[5]) ? 4'b0000 : 4'b0100;
												assign node10291 = (inp[1]) ? node10297 : node10292;
													assign node10292 = (inp[5]) ? node10294 : 4'b0000;
														assign node10294 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node10297 = (inp[9]) ? node10301 : node10298;
														assign node10298 = (inp[10]) ? 4'b0101 : 4'b0000;
														assign node10301 = (inp[7]) ? 4'b0101 : 4'b0000;
											assign node10304 = (inp[9]) ? node10318 : node10305;
												assign node10305 = (inp[1]) ? node10313 : node10306;
													assign node10306 = (inp[5]) ? 4'b0101 : node10307;
														assign node10307 = (inp[7]) ? node10309 : 4'b0001;
															assign node10309 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node10313 = (inp[10]) ? node10315 : 4'b0001;
														assign node10315 = (inp[12]) ? 4'b0100 : 4'b0001;
												assign node10318 = (inp[5]) ? node10326 : node10319;
													assign node10319 = (inp[1]) ? node10321 : 4'b0001;
														assign node10321 = (inp[12]) ? node10323 : 4'b0101;
															assign node10323 = (inp[7]) ? 4'b0001 : 4'b0100;
													assign node10326 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node10329 = (inp[2]) ? node10351 : node10330;
											assign node10330 = (inp[10]) ? node10346 : node10331;
												assign node10331 = (inp[9]) ? node10335 : node10332;
													assign node10332 = (inp[5]) ? 4'b0111 : 4'b0010;
													assign node10335 = (inp[5]) ? node10341 : node10336;
														assign node10336 = (inp[1]) ? node10338 : 4'b0111;
															assign node10338 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node10341 = (inp[1]) ? node10343 : 4'b0111;
															assign node10343 = (inp[7]) ? 4'b0111 : 4'b0011;
												assign node10346 = (inp[7]) ? node10348 : 4'b0011;
													assign node10348 = (inp[1]) ? 4'b0011 : 4'b0111;
											assign node10351 = (inp[5]) ? node10365 : node10352;
												assign node10352 = (inp[10]) ? node10358 : node10353;
													assign node10353 = (inp[7]) ? 4'b0011 : node10354;
														assign node10354 = (inp[12]) ? 4'b0111 : 4'b0110;
													assign node10358 = (inp[7]) ? node10360 : 4'b0010;
														assign node10360 = (inp[9]) ? node10362 : 4'b0110;
															assign node10362 = (inp[1]) ? 4'b0110 : 4'b0011;
												assign node10365 = (inp[12]) ? node10379 : node10366;
													assign node10366 = (inp[10]) ? node10372 : node10367;
														assign node10367 = (inp[1]) ? 4'b0110 : node10368;
															assign node10368 = (inp[7]) ? 4'b0011 : 4'b0110;
														assign node10372 = (inp[1]) ? node10376 : node10373;
															assign node10373 = (inp[9]) ? 4'b0110 : 4'b0011;
															assign node10376 = (inp[9]) ? 4'b0011 : 4'b0110;
													assign node10379 = (inp[1]) ? 4'b0010 : 4'b0110;
									assign node10382 = (inp[15]) ? node10418 : node10383;
										assign node10383 = (inp[5]) ? node10397 : node10384;
											assign node10384 = (inp[1]) ? node10392 : node10385;
												assign node10385 = (inp[7]) ? node10389 : node10386;
													assign node10386 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node10389 = (inp[12]) ? 4'b0011 : 4'b0010;
												assign node10392 = (inp[12]) ? node10394 : 4'b0110;
													assign node10394 = (inp[2]) ? 4'b0011 : 4'b0110;
											assign node10397 = (inp[1]) ? node10411 : node10398;
												assign node10398 = (inp[9]) ? 4'b0111 : node10399;
													assign node10399 = (inp[12]) ? node10405 : node10400;
														assign node10400 = (inp[10]) ? 4'b0110 : node10401;
															assign node10401 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node10405 = (inp[7]) ? node10407 : 4'b0011;
															assign node10407 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node10411 = (inp[12]) ? node10415 : node10412;
													assign node10412 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node10415 = (inp[7]) ? 4'b0010 : 4'b0110;
										assign node10418 = (inp[2]) ? node10442 : node10419;
											assign node10419 = (inp[1]) ? node10431 : node10420;
												assign node10420 = (inp[5]) ? node10426 : node10421;
													assign node10421 = (inp[7]) ? node10423 : 4'b0101;
														assign node10423 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node10426 = (inp[7]) ? 4'b0101 : node10427;
														assign node10427 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node10431 = (inp[5]) ? node10439 : node10432;
													assign node10432 = (inp[12]) ? node10436 : node10433;
														assign node10433 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node10436 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node10439 = (inp[12]) ? 4'b0000 : 4'b0101;
											assign node10442 = (inp[5]) ? node10454 : node10443;
												assign node10443 = (inp[1]) ? node10449 : node10444;
													assign node10444 = (inp[12]) ? 4'b0000 : node10445;
														assign node10445 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node10449 = (inp[7]) ? 4'b0100 : node10450;
														assign node10450 = (inp[12]) ? 4'b0101 : 4'b0000;
												assign node10454 = (inp[1]) ? 4'b0000 : node10455;
													assign node10455 = (inp[7]) ? node10459 : node10456;
														assign node10456 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node10459 = (inp[9]) ? 4'b0101 : 4'b0100;
				assign node10463 = (inp[4]) ? node12049 : node10464;
					assign node10464 = (inp[7]) ? node11166 : node10465;
						assign node10465 = (inp[8]) ? node10891 : node10466;
							assign node10466 = (inp[11]) ? node10700 : node10467;
								assign node10467 = (inp[2]) ? node10585 : node10468;
									assign node10468 = (inp[10]) ? node10526 : node10469;
										assign node10469 = (inp[9]) ? node10495 : node10470;
											assign node10470 = (inp[13]) ? node10480 : node10471;
												assign node10471 = (inp[12]) ? node10475 : node10472;
													assign node10472 = (inp[15]) ? 4'b0101 : 4'b0000;
													assign node10475 = (inp[5]) ? 4'b0100 : node10476;
														assign node10476 = (inp[15]) ? 4'b0000 : 4'b0100;
												assign node10480 = (inp[12]) ? node10486 : node10481;
													assign node10481 = (inp[1]) ? 4'b0000 : node10482;
														assign node10482 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node10486 = (inp[15]) ? node10492 : node10487;
														assign node10487 = (inp[0]) ? 4'b0001 : node10488;
															assign node10488 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node10492 = (inp[0]) ? 4'b0000 : 4'b0101;
											assign node10495 = (inp[1]) ? node10511 : node10496;
												assign node10496 = (inp[0]) ? node10508 : node10497;
													assign node10497 = (inp[15]) ? node10503 : node10498;
														assign node10498 = (inp[12]) ? 4'b0101 : node10499;
															assign node10499 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node10503 = (inp[13]) ? node10505 : 4'b0001;
															assign node10505 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node10508 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node10511 = (inp[0]) ? node10513 : 4'b0100;
													assign node10513 = (inp[15]) ? node10521 : node10514;
														assign node10514 = (inp[13]) ? node10518 : node10515;
															assign node10515 = (inp[5]) ? 4'b0101 : 4'b0001;
															assign node10518 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node10521 = (inp[13]) ? 4'b0101 : node10522;
															assign node10522 = (inp[12]) ? 4'b0000 : 4'b0100;
										assign node10526 = (inp[1]) ? node10558 : node10527;
											assign node10527 = (inp[12]) ? node10541 : node10528;
												assign node10528 = (inp[13]) ? node10534 : node10529;
													assign node10529 = (inp[9]) ? node10531 : 4'b0000;
														assign node10531 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node10534 = (inp[5]) ? node10536 : 4'b0101;
														assign node10536 = (inp[9]) ? 4'b0100 : node10537;
															assign node10537 = (inp[15]) ? 4'b0100 : 4'b0100;
												assign node10541 = (inp[13]) ? node10545 : node10542;
													assign node10542 = (inp[15]) ? 4'b0100 : 4'b0101;
													assign node10545 = (inp[9]) ? node10553 : node10546;
														assign node10546 = (inp[15]) ? node10550 : node10547;
															assign node10547 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node10550 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node10553 = (inp[15]) ? 4'b0001 : node10554;
															assign node10554 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node10558 = (inp[0]) ? node10572 : node10559;
												assign node10559 = (inp[9]) ? node10565 : node10560;
													assign node10560 = (inp[15]) ? node10562 : 4'b0000;
														assign node10562 = (inp[5]) ? 4'b0101 : 4'b0000;
													assign node10565 = (inp[12]) ? node10567 : 4'b0001;
														assign node10567 = (inp[15]) ? 4'b0001 : node10568;
															assign node10568 = (inp[13]) ? 4'b0001 : 4'b0100;
												assign node10572 = (inp[15]) ? node10578 : node10573;
													assign node10573 = (inp[12]) ? node10575 : 4'b0101;
														assign node10575 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node10578 = (inp[12]) ? node10580 : 4'b0000;
														assign node10580 = (inp[13]) ? 4'b0101 : node10581;
															assign node10581 = (inp[5]) ? 4'b0001 : 4'b0000;
									assign node10585 = (inp[1]) ? node10633 : node10586;
										assign node10586 = (inp[13]) ? node10606 : node10587;
											assign node10587 = (inp[12]) ? node10601 : node10588;
												assign node10588 = (inp[15]) ? 4'b0001 : node10589;
													assign node10589 = (inp[9]) ? node10595 : node10590;
														assign node10590 = (inp[0]) ? node10592 : 4'b0001;
															assign node10592 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node10595 = (inp[10]) ? 4'b0001 : node10596;
															assign node10596 = (inp[0]) ? 4'b0000 : 4'b0000;
												assign node10601 = (inp[9]) ? node10603 : 4'b0101;
													assign node10603 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node10606 = (inp[12]) ? node10616 : node10607;
												assign node10607 = (inp[5]) ? 4'b0101 : node10608;
													assign node10608 = (inp[9]) ? node10612 : node10609;
														assign node10609 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node10612 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node10616 = (inp[10]) ? node10626 : node10617;
													assign node10617 = (inp[0]) ? node10621 : node10618;
														assign node10618 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node10621 = (inp[9]) ? 4'b0001 : node10622;
															assign node10622 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node10626 = (inp[15]) ? node10628 : 4'b0000;
														assign node10628 = (inp[0]) ? 4'b0001 : node10629;
															assign node10629 = (inp[5]) ? 4'b0000 : 4'b0001;
										assign node10633 = (inp[13]) ? node10675 : node10634;
											assign node10634 = (inp[10]) ? node10650 : node10635;
												assign node10635 = (inp[0]) ? node10643 : node10636;
													assign node10636 = (inp[5]) ? 4'b0000 : node10637;
														assign node10637 = (inp[12]) ? 4'b0100 : node10638;
															assign node10638 = (inp[15]) ? 4'b0100 : 4'b0000;
													assign node10643 = (inp[12]) ? 4'b0000 : node10644;
														assign node10644 = (inp[15]) ? node10646 : 4'b0001;
															assign node10646 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node10650 = (inp[5]) ? node10662 : node10651;
													assign node10651 = (inp[12]) ? node10659 : node10652;
														assign node10652 = (inp[15]) ? node10656 : node10653;
															assign node10653 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node10656 = (inp[9]) ? 4'b0100 : 4'b0100;
														assign node10659 = (inp[15]) ? 4'b0001 : 4'b0101;
													assign node10662 = (inp[15]) ? node10670 : node10663;
														assign node10663 = (inp[12]) ? node10667 : node10664;
															assign node10664 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node10667 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node10670 = (inp[9]) ? node10672 : 4'b0000;
															assign node10672 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node10675 = (inp[9]) ? node10689 : node10676;
												assign node10676 = (inp[12]) ? node10682 : node10677;
													assign node10677 = (inp[15]) ? 4'b0001 : node10678;
														assign node10678 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node10682 = (inp[15]) ? 4'b0100 : node10683;
														assign node10683 = (inp[5]) ? 4'b0001 : node10684;
															assign node10684 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node10689 = (inp[15]) ? node10697 : node10690;
													assign node10690 = (inp[12]) ? node10694 : node10691;
														assign node10691 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node10694 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node10697 = (inp[12]) ? 4'b0101 : 4'b0001;
								assign node10700 = (inp[2]) ? node10786 : node10701;
									assign node10701 = (inp[9]) ? node10749 : node10702;
										assign node10702 = (inp[1]) ? node10722 : node10703;
											assign node10703 = (inp[0]) ? node10711 : node10704;
												assign node10704 = (inp[5]) ? node10708 : node10705;
													assign node10705 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node10708 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node10711 = (inp[5]) ? node10717 : node10712;
													assign node10712 = (inp[15]) ? node10714 : 4'b0100;
														assign node10714 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node10717 = (inp[12]) ? 4'b0101 : node10718;
														assign node10718 = (inp[15]) ? 4'b0001 : 4'b0101;
											assign node10722 = (inp[12]) ? node10734 : node10723;
												assign node10723 = (inp[15]) ? node10731 : node10724;
													assign node10724 = (inp[13]) ? node10726 : 4'b0000;
														assign node10726 = (inp[5]) ? node10728 : 4'b0100;
															assign node10728 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node10731 = (inp[13]) ? 4'b0000 : 4'b0101;
												assign node10734 = (inp[5]) ? node10744 : node10735;
													assign node10735 = (inp[13]) ? node10739 : node10736;
														assign node10736 = (inp[15]) ? 4'b0000 : 4'b0101;
														assign node10739 = (inp[15]) ? 4'b0101 : node10740;
															assign node10740 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node10744 = (inp[13]) ? 4'b0100 : node10745;
														assign node10745 = (inp[15]) ? 4'b0001 : 4'b0100;
										assign node10749 = (inp[12]) ? node10765 : node10750;
											assign node10750 = (inp[13]) ? node10756 : node10751;
												assign node10751 = (inp[0]) ? node10753 : 4'b0001;
													assign node10753 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node10756 = (inp[15]) ? node10758 : 4'b0101;
													assign node10758 = (inp[1]) ? node10762 : node10759;
														assign node10759 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node10762 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node10765 = (inp[13]) ? node10773 : node10766;
												assign node10766 = (inp[1]) ? 4'b0100 : node10767;
													assign node10767 = (inp[5]) ? node10769 : 4'b0101;
														assign node10769 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node10773 = (inp[15]) ? node10779 : node10774;
													assign node10774 = (inp[0]) ? 4'b0000 : node10775;
														assign node10775 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node10779 = (inp[1]) ? node10781 : 4'b0001;
														assign node10781 = (inp[0]) ? node10783 : 4'b0100;
															assign node10783 = (inp[5]) ? 4'b0101 : 4'b0100;
									assign node10786 = (inp[9]) ? node10842 : node10787;
										assign node10787 = (inp[0]) ? node10813 : node10788;
											assign node10788 = (inp[13]) ? node10798 : node10789;
												assign node10789 = (inp[1]) ? node10793 : node10790;
													assign node10790 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node10793 = (inp[10]) ? 4'b0100 : node10794;
														assign node10794 = (inp[5]) ? 4'b0001 : 4'b0101;
												assign node10798 = (inp[12]) ? node10804 : node10799;
													assign node10799 = (inp[15]) ? node10801 : 4'b0101;
														assign node10801 = (inp[1]) ? 4'b0001 : 4'b0100;
													assign node10804 = (inp[15]) ? node10810 : node10805;
														assign node10805 = (inp[1]) ? 4'b0000 : node10806;
															assign node10806 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node10810 = (inp[1]) ? 4'b0100 : 4'b0000;
											assign node10813 = (inp[12]) ? node10825 : node10814;
												assign node10814 = (inp[15]) ? node10820 : node10815;
													assign node10815 = (inp[5]) ? node10817 : 4'b0001;
														assign node10817 = (inp[13]) ? 4'b0100 : 4'b0000;
													assign node10820 = (inp[1]) ? 4'b0100 : node10821;
														assign node10821 = (inp[13]) ? 4'b0100 : 4'b0001;
												assign node10825 = (inp[5]) ? node10835 : node10826;
													assign node10826 = (inp[1]) ? node10828 : 4'b0101;
														assign node10828 = (inp[15]) ? node10832 : node10829;
															assign node10829 = (inp[13]) ? 4'b0001 : 4'b0100;
															assign node10832 = (inp[13]) ? 4'b0100 : 4'b0001;
													assign node10835 = (inp[13]) ? node10837 : 4'b0000;
														assign node10837 = (inp[1]) ? node10839 : 4'b0000;
															assign node10839 = (inp[15]) ? 4'b0101 : 4'b0001;
										assign node10842 = (inp[5]) ? node10868 : node10843;
											assign node10843 = (inp[12]) ? node10855 : node10844;
												assign node10844 = (inp[13]) ? node10852 : node10845;
													assign node10845 = (inp[1]) ? node10847 : 4'b0000;
														assign node10847 = (inp[0]) ? 4'b0101 : node10848;
															assign node10848 = (inp[15]) ? 4'b0100 : 4'b0000;
													assign node10852 = (inp[15]) ? 4'b0000 : 4'b0100;
												assign node10855 = (inp[13]) ? node10861 : node10856;
													assign node10856 = (inp[15]) ? node10858 : 4'b0101;
														assign node10858 = (inp[1]) ? 4'b0000 : 4'b0100;
													assign node10861 = (inp[10]) ? 4'b0001 : node10862;
														assign node10862 = (inp[15]) ? node10864 : 4'b0000;
															assign node10864 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node10868 = (inp[13]) ? node10882 : node10869;
												assign node10869 = (inp[0]) ? 4'b0001 : node10870;
													assign node10870 = (inp[1]) ? node10874 : node10871;
														assign node10871 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node10874 = (inp[12]) ? node10878 : node10875;
															assign node10875 = (inp[15]) ? 4'b0101 : 4'b0000;
															assign node10878 = (inp[15]) ? 4'b0000 : 4'b0101;
												assign node10882 = (inp[1]) ? node10886 : node10883;
													assign node10883 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node10886 = (inp[15]) ? 4'b0100 : node10887;
														assign node10887 = (inp[0]) ? 4'b0000 : 4'b0100;
							assign node10891 = (inp[0]) ? node10991 : node10892;
								assign node10892 = (inp[2]) ? node10944 : node10893;
									assign node10893 = (inp[13]) ? node10909 : node10894;
										assign node10894 = (inp[1]) ? node10898 : node10895;
											assign node10895 = (inp[12]) ? 4'b0110 : 4'b0010;
											assign node10898 = (inp[12]) ? node10904 : node10899;
												assign node10899 = (inp[15]) ? node10901 : 4'b0110;
													assign node10901 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node10904 = (inp[15]) ? 4'b0010 : node10905;
													assign node10905 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node10909 = (inp[1]) ? node10933 : node10910;
											assign node10910 = (inp[12]) ? node10918 : node10911;
												assign node10911 = (inp[15]) ? node10915 : node10912;
													assign node10912 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node10915 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node10918 = (inp[11]) ? node10928 : node10919;
													assign node10919 = (inp[9]) ? node10921 : 4'b0110;
														assign node10921 = (inp[15]) ? node10925 : node10922;
															assign node10922 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node10925 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node10928 = (inp[9]) ? node10930 : 4'b0111;
														assign node10930 = (inp[15]) ? 4'b0111 : 4'b0110;
											assign node10933 = (inp[12]) ? node10939 : node10934;
												assign node10934 = (inp[15]) ? 4'b0110 : node10935;
													assign node10935 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node10939 = (inp[15]) ? node10941 : 4'b0010;
													assign node10941 = (inp[5]) ? 4'b0010 : 4'b0011;
									assign node10944 = (inp[13]) ? node10960 : node10945;
										assign node10945 = (inp[1]) ? node10949 : node10946;
											assign node10946 = (inp[12]) ? 4'b0111 : 4'b0011;
											assign node10949 = (inp[12]) ? node10955 : node10950;
												assign node10950 = (inp[15]) ? node10952 : 4'b0111;
													assign node10952 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node10955 = (inp[15]) ? 4'b0011 : node10956;
													assign node10956 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node10960 = (inp[1]) ? node10980 : node10961;
											assign node10961 = (inp[12]) ? node10971 : node10962;
												assign node10962 = (inp[9]) ? node10968 : node10963;
													assign node10963 = (inp[10]) ? node10965 : 4'b0011;
														assign node10965 = (inp[15]) ? 4'b0010 : 4'b0011;
													assign node10968 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node10971 = (inp[9]) ? node10977 : node10972;
													assign node10972 = (inp[5]) ? node10974 : 4'b0111;
														assign node10974 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node10977 = (inp[15]) ? 4'b0110 : 4'b0111;
											assign node10980 = (inp[12]) ? node10986 : node10981;
												assign node10981 = (inp[15]) ? 4'b0111 : node10982;
													assign node10982 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node10986 = (inp[15]) ? node10988 : 4'b0011;
													assign node10988 = (inp[5]) ? 4'b0011 : 4'b0010;
								assign node10991 = (inp[2]) ? node11085 : node10992;
									assign node10992 = (inp[11]) ? node11044 : node10993;
										assign node10993 = (inp[10]) ? node11025 : node10994;
											assign node10994 = (inp[9]) ? node11008 : node10995;
												assign node10995 = (inp[12]) ? node11001 : node10996;
													assign node10996 = (inp[1]) ? 4'b0111 : node10997;
														assign node10997 = (inp[15]) ? 4'b0010 : 4'b0011;
													assign node11001 = (inp[5]) ? 4'b0011 : node11002;
														assign node11002 = (inp[15]) ? 4'b0010 : node11003;
															assign node11003 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node11008 = (inp[15]) ? node11016 : node11009;
													assign node11009 = (inp[12]) ? node11013 : node11010;
														assign node11010 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node11013 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node11016 = (inp[5]) ? node11020 : node11017;
														assign node11017 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node11020 = (inp[12]) ? 4'b0111 : node11021;
															assign node11021 = (inp[1]) ? 4'b0111 : 4'b0011;
											assign node11025 = (inp[15]) ? node11033 : node11026;
												assign node11026 = (inp[13]) ? node11028 : 4'b0011;
													assign node11028 = (inp[5]) ? node11030 : 4'b0011;
														assign node11030 = (inp[12]) ? 4'b0011 : 4'b0010;
												assign node11033 = (inp[9]) ? 4'b0011 : node11034;
													assign node11034 = (inp[12]) ? node11040 : node11035;
														assign node11035 = (inp[13]) ? 4'b0111 : node11036;
															assign node11036 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node11040 = (inp[1]) ? 4'b0011 : 4'b0111;
										assign node11044 = (inp[13]) ? node11062 : node11045;
											assign node11045 = (inp[9]) ? node11053 : node11046;
												assign node11046 = (inp[1]) ? node11050 : node11047;
													assign node11047 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node11050 = (inp[15]) ? 4'b0011 : 4'b0010;
												assign node11053 = (inp[12]) ? node11059 : node11054;
													assign node11054 = (inp[5]) ? node11056 : 4'b0111;
														assign node11056 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node11059 = (inp[1]) ? 4'b0011 : 4'b0111;
											assign node11062 = (inp[1]) ? node11074 : node11063;
												assign node11063 = (inp[12]) ? node11067 : node11064;
													assign node11064 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node11067 = (inp[9]) ? 4'b0110 : node11068;
														assign node11068 = (inp[10]) ? node11070 : 4'b0111;
															assign node11070 = (inp[15]) ? 4'b0111 : 4'b0110;
												assign node11074 = (inp[12]) ? node11080 : node11075;
													assign node11075 = (inp[5]) ? node11077 : 4'b0111;
														assign node11077 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node11080 = (inp[10]) ? node11082 : 4'b0011;
														assign node11082 = (inp[15]) ? 4'b0010 : 4'b0011;
									assign node11085 = (inp[13]) ? node11135 : node11086;
										assign node11086 = (inp[11]) ? node11108 : node11087;
											assign node11087 = (inp[10]) ? node11101 : node11088;
												assign node11088 = (inp[9]) ? node11092 : node11089;
													assign node11089 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node11092 = (inp[5]) ? node11096 : node11093;
														assign node11093 = (inp[12]) ? 4'b0011 : 4'b0110;
														assign node11096 = (inp[12]) ? node11098 : 4'b0010;
															assign node11098 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node11101 = (inp[1]) ? node11103 : 4'b0110;
													assign node11103 = (inp[5]) ? node11105 : 4'b0110;
														assign node11105 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node11108 = (inp[5]) ? node11128 : node11109;
												assign node11109 = (inp[9]) ? node11119 : node11110;
													assign node11110 = (inp[10]) ? node11112 : 4'b0110;
														assign node11112 = (inp[1]) ? node11116 : node11113;
															assign node11113 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node11116 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node11119 = (inp[10]) ? node11125 : node11120;
														assign node11120 = (inp[1]) ? node11122 : 4'b0010;
															assign node11122 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node11125 = (inp[1]) ? 4'b0011 : 4'b0110;
												assign node11128 = (inp[12]) ? node11132 : node11129;
													assign node11129 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node11132 = (inp[1]) ? 4'b0010 : 4'b0110;
										assign node11135 = (inp[1]) ? node11155 : node11136;
											assign node11136 = (inp[12]) ? node11144 : node11137;
												assign node11137 = (inp[15]) ? node11141 : node11138;
													assign node11138 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node11141 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node11144 = (inp[9]) ? node11150 : node11145;
													assign node11145 = (inp[5]) ? 4'b0110 : node11146;
														assign node11146 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node11150 = (inp[5]) ? 4'b0111 : node11151;
														assign node11151 = (inp[15]) ? 4'b0111 : 4'b0110;
											assign node11155 = (inp[12]) ? node11161 : node11156;
												assign node11156 = (inp[5]) ? node11158 : 4'b0110;
													assign node11158 = (inp[15]) ? 4'b0110 : 4'b0111;
												assign node11161 = (inp[15]) ? node11163 : 4'b0010;
													assign node11163 = (inp[5]) ? 4'b0010 : 4'b0011;
						assign node11166 = (inp[11]) ? node11610 : node11167;
							assign node11167 = (inp[2]) ? node11389 : node11168;
								assign node11168 = (inp[0]) ? node11288 : node11169;
									assign node11169 = (inp[8]) ? node11239 : node11170;
										assign node11170 = (inp[1]) ? node11196 : node11171;
											assign node11171 = (inp[5]) ? node11189 : node11172;
												assign node11172 = (inp[12]) ? node11182 : node11173;
													assign node11173 = (inp[9]) ? 4'b0011 : node11174;
														assign node11174 = (inp[13]) ? node11178 : node11175;
															assign node11175 = (inp[15]) ? 4'b0110 : 4'b0010;
															assign node11178 = (inp[10]) ? 4'b0011 : 4'b0110;
													assign node11182 = (inp[9]) ? node11184 : 4'b0011;
														assign node11184 = (inp[15]) ? 4'b0010 : node11185;
															assign node11185 = (inp[13]) ? 4'b0010 : 4'b0111;
												assign node11189 = (inp[13]) ? node11193 : node11190;
													assign node11190 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node11193 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node11196 = (inp[15]) ? node11220 : node11197;
												assign node11197 = (inp[5]) ? node11213 : node11198;
													assign node11198 = (inp[9]) ? node11206 : node11199;
														assign node11199 = (inp[10]) ? node11203 : node11200;
															assign node11200 = (inp[12]) ? 4'b0010 : 4'b0010;
															assign node11203 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node11206 = (inp[13]) ? node11210 : node11207;
															assign node11207 = (inp[12]) ? 4'b0110 : 4'b0011;
															assign node11210 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node11213 = (inp[9]) ? node11215 : 4'b0011;
														assign node11215 = (inp[13]) ? 4'b0010 : node11216;
															assign node11216 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node11220 = (inp[5]) ? node11232 : node11221;
													assign node11221 = (inp[10]) ? node11227 : node11222;
														assign node11222 = (inp[12]) ? 4'b0011 : node11223;
															assign node11223 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node11227 = (inp[12]) ? 4'b0110 : node11228;
															assign node11228 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node11232 = (inp[9]) ? node11236 : node11233;
														assign node11233 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node11236 = (inp[13]) ? 4'b0110 : 4'b0111;
										assign node11239 = (inp[15]) ? node11265 : node11240;
											assign node11240 = (inp[10]) ? node11254 : node11241;
												assign node11241 = (inp[5]) ? node11249 : node11242;
													assign node11242 = (inp[1]) ? 4'b0010 : node11243;
														assign node11243 = (inp[12]) ? node11245 : 4'b0010;
															assign node11245 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node11249 = (inp[1]) ? node11251 : 4'b0110;
														assign node11251 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node11254 = (inp[12]) ? node11260 : node11255;
													assign node11255 = (inp[5]) ? node11257 : 4'b0110;
														assign node11257 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node11260 = (inp[5]) ? node11262 : 4'b0111;
														assign node11262 = (inp[13]) ? 4'b0010 : 4'b0011;
											assign node11265 = (inp[10]) ? node11275 : node11266;
												assign node11266 = (inp[12]) ? node11272 : node11267;
													assign node11267 = (inp[1]) ? 4'b0110 : node11268;
														assign node11268 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node11272 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node11275 = (inp[9]) ? node11277 : 4'b0010;
													assign node11277 = (inp[5]) ? node11283 : node11278;
														assign node11278 = (inp[13]) ? 4'b0010 : node11279;
															assign node11279 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node11283 = (inp[13]) ? 4'b0110 : node11284;
															assign node11284 = (inp[12]) ? 4'b0010 : 4'b0010;
									assign node11288 = (inp[13]) ? node11346 : node11289;
										assign node11289 = (inp[12]) ? node11319 : node11290;
											assign node11290 = (inp[1]) ? node11304 : node11291;
												assign node11291 = (inp[5]) ? node11297 : node11292;
													assign node11292 = (inp[8]) ? 4'b0011 : node11293;
														assign node11293 = (inp[15]) ? 4'b0111 : 4'b0011;
													assign node11297 = (inp[15]) ? node11301 : node11298;
														assign node11298 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node11301 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node11304 = (inp[8]) ? node11312 : node11305;
													assign node11305 = (inp[10]) ? 4'b0011 : node11306;
														assign node11306 = (inp[15]) ? node11308 : 4'b0010;
															assign node11308 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node11312 = (inp[15]) ? node11316 : node11313;
														assign node11313 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node11316 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node11319 = (inp[15]) ? node11331 : node11320;
												assign node11320 = (inp[8]) ? node11328 : node11321;
													assign node11321 = (inp[1]) ? node11323 : 4'b0111;
														assign node11323 = (inp[10]) ? node11325 : 4'b0111;
															assign node11325 = (inp[5]) ? 4'b0110 : 4'b0110;
													assign node11328 = (inp[1]) ? 4'b0011 : 4'b0111;
												assign node11331 = (inp[5]) ? node11341 : node11332;
													assign node11332 = (inp[9]) ? node11334 : 4'b0110;
														assign node11334 = (inp[1]) ? node11338 : node11335;
															assign node11335 = (inp[8]) ? 4'b0110 : 4'b0010;
															assign node11338 = (inp[8]) ? 4'b0010 : 4'b0110;
													assign node11341 = (inp[8]) ? node11343 : 4'b0010;
														assign node11343 = (inp[1]) ? 4'b0011 : 4'b0111;
										assign node11346 = (inp[9]) ? node11370 : node11347;
											assign node11347 = (inp[8]) ? node11357 : node11348;
												assign node11348 = (inp[5]) ? node11350 : 4'b0011;
													assign node11350 = (inp[15]) ? node11352 : 4'b0110;
														assign node11352 = (inp[12]) ? node11354 : 4'b0011;
															assign node11354 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node11357 = (inp[12]) ? node11365 : node11358;
													assign node11358 = (inp[1]) ? 4'b0111 : node11359;
														assign node11359 = (inp[15]) ? node11361 : 4'b0011;
															assign node11361 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node11365 = (inp[1]) ? 4'b0011 : node11366;
														assign node11366 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node11370 = (inp[15]) ? node11384 : node11371;
												assign node11371 = (inp[8]) ? node11375 : node11372;
													assign node11372 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node11375 = (inp[10]) ? node11377 : 4'b0011;
														assign node11377 = (inp[12]) ? node11381 : node11378;
															assign node11378 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node11381 = (inp[1]) ? 4'b0011 : 4'b0110;
												assign node11384 = (inp[12]) ? 4'b0111 : node11385;
													assign node11385 = (inp[1]) ? 4'b0111 : 4'b0011;
								assign node11389 = (inp[0]) ? node11493 : node11390;
									assign node11390 = (inp[8]) ? node11466 : node11391;
										assign node11391 = (inp[1]) ? node11423 : node11392;
											assign node11392 = (inp[10]) ? node11404 : node11393;
												assign node11393 = (inp[13]) ? node11395 : 4'b0010;
													assign node11395 = (inp[5]) ? node11401 : node11396;
														assign node11396 = (inp[9]) ? 4'b0110 : node11397;
															assign node11397 = (inp[15]) ? 4'b0010 : 4'b0010;
														assign node11401 = (inp[15]) ? 4'b0110 : 4'b0111;
												assign node11404 = (inp[12]) ? node11414 : node11405;
													assign node11405 = (inp[13]) ? node11411 : node11406;
														assign node11406 = (inp[9]) ? 4'b0110 : node11407;
															assign node11407 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node11411 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node11414 = (inp[13]) ? node11418 : node11415;
														assign node11415 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node11418 = (inp[15]) ? node11420 : 4'b0011;
															assign node11420 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node11423 = (inp[5]) ? node11441 : node11424;
												assign node11424 = (inp[9]) ? node11428 : node11425;
													assign node11425 = (inp[13]) ? 4'b0011 : 4'b0110;
													assign node11428 = (inp[10]) ? node11436 : node11429;
														assign node11429 = (inp[13]) ? node11433 : node11430;
															assign node11430 = (inp[12]) ? 4'b0110 : 4'b0011;
															assign node11433 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node11436 = (inp[12]) ? 4'b0010 : node11437;
															assign node11437 = (inp[15]) ? 4'b0011 : 4'b0010;
												assign node11441 = (inp[9]) ? node11455 : node11442;
													assign node11442 = (inp[15]) ? node11448 : node11443;
														assign node11443 = (inp[13]) ? 4'b0010 : node11444;
															assign node11444 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node11448 = (inp[13]) ? node11452 : node11449;
															assign node11449 = (inp[10]) ? 4'b0111 : 4'b0011;
															assign node11452 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node11455 = (inp[15]) ? node11461 : node11456;
														assign node11456 = (inp[10]) ? node11458 : 4'b0011;
															assign node11458 = (inp[13]) ? 4'b0111 : 4'b0011;
														assign node11461 = (inp[13]) ? 4'b0111 : node11462;
															assign node11462 = (inp[10]) ? 4'b0110 : 4'b0010;
										assign node11466 = (inp[12]) ? node11484 : node11467;
											assign node11467 = (inp[1]) ? node11473 : node11468;
												assign node11468 = (inp[13]) ? node11470 : 4'b0011;
													assign node11470 = (inp[15]) ? 4'b0010 : 4'b0011;
												assign node11473 = (inp[13]) ? 4'b0111 : node11474;
													assign node11474 = (inp[9]) ? 4'b0110 : node11475;
														assign node11475 = (inp[15]) ? node11479 : node11476;
															assign node11476 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node11479 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node11484 = (inp[1]) ? 4'b0011 : node11485;
												assign node11485 = (inp[5]) ? 4'b0111 : node11486;
													assign node11486 = (inp[13]) ? node11488 : 4'b0111;
														assign node11488 = (inp[10]) ? 4'b0111 : 4'b0110;
									assign node11493 = (inp[9]) ? node11557 : node11494;
										assign node11494 = (inp[8]) ? node11526 : node11495;
											assign node11495 = (inp[12]) ? node11507 : node11496;
												assign node11496 = (inp[5]) ? node11502 : node11497;
													assign node11497 = (inp[15]) ? 4'b0111 : node11498;
														assign node11498 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node11502 = (inp[15]) ? 4'b0010 : node11503;
														assign node11503 = (inp[13]) ? 4'b0111 : 4'b0011;
												assign node11507 = (inp[13]) ? node11521 : node11508;
													assign node11508 = (inp[5]) ? node11516 : node11509;
														assign node11509 = (inp[15]) ? node11513 : node11510;
															assign node11510 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node11513 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node11516 = (inp[1]) ? node11518 : 4'b0111;
															assign node11518 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node11521 = (inp[1]) ? 4'b0011 : node11522;
														assign node11522 = (inp[15]) ? 4'b0111 : 4'b0010;
											assign node11526 = (inp[13]) ? node11544 : node11527;
												assign node11527 = (inp[5]) ? node11539 : node11528;
													assign node11528 = (inp[15]) ? node11532 : node11529;
														assign node11529 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node11532 = (inp[12]) ? node11536 : node11533;
															assign node11533 = (inp[1]) ? 4'b0111 : 4'b0010;
															assign node11536 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node11539 = (inp[15]) ? 4'b0110 : node11540;
														assign node11540 = (inp[10]) ? 4'b0111 : 4'b0011;
												assign node11544 = (inp[15]) ? node11552 : node11545;
													assign node11545 = (inp[1]) ? node11549 : node11546;
														assign node11546 = (inp[12]) ? 4'b0111 : 4'b0010;
														assign node11549 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node11552 = (inp[12]) ? node11554 : 4'b0110;
														assign node11554 = (inp[1]) ? 4'b0010 : 4'b0110;
										assign node11557 = (inp[12]) ? node11581 : node11558;
											assign node11558 = (inp[1]) ? node11572 : node11559;
												assign node11559 = (inp[8]) ? node11567 : node11560;
													assign node11560 = (inp[13]) ? node11564 : node11561;
														assign node11561 = (inp[15]) ? 4'b0110 : 4'b0010;
														assign node11564 = (inp[5]) ? 4'b0011 : 4'b0110;
													assign node11567 = (inp[13]) ? 4'b0010 : node11568;
														assign node11568 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node11572 = (inp[13]) ? 4'b0110 : node11573;
													assign node11573 = (inp[8]) ? node11577 : node11574;
														assign node11574 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node11577 = (inp[10]) ? 4'b0111 : 4'b0110;
											assign node11581 = (inp[1]) ? node11601 : node11582;
												assign node11582 = (inp[8]) ? node11592 : node11583;
													assign node11583 = (inp[5]) ? node11589 : node11584;
														assign node11584 = (inp[10]) ? node11586 : 4'b0011;
															assign node11586 = (inp[15]) ? 4'b0110 : 4'b0011;
														assign node11589 = (inp[10]) ? 4'b0011 : 4'b0110;
													assign node11592 = (inp[5]) ? 4'b0110 : node11593;
														assign node11593 = (inp[10]) ? node11597 : node11594;
															assign node11594 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node11597 = (inp[15]) ? 4'b0110 : 4'b0111;
												assign node11601 = (inp[13]) ? 4'b0010 : node11602;
													assign node11602 = (inp[5]) ? node11606 : node11603;
														assign node11603 = (inp[8]) ? 4'b0010 : 4'b0110;
														assign node11606 = (inp[8]) ? 4'b0011 : 4'b0111;
							assign node11610 = (inp[9]) ? node11854 : node11611;
								assign node11611 = (inp[2]) ? node11733 : node11612;
									assign node11612 = (inp[10]) ? node11674 : node11613;
										assign node11613 = (inp[1]) ? node11651 : node11614;
											assign node11614 = (inp[12]) ? node11632 : node11615;
												assign node11615 = (inp[8]) ? node11625 : node11616;
													assign node11616 = (inp[13]) ? node11622 : node11617;
														assign node11617 = (inp[15]) ? 4'b0110 : node11618;
															assign node11618 = (inp[5]) ? 4'b0010 : 4'b0010;
														assign node11622 = (inp[15]) ? 4'b0011 : 4'b0111;
													assign node11625 = (inp[13]) ? 4'b0010 : node11626;
														assign node11626 = (inp[0]) ? 4'b0011 : node11627;
															assign node11627 = (inp[15]) ? 4'b0010 : 4'b0011;
												assign node11632 = (inp[5]) ? node11644 : node11633;
													assign node11633 = (inp[8]) ? node11639 : node11634;
														assign node11634 = (inp[0]) ? node11636 : 4'b0011;
															assign node11636 = (inp[15]) ? 4'b0011 : 4'b0111;
														assign node11639 = (inp[0]) ? 4'b0111 : node11640;
															assign node11640 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node11644 = (inp[15]) ? node11648 : node11645;
														assign node11645 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node11648 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node11651 = (inp[12]) ? node11665 : node11652;
												assign node11652 = (inp[15]) ? node11658 : node11653;
													assign node11653 = (inp[8]) ? 4'b0110 : node11654;
														assign node11654 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node11658 = (inp[0]) ? 4'b0110 : node11659;
														assign node11659 = (inp[8]) ? node11661 : 4'b0111;
															assign node11661 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node11665 = (inp[15]) ? node11669 : node11666;
													assign node11666 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node11669 = (inp[13]) ? 4'b0010 : node11670;
														assign node11670 = (inp[8]) ? 4'b0010 : 4'b0110;
										assign node11674 = (inp[13]) ? node11706 : node11675;
											assign node11675 = (inp[8]) ? node11689 : node11676;
												assign node11676 = (inp[1]) ? node11686 : node11677;
													assign node11677 = (inp[15]) ? node11683 : node11678;
														assign node11678 = (inp[5]) ? 4'b0110 : node11679;
															assign node11679 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node11683 = (inp[12]) ? 4'b0011 : 4'b0110;
													assign node11686 = (inp[15]) ? 4'b0110 : 4'b0111;
												assign node11689 = (inp[5]) ? node11697 : node11690;
													assign node11690 = (inp[12]) ? 4'b0111 : node11691;
														assign node11691 = (inp[0]) ? 4'b0110 : node11692;
															assign node11692 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node11697 = (inp[12]) ? node11703 : node11698;
														assign node11698 = (inp[1]) ? 4'b0111 : node11699;
															assign node11699 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node11703 = (inp[1]) ? 4'b0010 : 4'b0111;
											assign node11706 = (inp[12]) ? node11722 : node11707;
												assign node11707 = (inp[1]) ? node11713 : node11708;
													assign node11708 = (inp[5]) ? node11710 : 4'b0110;
														assign node11710 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node11713 = (inp[15]) ? node11715 : 4'b0110;
														assign node11715 = (inp[8]) ? node11719 : node11716;
															assign node11716 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node11719 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node11722 = (inp[1]) ? node11728 : node11723;
													assign node11723 = (inp[8]) ? node11725 : 4'b0011;
														assign node11725 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node11728 = (inp[8]) ? node11730 : 4'b0010;
														assign node11730 = (inp[0]) ? 4'b0011 : 4'b0010;
									assign node11733 = (inp[0]) ? node11791 : node11734;
										assign node11734 = (inp[5]) ? node11762 : node11735;
											assign node11735 = (inp[12]) ? node11749 : node11736;
												assign node11736 = (inp[1]) ? node11744 : node11737;
													assign node11737 = (inp[8]) ? 4'b0011 : node11738;
														assign node11738 = (inp[13]) ? 4'b0111 : node11739;
															assign node11739 = (inp[15]) ? 4'b0111 : 4'b0011;
													assign node11744 = (inp[13]) ? 4'b0111 : node11745;
														assign node11745 = (inp[15]) ? 4'b0110 : 4'b0111;
												assign node11749 = (inp[1]) ? node11755 : node11750;
													assign node11750 = (inp[10]) ? node11752 : 4'b0111;
														assign node11752 = (inp[15]) ? 4'b0010 : 4'b0111;
													assign node11755 = (inp[15]) ? node11757 : 4'b0011;
														assign node11757 = (inp[8]) ? node11759 : 4'b0111;
															assign node11759 = (inp[13]) ? 4'b0011 : 4'b0010;
											assign node11762 = (inp[12]) ? node11776 : node11763;
												assign node11763 = (inp[1]) ? node11769 : node11764;
													assign node11764 = (inp[15]) ? 4'b0010 : node11765;
														assign node11765 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node11769 = (inp[13]) ? node11773 : node11770;
														assign node11770 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node11773 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node11776 = (inp[1]) ? node11784 : node11777;
													assign node11777 = (inp[8]) ? 4'b0111 : node11778;
														assign node11778 = (inp[15]) ? 4'b0110 : node11779;
															assign node11779 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node11784 = (inp[13]) ? 4'b0010 : node11785;
														assign node11785 = (inp[8]) ? node11787 : 4'b0111;
															assign node11787 = (inp[15]) ? 4'b0011 : 4'b0010;
										assign node11791 = (inp[8]) ? node11817 : node11792;
											assign node11792 = (inp[13]) ? node11806 : node11793;
												assign node11793 = (inp[12]) ? node11797 : node11794;
													assign node11794 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node11797 = (inp[5]) ? node11801 : node11798;
														assign node11798 = (inp[15]) ? 4'b0010 : 4'b0111;
														assign node11801 = (inp[15]) ? 4'b0111 : node11802;
															assign node11802 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node11806 = (inp[15]) ? node11812 : node11807;
													assign node11807 = (inp[1]) ? node11809 : 4'b0010;
														assign node11809 = (inp[5]) ? 4'b0011 : 4'b0111;
													assign node11812 = (inp[1]) ? 4'b0111 : node11813;
														assign node11813 = (inp[12]) ? 4'b0111 : 4'b0011;
											assign node11817 = (inp[10]) ? node11837 : node11818;
												assign node11818 = (inp[5]) ? node11828 : node11819;
													assign node11819 = (inp[13]) ? node11825 : node11820;
														assign node11820 = (inp[1]) ? node11822 : 4'b0010;
															assign node11822 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node11825 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node11828 = (inp[15]) ? node11830 : 4'b0110;
														assign node11830 = (inp[13]) ? node11834 : node11831;
															assign node11831 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node11834 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node11837 = (inp[13]) ? node11849 : node11838;
													assign node11838 = (inp[1]) ? node11842 : node11839;
														assign node11839 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node11842 = (inp[12]) ? node11846 : node11843;
															assign node11843 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node11846 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node11849 = (inp[1]) ? 4'b0010 : node11850;
														assign node11850 = (inp[15]) ? 4'b0011 : 4'b0010;
								assign node11854 = (inp[2]) ? node11964 : node11855;
									assign node11855 = (inp[0]) ? node11911 : node11856;
										assign node11856 = (inp[10]) ? node11888 : node11857;
											assign node11857 = (inp[12]) ? node11871 : node11858;
												assign node11858 = (inp[13]) ? node11868 : node11859;
													assign node11859 = (inp[1]) ? node11863 : node11860;
														assign node11860 = (inp[8]) ? 4'b0010 : 4'b0111;
														assign node11863 = (inp[8]) ? node11865 : 4'b0010;
															assign node11865 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node11868 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node11871 = (inp[1]) ? node11881 : node11872;
													assign node11872 = (inp[8]) ? node11878 : node11873;
														assign node11873 = (inp[13]) ? node11875 : 4'b0011;
															assign node11875 = (inp[15]) ? 4'b0110 : 4'b0010;
														assign node11878 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node11881 = (inp[8]) ? node11883 : 4'b0110;
														assign node11883 = (inp[15]) ? 4'b0010 : node11884;
															assign node11884 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node11888 = (inp[5]) ? node11900 : node11889;
												assign node11889 = (inp[8]) ? node11891 : 4'b0010;
													assign node11891 = (inp[15]) ? node11897 : node11892;
														assign node11892 = (inp[12]) ? node11894 : 4'b0010;
															assign node11894 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node11897 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node11900 = (inp[13]) ? node11908 : node11901;
													assign node11901 = (inp[8]) ? node11903 : 4'b0010;
														assign node11903 = (inp[12]) ? node11905 : 4'b0011;
															assign node11905 = (inp[1]) ? 4'b0011 : 4'b0110;
													assign node11908 = (inp[12]) ? 4'b0010 : 4'b0110;
										assign node11911 = (inp[15]) ? node11933 : node11912;
											assign node11912 = (inp[12]) ? node11916 : node11913;
												assign node11913 = (inp[13]) ? 4'b0111 : 4'b0011;
												assign node11916 = (inp[13]) ? node11926 : node11917;
													assign node11917 = (inp[10]) ? node11923 : node11918;
														assign node11918 = (inp[1]) ? node11920 : 4'b0111;
															assign node11920 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node11923 = (inp[8]) ? 4'b0010 : 4'b0110;
													assign node11926 = (inp[5]) ? node11930 : node11927;
														assign node11927 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node11930 = (inp[8]) ? 4'b0111 : 4'b0011;
											assign node11933 = (inp[8]) ? node11951 : node11934;
												assign node11934 = (inp[10]) ? node11946 : node11935;
													assign node11935 = (inp[1]) ? node11941 : node11936;
														assign node11936 = (inp[13]) ? node11938 : 4'b0111;
															assign node11938 = (inp[12]) ? 4'b0111 : 4'b0010;
														assign node11941 = (inp[12]) ? node11943 : 4'b0010;
															assign node11943 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node11946 = (inp[13]) ? 4'b0111 : node11947;
														assign node11947 = (inp[1]) ? 4'b0111 : 4'b0010;
												assign node11951 = (inp[5]) ? node11957 : node11952;
													assign node11952 = (inp[1]) ? node11954 : 4'b0011;
														assign node11954 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node11957 = (inp[12]) ? node11961 : node11958;
														assign node11958 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node11961 = (inp[1]) ? 4'b0011 : 4'b0111;
									assign node11964 = (inp[5]) ? node12002 : node11965;
										assign node11965 = (inp[13]) ? node11985 : node11966;
											assign node11966 = (inp[12]) ? node11974 : node11967;
												assign node11967 = (inp[8]) ? node11971 : node11968;
													assign node11968 = (inp[15]) ? 4'b0110 : 4'b0010;
													assign node11971 = (inp[1]) ? 4'b0110 : 4'b0011;
												assign node11974 = (inp[0]) ? node11978 : node11975;
													assign node11975 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node11978 = (inp[15]) ? node11980 : 4'b0010;
														assign node11980 = (inp[10]) ? 4'b0111 : node11981;
															assign node11981 = (inp[1]) ? 4'b0011 : 4'b0011;
											assign node11985 = (inp[12]) ? node11993 : node11986;
												assign node11986 = (inp[8]) ? 4'b0010 : node11987;
													assign node11987 = (inp[15]) ? node11989 : 4'b0110;
														assign node11989 = (inp[1]) ? 4'b0110 : 4'b0010;
												assign node11993 = (inp[1]) ? 4'b0010 : node11994;
													assign node11994 = (inp[15]) ? node11996 : 4'b0011;
														assign node11996 = (inp[0]) ? 4'b0110 : node11997;
															assign node11997 = (inp[8]) ? 4'b0111 : 4'b0110;
										assign node12002 = (inp[13]) ? node12026 : node12003;
											assign node12003 = (inp[12]) ? node12013 : node12004;
												assign node12004 = (inp[1]) ? node12006 : 4'b0010;
													assign node12006 = (inp[8]) ? node12008 : 4'b0010;
														assign node12008 = (inp[15]) ? 4'b0111 : node12009;
															assign node12009 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node12013 = (inp[8]) ? node12019 : node12014;
													assign node12014 = (inp[15]) ? 4'b0110 : node12015;
														assign node12015 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node12019 = (inp[1]) ? node12023 : node12020;
														assign node12020 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node12023 = (inp[15]) ? 4'b0011 : 4'b0010;
											assign node12026 = (inp[1]) ? node12046 : node12027;
												assign node12027 = (inp[10]) ? node12037 : node12028;
													assign node12028 = (inp[0]) ? 4'b0011 : node12029;
														assign node12029 = (inp[15]) ? node12033 : node12030;
															assign node12030 = (inp[12]) ? 4'b0010 : 4'b0011;
															assign node12033 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node12037 = (inp[8]) ? 4'b0010 : node12038;
														assign node12038 = (inp[0]) ? node12042 : node12039;
															assign node12039 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node12042 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node12046 = (inp[0]) ? 4'b0010 : 4'b0011;
					assign node12049 = (inp[8]) ? node12413 : node12050;
						assign node12050 = (inp[7]) ? node12304 : node12051;
							assign node12051 = (inp[0]) ? node12173 : node12052;
								assign node12052 = (inp[9]) ? node12114 : node12053;
									assign node12053 = (inp[5]) ? node12087 : node12054;
										assign node12054 = (inp[1]) ? node12064 : node12055;
											assign node12055 = (inp[15]) ? node12059 : node12056;
												assign node12056 = (inp[13]) ? 4'b0110 : 4'b0010;
												assign node12059 = (inp[13]) ? node12061 : 4'b0110;
													assign node12061 = (inp[12]) ? 4'b0010 : 4'b0011;
											assign node12064 = (inp[12]) ? node12080 : node12065;
												assign node12065 = (inp[10]) ? node12075 : node12066;
													assign node12066 = (inp[11]) ? node12072 : node12067;
														assign node12067 = (inp[13]) ? 4'b0110 : node12068;
															assign node12068 = (inp[15]) ? 4'b0110 : 4'b0010;
														assign node12072 = (inp[15]) ? 4'b0010 : 4'b0110;
													assign node12075 = (inp[15]) ? node12077 : 4'b0010;
														assign node12077 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node12080 = (inp[13]) ? node12084 : node12081;
													assign node12081 = (inp[15]) ? 4'b0110 : 4'b0011;
													assign node12084 = (inp[15]) ? 4'b0011 : 4'b0111;
										assign node12087 = (inp[13]) ? node12095 : node12088;
											assign node12088 = (inp[15]) ? 4'b0111 : node12089;
												assign node12089 = (inp[12]) ? node12091 : 4'b0011;
													assign node12091 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node12095 = (inp[15]) ? node12099 : node12096;
												assign node12096 = (inp[12]) ? 4'b0110 : 4'b0111;
												assign node12099 = (inp[10]) ? node12107 : node12100;
													assign node12100 = (inp[1]) ? node12104 : node12101;
														assign node12101 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node12104 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node12107 = (inp[2]) ? node12109 : 4'b0010;
														assign node12109 = (inp[12]) ? node12111 : 4'b0010;
															assign node12111 = (inp[1]) ? 4'b0010 : 4'b0011;
									assign node12114 = (inp[5]) ? node12150 : node12115;
										assign node12115 = (inp[12]) ? node12129 : node12116;
											assign node12116 = (inp[1]) ? node12124 : node12117;
												assign node12117 = (inp[13]) ? node12121 : node12118;
													assign node12118 = (inp[15]) ? 4'b0111 : 4'b0011;
													assign node12121 = (inp[15]) ? 4'b0010 : 4'b0111;
												assign node12124 = (inp[15]) ? node12126 : 4'b0111;
													assign node12126 = (inp[13]) ? 4'b0011 : 4'b0111;
											assign node12129 = (inp[1]) ? node12143 : node12130;
												assign node12130 = (inp[2]) ? node12132 : 4'b0111;
													assign node12132 = (inp[11]) ? node12138 : node12133;
														assign node12133 = (inp[15]) ? 4'b0111 : node12134;
															assign node12134 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node12138 = (inp[10]) ? 4'b0011 : node12139;
															assign node12139 = (inp[13]) ? 4'b0111 : 4'b0011;
												assign node12143 = (inp[15]) ? node12147 : node12144;
													assign node12144 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node12147 = (inp[13]) ? 4'b0010 : 4'b0111;
										assign node12150 = (inp[13]) ? node12158 : node12151;
											assign node12151 = (inp[15]) ? 4'b0110 : node12152;
												assign node12152 = (inp[12]) ? node12154 : 4'b0010;
													assign node12154 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node12158 = (inp[15]) ? node12164 : node12159;
												assign node12159 = (inp[1]) ? node12161 : 4'b0110;
													assign node12161 = (inp[12]) ? 4'b0111 : 4'b0110;
												assign node12164 = (inp[2]) ? node12166 : 4'b0011;
													assign node12166 = (inp[11]) ? node12168 : 4'b0010;
														assign node12168 = (inp[1]) ? 4'b0011 : node12169;
															assign node12169 = (inp[12]) ? 4'b0010 : 4'b0011;
								assign node12173 = (inp[9]) ? node12233 : node12174;
									assign node12174 = (inp[5]) ? node12198 : node12175;
										assign node12175 = (inp[13]) ? node12191 : node12176;
											assign node12176 = (inp[15]) ? node12182 : node12177;
												assign node12177 = (inp[12]) ? node12179 : 4'b0010;
													assign node12179 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node12182 = (inp[2]) ? node12184 : 4'b0111;
													assign node12184 = (inp[10]) ? 4'b0111 : node12185;
														assign node12185 = (inp[11]) ? 4'b0110 : node12186;
															assign node12186 = (inp[1]) ? 4'b0110 : 4'b0110;
											assign node12191 = (inp[15]) ? 4'b0010 : node12192;
												assign node12192 = (inp[12]) ? node12194 : 4'b0110;
													assign node12194 = (inp[1]) ? 4'b0110 : 4'b0111;
										assign node12198 = (inp[1]) ? node12220 : node12199;
											assign node12199 = (inp[12]) ? node12213 : node12200;
												assign node12200 = (inp[11]) ? node12206 : node12201;
													assign node12201 = (inp[13]) ? 4'b0011 : node12202;
														assign node12202 = (inp[15]) ? 4'b0111 : 4'b0011;
													assign node12206 = (inp[2]) ? node12208 : 4'b0011;
														assign node12208 = (inp[15]) ? 4'b0011 : node12209;
															assign node12209 = (inp[13]) ? 4'b0111 : 4'b0011;
												assign node12213 = (inp[15]) ? node12217 : node12214;
													assign node12214 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node12217 = (inp[13]) ? 4'b0011 : 4'b0110;
											assign node12220 = (inp[2]) ? node12226 : node12221;
												assign node12221 = (inp[15]) ? 4'b0011 : node12222;
													assign node12222 = (inp[13]) ? 4'b0111 : 4'b0011;
												assign node12226 = (inp[15]) ? node12230 : node12227;
													assign node12227 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node12230 = (inp[13]) ? 4'b0011 : 4'b0111;
									assign node12233 = (inp[5]) ? node12275 : node12234;
										assign node12234 = (inp[2]) ? node12258 : node12235;
											assign node12235 = (inp[13]) ? node12251 : node12236;
												assign node12236 = (inp[15]) ? node12240 : node12237;
													assign node12237 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node12240 = (inp[10]) ? node12246 : node12241;
														assign node12241 = (inp[1]) ? 4'b0110 : node12242;
															assign node12242 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node12246 = (inp[12]) ? node12248 : 4'b0111;
															assign node12248 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node12251 = (inp[15]) ? 4'b0011 : node12252;
													assign node12252 = (inp[12]) ? node12254 : 4'b0111;
														assign node12254 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node12258 = (inp[12]) ? node12266 : node12259;
												assign node12259 = (inp[11]) ? 4'b0011 : node12260;
													assign node12260 = (inp[15]) ? node12262 : 4'b0011;
														assign node12262 = (inp[1]) ? 4'b0110 : 4'b0011;
												assign node12266 = (inp[15]) ? node12272 : node12267;
													assign node12267 = (inp[1]) ? 4'b0111 : node12268;
														assign node12268 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node12272 = (inp[13]) ? 4'b0011 : 4'b0111;
										assign node12275 = (inp[13]) ? node12297 : node12276;
											assign node12276 = (inp[15]) ? node12280 : node12277;
												assign node12277 = (inp[12]) ? 4'b0011 : 4'b0010;
												assign node12280 = (inp[10]) ? node12290 : node12281;
													assign node12281 = (inp[2]) ? 4'b0111 : node12282;
														assign node12282 = (inp[12]) ? node12286 : node12283;
															assign node12283 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node12286 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node12290 = (inp[1]) ? node12294 : node12291;
														assign node12291 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node12294 = (inp[12]) ? 4'b0110 : 4'b0111;
											assign node12297 = (inp[15]) ? 4'b0010 : node12298;
												assign node12298 = (inp[1]) ? 4'b0110 : node12299;
													assign node12299 = (inp[10]) ? 4'b0111 : 4'b0110;
							assign node12304 = (inp[0]) ? node12362 : node12305;
								assign node12305 = (inp[9]) ? node12337 : node12306;
									assign node12306 = (inp[12]) ? node12326 : node12307;
										assign node12307 = (inp[15]) ? node12315 : node12308;
											assign node12308 = (inp[13]) ? node12312 : node12309;
												assign node12309 = (inp[1]) ? 4'b0100 : 4'b0000;
												assign node12312 = (inp[1]) ? 4'b0000 : 4'b0100;
											assign node12315 = (inp[2]) ? node12321 : node12316;
												assign node12316 = (inp[13]) ? node12318 : 4'b0000;
													assign node12318 = (inp[1]) ? 4'b0000 : 4'b0101;
												assign node12321 = (inp[13]) ? 4'b0000 : node12322;
													assign node12322 = (inp[1]) ? 4'b0101 : 4'b0000;
										assign node12326 = (inp[13]) ? node12332 : node12327;
											assign node12327 = (inp[1]) ? node12329 : 4'b0001;
												assign node12329 = (inp[15]) ? 4'b0101 : 4'b0100;
											assign node12332 = (inp[1]) ? 4'b0000 : node12333;
												assign node12333 = (inp[15]) ? 4'b0100 : 4'b0101;
									assign node12337 = (inp[1]) ? node12357 : node12338;
										assign node12338 = (inp[13]) ? node12342 : node12339;
											assign node12339 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node12342 = (inp[2]) ? node12352 : node12343;
												assign node12343 = (inp[11]) ? node12345 : 4'b0100;
													assign node12345 = (inp[15]) ? node12349 : node12346;
														assign node12346 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node12349 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node12352 = (inp[15]) ? node12354 : 4'b0101;
													assign node12354 = (inp[12]) ? 4'b0101 : 4'b0100;
										assign node12357 = (inp[13]) ? 4'b0001 : node12358;
											assign node12358 = (inp[15]) ? 4'b0100 : 4'b0101;
								assign node12362 = (inp[9]) ? node12386 : node12363;
									assign node12363 = (inp[15]) ? node12375 : node12364;
										assign node12364 = (inp[13]) ? node12370 : node12365;
											assign node12365 = (inp[1]) ? 4'b0100 : node12366;
												assign node12366 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node12370 = (inp[1]) ? 4'b0001 : node12371;
												assign node12371 = (inp[12]) ? 4'b0101 : 4'b0100;
										assign node12375 = (inp[1]) ? node12383 : node12376;
											assign node12376 = (inp[13]) ? node12380 : node12377;
												assign node12377 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node12380 = (inp[12]) ? 4'b0101 : 4'b0100;
											assign node12383 = (inp[13]) ? 4'b0001 : 4'b0101;
									assign node12386 = (inp[15]) ? node12402 : node12387;
										assign node12387 = (inp[12]) ? node12395 : node12388;
											assign node12388 = (inp[13]) ? node12392 : node12389;
												assign node12389 = (inp[1]) ? 4'b0101 : 4'b0001;
												assign node12392 = (inp[1]) ? 4'b0000 : 4'b0101;
											assign node12395 = (inp[1]) ? node12399 : node12396;
												assign node12396 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node12399 = (inp[13]) ? 4'b0000 : 4'b0101;
										assign node12402 = (inp[1]) ? node12410 : node12403;
											assign node12403 = (inp[13]) ? node12407 : node12404;
												assign node12404 = (inp[12]) ? 4'b0001 : 4'b0000;
												assign node12407 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node12410 = (inp[13]) ? 4'b0000 : 4'b0100;
						assign node12413 = (inp[1]) ? node12521 : node12414;
							assign node12414 = (inp[7]) ? node12498 : node12415;
								assign node12415 = (inp[15]) ? node12475 : node12416;
									assign node12416 = (inp[10]) ? node12440 : node12417;
										assign node12417 = (inp[0]) ? node12429 : node12418;
											assign node12418 = (inp[5]) ? node12424 : node12419;
												assign node12419 = (inp[12]) ? node12421 : 4'b0000;
													assign node12421 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node12424 = (inp[12]) ? node12426 : 4'b0001;
													assign node12426 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node12429 = (inp[5]) ? node12435 : node12430;
												assign node12430 = (inp[12]) ? node12432 : 4'b0001;
													assign node12432 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node12435 = (inp[12]) ? node12437 : 4'b0000;
													assign node12437 = (inp[13]) ? 4'b0001 : 4'b0000;
										assign node12440 = (inp[9]) ? node12460 : node12441;
											assign node12441 = (inp[12]) ? node12449 : node12442;
												assign node12442 = (inp[0]) ? node12446 : node12443;
													assign node12443 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node12446 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node12449 = (inp[13]) ? 4'b0001 : node12450;
													assign node12450 = (inp[2]) ? 4'b0001 : node12451;
														assign node12451 = (inp[5]) ? node12455 : node12452;
															assign node12452 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node12455 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node12460 = (inp[12]) ? node12468 : node12461;
												assign node12461 = (inp[5]) ? node12465 : node12462;
													assign node12462 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node12465 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node12468 = (inp[5]) ? node12470 : 4'b0000;
													assign node12470 = (inp[0]) ? 4'b0001 : node12471;
														assign node12471 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node12475 = (inp[0]) ? node12487 : node12476;
										assign node12476 = (inp[5]) ? node12482 : node12477;
											assign node12477 = (inp[13]) ? node12479 : 4'b0100;
												assign node12479 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node12482 = (inp[13]) ? node12484 : 4'b0101;
												assign node12484 = (inp[12]) ? 4'b0101 : 4'b0100;
										assign node12487 = (inp[5]) ? node12493 : node12488;
											assign node12488 = (inp[12]) ? 4'b0101 : node12489;
												assign node12489 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node12493 = (inp[13]) ? node12495 : 4'b0100;
												assign node12495 = (inp[12]) ? 4'b0100 : 4'b0101;
								assign node12498 = (inp[15]) ? node12514 : node12499;
									assign node12499 = (inp[10]) ? node12507 : node12500;
										assign node12500 = (inp[12]) ? node12504 : node12501;
											assign node12501 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node12504 = (inp[0]) ? 4'b0100 : 4'b0101;
										assign node12507 = (inp[12]) ? node12511 : node12508;
											assign node12508 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node12511 = (inp[0]) ? 4'b0100 : 4'b0101;
									assign node12514 = (inp[0]) ? node12518 : node12515;
										assign node12515 = (inp[12]) ? 4'b0101 : 4'b0100;
										assign node12518 = (inp[12]) ? 4'b0100 : 4'b0101;
							assign node12521 = (inp[15]) ? node12629 : node12522;
								assign node12522 = (inp[7]) ? node12622 : node12523;
									assign node12523 = (inp[2]) ? node12583 : node12524;
										assign node12524 = (inp[11]) ? node12550 : node12525;
											assign node12525 = (inp[9]) ? node12533 : node12526;
												assign node12526 = (inp[10]) ? node12528 : 4'b0101;
													assign node12528 = (inp[5]) ? 4'b0101 : node12529;
														assign node12529 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node12533 = (inp[0]) ? node12543 : node12534;
													assign node12534 = (inp[12]) ? node12536 : 4'b0101;
														assign node12536 = (inp[10]) ? node12540 : node12537;
															assign node12537 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node12540 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node12543 = (inp[12]) ? node12547 : node12544;
														assign node12544 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node12547 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node12550 = (inp[9]) ? node12564 : node12551;
												assign node12551 = (inp[10]) ? node12557 : node12552;
													assign node12552 = (inp[12]) ? node12554 : 4'b0100;
														assign node12554 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node12557 = (inp[12]) ? 4'b0100 : node12558;
														assign node12558 = (inp[0]) ? 4'b0101 : node12559;
															assign node12559 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node12564 = (inp[12]) ? node12576 : node12565;
													assign node12565 = (inp[13]) ? node12571 : node12566;
														assign node12566 = (inp[10]) ? node12568 : 4'b0100;
															assign node12568 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node12571 = (inp[0]) ? 4'b0101 : node12572;
															assign node12572 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node12576 = (inp[5]) ? node12578 : 4'b0101;
														assign node12578 = (inp[13]) ? node12580 : 4'b0101;
															assign node12580 = (inp[0]) ? 4'b0100 : 4'b0101;
										assign node12583 = (inp[11]) ? node12603 : node12584;
											assign node12584 = (inp[0]) ? node12596 : node12585;
												assign node12585 = (inp[9]) ? node12591 : node12586;
													assign node12586 = (inp[5]) ? 4'b0100 : node12587;
														assign node12587 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node12591 = (inp[12]) ? 4'b0101 : node12592;
														assign node12592 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node12596 = (inp[5]) ? 4'b0100 : node12597;
													assign node12597 = (inp[13]) ? 4'b0101 : node12598;
														assign node12598 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node12603 = (inp[9]) ? node12613 : node12604;
												assign node12604 = (inp[0]) ? node12606 : 4'b0101;
													assign node12606 = (inp[5]) ? node12610 : node12607;
														assign node12607 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node12610 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node12613 = (inp[12]) ? node12615 : 4'b0101;
													assign node12615 = (inp[10]) ? 4'b0101 : node12616;
														assign node12616 = (inp[13]) ? node12618 : 4'b0100;
															assign node12618 = (inp[5]) ? 4'b0101 : 4'b0100;
									assign node12622 = (inp[0]) ? node12626 : node12623;
										assign node12623 = (inp[13]) ? 4'b0001 : 4'b0000;
										assign node12626 = (inp[13]) ? 4'b0000 : 4'b0001;
								assign node12629 = (inp[0]) ? node12643 : node12630;
									assign node12630 = (inp[7]) ? 4'b0001 : node12631;
										assign node12631 = (inp[5]) ? node12637 : node12632;
											assign node12632 = (inp[12]) ? 4'b0000 : node12633;
												assign node12633 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node12637 = (inp[13]) ? 4'b0001 : node12638;
												assign node12638 = (inp[12]) ? 4'b0001 : 4'b0000;
									assign node12643 = (inp[7]) ? 4'b0000 : node12644;
										assign node12644 = (inp[5]) ? node12650 : node12645;
											assign node12645 = (inp[13]) ? 4'b0001 : node12646;
												assign node12646 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node12650 = (inp[13]) ? 4'b0000 : node12651;
												assign node12651 = (inp[12]) ? 4'b0000 : 4'b0001;
		assign node12656 = (inp[8]) ? node19402 : node12657;
			assign node12657 = (inp[14]) ? node16315 : node12658;
				assign node12658 = (inp[7]) ? node14472 : node12659;
					assign node12659 = (inp[15]) ? node13549 : node12660;
						assign node12660 = (inp[6]) ? node13090 : node12661;
							assign node12661 = (inp[2]) ? node12865 : node12662;
								assign node12662 = (inp[13]) ? node12760 : node12663;
									assign node12663 = (inp[1]) ? node12715 : node12664;
										assign node12664 = (inp[4]) ? node12694 : node12665;
											assign node12665 = (inp[12]) ? node12683 : node12666;
												assign node12666 = (inp[9]) ? node12674 : node12667;
													assign node12667 = (inp[11]) ? 4'b1001 : node12668;
														assign node12668 = (inp[0]) ? node12670 : 4'b1001;
															assign node12670 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node12674 = (inp[0]) ? node12676 : 4'b1000;
														assign node12676 = (inp[10]) ? node12680 : node12677;
															assign node12677 = (inp[5]) ? 4'b1000 : 4'b1001;
															assign node12680 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node12683 = (inp[0]) ? node12689 : node12684;
													assign node12684 = (inp[10]) ? 4'b1010 : node12685;
														assign node12685 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node12689 = (inp[10]) ? 4'b1011 : node12690;
														assign node12690 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node12694 = (inp[12]) ? node12706 : node12695;
												assign node12695 = (inp[10]) ? node12703 : node12696;
													assign node12696 = (inp[9]) ? 4'b1011 : node12697;
														assign node12697 = (inp[5]) ? node12699 : 4'b1010;
															assign node12699 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node12703 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node12706 = (inp[5]) ? node12712 : node12707;
													assign node12707 = (inp[0]) ? 4'b1100 : node12708;
														assign node12708 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node12712 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node12715 = (inp[5]) ? node12743 : node12716;
											assign node12716 = (inp[10]) ? node12730 : node12717;
												assign node12717 = (inp[9]) ? node12723 : node12718;
													assign node12718 = (inp[12]) ? node12720 : 4'b1100;
														assign node12720 = (inp[4]) ? 4'b1101 : 4'b1111;
													assign node12723 = (inp[12]) ? node12727 : node12724;
														assign node12724 = (inp[4]) ? 4'b1111 : 4'b1101;
														assign node12727 = (inp[4]) ? 4'b1100 : 4'b1110;
												assign node12730 = (inp[11]) ? node12736 : node12731;
													assign node12731 = (inp[0]) ? 4'b1101 : node12732;
														assign node12732 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node12736 = (inp[9]) ? node12738 : 4'b1101;
														assign node12738 = (inp[12]) ? node12740 : 4'b1110;
															assign node12740 = (inp[4]) ? 4'b1101 : 4'b1111;
											assign node12743 = (inp[12]) ? node12749 : node12744;
												assign node12744 = (inp[4]) ? 4'b1011 : node12745;
													assign node12745 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node12749 = (inp[4]) ? node12751 : 4'b1010;
													assign node12751 = (inp[0]) ? node12757 : node12752;
														assign node12752 = (inp[11]) ? 4'b1101 : node12753;
															assign node12753 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node12757 = (inp[10]) ? 4'b1101 : 4'b1100;
									assign node12760 = (inp[5]) ? node12812 : node12761;
										assign node12761 = (inp[1]) ? node12785 : node12762;
											assign node12762 = (inp[12]) ? node12774 : node12763;
												assign node12763 = (inp[4]) ? node12769 : node12764;
													assign node12764 = (inp[9]) ? node12766 : 4'b1101;
														assign node12766 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node12769 = (inp[0]) ? 4'b1111 : node12770;
														assign node12770 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node12774 = (inp[4]) ? node12778 : node12775;
													assign node12775 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node12778 = (inp[0]) ? node12780 : 4'b1001;
														assign node12780 = (inp[10]) ? node12782 : 4'b1000;
															assign node12782 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node12785 = (inp[12]) ? node12799 : node12786;
												assign node12786 = (inp[4]) ? node12792 : node12787;
													assign node12787 = (inp[11]) ? 4'b1001 : node12788;
														assign node12788 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node12792 = (inp[10]) ? 4'b1011 : node12793;
														assign node12793 = (inp[0]) ? node12795 : 4'b1010;
															assign node12795 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node12799 = (inp[4]) ? node12803 : node12800;
													assign node12800 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node12803 = (inp[9]) ? 4'b1000 : node12804;
														assign node12804 = (inp[0]) ? node12808 : node12805;
															assign node12805 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node12808 = (inp[10]) ? 4'b1001 : 4'b1000;
										assign node12812 = (inp[12]) ? node12840 : node12813;
											assign node12813 = (inp[4]) ? node12827 : node12814;
												assign node12814 = (inp[10]) ? node12822 : node12815;
													assign node12815 = (inp[0]) ? 4'b1100 : node12816;
														assign node12816 = (inp[11]) ? node12818 : 4'b1100;
															assign node12818 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node12822 = (inp[9]) ? 4'b1101 : node12823;
														assign node12823 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node12827 = (inp[0]) ? node12833 : node12828;
													assign node12828 = (inp[1]) ? 4'b1110 : node12829;
														assign node12829 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node12833 = (inp[10]) ? 4'b1111 : node12834;
														assign node12834 = (inp[9]) ? node12836 : 4'b1111;
															assign node12836 = (inp[1]) ? 4'b1110 : 4'b1111;
											assign node12840 = (inp[4]) ? node12848 : node12841;
												assign node12841 = (inp[11]) ? 4'b1110 : node12842;
													assign node12842 = (inp[1]) ? node12844 : 4'b1111;
														assign node12844 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node12848 = (inp[1]) ? node12856 : node12849;
													assign node12849 = (inp[9]) ? node12851 : 4'b1101;
														assign node12851 = (inp[11]) ? 4'b1101 : node12852;
															assign node12852 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node12856 = (inp[9]) ? 4'b1001 : node12857;
														assign node12857 = (inp[10]) ? node12861 : node12858;
															assign node12858 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node12861 = (inp[0]) ? 4'b1001 : 4'b1000;
								assign node12865 = (inp[13]) ? node12963 : node12866;
									assign node12866 = (inp[1]) ? node12920 : node12867;
										assign node12867 = (inp[12]) ? node12895 : node12868;
											assign node12868 = (inp[4]) ? node12876 : node12869;
												assign node12869 = (inp[11]) ? node12871 : 4'b1101;
													assign node12871 = (inp[10]) ? node12873 : 4'b1100;
														assign node12873 = (inp[5]) ? 4'b1101 : 4'b1100;
												assign node12876 = (inp[0]) ? node12890 : node12877;
													assign node12877 = (inp[10]) ? node12885 : node12878;
														assign node12878 = (inp[11]) ? node12882 : node12879;
															assign node12879 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node12882 = (inp[9]) ? 4'b1110 : 4'b1110;
														assign node12885 = (inp[9]) ? 4'b1111 : node12886;
															assign node12886 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node12890 = (inp[10]) ? node12892 : 4'b1111;
														assign node12892 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node12895 = (inp[4]) ? node12905 : node12896;
												assign node12896 = (inp[0]) ? 4'b1111 : node12897;
													assign node12897 = (inp[5]) ? node12899 : 4'b1111;
														assign node12899 = (inp[10]) ? 4'b1110 : node12900;
															assign node12900 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node12905 = (inp[5]) ? node12913 : node12906;
													assign node12906 = (inp[11]) ? 4'b1000 : node12907;
														assign node12907 = (inp[9]) ? 4'b1000 : node12908;
															assign node12908 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node12913 = (inp[11]) ? node12915 : 4'b1100;
														assign node12915 = (inp[9]) ? 4'b1101 : node12916;
															assign node12916 = (inp[10]) ? 4'b1101 : 4'b1100;
										assign node12920 = (inp[5]) ? node12946 : node12921;
											assign node12921 = (inp[9]) ? node12935 : node12922;
												assign node12922 = (inp[11]) ? node12926 : node12923;
													assign node12923 = (inp[10]) ? 4'b1001 : 4'b1011;
													assign node12926 = (inp[10]) ? node12928 : 4'b1001;
														assign node12928 = (inp[12]) ? node12932 : node12929;
															assign node12929 = (inp[4]) ? 4'b1011 : 4'b1000;
															assign node12932 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node12935 = (inp[0]) ? node12943 : node12936;
													assign node12936 = (inp[10]) ? node12940 : node12937;
														assign node12937 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node12940 = (inp[12]) ? 4'b1010 : 4'b1000;
													assign node12943 = (inp[10]) ? 4'b1011 : 4'b1010;
											assign node12946 = (inp[4]) ? node12956 : node12947;
												assign node12947 = (inp[12]) ? 4'b1111 : node12948;
													assign node12948 = (inp[11]) ? node12950 : 4'b1100;
														assign node12950 = (inp[0]) ? 4'b1100 : node12951;
															assign node12951 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node12956 = (inp[12]) ? node12958 : 4'b1111;
													assign node12958 = (inp[11]) ? node12960 : 4'b1000;
														assign node12960 = (inp[10]) ? 4'b1001 : 4'b1000;
									assign node12963 = (inp[5]) ? node13031 : node12964;
										assign node12964 = (inp[1]) ? node12992 : node12965;
											assign node12965 = (inp[4]) ? node12981 : node12966;
												assign node12966 = (inp[12]) ? node12974 : node12967;
													assign node12967 = (inp[10]) ? node12969 : 4'b1000;
														assign node12969 = (inp[9]) ? 4'b1001 : node12970;
															assign node12970 = (inp[0]) ? 4'b1000 : 4'b1000;
													assign node12974 = (inp[10]) ? 4'b1010 : node12975;
														assign node12975 = (inp[0]) ? node12977 : 4'b1011;
															assign node12977 = (inp[9]) ? 4'b1010 : 4'b1010;
												assign node12981 = (inp[12]) ? node12985 : node12982;
													assign node12982 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node12985 = (inp[0]) ? node12987 : 4'b1100;
														assign node12987 = (inp[10]) ? node12989 : 4'b1101;
															assign node12989 = (inp[9]) ? 4'b1101 : 4'b1100;
											assign node12992 = (inp[9]) ? node13014 : node12993;
												assign node12993 = (inp[11]) ? node13005 : node12994;
													assign node12994 = (inp[4]) ? node12998 : node12995;
														assign node12995 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node12998 = (inp[10]) ? node13002 : node12999;
															assign node12999 = (inp[12]) ? 4'b1101 : 4'b1111;
															assign node13002 = (inp[12]) ? 4'b1100 : 4'b1110;
													assign node13005 = (inp[10]) ? node13007 : 4'b1110;
														assign node13007 = (inp[12]) ? node13011 : node13008;
															assign node13008 = (inp[4]) ? 4'b1111 : 4'b1100;
															assign node13011 = (inp[0]) ? 4'b1100 : 4'b1111;
												assign node13014 = (inp[10]) ? node13026 : node13015;
													assign node13015 = (inp[0]) ? node13023 : node13016;
														assign node13016 = (inp[12]) ? node13020 : node13017;
															assign node13017 = (inp[4]) ? 4'b1111 : 4'b1100;
															assign node13020 = (inp[4]) ? 4'b1101 : 4'b1111;
														assign node13023 = (inp[4]) ? 4'b1100 : 4'b1110;
													assign node13026 = (inp[0]) ? node13028 : 4'b1110;
														assign node13028 = (inp[11]) ? 4'b1110 : 4'b1111;
										assign node13031 = (inp[11]) ? node13057 : node13032;
											assign node13032 = (inp[12]) ? node13050 : node13033;
												assign node13033 = (inp[4]) ? node13045 : node13034;
													assign node13034 = (inp[1]) ? node13040 : node13035;
														assign node13035 = (inp[9]) ? node13037 : 4'b1001;
															assign node13037 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node13040 = (inp[0]) ? node13042 : 4'b1000;
															assign node13042 = (inp[10]) ? 4'b1000 : 4'b1000;
													assign node13045 = (inp[1]) ? 4'b1011 : node13046;
														assign node13046 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node13050 = (inp[4]) ? node13052 : 4'b1010;
													assign node13052 = (inp[1]) ? node13054 : 4'b1000;
														assign node13054 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node13057 = (inp[10]) ? node13073 : node13058;
												assign node13058 = (inp[9]) ? node13064 : node13059;
													assign node13059 = (inp[4]) ? node13061 : 4'b1011;
														assign node13061 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node13064 = (inp[0]) ? node13066 : 4'b1010;
														assign node13066 = (inp[1]) ? node13070 : node13067;
															assign node13067 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node13070 = (inp[4]) ? 4'b1010 : 4'b1011;
												assign node13073 = (inp[0]) ? node13079 : node13074;
													assign node13074 = (inp[1]) ? node13076 : 4'b1011;
														assign node13076 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node13079 = (inp[1]) ? node13083 : node13080;
														assign node13080 = (inp[9]) ? 4'b1011 : 4'b1000;
														assign node13083 = (inp[12]) ? node13087 : node13084;
															assign node13084 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node13087 = (inp[9]) ? 4'b1010 : 4'b1011;
							assign node13090 = (inp[1]) ? node13296 : node13091;
								assign node13091 = (inp[2]) ? node13179 : node13092;
									assign node13092 = (inp[11]) ? node13130 : node13093;
										assign node13093 = (inp[5]) ? node13111 : node13094;
											assign node13094 = (inp[13]) ? node13106 : node13095;
												assign node13095 = (inp[12]) ? node13101 : node13096;
													assign node13096 = (inp[10]) ? 4'b1000 : node13097;
														assign node13097 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node13101 = (inp[9]) ? 4'b1001 : node13102;
														assign node13102 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node13106 = (inp[9]) ? 4'b1101 : node13107;
													assign node13107 = (inp[12]) ? 4'b1101 : 4'b1100;
											assign node13111 = (inp[13]) ? node13117 : node13112;
												assign node13112 = (inp[12]) ? 4'b1101 : node13113;
													assign node13113 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node13117 = (inp[4]) ? node13123 : node13118;
													assign node13118 = (inp[0]) ? node13120 : 4'b1001;
														assign node13120 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node13123 = (inp[9]) ? 4'b1000 : node13124;
														assign node13124 = (inp[12]) ? node13126 : 4'b1001;
															assign node13126 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node13130 = (inp[12]) ? node13158 : node13131;
											assign node13131 = (inp[9]) ? node13151 : node13132;
												assign node13132 = (inp[4]) ? node13144 : node13133;
													assign node13133 = (inp[0]) ? node13141 : node13134;
														assign node13134 = (inp[13]) ? node13138 : node13135;
															assign node13135 = (inp[5]) ? 4'b1101 : 4'b1001;
															assign node13138 = (inp[5]) ? 4'b1000 : 4'b1101;
														assign node13141 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node13144 = (inp[0]) ? node13146 : 4'b1000;
														assign node13146 = (inp[5]) ? 4'b1101 : node13147;
															assign node13147 = (inp[13]) ? 4'b1101 : 4'b1000;
												assign node13151 = (inp[5]) ? 4'b1001 : node13152;
													assign node13152 = (inp[13]) ? 4'b1100 : node13153;
														assign node13153 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node13158 = (inp[13]) ? node13172 : node13159;
												assign node13159 = (inp[5]) ? node13169 : node13160;
													assign node13160 = (inp[4]) ? 4'b1000 : node13161;
														assign node13161 = (inp[10]) ? node13165 : node13162;
															assign node13162 = (inp[0]) ? 4'b1000 : 4'b1000;
															assign node13165 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node13169 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node13172 = (inp[5]) ? node13176 : node13173;
													assign node13173 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node13176 = (inp[0]) ? 4'b1001 : 4'b1000;
									assign node13179 = (inp[10]) ? node13233 : node13180;
										assign node13180 = (inp[11]) ? node13206 : node13181;
											assign node13181 = (inp[5]) ? node13195 : node13182;
												assign node13182 = (inp[13]) ? node13184 : 4'b1000;
													assign node13184 = (inp[12]) ? node13190 : node13185;
														assign node13185 = (inp[9]) ? 4'b1100 : node13186;
															assign node13186 = (inp[4]) ? 4'b1100 : 4'b1100;
														assign node13190 = (inp[9]) ? node13192 : 4'b1100;
															assign node13192 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node13195 = (inp[13]) ? node13199 : node13196;
													assign node13196 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node13199 = (inp[9]) ? 4'b1000 : node13200;
														assign node13200 = (inp[12]) ? 4'b1001 : node13201;
															assign node13201 = (inp[4]) ? 4'b1000 : 4'b1001;
											assign node13206 = (inp[12]) ? node13218 : node13207;
												assign node13207 = (inp[0]) ? node13211 : node13208;
													assign node13208 = (inp[5]) ? 4'b1001 : 4'b1101;
													assign node13211 = (inp[4]) ? 4'b1101 : node13212;
														assign node13212 = (inp[13]) ? 4'b1000 : node13213;
															assign node13213 = (inp[5]) ? 4'b1101 : 4'b1000;
												assign node13218 = (inp[9]) ? node13228 : node13219;
													assign node13219 = (inp[13]) ? node13223 : node13220;
														assign node13220 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node13223 = (inp[4]) ? 4'b1101 : node13224;
															assign node13224 = (inp[5]) ? 4'b1000 : 4'b1100;
													assign node13228 = (inp[13]) ? 4'b1001 : node13229;
														assign node13229 = (inp[5]) ? 4'b1100 : 4'b1000;
										assign node13233 = (inp[0]) ? node13271 : node13234;
											assign node13234 = (inp[13]) ? node13254 : node13235;
												assign node13235 = (inp[5]) ? node13243 : node13236;
													assign node13236 = (inp[4]) ? 4'b1001 : node13237;
														assign node13237 = (inp[11]) ? node13239 : 4'b1000;
															assign node13239 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node13243 = (inp[12]) ? node13249 : node13244;
														assign node13244 = (inp[11]) ? 4'b1100 : node13245;
															assign node13245 = (inp[4]) ? 4'b1100 : 4'b1101;
														assign node13249 = (inp[4]) ? node13251 : 4'b1101;
															assign node13251 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node13254 = (inp[5]) ? node13264 : node13255;
													assign node13255 = (inp[11]) ? 4'b1101 : node13256;
														assign node13256 = (inp[12]) ? node13260 : node13257;
															assign node13257 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node13260 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node13264 = (inp[12]) ? node13266 : 4'b1001;
														assign node13266 = (inp[4]) ? node13268 : 4'b1001;
															assign node13268 = (inp[9]) ? 4'b1000 : 4'b1000;
											assign node13271 = (inp[12]) ? node13281 : node13272;
												assign node13272 = (inp[11]) ? node13278 : node13273;
													assign node13273 = (inp[13]) ? node13275 : 4'b1101;
														assign node13275 = (inp[5]) ? 4'b1001 : 4'b1101;
													assign node13278 = (inp[4]) ? 4'b1000 : 4'b1101;
												assign node13281 = (inp[4]) ? node13289 : node13282;
													assign node13282 = (inp[11]) ? node13284 : 4'b1000;
														assign node13284 = (inp[5]) ? node13286 : 4'b1100;
															assign node13286 = (inp[13]) ? 4'b1001 : 4'b1100;
													assign node13289 = (inp[13]) ? 4'b1000 : node13290;
														assign node13290 = (inp[5]) ? 4'b1101 : node13291;
															assign node13291 = (inp[11]) ? 4'b1000 : 4'b1001;
								assign node13296 = (inp[9]) ? node13406 : node13297;
									assign node13297 = (inp[0]) ? node13347 : node13298;
										assign node13298 = (inp[13]) ? node13332 : node13299;
											assign node13299 = (inp[12]) ? node13319 : node13300;
												assign node13300 = (inp[2]) ? node13310 : node13301;
													assign node13301 = (inp[11]) ? node13305 : node13302;
														assign node13302 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node13305 = (inp[4]) ? node13307 : 4'b1001;
															assign node13307 = (inp[5]) ? 4'b1100 : 4'b1001;
													assign node13310 = (inp[5]) ? node13316 : node13311;
														assign node13311 = (inp[4]) ? node13313 : 4'b1100;
															assign node13313 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node13316 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node13319 = (inp[5]) ? node13325 : node13320;
													assign node13320 = (inp[10]) ? node13322 : 4'b1001;
														assign node13322 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node13325 = (inp[2]) ? node13329 : node13326;
														assign node13326 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node13329 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node13332 = (inp[5]) ? node13340 : node13333;
												assign node13333 = (inp[11]) ? node13335 : 4'b1100;
													assign node13335 = (inp[12]) ? node13337 : 4'b1101;
														assign node13337 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node13340 = (inp[11]) ? 4'b1100 : node13341;
													assign node13341 = (inp[4]) ? node13343 : 4'b1101;
														assign node13343 = (inp[2]) ? 4'b1100 : 4'b1101;
										assign node13347 = (inp[11]) ? node13377 : node13348;
											assign node13348 = (inp[12]) ? node13360 : node13349;
												assign node13349 = (inp[10]) ? node13355 : node13350;
													assign node13350 = (inp[4]) ? 4'b1001 : node13351;
														assign node13351 = (inp[5]) ? 4'b1101 : 4'b1001;
													assign node13355 = (inp[5]) ? 4'b1000 : node13356;
														assign node13356 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node13360 = (inp[2]) ? node13368 : node13361;
													assign node13361 = (inp[13]) ? 4'b1101 : node13362;
														assign node13362 = (inp[10]) ? 4'b1101 : node13363;
															assign node13363 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node13368 = (inp[10]) ? node13374 : node13369;
														assign node13369 = (inp[4]) ? 4'b1100 : node13370;
															assign node13370 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node13374 = (inp[4]) ? 4'b1001 : 4'b1000;
											assign node13377 = (inp[5]) ? node13387 : node13378;
												assign node13378 = (inp[13]) ? node13382 : node13379;
													assign node13379 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node13382 = (inp[12]) ? node13384 : 4'b1101;
														assign node13384 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node13387 = (inp[10]) ? node13397 : node13388;
													assign node13388 = (inp[12]) ? node13394 : node13389;
														assign node13389 = (inp[13]) ? node13391 : 4'b1001;
															assign node13391 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node13394 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node13397 = (inp[13]) ? node13401 : node13398;
														assign node13398 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node13401 = (inp[4]) ? 4'b1101 : node13402;
															assign node13402 = (inp[12]) ? 4'b1001 : 4'b1101;
									assign node13406 = (inp[10]) ? node13490 : node13407;
										assign node13407 = (inp[13]) ? node13449 : node13408;
											assign node13408 = (inp[2]) ? node13424 : node13409;
												assign node13409 = (inp[12]) ? node13413 : node13410;
													assign node13410 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node13413 = (inp[11]) ? node13419 : node13414;
														assign node13414 = (inp[4]) ? 4'b1001 : node13415;
															assign node13415 = (inp[0]) ? 4'b1000 : 4'b1100;
														assign node13419 = (inp[5]) ? 4'b1101 : node13420;
															assign node13420 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node13424 = (inp[11]) ? node13436 : node13425;
													assign node13425 = (inp[12]) ? node13433 : node13426;
														assign node13426 = (inp[5]) ? node13430 : node13427;
															assign node13427 = (inp[4]) ? 4'b1000 : 4'b1101;
															assign node13430 = (inp[4]) ? 4'b1101 : 4'b1000;
														assign node13433 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node13436 = (inp[0]) ? node13444 : node13437;
														assign node13437 = (inp[5]) ? node13441 : node13438;
															assign node13438 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node13441 = (inp[12]) ? 4'b1000 : 4'b1001;
														assign node13444 = (inp[5]) ? node13446 : 4'b1001;
															assign node13446 = (inp[12]) ? 4'b1001 : 4'b1100;
											assign node13449 = (inp[0]) ? node13467 : node13450;
												assign node13450 = (inp[5]) ? node13460 : node13451;
													assign node13451 = (inp[11]) ? node13455 : node13452;
														assign node13452 = (inp[12]) ? 4'b1001 : 4'b1000;
														assign node13455 = (inp[2]) ? 4'b1100 : node13456;
															assign node13456 = (inp[12]) ? 4'b1000 : 4'b1001;
													assign node13460 = (inp[11]) ? node13464 : node13461;
														assign node13461 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node13464 = (inp[12]) ? 4'b1100 : 4'b1000;
												assign node13467 = (inp[11]) ? node13479 : node13468;
													assign node13468 = (inp[4]) ? node13474 : node13469;
														assign node13469 = (inp[12]) ? node13471 : 4'b1100;
															assign node13471 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node13474 = (inp[2]) ? node13476 : 4'b1101;
															assign node13476 = (inp[12]) ? 4'b1000 : 4'b1101;
													assign node13479 = (inp[2]) ? node13483 : node13480;
														assign node13480 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node13483 = (inp[12]) ? node13487 : node13484;
															assign node13484 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node13487 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node13490 = (inp[12]) ? node13520 : node13491;
											assign node13491 = (inp[5]) ? node13501 : node13492;
												assign node13492 = (inp[13]) ? node13498 : node13493;
													assign node13493 = (inp[4]) ? 4'b1001 : node13494;
														assign node13494 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node13498 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node13501 = (inp[11]) ? node13509 : node13502;
													assign node13502 = (inp[4]) ? node13506 : node13503;
														assign node13503 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node13506 = (inp[13]) ? 4'b1000 : 4'b1101;
													assign node13509 = (inp[13]) ? node13515 : node13510;
														assign node13510 = (inp[4]) ? node13512 : 4'b1000;
															assign node13512 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node13515 = (inp[4]) ? 4'b1001 : node13516;
															assign node13516 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node13520 = (inp[2]) ? node13546 : node13521;
												assign node13521 = (inp[0]) ? node13535 : node13522;
													assign node13522 = (inp[13]) ? node13530 : node13523;
														assign node13523 = (inp[5]) ? node13527 : node13524;
															assign node13524 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node13527 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node13530 = (inp[5]) ? node13532 : 4'b1101;
															assign node13532 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node13535 = (inp[4]) ? node13541 : node13536;
														assign node13536 = (inp[5]) ? node13538 : 4'b1101;
															assign node13538 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node13541 = (inp[11]) ? 4'b1101 : node13542;
															assign node13542 = (inp[13]) ? 4'b1101 : 4'b1100;
												assign node13546 = (inp[4]) ? 4'b1000 : 4'b1100;
						assign node13549 = (inp[6]) ? node14009 : node13550;
							assign node13550 = (inp[12]) ? node13760 : node13551;
								assign node13551 = (inp[4]) ? node13661 : node13552;
									assign node13552 = (inp[13]) ? node13602 : node13553;
										assign node13553 = (inp[2]) ? node13581 : node13554;
											assign node13554 = (inp[1]) ? node13570 : node13555;
												assign node13555 = (inp[11]) ? node13563 : node13556;
													assign node13556 = (inp[9]) ? 4'b1001 : node13557;
														assign node13557 = (inp[0]) ? node13559 : 4'b1000;
															assign node13559 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node13563 = (inp[0]) ? 4'b1000 : node13564;
														assign node13564 = (inp[5]) ? node13566 : 4'b1000;
															assign node13566 = (inp[10]) ? 4'b1000 : 4'b1000;
												assign node13570 = (inp[5]) ? node13578 : node13571;
													assign node13571 = (inp[0]) ? node13573 : 4'b1101;
														assign node13573 = (inp[9]) ? 4'b1100 : node13574;
															assign node13574 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node13578 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node13581 = (inp[1]) ? node13595 : node13582;
												assign node13582 = (inp[0]) ? node13588 : node13583;
													assign node13583 = (inp[10]) ? node13585 : 4'b1100;
														assign node13585 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node13588 = (inp[5]) ? 4'b1101 : node13589;
														assign node13589 = (inp[9]) ? node13591 : 4'b1101;
															assign node13591 = (inp[10]) ? 4'b1100 : 4'b1100;
												assign node13595 = (inp[5]) ? 4'b1101 : node13596;
													assign node13596 = (inp[10]) ? 4'b1000 : node13597;
														assign node13597 = (inp[9]) ? 4'b1000 : 4'b1001;
										assign node13602 = (inp[2]) ? node13632 : node13603;
											assign node13603 = (inp[1]) ? node13613 : node13604;
												assign node13604 = (inp[11]) ? 4'b1101 : node13605;
													assign node13605 = (inp[9]) ? node13609 : node13606;
														assign node13606 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node13609 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node13613 = (inp[5]) ? node13625 : node13614;
													assign node13614 = (inp[11]) ? node13620 : node13615;
														assign node13615 = (inp[10]) ? 4'b1000 : node13616;
															assign node13616 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node13620 = (inp[10]) ? 4'b1001 : node13621;
															assign node13621 = (inp[9]) ? 4'b1000 : 4'b1000;
													assign node13625 = (inp[9]) ? 4'b1100 : node13626;
														assign node13626 = (inp[11]) ? 4'b1101 : node13627;
															assign node13627 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node13632 = (inp[0]) ? node13648 : node13633;
												assign node13633 = (inp[5]) ? node13641 : node13634;
													assign node13634 = (inp[1]) ? node13636 : 4'b1000;
														assign node13636 = (inp[11]) ? 4'b1101 : node13637;
															assign node13637 = (inp[9]) ? 4'b1100 : 4'b1100;
													assign node13641 = (inp[1]) ? node13643 : 4'b1000;
														assign node13643 = (inp[10]) ? node13645 : 4'b1001;
															assign node13645 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node13648 = (inp[5]) ? node13656 : node13649;
													assign node13649 = (inp[10]) ? node13653 : node13650;
														assign node13650 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node13653 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node13656 = (inp[9]) ? 4'b1001 : node13657;
														assign node13657 = (inp[1]) ? 4'b1000 : 4'b1001;
									assign node13661 = (inp[9]) ? node13701 : node13662;
										assign node13662 = (inp[13]) ? node13682 : node13663;
											assign node13663 = (inp[2]) ? node13673 : node13664;
												assign node13664 = (inp[5]) ? 4'b1101 : node13665;
													assign node13665 = (inp[1]) ? node13669 : node13666;
														assign node13666 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node13669 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node13673 = (inp[11]) ? node13677 : node13674;
													assign node13674 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node13677 = (inp[5]) ? 4'b1000 : node13678;
														assign node13678 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node13682 = (inp[2]) ? node13690 : node13683;
												assign node13683 = (inp[11]) ? 4'b1001 : node13684;
													assign node13684 = (inp[10]) ? 4'b1000 : node13685;
														assign node13685 = (inp[1]) ? 4'b1100 : 4'b1000;
												assign node13690 = (inp[5]) ? node13696 : node13691;
													assign node13691 = (inp[10]) ? 4'b1100 : node13692;
														assign node13692 = (inp[0]) ? 4'b1001 : 4'b1101;
													assign node13696 = (inp[0]) ? node13698 : 4'b1100;
														assign node13698 = (inp[1]) ? 4'b1100 : 4'b1101;
										assign node13701 = (inp[1]) ? node13735 : node13702;
											assign node13702 = (inp[0]) ? node13720 : node13703;
												assign node13703 = (inp[13]) ? node13711 : node13704;
													assign node13704 = (inp[2]) ? node13706 : 4'b1100;
														assign node13706 = (inp[10]) ? node13708 : 4'b1001;
															assign node13708 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node13711 = (inp[2]) ? node13715 : node13712;
														assign node13712 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node13715 = (inp[10]) ? 4'b1101 : node13716;
															assign node13716 = (inp[11]) ? 4'b1100 : 4'b1100;
												assign node13720 = (inp[5]) ? node13730 : node13721;
													assign node13721 = (inp[13]) ? node13727 : node13722;
														assign node13722 = (inp[11]) ? node13724 : 4'b1101;
															assign node13724 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node13727 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node13730 = (inp[2]) ? 4'b1000 : node13731;
														assign node13731 = (inp[13]) ? 4'b1001 : 4'b1101;
											assign node13735 = (inp[10]) ? node13743 : node13736;
												assign node13736 = (inp[13]) ? node13738 : 4'b1101;
													assign node13738 = (inp[0]) ? node13740 : 4'b1101;
														assign node13740 = (inp[5]) ? 4'b1101 : 4'b1001;
												assign node13743 = (inp[13]) ? node13755 : node13744;
													assign node13744 = (inp[5]) ? node13750 : node13745;
														assign node13745 = (inp[2]) ? 4'b1101 : node13746;
															assign node13746 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node13750 = (inp[2]) ? 4'b1001 : node13751;
															assign node13751 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node13755 = (inp[11]) ? node13757 : 4'b1001;
														assign node13757 = (inp[2]) ? 4'b1100 : 4'b1001;
								assign node13760 = (inp[5]) ? node13894 : node13761;
									assign node13761 = (inp[4]) ? node13827 : node13762;
										assign node13762 = (inp[0]) ? node13802 : node13763;
											assign node13763 = (inp[2]) ? node13783 : node13764;
												assign node13764 = (inp[10]) ? node13778 : node13765;
													assign node13765 = (inp[9]) ? node13771 : node13766;
														assign node13766 = (inp[13]) ? node13768 : 4'b1010;
															assign node13768 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node13771 = (inp[11]) ? node13775 : node13772;
															assign node13772 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node13775 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node13778 = (inp[13]) ? node13780 : 4'b1110;
														assign node13780 = (inp[1]) ? 4'b1011 : 4'b1111;
												assign node13783 = (inp[11]) ? node13795 : node13784;
													assign node13784 = (inp[1]) ? node13790 : node13785;
														assign node13785 = (inp[13]) ? node13787 : 4'b1111;
															assign node13787 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node13790 = (inp[13]) ? 4'b1111 : node13791;
															assign node13791 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node13795 = (inp[13]) ? node13797 : 4'b1010;
														assign node13797 = (inp[9]) ? node13799 : 4'b1011;
															assign node13799 = (inp[10]) ? 4'b1010 : 4'b1011;
											assign node13802 = (inp[2]) ? node13814 : node13803;
												assign node13803 = (inp[13]) ? 4'b1011 : node13804;
													assign node13804 = (inp[1]) ? node13810 : node13805;
														assign node13805 = (inp[11]) ? 4'b1011 : node13806;
															assign node13806 = (inp[9]) ? 4'b1010 : 4'b1010;
														assign node13810 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node13814 = (inp[1]) ? node13822 : node13815;
													assign node13815 = (inp[13]) ? node13817 : 4'b1110;
														assign node13817 = (inp[11]) ? 4'b1010 : node13818;
															assign node13818 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node13822 = (inp[10]) ? node13824 : 4'b1010;
														assign node13824 = (inp[11]) ? 4'b1011 : 4'b1010;
										assign node13827 = (inp[11]) ? node13851 : node13828;
											assign node13828 = (inp[9]) ? node13840 : node13829;
												assign node13829 = (inp[2]) ? node13835 : node13830;
													assign node13830 = (inp[1]) ? 4'b1111 : node13831;
														assign node13831 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node13835 = (inp[0]) ? node13837 : 4'b1110;
														assign node13837 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node13840 = (inp[2]) ? node13844 : node13841;
													assign node13841 = (inp[13]) ? 4'b1110 : 4'b1010;
													assign node13844 = (inp[1]) ? node13848 : node13845;
														assign node13845 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node13848 = (inp[10]) ? 4'b1110 : 4'b1111;
											assign node13851 = (inp[9]) ? node13875 : node13852;
												assign node13852 = (inp[0]) ? node13862 : node13853;
													assign node13853 = (inp[2]) ? node13857 : node13854;
														assign node13854 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node13857 = (inp[1]) ? 4'b1111 : node13858;
															assign node13858 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node13862 = (inp[1]) ? node13868 : node13863;
														assign node13863 = (inp[13]) ? 4'b1011 : node13864;
															assign node13864 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node13868 = (inp[2]) ? node13872 : node13869;
															assign node13869 = (inp[13]) ? 4'b1011 : 4'b1111;
															assign node13872 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node13875 = (inp[10]) ? node13881 : node13876;
													assign node13876 = (inp[2]) ? node13878 : 4'b1111;
														assign node13878 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node13881 = (inp[0]) ? node13889 : node13882;
														assign node13882 = (inp[1]) ? node13886 : node13883;
															assign node13883 = (inp[2]) ? 4'b1010 : 4'b1010;
															assign node13886 = (inp[13]) ? 4'b1010 : 4'b1010;
														assign node13889 = (inp[13]) ? node13891 : 4'b1111;
															assign node13891 = (inp[2]) ? 4'b1011 : 4'b1010;
									assign node13894 = (inp[1]) ? node13954 : node13895;
										assign node13895 = (inp[9]) ? node13923 : node13896;
											assign node13896 = (inp[2]) ? node13912 : node13897;
												assign node13897 = (inp[13]) ? node13899 : 4'b1011;
													assign node13899 = (inp[10]) ? node13907 : node13900;
														assign node13900 = (inp[4]) ? node13904 : node13901;
															assign node13901 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node13904 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node13907 = (inp[11]) ? 4'b1110 : node13908;
															assign node13908 = (inp[4]) ? 4'b1111 : 4'b1110;
												assign node13912 = (inp[13]) ? node13918 : node13913;
													assign node13913 = (inp[10]) ? node13915 : 4'b1110;
														assign node13915 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node13918 = (inp[0]) ? node13920 : 4'b1010;
														assign node13920 = (inp[10]) ? 4'b1010 : 4'b1011;
											assign node13923 = (inp[10]) ? node13939 : node13924;
												assign node13924 = (inp[11]) ? node13934 : node13925;
													assign node13925 = (inp[13]) ? node13931 : node13926;
														assign node13926 = (inp[2]) ? 4'b1111 : node13927;
															assign node13927 = (inp[4]) ? 4'b1010 : 4'b1011;
														assign node13931 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node13934 = (inp[13]) ? node13936 : 4'b1111;
														assign node13936 = (inp[2]) ? 4'b1011 : 4'b1111;
												assign node13939 = (inp[4]) ? node13945 : node13940;
													assign node13940 = (inp[2]) ? node13942 : 4'b1010;
														assign node13942 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node13945 = (inp[11]) ? node13949 : node13946;
														assign node13946 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node13949 = (inp[2]) ? 4'b1010 : node13950;
															assign node13950 = (inp[13]) ? 4'b1111 : 4'b1011;
										assign node13954 = (inp[13]) ? node13988 : node13955;
											assign node13955 = (inp[2]) ? node13975 : node13956;
												assign node13956 = (inp[0]) ? node13964 : node13957;
													assign node13957 = (inp[11]) ? 4'b1010 : node13958;
														assign node13958 = (inp[9]) ? 4'b1010 : node13959;
															assign node13959 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node13964 = (inp[11]) ? node13970 : node13965;
														assign node13965 = (inp[4]) ? 4'b1010 : node13966;
															assign node13966 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node13970 = (inp[4]) ? 4'b1011 : node13971;
															assign node13971 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node13975 = (inp[9]) ? node13981 : node13976;
													assign node13976 = (inp[11]) ? node13978 : 4'b1110;
														assign node13978 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node13981 = (inp[10]) ? node13983 : 4'b1111;
														assign node13983 = (inp[4]) ? node13985 : 4'b1110;
															assign node13985 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node13988 = (inp[2]) ? node14000 : node13989;
												assign node13989 = (inp[11]) ? node13991 : 4'b1111;
													assign node13991 = (inp[10]) ? 4'b1111 : node13992;
														assign node13992 = (inp[0]) ? node13996 : node13993;
															assign node13993 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node13996 = (inp[4]) ? 4'b1111 : 4'b1110;
												assign node14000 = (inp[10]) ? 4'b1010 : node14001;
													assign node14001 = (inp[4]) ? node14003 : 4'b1011;
														assign node14003 = (inp[11]) ? 4'b1011 : node14004;
															assign node14004 = (inp[9]) ? 4'b1010 : 4'b1010;
							assign node14009 = (inp[0]) ? node14221 : node14010;
								assign node14010 = (inp[12]) ? node14148 : node14011;
									assign node14011 = (inp[9]) ? node14091 : node14012;
										assign node14012 = (inp[11]) ? node14054 : node14013;
											assign node14013 = (inp[1]) ? node14039 : node14014;
												assign node14014 = (inp[5]) ? node14026 : node14015;
													assign node14015 = (inp[10]) ? node14021 : node14016;
														assign node14016 = (inp[2]) ? 4'b1010 : node14017;
															assign node14017 = (inp[4]) ? 4'b1010 : 4'b1111;
														assign node14021 = (inp[4]) ? node14023 : 4'b1111;
															assign node14023 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node14026 = (inp[10]) ? node14032 : node14027;
														assign node14027 = (inp[4]) ? node14029 : 4'b1110;
															assign node14029 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node14032 = (inp[4]) ? node14036 : node14033;
															assign node14033 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node14036 = (inp[13]) ? 4'b1110 : 4'b1010;
												assign node14039 = (inp[5]) ? node14049 : node14040;
													assign node14040 = (inp[4]) ? node14046 : node14041;
														assign node14041 = (inp[10]) ? 4'b1111 : node14042;
															assign node14042 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node14046 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node14049 = (inp[13]) ? 4'b1011 : node14050;
														assign node14050 = (inp[4]) ? 4'b1111 : 4'b1011;
											assign node14054 = (inp[1]) ? node14074 : node14055;
												assign node14055 = (inp[2]) ? node14065 : node14056;
													assign node14056 = (inp[5]) ? node14060 : node14057;
														assign node14057 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node14060 = (inp[13]) ? node14062 : 4'b1010;
															assign node14062 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node14065 = (inp[5]) ? node14067 : 4'b1011;
														assign node14067 = (inp[4]) ? node14071 : node14068;
															assign node14068 = (inp[13]) ? 4'b1011 : 4'b1111;
															assign node14071 = (inp[13]) ? 4'b1111 : 4'b1011;
												assign node14074 = (inp[5]) ? node14084 : node14075;
													assign node14075 = (inp[4]) ? 4'b1011 : node14076;
														assign node14076 = (inp[2]) ? node14080 : node14077;
															assign node14077 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node14080 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node14084 = (inp[10]) ? node14088 : node14085;
														assign node14085 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node14088 = (inp[13]) ? 4'b1111 : 4'b1110;
										assign node14091 = (inp[5]) ? node14113 : node14092;
											assign node14092 = (inp[4]) ? node14100 : node14093;
												assign node14093 = (inp[10]) ? 4'b1110 : node14094;
													assign node14094 = (inp[1]) ? node14096 : 4'b1110;
														assign node14096 = (inp[13]) ? 4'b1011 : 4'b1111;
												assign node14100 = (inp[1]) ? node14110 : node14101;
													assign node14101 = (inp[13]) ? node14105 : node14102;
														assign node14102 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node14105 = (inp[10]) ? 4'b1010 : node14106;
															assign node14106 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node14110 = (inp[13]) ? 4'b1110 : 4'b1010;
											assign node14113 = (inp[1]) ? node14129 : node14114;
												assign node14114 = (inp[11]) ? node14122 : node14115;
													assign node14115 = (inp[10]) ? 4'b1111 : node14116;
														assign node14116 = (inp[13]) ? node14118 : 4'b1010;
															assign node14118 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node14122 = (inp[13]) ? node14126 : node14123;
														assign node14123 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node14126 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node14129 = (inp[11]) ? node14137 : node14130;
													assign node14130 = (inp[10]) ? 4'b1010 : node14131;
														assign node14131 = (inp[2]) ? 4'b1010 : node14132;
															assign node14132 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node14137 = (inp[2]) ? node14143 : node14138;
														assign node14138 = (inp[4]) ? 4'b1011 : node14139;
															assign node14139 = (inp[10]) ? 4'b1110 : 4'b1011;
														assign node14143 = (inp[10]) ? node14145 : 4'b1111;
															assign node14145 = (inp[13]) ? 4'b1111 : 4'b1011;
									assign node14148 = (inp[10]) ? node14182 : node14149;
										assign node14149 = (inp[5]) ? node14163 : node14150;
											assign node14150 = (inp[13]) ? 4'b1111 : node14151;
												assign node14151 = (inp[4]) ? node14157 : node14152;
													assign node14152 = (inp[1]) ? 4'b1010 : node14153;
														assign node14153 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node14157 = (inp[9]) ? node14159 : 4'b1011;
														assign node14159 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node14163 = (inp[13]) ? node14171 : node14164;
												assign node14164 = (inp[2]) ? 4'b1111 : node14165;
													assign node14165 = (inp[4]) ? 4'b1110 : node14166;
														assign node14166 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node14171 = (inp[9]) ? node14177 : node14172;
													assign node14172 = (inp[11]) ? node14174 : 4'b1010;
														assign node14174 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node14177 = (inp[11]) ? node14179 : 4'b1011;
														assign node14179 = (inp[2]) ? 4'b1010 : 4'b1011;
										assign node14182 = (inp[5]) ? node14198 : node14183;
											assign node14183 = (inp[13]) ? node14191 : node14184;
												assign node14184 = (inp[9]) ? node14188 : node14185;
													assign node14185 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node14188 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node14191 = (inp[11]) ? 4'b1110 : node14192;
													assign node14192 = (inp[1]) ? 4'b1111 : node14193;
														assign node14193 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node14198 = (inp[13]) ? node14210 : node14199;
												assign node14199 = (inp[11]) ? node14205 : node14200;
													assign node14200 = (inp[9]) ? node14202 : 4'b1110;
														assign node14202 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node14205 = (inp[9]) ? node14207 : 4'b1111;
														assign node14207 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node14210 = (inp[9]) ? node14216 : node14211;
													assign node14211 = (inp[11]) ? 4'b1011 : node14212;
														assign node14212 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node14216 = (inp[2]) ? node14218 : 4'b1010;
														assign node14218 = (inp[11]) ? 4'b1010 : 4'b1011;
								assign node14221 = (inp[1]) ? node14339 : node14222;
									assign node14222 = (inp[4]) ? node14280 : node14223;
										assign node14223 = (inp[2]) ? node14263 : node14224;
											assign node14224 = (inp[12]) ? node14242 : node14225;
												assign node14225 = (inp[10]) ? node14233 : node14226;
													assign node14226 = (inp[13]) ? node14228 : 4'b1110;
														assign node14228 = (inp[9]) ? node14230 : 4'b1011;
															assign node14230 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node14233 = (inp[9]) ? node14237 : node14234;
														assign node14234 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node14237 = (inp[5]) ? 4'b1011 : node14238;
															assign node14238 = (inp[13]) ? 4'b1111 : 4'b1011;
												assign node14242 = (inp[13]) ? node14252 : node14243;
													assign node14243 = (inp[5]) ? node14249 : node14244;
														assign node14244 = (inp[11]) ? 4'b1011 : node14245;
															assign node14245 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node14249 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node14252 = (inp[10]) ? node14258 : node14253;
														assign node14253 = (inp[9]) ? 4'b1110 : node14254;
															assign node14254 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node14258 = (inp[11]) ? node14260 : 4'b1110;
															assign node14260 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node14263 = (inp[5]) ? node14271 : node14264;
												assign node14264 = (inp[13]) ? node14266 : 4'b1010;
													assign node14266 = (inp[11]) ? 4'b1110 : node14267;
														assign node14267 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node14271 = (inp[13]) ? 4'b1010 : node14272;
													assign node14272 = (inp[9]) ? node14276 : node14273;
														assign node14273 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node14276 = (inp[11]) ? 4'b1110 : 4'b1111;
										assign node14280 = (inp[12]) ? node14308 : node14281;
											assign node14281 = (inp[11]) ? node14291 : node14282;
												assign node14282 = (inp[9]) ? node14284 : 4'b1111;
													assign node14284 = (inp[5]) ? node14288 : node14285;
														assign node14285 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node14288 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node14291 = (inp[2]) ? node14297 : node14292;
													assign node14292 = (inp[13]) ? node14294 : 4'b1111;
														assign node14294 = (inp[5]) ? 4'b1111 : 4'b1010;
													assign node14297 = (inp[10]) ? node14303 : node14298;
														assign node14298 = (inp[13]) ? node14300 : 4'b1011;
															assign node14300 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node14303 = (inp[9]) ? node14305 : 4'b1010;
															assign node14305 = (inp[13]) ? 4'b1011 : 4'b1010;
											assign node14308 = (inp[10]) ? node14334 : node14309;
												assign node14309 = (inp[11]) ? node14319 : node14310;
													assign node14310 = (inp[13]) ? node14316 : node14311;
														assign node14311 = (inp[5]) ? 4'b1111 : node14312;
															assign node14312 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node14316 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node14319 = (inp[2]) ? node14327 : node14320;
														assign node14320 = (inp[5]) ? node14324 : node14321;
															assign node14321 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node14324 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node14327 = (inp[9]) ? node14331 : node14328;
															assign node14328 = (inp[13]) ? 4'b1011 : 4'b1111;
															assign node14331 = (inp[5]) ? 4'b1110 : 4'b1011;
												assign node14334 = (inp[5]) ? 4'b1111 : node14335;
													assign node14335 = (inp[11]) ? 4'b1011 : 4'b1010;
									assign node14339 = (inp[10]) ? node14405 : node14340;
										assign node14340 = (inp[4]) ? node14380 : node14341;
											assign node14341 = (inp[2]) ? node14361 : node14342;
												assign node14342 = (inp[13]) ? node14348 : node14343;
													assign node14343 = (inp[11]) ? node14345 : 4'b1010;
														assign node14345 = (inp[5]) ? 4'b1010 : 4'b1011;
													assign node14348 = (inp[11]) ? node14356 : node14349;
														assign node14349 = (inp[12]) ? node14353 : node14350;
															assign node14350 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node14353 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node14356 = (inp[12]) ? 4'b1110 : node14357;
															assign node14357 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node14361 = (inp[9]) ? node14369 : node14362;
													assign node14362 = (inp[13]) ? node14364 : 4'b1110;
														assign node14364 = (inp[11]) ? node14366 : 4'b1111;
															assign node14366 = (inp[5]) ? 4'b1111 : 4'b1110;
													assign node14369 = (inp[12]) ? node14375 : node14370;
														assign node14370 = (inp[5]) ? node14372 : 4'b1011;
															assign node14372 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node14375 = (inp[13]) ? 4'b1111 : node14376;
															assign node14376 = (inp[5]) ? 4'b1111 : 4'b1011;
											assign node14380 = (inp[13]) ? node14392 : node14381;
												assign node14381 = (inp[12]) ? node14387 : node14382;
													assign node14382 = (inp[2]) ? node14384 : 4'b1111;
														assign node14384 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node14387 = (inp[11]) ? 4'b1110 : node14388;
														assign node14388 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node14392 = (inp[5]) ? node14398 : node14393;
													assign node14393 = (inp[2]) ? 4'b1110 : node14394;
														assign node14394 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node14398 = (inp[2]) ? 4'b1010 : node14399;
														assign node14399 = (inp[11]) ? 4'b1011 : node14400;
															assign node14400 = (inp[12]) ? 4'b1010 : 4'b1011;
										assign node14405 = (inp[12]) ? node14443 : node14406;
											assign node14406 = (inp[5]) ? node14420 : node14407;
												assign node14407 = (inp[2]) ? node14415 : node14408;
													assign node14408 = (inp[4]) ? node14412 : node14409;
														assign node14409 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node14412 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node14415 = (inp[13]) ? 4'b1111 : node14416;
														assign node14416 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node14420 = (inp[2]) ? node14436 : node14421;
													assign node14421 = (inp[9]) ? node14429 : node14422;
														assign node14422 = (inp[13]) ? node14426 : node14423;
															assign node14423 = (inp[4]) ? 4'b1111 : 4'b1010;
															assign node14426 = (inp[4]) ? 4'b1010 : 4'b1111;
														assign node14429 = (inp[13]) ? node14433 : node14430;
															assign node14430 = (inp[4]) ? 4'b1110 : 4'b1011;
															assign node14433 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node14436 = (inp[9]) ? 4'b1011 : node14437;
														assign node14437 = (inp[13]) ? node14439 : 4'b1010;
															assign node14439 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node14443 = (inp[2]) ? node14453 : node14444;
												assign node14444 = (inp[5]) ? node14446 : 4'b1010;
													assign node14446 = (inp[13]) ? node14448 : 4'b1111;
														assign node14448 = (inp[9]) ? node14450 : 4'b1011;
															assign node14450 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node14453 = (inp[13]) ? node14461 : node14454;
													assign node14454 = (inp[5]) ? 4'b1111 : node14455;
														assign node14455 = (inp[9]) ? 4'b1011 : node14456;
															assign node14456 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node14461 = (inp[5]) ? node14467 : node14462;
														assign node14462 = (inp[4]) ? node14464 : 4'b1111;
															assign node14464 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node14467 = (inp[9]) ? node14469 : 4'b1010;
															assign node14469 = (inp[11]) ? 4'b1010 : 4'b1011;
					assign node14472 = (inp[15]) ? node15420 : node14473;
						assign node14473 = (inp[6]) ? node14969 : node14474;
							assign node14474 = (inp[4]) ? node14726 : node14475;
								assign node14475 = (inp[12]) ? node14589 : node14476;
									assign node14476 = (inp[1]) ? node14530 : node14477;
										assign node14477 = (inp[13]) ? node14493 : node14478;
											assign node14478 = (inp[0]) ? node14484 : node14479;
												assign node14479 = (inp[5]) ? 4'b1110 : node14480;
													assign node14480 = (inp[2]) ? 4'b1110 : 4'b1010;
												assign node14484 = (inp[5]) ? node14488 : node14485;
													assign node14485 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node14488 = (inp[2]) ? node14490 : 4'b1110;
														assign node14490 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node14493 = (inp[0]) ? node14509 : node14494;
												assign node14494 = (inp[11]) ? node14502 : node14495;
													assign node14495 = (inp[9]) ? node14497 : 4'b1011;
														assign node14497 = (inp[5]) ? node14499 : 4'b1011;
															assign node14499 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node14502 = (inp[10]) ? node14504 : 4'b1010;
														assign node14504 = (inp[9]) ? node14506 : 4'b1110;
															assign node14506 = (inp[2]) ? 4'b1110 : 4'b1010;
												assign node14509 = (inp[11]) ? node14519 : node14510;
													assign node14510 = (inp[5]) ? 4'b1110 : node14511;
														assign node14511 = (inp[2]) ? node14515 : node14512;
															assign node14512 = (inp[10]) ? 4'b1110 : 4'b1110;
															assign node14515 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node14519 = (inp[9]) ? node14525 : node14520;
														assign node14520 = (inp[5]) ? 4'b1111 : node14521;
															assign node14521 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node14525 = (inp[5]) ? node14527 : 4'b1011;
															assign node14527 = (inp[2]) ? 4'b1110 : 4'b1010;
										assign node14530 = (inp[5]) ? node14558 : node14531;
											assign node14531 = (inp[11]) ? node14547 : node14532;
												assign node14532 = (inp[0]) ? node14536 : node14533;
													assign node14533 = (inp[13]) ? 4'b1011 : 4'b1110;
													assign node14536 = (inp[9]) ? node14542 : node14537;
														assign node14537 = (inp[13]) ? node14539 : 4'b1010;
															assign node14539 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node14542 = (inp[2]) ? node14544 : 4'b1011;
															assign node14544 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node14547 = (inp[9]) ? node14555 : node14548;
													assign node14548 = (inp[2]) ? node14552 : node14549;
														assign node14549 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node14552 = (inp[0]) ? 4'b1111 : 4'b1010;
													assign node14555 = (inp[0]) ? 4'b1110 : 4'b1010;
											assign node14558 = (inp[2]) ? node14572 : node14559;
												assign node14559 = (inp[13]) ? node14565 : node14560;
													assign node14560 = (inp[0]) ? 4'b1011 : node14561;
														assign node14561 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node14565 = (inp[11]) ? node14567 : 4'b1111;
														assign node14567 = (inp[10]) ? 4'b1110 : node14568;
															assign node14568 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node14572 = (inp[13]) ? node14584 : node14573;
													assign node14573 = (inp[11]) ? node14579 : node14574;
														assign node14574 = (inp[9]) ? node14576 : 4'b1110;
															assign node14576 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node14579 = (inp[0]) ? node14581 : 4'b1110;
															assign node14581 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node14584 = (inp[0]) ? 4'b1011 : node14585;
														assign node14585 = (inp[9]) ? 4'b1011 : 4'b1010;
									assign node14589 = (inp[5]) ? node14667 : node14590;
										assign node14590 = (inp[0]) ? node14624 : node14591;
											assign node14591 = (inp[9]) ? node14609 : node14592;
												assign node14592 = (inp[1]) ? node14598 : node14593;
													assign node14593 = (inp[13]) ? node14595 : 4'b1101;
														assign node14595 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node14598 = (inp[2]) ? node14604 : node14599;
														assign node14599 = (inp[13]) ? node14601 : 4'b1000;
															assign node14601 = (inp[10]) ? 4'b1100 : 4'b1100;
														assign node14604 = (inp[13]) ? node14606 : 4'b1101;
															assign node14606 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node14609 = (inp[1]) ? node14617 : node14610;
													assign node14610 = (inp[11]) ? node14612 : 4'b1101;
														assign node14612 = (inp[10]) ? 4'b1000 : node14613;
															assign node14613 = (inp[13]) ? 4'b1101 : 4'b1000;
													assign node14617 = (inp[13]) ? node14621 : node14618;
														assign node14618 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node14621 = (inp[2]) ? 4'b1000 : 4'b1100;
											assign node14624 = (inp[1]) ? node14644 : node14625;
												assign node14625 = (inp[11]) ? node14637 : node14626;
													assign node14626 = (inp[10]) ? node14630 : node14627;
														assign node14627 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node14630 = (inp[13]) ? node14634 : node14631;
															assign node14631 = (inp[2]) ? 4'b1001 : 4'b1100;
															assign node14634 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node14637 = (inp[2]) ? node14641 : node14638;
														assign node14638 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node14641 = (inp[13]) ? 4'b1100 : 4'b1000;
												assign node14644 = (inp[11]) ? node14658 : node14645;
													assign node14645 = (inp[9]) ? node14653 : node14646;
														assign node14646 = (inp[2]) ? node14650 : node14647;
															assign node14647 = (inp[10]) ? 4'b1000 : 4'b1100;
															assign node14650 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node14653 = (inp[10]) ? node14655 : 4'b1001;
															assign node14655 = (inp[13]) ? 4'b1000 : 4'b1101;
													assign node14658 = (inp[9]) ? 4'b1000 : node14659;
														assign node14659 = (inp[13]) ? node14663 : node14660;
															assign node14660 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node14663 = (inp[10]) ? 4'b1101 : 4'b1001;
										assign node14667 = (inp[11]) ? node14705 : node14668;
											assign node14668 = (inp[1]) ? node14688 : node14669;
												assign node14669 = (inp[0]) ? node14681 : node14670;
													assign node14670 = (inp[13]) ? node14678 : node14671;
														assign node14671 = (inp[2]) ? node14675 : node14672;
															assign node14672 = (inp[9]) ? 4'b1100 : 4'b1100;
															assign node14675 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node14678 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node14681 = (inp[9]) ? 4'b1101 : node14682;
														assign node14682 = (inp[2]) ? node14684 : 4'b1101;
															assign node14684 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node14688 = (inp[9]) ? node14700 : node14689;
													assign node14689 = (inp[13]) ? node14695 : node14690;
														assign node14690 = (inp[2]) ? node14692 : 4'b1100;
															assign node14692 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node14695 = (inp[2]) ? 4'b1101 : node14696;
															assign node14696 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node14700 = (inp[2]) ? 4'b1100 : node14701;
														assign node14701 = (inp[13]) ? 4'b1001 : 4'b1100;
											assign node14705 = (inp[1]) ? node14715 : node14706;
												assign node14706 = (inp[9]) ? node14708 : 4'b1000;
													assign node14708 = (inp[2]) ? node14712 : node14709;
														assign node14709 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node14712 = (inp[13]) ? 4'b1100 : 4'b1001;
												assign node14715 = (inp[9]) ? node14721 : node14716;
													assign node14716 = (inp[13]) ? 4'b1100 : node14717;
														assign node14717 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node14721 = (inp[13]) ? node14723 : 4'b1000;
														assign node14723 = (inp[2]) ? 4'b1100 : 4'b1000;
								assign node14726 = (inp[12]) ? node14848 : node14727;
									assign node14727 = (inp[1]) ? node14775 : node14728;
										assign node14728 = (inp[10]) ? node14752 : node14729;
											assign node14729 = (inp[5]) ? node14739 : node14730;
												assign node14730 = (inp[9]) ? node14732 : 4'b1100;
													assign node14732 = (inp[2]) ? node14736 : node14733;
														assign node14733 = (inp[0]) ? 4'b1001 : 4'b1101;
														assign node14736 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node14739 = (inp[9]) ? node14749 : node14740;
													assign node14740 = (inp[13]) ? node14744 : node14741;
														assign node14741 = (inp[0]) ? 4'b1101 : 4'b1001;
														assign node14744 = (inp[2]) ? node14746 : 4'b1000;
															assign node14746 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node14749 = (inp[11]) ? 4'b1000 : 4'b1100;
											assign node14752 = (inp[9]) ? node14764 : node14753;
												assign node14753 = (inp[13]) ? node14757 : node14754;
													assign node14754 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node14757 = (inp[11]) ? 4'b1000 : node14758;
														assign node14758 = (inp[5]) ? 4'b1001 : node14759;
															assign node14759 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node14764 = (inp[0]) ? node14772 : node14765;
													assign node14765 = (inp[11]) ? 4'b1100 : node14766;
														assign node14766 = (inp[5]) ? node14768 : 4'b1100;
															assign node14768 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node14772 = (inp[2]) ? 4'b1100 : 4'b1000;
										assign node14775 = (inp[9]) ? node14813 : node14776;
											assign node14776 = (inp[10]) ? node14794 : node14777;
												assign node14777 = (inp[5]) ? node14783 : node14778;
													assign node14778 = (inp[13]) ? node14780 : 4'b1101;
														assign node14780 = (inp[0]) ? 4'b1101 : 4'b1000;
													assign node14783 = (inp[11]) ? node14789 : node14784;
														assign node14784 = (inp[2]) ? 4'b1001 : node14785;
															assign node14785 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node14789 = (inp[13]) ? 4'b1100 : node14790;
															assign node14790 = (inp[2]) ? 4'b1000 : 4'b1100;
												assign node14794 = (inp[2]) ? node14802 : node14795;
													assign node14795 = (inp[13]) ? node14799 : node14796;
														assign node14796 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node14799 = (inp[11]) ? 4'b1000 : 4'b1101;
													assign node14802 = (inp[13]) ? node14808 : node14803;
														assign node14803 = (inp[5]) ? node14805 : 4'b1100;
															assign node14805 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node14808 = (inp[5]) ? node14810 : 4'b1001;
															assign node14810 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node14813 = (inp[10]) ? node14829 : node14814;
												assign node14814 = (inp[0]) ? node14824 : node14815;
													assign node14815 = (inp[13]) ? node14817 : 4'b1101;
														assign node14817 = (inp[5]) ? node14821 : node14818;
															assign node14818 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node14821 = (inp[2]) ? 4'b1101 : 4'b1000;
													assign node14824 = (inp[11]) ? 4'b1101 : node14825;
														assign node14825 = (inp[5]) ? 4'b1000 : 4'b1001;
												assign node14829 = (inp[0]) ? node14839 : node14830;
													assign node14830 = (inp[2]) ? node14832 : 4'b1001;
														assign node14832 = (inp[5]) ? node14836 : node14833;
															assign node14833 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node14836 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node14839 = (inp[2]) ? 4'b1000 : node14840;
														assign node14840 = (inp[5]) ? node14844 : node14841;
															assign node14841 = (inp[13]) ? 4'b1101 : 4'b1000;
															assign node14844 = (inp[13]) ? 4'b1000 : 4'b1101;
									assign node14848 = (inp[1]) ? node14910 : node14849;
										assign node14849 = (inp[10]) ? node14875 : node14850;
											assign node14850 = (inp[9]) ? node14864 : node14851;
												assign node14851 = (inp[5]) ? node14857 : node14852;
													assign node14852 = (inp[2]) ? node14854 : 4'b1111;
														assign node14854 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node14857 = (inp[0]) ? 4'b1010 : node14858;
														assign node14858 = (inp[2]) ? node14860 : 4'b1011;
															assign node14860 = (inp[13]) ? 4'b1010 : 4'b1110;
												assign node14864 = (inp[2]) ? node14868 : node14865;
													assign node14865 = (inp[13]) ? 4'b1110 : 4'b1010;
													assign node14868 = (inp[13]) ? node14872 : node14869;
														assign node14869 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node14872 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node14875 = (inp[11]) ? node14893 : node14876;
												assign node14876 = (inp[2]) ? node14882 : node14877;
													assign node14877 = (inp[13]) ? 4'b1110 : node14878;
														assign node14878 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node14882 = (inp[13]) ? node14886 : node14883;
														assign node14883 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node14886 = (inp[9]) ? node14890 : node14887;
															assign node14887 = (inp[5]) ? 4'b1011 : 4'b1010;
															assign node14890 = (inp[5]) ? 4'b1010 : 4'b1011;
												assign node14893 = (inp[2]) ? node14901 : node14894;
													assign node14894 = (inp[13]) ? node14896 : 4'b1011;
														assign node14896 = (inp[0]) ? node14898 : 4'b1111;
															assign node14898 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node14901 = (inp[0]) ? node14903 : 4'b1110;
														assign node14903 = (inp[9]) ? node14907 : node14904;
															assign node14904 = (inp[5]) ? 4'b1110 : 4'b1111;
															assign node14907 = (inp[5]) ? 4'b1111 : 4'b1110;
										assign node14910 = (inp[10]) ? node14940 : node14911;
											assign node14911 = (inp[11]) ? node14929 : node14912;
												assign node14912 = (inp[13]) ? node14924 : node14913;
													assign node14913 = (inp[2]) ? node14919 : node14914;
														assign node14914 = (inp[5]) ? node14916 : 4'b1110;
															assign node14916 = (inp[9]) ? 4'b1010 : 4'b1010;
														assign node14919 = (inp[5]) ? 4'b1110 : node14920;
															assign node14920 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node14924 = (inp[9]) ? node14926 : 4'b1010;
														assign node14926 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node14929 = (inp[9]) ? node14933 : node14930;
													assign node14930 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node14933 = (inp[2]) ? 4'b1011 : node14934;
														assign node14934 = (inp[13]) ? 4'b1111 : node14935;
															assign node14935 = (inp[5]) ? 4'b1011 : 4'b1111;
											assign node14940 = (inp[13]) ? node14952 : node14941;
												assign node14941 = (inp[2]) ? node14943 : 4'b1010;
													assign node14943 = (inp[11]) ? node14947 : node14944;
														assign node14944 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node14947 = (inp[0]) ? 4'b1011 : node14948;
															assign node14948 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node14952 = (inp[11]) ? node14960 : node14953;
													assign node14953 = (inp[0]) ? 4'b1010 : node14954;
														assign node14954 = (inp[2]) ? 4'b1011 : node14955;
															assign node14955 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node14960 = (inp[2]) ? node14966 : node14961;
														assign node14961 = (inp[0]) ? node14963 : 4'b1010;
															assign node14963 = (inp[5]) ? 4'b1111 : 4'b1011;
														assign node14966 = (inp[5]) ? 4'b1010 : 4'b1110;
							assign node14969 = (inp[9]) ? node15189 : node14970;
								assign node14970 = (inp[0]) ? node15084 : node14971;
									assign node14971 = (inp[13]) ? node15023 : node14972;
										assign node14972 = (inp[5]) ? node14992 : node14973;
											assign node14973 = (inp[1]) ? node14987 : node14974;
												assign node14974 = (inp[12]) ? node14980 : node14975;
													assign node14975 = (inp[10]) ? node14977 : 4'b1011;
														assign node14977 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node14980 = (inp[4]) ? 4'b1010 : node14981;
														assign node14981 = (inp[10]) ? node14983 : 4'b1110;
															assign node14983 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node14987 = (inp[12]) ? node14989 : 4'b1011;
													assign node14989 = (inp[11]) ? 4'b1011 : 4'b1010;
											assign node14992 = (inp[1]) ? node15010 : node14993;
												assign node14993 = (inp[2]) ? node15003 : node14994;
													assign node14994 = (inp[11]) ? node15000 : node14995;
														assign node14995 = (inp[12]) ? node14997 : 4'b1010;
															assign node14997 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node15000 = (inp[12]) ? 4'b1011 : 4'b1110;
													assign node15003 = (inp[10]) ? 4'b1111 : node15004;
														assign node15004 = (inp[12]) ? 4'b1011 : node15005;
															assign node15005 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node15010 = (inp[2]) ? node15016 : node15011;
													assign node15011 = (inp[4]) ? node15013 : 4'b1111;
														assign node15013 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node15016 = (inp[4]) ? 4'b1110 : node15017;
														assign node15017 = (inp[12]) ? 4'b1110 : node15018;
															assign node15018 = (inp[11]) ? 4'b1111 : 4'b1110;
										assign node15023 = (inp[5]) ? node15051 : node15024;
											assign node15024 = (inp[1]) ? node15042 : node15025;
												assign node15025 = (inp[2]) ? node15035 : node15026;
													assign node15026 = (inp[4]) ? node15032 : node15027;
														assign node15027 = (inp[12]) ? node15029 : 4'b1110;
															assign node15029 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node15032 = (inp[12]) ? 4'b1110 : 4'b1010;
													assign node15035 = (inp[11]) ? 4'b1011 : node15036;
														assign node15036 = (inp[12]) ? 4'b1111 : node15037;
															assign node15037 = (inp[4]) ? 4'b1010 : 4'b1111;
												assign node15042 = (inp[2]) ? 4'b1110 : node15043;
													assign node15043 = (inp[11]) ? node15045 : 4'b1111;
														assign node15045 = (inp[12]) ? node15047 : 4'b1110;
															assign node15047 = (inp[4]) ? 4'b1110 : 4'b1111;
											assign node15051 = (inp[1]) ? node15071 : node15052;
												assign node15052 = (inp[11]) ? node15062 : node15053;
													assign node15053 = (inp[12]) ? node15057 : node15054;
														assign node15054 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node15057 = (inp[4]) ? 4'b1011 : node15058;
															assign node15058 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node15062 = (inp[12]) ? node15066 : node15063;
														assign node15063 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node15066 = (inp[10]) ? node15068 : 4'b1010;
															assign node15068 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node15071 = (inp[12]) ? node15079 : node15072;
													assign node15072 = (inp[10]) ? node15074 : 4'b1011;
														assign node15074 = (inp[2]) ? node15076 : 4'b1011;
															assign node15076 = (inp[4]) ? 4'b1010 : 4'b1010;
													assign node15079 = (inp[11]) ? node15081 : 4'b1010;
														assign node15081 = (inp[4]) ? 4'b1010 : 4'b1011;
									assign node15084 = (inp[11]) ? node15144 : node15085;
										assign node15085 = (inp[13]) ? node15113 : node15086;
											assign node15086 = (inp[5]) ? node15100 : node15087;
												assign node15087 = (inp[1]) ? node15093 : node15088;
													assign node15088 = (inp[4]) ? 4'b1111 : node15089;
														assign node15089 = (inp[12]) ? 4'b1110 : 4'b1010;
													assign node15093 = (inp[10]) ? node15095 : 4'b1011;
														assign node15095 = (inp[12]) ? 4'b1011 : node15096;
															assign node15096 = (inp[4]) ? 4'b1010 : 4'b1010;
												assign node15100 = (inp[1]) ? node15108 : node15101;
													assign node15101 = (inp[10]) ? node15103 : 4'b1011;
														assign node15103 = (inp[2]) ? 4'b1111 : node15104;
															assign node15104 = (inp[12]) ? 4'b1010 : 4'b1010;
													assign node15108 = (inp[2]) ? 4'b1111 : node15109;
														assign node15109 = (inp[10]) ? 4'b1111 : 4'b1110;
											assign node15113 = (inp[4]) ? node15125 : node15114;
												assign node15114 = (inp[2]) ? node15122 : node15115;
													assign node15115 = (inp[5]) ? node15117 : 4'b1110;
														assign node15117 = (inp[10]) ? 4'b1010 : node15118;
															assign node15118 = (inp[12]) ? 4'b1010 : 4'b1011;
													assign node15122 = (inp[5]) ? 4'b1010 : 4'b1011;
												assign node15125 = (inp[2]) ? node15133 : node15126;
													assign node15126 = (inp[12]) ? node15130 : node15127;
														assign node15127 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node15130 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node15133 = (inp[5]) ? node15139 : node15134;
														assign node15134 = (inp[12]) ? 4'b1110 : node15135;
															assign node15135 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node15139 = (inp[12]) ? 4'b1010 : node15140;
															assign node15140 = (inp[10]) ? 4'b1111 : 4'b1010;
										assign node15144 = (inp[13]) ? node15164 : node15145;
											assign node15145 = (inp[5]) ? node15157 : node15146;
												assign node15146 = (inp[2]) ? node15152 : node15147;
													assign node15147 = (inp[4]) ? 4'b1011 : node15148;
														assign node15148 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node15152 = (inp[4]) ? node15154 : 4'b1011;
														assign node15154 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node15157 = (inp[1]) ? 4'b1110 : node15158;
													assign node15158 = (inp[12]) ? node15160 : 4'b1111;
														assign node15160 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node15164 = (inp[5]) ? node15174 : node15165;
												assign node15165 = (inp[4]) ? node15171 : node15166;
													assign node15166 = (inp[12]) ? 4'b1010 : node15167;
														assign node15167 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node15171 = (inp[10]) ? 4'b1111 : 4'b1011;
												assign node15174 = (inp[1]) ? node15184 : node15175;
													assign node15175 = (inp[12]) ? node15181 : node15176;
														assign node15176 = (inp[4]) ? 4'b1110 : node15177;
															assign node15177 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node15181 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node15184 = (inp[12]) ? node15186 : 4'b1011;
														assign node15186 = (inp[2]) ? 4'b1011 : 4'b1010;
								assign node15189 = (inp[11]) ? node15315 : node15190;
									assign node15190 = (inp[10]) ? node15254 : node15191;
										assign node15191 = (inp[1]) ? node15223 : node15192;
											assign node15192 = (inp[12]) ? node15214 : node15193;
												assign node15193 = (inp[2]) ? node15207 : node15194;
													assign node15194 = (inp[0]) ? node15202 : node15195;
														assign node15195 = (inp[5]) ? node15199 : node15196;
															assign node15196 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node15199 = (inp[4]) ? 4'b1011 : 4'b1110;
														assign node15202 = (inp[5]) ? 4'b1010 : node15203;
															assign node15203 = (inp[13]) ? 4'b1111 : 4'b1010;
													assign node15207 = (inp[13]) ? node15209 : 4'b1110;
														assign node15209 = (inp[0]) ? 4'b1110 : node15210;
															assign node15210 = (inp[5]) ? 4'b1011 : 4'b1110;
												assign node15214 = (inp[2]) ? node15220 : node15215;
													assign node15215 = (inp[4]) ? node15217 : 4'b1111;
														assign node15217 = (inp[13]) ? 4'b1110 : 4'b1011;
													assign node15220 = (inp[5]) ? 4'b1011 : 4'b1010;
											assign node15223 = (inp[0]) ? node15247 : node15224;
												assign node15224 = (inp[4]) ? node15234 : node15225;
													assign node15225 = (inp[13]) ? node15231 : node15226;
														assign node15226 = (inp[5]) ? node15228 : 4'b1011;
															assign node15228 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node15231 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node15234 = (inp[13]) ? node15240 : node15235;
														assign node15235 = (inp[5]) ? node15237 : 4'b1011;
															assign node15237 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node15240 = (inp[5]) ? node15244 : node15241;
															assign node15241 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node15244 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node15247 = (inp[5]) ? 4'b1110 : node15248;
													assign node15248 = (inp[13]) ? node15250 : 4'b1010;
														assign node15250 = (inp[4]) ? 4'b1111 : 4'b1110;
										assign node15254 = (inp[2]) ? node15286 : node15255;
											assign node15255 = (inp[1]) ? node15273 : node15256;
												assign node15256 = (inp[4]) ? node15270 : node15257;
													assign node15257 = (inp[0]) ? node15265 : node15258;
														assign node15258 = (inp[5]) ? node15262 : node15259;
															assign node15259 = (inp[12]) ? 4'b1111 : 4'b1011;
															assign node15262 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node15265 = (inp[12]) ? node15267 : 4'b1010;
															assign node15267 = (inp[5]) ? 4'b1010 : 4'b1010;
													assign node15270 = (inp[13]) ? 4'b1010 : 4'b1011;
												assign node15273 = (inp[0]) ? node15275 : 4'b1011;
													assign node15275 = (inp[4]) ? node15283 : node15276;
														assign node15276 = (inp[13]) ? node15280 : node15277;
															assign node15277 = (inp[12]) ? 4'b1111 : 4'b1110;
															assign node15280 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node15283 = (inp[13]) ? 4'b1111 : 4'b1011;
											assign node15286 = (inp[4]) ? node15298 : node15287;
												assign node15287 = (inp[12]) ? node15293 : node15288;
													assign node15288 = (inp[13]) ? node15290 : 4'b1010;
														assign node15290 = (inp[5]) ? 4'b1010 : 4'b1110;
													assign node15293 = (inp[13]) ? node15295 : 4'b1011;
														assign node15295 = (inp[5]) ? 4'b1011 : 4'b1010;
												assign node15298 = (inp[13]) ? node15306 : node15299;
													assign node15299 = (inp[12]) ? 4'b1110 : node15300;
														assign node15300 = (inp[5]) ? 4'b1010 : node15301;
															assign node15301 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node15306 = (inp[5]) ? node15310 : node15307;
														assign node15307 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node15310 = (inp[0]) ? 4'b1011 : node15311;
															assign node15311 = (inp[1]) ? 4'b1011 : 4'b1111;
									assign node15315 = (inp[1]) ? node15373 : node15316;
										assign node15316 = (inp[10]) ? node15352 : node15317;
											assign node15317 = (inp[2]) ? node15331 : node15318;
												assign node15318 = (inp[13]) ? node15324 : node15319;
													assign node15319 = (inp[4]) ? node15321 : 4'b1010;
														assign node15321 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node15324 = (inp[0]) ? node15326 : 4'b1011;
														assign node15326 = (inp[4]) ? node15328 : 4'b1011;
															assign node15328 = (inp[12]) ? 4'b1011 : 4'b1110;
												assign node15331 = (inp[5]) ? node15341 : node15332;
													assign node15332 = (inp[13]) ? node15336 : node15333;
														assign node15333 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node15336 = (inp[4]) ? 4'b1110 : node15337;
															assign node15337 = (inp[0]) ? 4'b1011 : 4'b1111;
													assign node15341 = (inp[13]) ? node15345 : node15342;
														assign node15342 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node15345 = (inp[0]) ? node15349 : node15346;
															assign node15346 = (inp[12]) ? 4'b1111 : 4'b1110;
															assign node15349 = (inp[4]) ? 4'b1111 : 4'b1110;
											assign node15352 = (inp[2]) ? node15368 : node15353;
												assign node15353 = (inp[4]) ? node15361 : node15354;
													assign node15354 = (inp[12]) ? node15356 : 4'b1010;
														assign node15356 = (inp[0]) ? node15358 : 4'b1110;
															assign node15358 = (inp[5]) ? 4'b1110 : 4'b1011;
													assign node15361 = (inp[12]) ? node15363 : 4'b1011;
														assign node15363 = (inp[0]) ? 4'b1110 : node15364;
															assign node15364 = (inp[13]) ? 4'b1011 : 4'b1011;
												assign node15368 = (inp[4]) ? node15370 : 4'b1010;
													assign node15370 = (inp[0]) ? 4'b1010 : 4'b1110;
										assign node15373 = (inp[2]) ? node15401 : node15374;
											assign node15374 = (inp[4]) ? node15388 : node15375;
												assign node15375 = (inp[13]) ? node15385 : node15376;
													assign node15376 = (inp[5]) ? node15382 : node15377;
														assign node15377 = (inp[0]) ? node15379 : 4'b1010;
															assign node15379 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node15382 = (inp[12]) ? 4'b1110 : 4'b1111;
													assign node15385 = (inp[5]) ? 4'b1010 : 4'b1110;
												assign node15388 = (inp[13]) ? node15394 : node15389;
													assign node15389 = (inp[5]) ? node15391 : 4'b1010;
														assign node15391 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node15394 = (inp[0]) ? node15398 : node15395;
														assign node15395 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node15398 = (inp[12]) ? 4'b1110 : 4'b1010;
											assign node15401 = (inp[13]) ? node15415 : node15402;
												assign node15402 = (inp[5]) ? node15412 : node15403;
													assign node15403 = (inp[12]) ? node15407 : node15404;
														assign node15404 = (inp[4]) ? 4'b1010 : 4'b1011;
														assign node15407 = (inp[0]) ? node15409 : 4'b1010;
															assign node15409 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node15412 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node15415 = (inp[5]) ? 4'b1010 : node15416;
													assign node15416 = (inp[4]) ? 4'b1110 : 4'b1111;
						assign node15420 = (inp[6]) ? node15896 : node15421;
							assign node15421 = (inp[12]) ? node15655 : node15422;
								assign node15422 = (inp[5]) ? node15550 : node15423;
									assign node15423 = (inp[11]) ? node15489 : node15424;
										assign node15424 = (inp[0]) ? node15446 : node15425;
											assign node15425 = (inp[10]) ? node15429 : node15426;
												assign node15426 = (inp[2]) ? 4'b1110 : 4'b1010;
												assign node15429 = (inp[1]) ? node15437 : node15430;
													assign node15430 = (inp[9]) ? 4'b1110 : node15431;
														assign node15431 = (inp[4]) ? node15433 : 4'b1011;
															assign node15433 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node15437 = (inp[9]) ? node15443 : node15438;
														assign node15438 = (inp[13]) ? node15440 : 4'b1110;
															assign node15440 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node15443 = (inp[13]) ? 4'b1010 : 4'b1011;
											assign node15446 = (inp[13]) ? node15468 : node15447;
												assign node15447 = (inp[9]) ? node15459 : node15448;
													assign node15448 = (inp[2]) ? node15452 : node15449;
														assign node15449 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node15452 = (inp[10]) ? node15456 : node15453;
															assign node15453 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node15456 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node15459 = (inp[10]) ? node15465 : node15460;
														assign node15460 = (inp[1]) ? 4'b1111 : node15461;
															assign node15461 = (inp[2]) ? 4'b1110 : 4'b1011;
														assign node15465 = (inp[4]) ? 4'b1111 : 4'b1110;
												assign node15468 = (inp[9]) ? node15478 : node15469;
													assign node15469 = (inp[2]) ? node15475 : node15470;
														assign node15470 = (inp[4]) ? node15472 : 4'b1011;
															assign node15472 = (inp[1]) ? 4'b1110 : 4'b1110;
														assign node15475 = (inp[10]) ? 4'b1011 : 4'b1110;
													assign node15478 = (inp[2]) ? node15482 : node15479;
														assign node15479 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node15482 = (inp[1]) ? node15486 : node15483;
															assign node15483 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node15486 = (inp[10]) ? 4'b1110 : 4'b1111;
										assign node15489 = (inp[10]) ? node15523 : node15490;
											assign node15490 = (inp[0]) ? node15510 : node15491;
												assign node15491 = (inp[13]) ? node15503 : node15492;
													assign node15492 = (inp[2]) ? node15498 : node15493;
														assign node15493 = (inp[4]) ? 4'b1011 : node15494;
															assign node15494 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node15498 = (inp[4]) ? node15500 : 4'b1011;
															assign node15500 = (inp[1]) ? 4'b1111 : 4'b1110;
													assign node15503 = (inp[4]) ? node15507 : node15504;
														assign node15504 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node15507 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node15510 = (inp[4]) ? node15516 : node15511;
													assign node15511 = (inp[9]) ? 4'b1110 : node15512;
														assign node15512 = (inp[1]) ? 4'b1011 : 4'b1110;
													assign node15516 = (inp[2]) ? 4'b1011 : node15517;
														assign node15517 = (inp[13]) ? 4'b1110 : node15518;
															assign node15518 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node15523 = (inp[1]) ? node15543 : node15524;
												assign node15524 = (inp[0]) ? node15530 : node15525;
													assign node15525 = (inp[2]) ? node15527 : 4'b1010;
														assign node15527 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node15530 = (inp[13]) ? node15536 : node15531;
														assign node15531 = (inp[4]) ? node15533 : 4'b1111;
															assign node15533 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node15536 = (inp[9]) ? node15540 : node15537;
															assign node15537 = (inp[4]) ? 4'b1010 : 4'b1111;
															assign node15540 = (inp[2]) ? 4'b1110 : 4'b1010;
												assign node15543 = (inp[13]) ? node15545 : 4'b1111;
													assign node15545 = (inp[2]) ? 4'b1011 : node15546;
														assign node15546 = (inp[4]) ? 4'b1111 : 4'b1011;
									assign node15550 = (inp[1]) ? node15610 : node15551;
										assign node15551 = (inp[0]) ? node15591 : node15552;
											assign node15552 = (inp[2]) ? node15568 : node15553;
												assign node15553 = (inp[9]) ? node15563 : node15554;
													assign node15554 = (inp[11]) ? 4'b1011 : node15555;
														assign node15555 = (inp[10]) ? node15559 : node15556;
															assign node15556 = (inp[4]) ? 4'b1010 : 4'b1011;
															assign node15559 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node15563 = (inp[10]) ? node15565 : 4'b1010;
														assign node15565 = (inp[4]) ? 4'b1010 : 4'b1111;
												assign node15568 = (inp[11]) ? node15580 : node15569;
													assign node15569 = (inp[4]) ? node15573 : node15570;
														assign node15570 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node15573 = (inp[13]) ? node15577 : node15574;
															assign node15574 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node15577 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node15580 = (inp[13]) ? node15586 : node15581;
														assign node15581 = (inp[4]) ? 4'b1011 : node15582;
															assign node15582 = (inp[10]) ? 4'b1110 : 4'b1110;
														assign node15586 = (inp[4]) ? 4'b1110 : node15587;
															assign node15587 = (inp[9]) ? 4'b1011 : 4'b1010;
											assign node15591 = (inp[2]) ? node15597 : node15592;
												assign node15592 = (inp[11]) ? 4'b1010 : node15593;
													assign node15593 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node15597 = (inp[11]) ? node15603 : node15598;
													assign node15598 = (inp[9]) ? node15600 : 4'b1010;
														assign node15600 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node15603 = (inp[4]) ? node15607 : node15604;
														assign node15604 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node15607 = (inp[13]) ? 4'b1111 : 4'b1011;
										assign node15610 = (inp[2]) ? node15632 : node15611;
											assign node15611 = (inp[9]) ? node15619 : node15612;
												assign node15612 = (inp[10]) ? 4'b1111 : node15613;
													assign node15613 = (inp[13]) ? node15615 : 4'b1110;
														assign node15615 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node15619 = (inp[4]) ? node15623 : node15620;
													assign node15620 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node15623 = (inp[13]) ? node15629 : node15624;
														assign node15624 = (inp[0]) ? 4'b1010 : node15625;
															assign node15625 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node15629 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node15632 = (inp[13]) ? node15640 : node15633;
												assign node15633 = (inp[4]) ? 4'b1111 : node15634;
													assign node15634 = (inp[10]) ? 4'b1011 : node15635;
														assign node15635 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node15640 = (inp[4]) ? node15648 : node15641;
													assign node15641 = (inp[9]) ? 4'b1111 : node15642;
														assign node15642 = (inp[11]) ? 4'b1110 : node15643;
															assign node15643 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node15648 = (inp[10]) ? 4'b1010 : node15649;
														assign node15649 = (inp[11]) ? 4'b1011 : node15650;
															assign node15650 = (inp[9]) ? 4'b1010 : 4'b1010;
								assign node15655 = (inp[10]) ? node15767 : node15656;
									assign node15656 = (inp[9]) ? node15714 : node15657;
										assign node15657 = (inp[11]) ? node15683 : node15658;
											assign node15658 = (inp[5]) ? node15674 : node15659;
												assign node15659 = (inp[0]) ? node15667 : node15660;
													assign node15660 = (inp[1]) ? node15662 : 4'b1101;
														assign node15662 = (inp[4]) ? node15664 : 4'b1100;
															assign node15664 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node15667 = (inp[4]) ? 4'b1100 : node15668;
														assign node15668 = (inp[1]) ? 4'b1100 : node15669;
															assign node15669 = (inp[13]) ? 4'b1000 : 4'b1000;
												assign node15674 = (inp[2]) ? node15680 : node15675;
													assign node15675 = (inp[13]) ? node15677 : 4'b1000;
														assign node15677 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node15680 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node15683 = (inp[2]) ? node15703 : node15684;
												assign node15684 = (inp[4]) ? node15694 : node15685;
													assign node15685 = (inp[13]) ? node15689 : node15686;
														assign node15686 = (inp[5]) ? 4'b1000 : 4'b1100;
														assign node15689 = (inp[0]) ? node15691 : 4'b1100;
															assign node15691 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node15694 = (inp[0]) ? node15700 : node15695;
														assign node15695 = (inp[5]) ? 4'b1101 : node15696;
															assign node15696 = (inp[1]) ? 4'b1001 : 4'b1101;
														assign node15700 = (inp[13]) ? 4'b1100 : 4'b1101;
												assign node15703 = (inp[13]) ? node15707 : node15704;
													assign node15704 = (inp[5]) ? 4'b1100 : 4'b1001;
													assign node15707 = (inp[5]) ? 4'b1000 : node15708;
														assign node15708 = (inp[1]) ? 4'b1100 : node15709;
															assign node15709 = (inp[4]) ? 4'b1000 : 4'b1001;
										assign node15714 = (inp[4]) ? node15738 : node15715;
											assign node15715 = (inp[1]) ? node15727 : node15716;
												assign node15716 = (inp[11]) ? node15720 : node15717;
													assign node15717 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node15720 = (inp[5]) ? 4'b1100 : node15721;
														assign node15721 = (inp[0]) ? 4'b1000 : node15722;
															assign node15722 = (inp[13]) ? 4'b1000 : 4'b1100;
												assign node15727 = (inp[5]) ? node15731 : node15728;
													assign node15728 = (inp[0]) ? 4'b1101 : 4'b1000;
													assign node15731 = (inp[11]) ? node15733 : 4'b1000;
														assign node15733 = (inp[13]) ? node15735 : 4'b1101;
															assign node15735 = (inp[2]) ? 4'b1001 : 4'b1101;
											assign node15738 = (inp[1]) ? node15750 : node15739;
												assign node15739 = (inp[13]) ? node15747 : node15740;
													assign node15740 = (inp[2]) ? node15742 : 4'b1001;
														assign node15742 = (inp[11]) ? node15744 : 4'b1101;
															assign node15744 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node15747 = (inp[2]) ? 4'b1001 : 4'b1101;
												assign node15750 = (inp[11]) ? node15760 : node15751;
													assign node15751 = (inp[13]) ? node15753 : 4'b1001;
														assign node15753 = (inp[2]) ? node15757 : node15754;
															assign node15754 = (inp[5]) ? 4'b1101 : 4'b1001;
															assign node15757 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node15760 = (inp[5]) ? node15762 : 4'b1000;
														assign node15762 = (inp[0]) ? node15764 : 4'b1000;
															assign node15764 = (inp[2]) ? 4'b1001 : 4'b1101;
									assign node15767 = (inp[1]) ? node15825 : node15768;
										assign node15768 = (inp[4]) ? node15792 : node15769;
											assign node15769 = (inp[0]) ? node15775 : node15770;
												assign node15770 = (inp[11]) ? 4'b1001 : node15771;
													assign node15771 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node15775 = (inp[9]) ? node15783 : node15776;
													assign node15776 = (inp[5]) ? 4'b1001 : node15777;
														assign node15777 = (inp[2]) ? node15779 : 4'b1101;
															assign node15779 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node15783 = (inp[11]) ? node15785 : 4'b1000;
														assign node15785 = (inp[2]) ? node15789 : node15786;
															assign node15786 = (inp[5]) ? 4'b1101 : 4'b1100;
															assign node15789 = (inp[5]) ? 4'b1100 : 4'b1101;
											assign node15792 = (inp[11]) ? node15812 : node15793;
												assign node15793 = (inp[13]) ? node15799 : node15794;
													assign node15794 = (inp[9]) ? 4'b1001 : node15795;
														assign node15795 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node15799 = (inp[2]) ? node15805 : node15800;
														assign node15800 = (inp[0]) ? 4'b1101 : node15801;
															assign node15801 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node15805 = (inp[9]) ? node15809 : node15806;
															assign node15806 = (inp[5]) ? 4'b1000 : 4'b1001;
															assign node15809 = (inp[5]) ? 4'b1001 : 4'b1000;
												assign node15812 = (inp[5]) ? node15820 : node15813;
													assign node15813 = (inp[9]) ? node15815 : 4'b1000;
														assign node15815 = (inp[2]) ? node15817 : 4'b1000;
															assign node15817 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node15820 = (inp[2]) ? 4'b1000 : node15821;
														assign node15821 = (inp[13]) ? 4'b1100 : 4'b1000;
										assign node15825 = (inp[5]) ? node15867 : node15826;
											assign node15826 = (inp[0]) ? node15848 : node15827;
												assign node15827 = (inp[11]) ? node15837 : node15828;
													assign node15828 = (inp[4]) ? node15830 : 4'b1001;
														assign node15830 = (inp[2]) ? node15834 : node15831;
															assign node15831 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node15834 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node15837 = (inp[9]) ? node15843 : node15838;
														assign node15838 = (inp[2]) ? 4'b1101 : node15839;
															assign node15839 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node15843 = (inp[2]) ? node15845 : 4'b1101;
															assign node15845 = (inp[13]) ? 4'b1101 : 4'b1001;
												assign node15848 = (inp[9]) ? node15856 : node15849;
													assign node15849 = (inp[11]) ? 4'b1001 : node15850;
														assign node15850 = (inp[2]) ? 4'b1100 : node15851;
															assign node15851 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node15856 = (inp[4]) ? node15862 : node15857;
														assign node15857 = (inp[2]) ? 4'b1100 : node15858;
															assign node15858 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node15862 = (inp[2]) ? 4'b1000 : node15863;
															assign node15863 = (inp[13]) ? 4'b1000 : 4'b1100;
											assign node15867 = (inp[2]) ? node15883 : node15868;
												assign node15868 = (inp[13]) ? node15876 : node15869;
													assign node15869 = (inp[0]) ? 4'b1001 : node15870;
														assign node15870 = (inp[9]) ? 4'b1001 : node15871;
															assign node15871 = (inp[4]) ? 4'b1000 : 4'b1001;
													assign node15876 = (inp[9]) ? 4'b1101 : node15877;
														assign node15877 = (inp[4]) ? node15879 : 4'b1100;
															assign node15879 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node15883 = (inp[13]) ? node15891 : node15884;
													assign node15884 = (inp[9]) ? 4'b1100 : node15885;
														assign node15885 = (inp[4]) ? 4'b1101 : node15886;
															assign node15886 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node15891 = (inp[11]) ? node15893 : 4'b1000;
														assign node15893 = (inp[9]) ? 4'b1000 : 4'b1001;
							assign node15896 = (inp[13]) ? node16120 : node15897;
								assign node15897 = (inp[5]) ? node16017 : node15898;
									assign node15898 = (inp[12]) ? node15972 : node15899;
										assign node15899 = (inp[10]) ? node15937 : node15900;
											assign node15900 = (inp[11]) ? node15918 : node15901;
												assign node15901 = (inp[0]) ? node15909 : node15902;
													assign node15902 = (inp[4]) ? node15904 : 4'b1001;
														assign node15904 = (inp[1]) ? node15906 : 4'b1100;
															assign node15906 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node15909 = (inp[9]) ? node15915 : node15910;
														assign node15910 = (inp[4]) ? node15912 : 4'b1000;
															assign node15912 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node15915 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node15918 = (inp[2]) ? node15924 : node15919;
													assign node15919 = (inp[0]) ? node15921 : 4'b1001;
														assign node15921 = (inp[1]) ? 4'b1100 : 4'b1001;
													assign node15924 = (inp[0]) ? node15930 : node15925;
														assign node15925 = (inp[1]) ? node15927 : 4'b1101;
															assign node15927 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node15930 = (inp[1]) ? node15934 : node15931;
															assign node15931 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node15934 = (inp[4]) ? 4'b1001 : 4'b1100;
											assign node15937 = (inp[11]) ? node15957 : node15938;
												assign node15938 = (inp[4]) ? node15948 : node15939;
													assign node15939 = (inp[1]) ? 4'b1100 : node15940;
														assign node15940 = (inp[0]) ? node15944 : node15941;
															assign node15941 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node15944 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node15948 = (inp[1]) ? node15952 : node15949;
														assign node15949 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node15952 = (inp[9]) ? node15954 : 4'b1001;
															assign node15954 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node15957 = (inp[1]) ? node15961 : node15958;
													assign node15958 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node15961 = (inp[4]) ? node15967 : node15962;
														assign node15962 = (inp[9]) ? 4'b1101 : node15963;
															assign node15963 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node15967 = (inp[0]) ? node15969 : 4'b1001;
															assign node15969 = (inp[9]) ? 4'b1000 : 4'b1001;
										assign node15972 = (inp[10]) ? node15994 : node15973;
											assign node15973 = (inp[9]) ? node15987 : node15974;
												assign node15974 = (inp[1]) ? node15980 : node15975;
													assign node15975 = (inp[11]) ? 4'b1000 : node15976;
														assign node15976 = (inp[4]) ? 4'b1001 : 4'b1000;
													assign node15980 = (inp[2]) ? 4'b1001 : node15981;
														assign node15981 = (inp[11]) ? node15983 : 4'b1000;
															assign node15983 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node15987 = (inp[11]) ? 4'b1001 : node15988;
													assign node15988 = (inp[1]) ? 4'b1000 : node15989;
														assign node15989 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node15994 = (inp[4]) ? node16008 : node15995;
												assign node15995 = (inp[0]) ? node16001 : node15996;
													assign node15996 = (inp[9]) ? node15998 : 4'b1001;
														assign node15998 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node16001 = (inp[1]) ? 4'b1001 : node16002;
														assign node16002 = (inp[9]) ? 4'b1000 : node16003;
															assign node16003 = (inp[11]) ? 4'b1000 : 4'b1000;
												assign node16008 = (inp[2]) ? node16010 : 4'b1000;
													assign node16010 = (inp[0]) ? 4'b1000 : node16011;
														assign node16011 = (inp[9]) ? 4'b1001 : node16012;
															assign node16012 = (inp[11]) ? 4'b1000 : 4'b1001;
									assign node16017 = (inp[12]) ? node16077 : node16018;
										assign node16018 = (inp[1]) ? node16052 : node16019;
											assign node16019 = (inp[4]) ? node16033 : node16020;
												assign node16020 = (inp[10]) ? 4'b1100 : node16021;
													assign node16021 = (inp[2]) ? node16029 : node16022;
														assign node16022 = (inp[9]) ? node16026 : node16023;
															assign node16023 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node16026 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node16029 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node16033 = (inp[10]) ? node16043 : node16034;
													assign node16034 = (inp[2]) ? 4'b1001 : node16035;
														assign node16035 = (inp[11]) ? node16039 : node16036;
															assign node16036 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node16039 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node16043 = (inp[2]) ? node16047 : node16044;
														assign node16044 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node16047 = (inp[0]) ? 4'b1000 : node16048;
															assign node16048 = (inp[9]) ? 4'b1001 : 4'b1000;
											assign node16052 = (inp[4]) ? node16068 : node16053;
												assign node16053 = (inp[11]) ? node16063 : node16054;
													assign node16054 = (inp[9]) ? node16058 : node16055;
														assign node16055 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node16058 = (inp[2]) ? node16060 : 4'b1001;
															assign node16060 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node16063 = (inp[0]) ? node16065 : 4'b1000;
														assign node16065 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node16068 = (inp[10]) ? node16070 : 4'b1101;
													assign node16070 = (inp[11]) ? 4'b1100 : node16071;
														assign node16071 = (inp[0]) ? node16073 : 4'b1101;
															assign node16073 = (inp[9]) ? 4'b1101 : 4'b1100;
										assign node16077 = (inp[0]) ? node16095 : node16078;
											assign node16078 = (inp[2]) ? node16088 : node16079;
												assign node16079 = (inp[4]) ? node16083 : node16080;
													assign node16080 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node16083 = (inp[9]) ? 4'b1100 : node16084;
														assign node16084 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node16088 = (inp[11]) ? node16092 : node16089;
													assign node16089 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node16092 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node16095 = (inp[2]) ? node16105 : node16096;
												assign node16096 = (inp[10]) ? node16100 : node16097;
													assign node16097 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node16100 = (inp[11]) ? node16102 : 4'b1101;
														assign node16102 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node16105 = (inp[10]) ? node16115 : node16106;
													assign node16106 = (inp[1]) ? 4'b1101 : node16107;
														assign node16107 = (inp[9]) ? node16111 : node16108;
															assign node16108 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node16111 = (inp[4]) ? 4'b1100 : 4'b1101;
													assign node16115 = (inp[11]) ? 4'b1100 : node16116;
														assign node16116 = (inp[9]) ? 4'b1101 : 4'b1100;
								assign node16120 = (inp[5]) ? node16236 : node16121;
									assign node16121 = (inp[12]) ? node16187 : node16122;
										assign node16122 = (inp[2]) ? node16160 : node16123;
											assign node16123 = (inp[9]) ? node16137 : node16124;
												assign node16124 = (inp[4]) ? node16134 : node16125;
													assign node16125 = (inp[1]) ? node16129 : node16126;
														assign node16126 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node16129 = (inp[0]) ? 4'b1001 : node16130;
															assign node16130 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node16134 = (inp[1]) ? 4'b1101 : 4'b1001;
												assign node16137 = (inp[0]) ? node16149 : node16138;
													assign node16138 = (inp[10]) ? node16146 : node16139;
														assign node16139 = (inp[11]) ? node16143 : node16140;
															assign node16140 = (inp[1]) ? 4'b1100 : 4'b1001;
															assign node16143 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node16146 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node16149 = (inp[11]) ? node16157 : node16150;
														assign node16150 = (inp[1]) ? node16154 : node16151;
															assign node16151 = (inp[10]) ? 4'b1001 : 4'b1100;
															assign node16154 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node16157 = (inp[4]) ? 4'b1100 : 4'b1101;
											assign node16160 = (inp[10]) ? node16170 : node16161;
												assign node16161 = (inp[1]) ? node16165 : node16162;
													assign node16162 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node16165 = (inp[4]) ? node16167 : 4'b1000;
														assign node16167 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node16170 = (inp[11]) ? node16182 : node16171;
													assign node16171 = (inp[1]) ? node16177 : node16172;
														assign node16172 = (inp[4]) ? 4'b1000 : node16173;
															assign node16173 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node16177 = (inp[4]) ? 4'b1101 : node16178;
															assign node16178 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node16182 = (inp[0]) ? node16184 : 4'b1000;
														assign node16184 = (inp[9]) ? 4'b1100 : 4'b1101;
										assign node16187 = (inp[1]) ? node16211 : node16188;
											assign node16188 = (inp[0]) ? node16204 : node16189;
												assign node16189 = (inp[10]) ? node16197 : node16190;
													assign node16190 = (inp[9]) ? 4'b1100 : node16191;
														assign node16191 = (inp[2]) ? node16193 : 4'b1100;
															assign node16193 = (inp[4]) ? 4'b1100 : 4'b1100;
													assign node16197 = (inp[9]) ? node16199 : 4'b1100;
														assign node16199 = (inp[11]) ? node16201 : 4'b1101;
															assign node16201 = (inp[2]) ? 4'b1100 : 4'b1100;
												assign node16204 = (inp[11]) ? node16208 : node16205;
													assign node16205 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node16208 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node16211 = (inp[11]) ? node16225 : node16212;
												assign node16212 = (inp[4]) ? node16220 : node16213;
													assign node16213 = (inp[9]) ? 4'b1100 : node16214;
														assign node16214 = (inp[2]) ? node16216 : 4'b1100;
															assign node16216 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node16220 = (inp[9]) ? 4'b1101 : node16221;
														assign node16221 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node16225 = (inp[9]) ? node16233 : node16226;
													assign node16226 = (inp[0]) ? 4'b1101 : node16227;
														assign node16227 = (inp[4]) ? 4'b1101 : node16228;
															assign node16228 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node16233 = (inp[2]) ? 4'b1101 : 4'b1100;
									assign node16236 = (inp[12]) ? node16288 : node16237;
										assign node16237 = (inp[1]) ? node16263 : node16238;
											assign node16238 = (inp[4]) ? node16248 : node16239;
												assign node16239 = (inp[2]) ? node16245 : node16240;
													assign node16240 = (inp[9]) ? node16242 : 4'b1001;
														assign node16242 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node16245 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node16248 = (inp[9]) ? node16260 : node16249;
													assign node16249 = (inp[0]) ? node16257 : node16250;
														assign node16250 = (inp[11]) ? node16254 : node16251;
															assign node16251 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node16254 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node16257 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node16260 = (inp[11]) ? 4'b1101 : 4'b1100;
											assign node16263 = (inp[4]) ? node16275 : node16264;
												assign node16264 = (inp[0]) ? node16266 : 4'b1101;
													assign node16266 = (inp[9]) ? 4'b1100 : node16267;
														assign node16267 = (inp[11]) ? node16271 : node16268;
															assign node16268 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node16271 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node16275 = (inp[0]) ? node16283 : node16276;
													assign node16276 = (inp[2]) ? node16278 : 4'b1001;
														assign node16278 = (inp[9]) ? node16280 : 4'b1000;
															assign node16280 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node16283 = (inp[11]) ? node16285 : 4'b1000;
														assign node16285 = (inp[9]) ? 4'b1000 : 4'b1001;
										assign node16288 = (inp[11]) ? node16306 : node16289;
											assign node16289 = (inp[0]) ? node16297 : node16290;
												assign node16290 = (inp[10]) ? node16292 : 4'b1000;
													assign node16292 = (inp[2]) ? 4'b1000 : node16293;
														assign node16293 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node16297 = (inp[9]) ? node16301 : node16298;
													assign node16298 = (inp[4]) ? 4'b1000 : 4'b1001;
													assign node16301 = (inp[4]) ? 4'b1001 : node16302;
														assign node16302 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node16306 = (inp[9]) ? node16310 : node16307;
												assign node16307 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node16310 = (inp[2]) ? 4'b1000 : node16311;
													assign node16311 = (inp[0]) ? 4'b1001 : 4'b1000;
				assign node16315 = (inp[7]) ? node17931 : node16316;
					assign node16316 = (inp[6]) ? node17254 : node16317;
						assign node16317 = (inp[12]) ? node16807 : node16318;
							assign node16318 = (inp[15]) ? node16550 : node16319;
								assign node16319 = (inp[4]) ? node16449 : node16320;
									assign node16320 = (inp[0]) ? node16392 : node16321;
										assign node16321 = (inp[5]) ? node16357 : node16322;
											assign node16322 = (inp[10]) ? node16336 : node16323;
												assign node16323 = (inp[1]) ? node16333 : node16324;
													assign node16324 = (inp[9]) ? node16328 : node16325;
														assign node16325 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node16328 = (inp[2]) ? node16330 : 4'b0111;
															assign node16330 = (inp[13]) ? 4'b0010 : 4'b0111;
													assign node16333 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node16336 = (inp[13]) ? node16342 : node16337;
													assign node16337 = (inp[11]) ? 4'b0010 : node16338;
														assign node16338 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node16342 = (inp[11]) ? node16350 : node16343;
														assign node16343 = (inp[1]) ? node16347 : node16344;
															assign node16344 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node16347 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node16350 = (inp[9]) ? node16354 : node16351;
															assign node16351 = (inp[2]) ? 4'b0010 : 4'b0111;
															assign node16354 = (inp[2]) ? 4'b0111 : 4'b0010;
											assign node16357 = (inp[11]) ? node16373 : node16358;
												assign node16358 = (inp[13]) ? node16368 : node16359;
													assign node16359 = (inp[2]) ? 4'b0011 : node16360;
														assign node16360 = (inp[9]) ? node16364 : node16361;
															assign node16361 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node16364 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node16368 = (inp[9]) ? node16370 : 4'b0011;
														assign node16370 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node16373 = (inp[10]) ? node16385 : node16374;
													assign node16374 = (inp[1]) ? node16378 : node16375;
														assign node16375 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node16378 = (inp[13]) ? node16382 : node16379;
															assign node16379 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node16382 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node16385 = (inp[1]) ? 4'b0010 : node16386;
														assign node16386 = (inp[9]) ? 4'b0010 : node16387;
															assign node16387 = (inp[2]) ? 4'b0010 : 4'b0110;
										assign node16392 = (inp[2]) ? node16424 : node16393;
											assign node16393 = (inp[13]) ? node16409 : node16394;
												assign node16394 = (inp[1]) ? node16400 : node16395;
													assign node16395 = (inp[5]) ? node16397 : 4'b0010;
														assign node16397 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node16400 = (inp[10]) ? node16406 : node16401;
														assign node16401 = (inp[11]) ? 4'b0110 : node16402;
															assign node16402 = (inp[5]) ? 4'b0110 : 4'b0110;
														assign node16406 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node16409 = (inp[5]) ? node16417 : node16410;
													assign node16410 = (inp[1]) ? 4'b0010 : node16411;
														assign node16411 = (inp[11]) ? 4'b0110 : node16412;
															assign node16412 = (inp[9]) ? 4'b0110 : 4'b0110;
													assign node16417 = (inp[1]) ? node16419 : 4'b0010;
														assign node16419 = (inp[10]) ? 4'b0010 : node16420;
															assign node16420 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node16424 = (inp[13]) ? node16434 : node16425;
												assign node16425 = (inp[9]) ? node16431 : node16426;
													assign node16426 = (inp[1]) ? node16428 : 4'b0110;
														assign node16428 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node16431 = (inp[11]) ? 4'b0011 : 4'b0111;
												assign node16434 = (inp[5]) ? node16444 : node16435;
													assign node16435 = (inp[1]) ? node16439 : node16436;
														assign node16436 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node16439 = (inp[10]) ? 4'b0111 : node16440;
															assign node16440 = (inp[11]) ? 4'b0110 : 4'b0110;
													assign node16444 = (inp[10]) ? 4'b0110 : node16445;
														assign node16445 = (inp[9]) ? 4'b0110 : 4'b0111;
									assign node16449 = (inp[9]) ? node16493 : node16450;
										assign node16450 = (inp[2]) ? node16466 : node16451;
											assign node16451 = (inp[13]) ? node16459 : node16452;
												assign node16452 = (inp[11]) ? node16454 : 4'b0000;
													assign node16454 = (inp[10]) ? node16456 : 4'b0001;
														assign node16456 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node16459 = (inp[5]) ? node16461 : 4'b0100;
													assign node16461 = (inp[1]) ? node16463 : 4'b0101;
														assign node16463 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node16466 = (inp[13]) ? node16482 : node16467;
												assign node16467 = (inp[5]) ? node16477 : node16468;
													assign node16468 = (inp[1]) ? 4'b0101 : node16469;
														assign node16469 = (inp[11]) ? node16473 : node16470;
															assign node16470 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node16473 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node16477 = (inp[1]) ? 4'b0000 : node16478;
														assign node16478 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node16482 = (inp[5]) ? node16486 : node16483;
													assign node16483 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node16486 = (inp[1]) ? node16490 : node16487;
														assign node16487 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node16490 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node16493 = (inp[2]) ? node16523 : node16494;
											assign node16494 = (inp[13]) ? node16510 : node16495;
												assign node16495 = (inp[1]) ? node16501 : node16496;
													assign node16496 = (inp[11]) ? 4'b0000 : node16497;
														assign node16497 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node16501 = (inp[5]) ? node16503 : 4'b0000;
														assign node16503 = (inp[11]) ? node16507 : node16504;
															assign node16504 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node16507 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node16510 = (inp[5]) ? node16520 : node16511;
													assign node16511 = (inp[0]) ? node16515 : node16512;
														assign node16512 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node16515 = (inp[1]) ? 4'b0100 : node16516;
															assign node16516 = (inp[11]) ? 4'b0100 : 4'b0100;
													assign node16520 = (inp[1]) ? 4'b0001 : 4'b0101;
											assign node16523 = (inp[13]) ? node16537 : node16524;
												assign node16524 = (inp[1]) ? node16532 : node16525;
													assign node16525 = (inp[10]) ? node16527 : 4'b0100;
														assign node16527 = (inp[0]) ? 4'b0101 : node16528;
															assign node16528 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node16532 = (inp[5]) ? node16534 : 4'b0101;
														assign node16534 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node16537 = (inp[1]) ? node16545 : node16538;
													assign node16538 = (inp[0]) ? 4'b0001 : node16539;
														assign node16539 = (inp[5]) ? 4'b0000 : node16540;
															assign node16540 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node16545 = (inp[10]) ? node16547 : 4'b0001;
														assign node16547 = (inp[11]) ? 4'b0100 : 4'b0101;
								assign node16550 = (inp[9]) ? node16670 : node16551;
									assign node16551 = (inp[10]) ? node16611 : node16552;
										assign node16552 = (inp[2]) ? node16584 : node16553;
											assign node16553 = (inp[1]) ? node16569 : node16554;
												assign node16554 = (inp[11]) ? node16562 : node16555;
													assign node16555 = (inp[0]) ? node16557 : 4'b0000;
														assign node16557 = (inp[4]) ? 4'b0101 : node16558;
															assign node16558 = (inp[13]) ? 4'b0101 : 4'b0000;
													assign node16562 = (inp[4]) ? node16566 : node16563;
														assign node16563 = (inp[5]) ? 4'b0101 : 4'b0001;
														assign node16566 = (inp[0]) ? 4'b0000 : 4'b0101;
												assign node16569 = (inp[11]) ? node16577 : node16570;
													assign node16570 = (inp[4]) ? node16572 : 4'b0000;
														assign node16572 = (inp[5]) ? node16574 : 4'b0000;
															assign node16574 = (inp[13]) ? 4'b0101 : 4'b0000;
													assign node16577 = (inp[13]) ? node16579 : 4'b0100;
														assign node16579 = (inp[5]) ? 4'b0000 : node16580;
															assign node16580 = (inp[4]) ? 4'b0000 : 4'b0101;
											assign node16584 = (inp[11]) ? node16598 : node16585;
												assign node16585 = (inp[1]) ? node16595 : node16586;
													assign node16586 = (inp[13]) ? node16592 : node16587;
														assign node16587 = (inp[4]) ? node16589 : 4'b0101;
															assign node16589 = (inp[5]) ? 4'b0000 : 4'b0000;
														assign node16592 = (inp[4]) ? 4'b0101 : 4'b0000;
													assign node16595 = (inp[13]) ? 4'b0001 : 4'b0101;
												assign node16598 = (inp[13]) ? node16608 : node16599;
													assign node16599 = (inp[5]) ? node16605 : node16600;
														assign node16600 = (inp[1]) ? 4'b0000 : node16601;
															assign node16601 = (inp[0]) ? 4'b0101 : 4'b0001;
														assign node16605 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node16608 = (inp[5]) ? 4'b0000 : 4'b0001;
										assign node16611 = (inp[11]) ? node16641 : node16612;
											assign node16612 = (inp[1]) ? node16622 : node16613;
												assign node16613 = (inp[4]) ? node16619 : node16614;
													assign node16614 = (inp[2]) ? node16616 : 4'b0001;
														assign node16616 = (inp[0]) ? 4'b0101 : 4'b0001;
													assign node16619 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node16622 = (inp[2]) ? node16634 : node16623;
													assign node16623 = (inp[13]) ? node16631 : node16624;
														assign node16624 = (inp[5]) ? node16628 : node16625;
															assign node16625 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node16628 = (inp[4]) ? 4'b0000 : 4'b0101;
														assign node16631 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node16634 = (inp[5]) ? 4'b0100 : node16635;
														assign node16635 = (inp[0]) ? 4'b0100 : node16636;
															assign node16636 = (inp[13]) ? 4'b0000 : 4'b0000;
											assign node16641 = (inp[1]) ? node16653 : node16642;
												assign node16642 = (inp[5]) ? node16646 : node16643;
													assign node16643 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node16646 = (inp[2]) ? node16650 : node16647;
														assign node16647 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node16650 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node16653 = (inp[4]) ? node16661 : node16654;
													assign node16654 = (inp[5]) ? node16658 : node16655;
														assign node16655 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node16658 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node16661 = (inp[5]) ? node16667 : node16662;
														assign node16662 = (inp[2]) ? 4'b0001 : node16663;
															assign node16663 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node16667 = (inp[13]) ? 4'b0001 : 4'b0000;
									assign node16670 = (inp[5]) ? node16752 : node16671;
										assign node16671 = (inp[11]) ? node16707 : node16672;
											assign node16672 = (inp[13]) ? node16686 : node16673;
												assign node16673 = (inp[10]) ? node16675 : 4'b0101;
													assign node16675 = (inp[0]) ? node16681 : node16676;
														assign node16676 = (inp[1]) ? node16678 : 4'b0100;
															assign node16678 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node16681 = (inp[4]) ? 4'b0001 : node16682;
															assign node16682 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node16686 = (inp[1]) ? node16696 : node16687;
													assign node16687 = (inp[2]) ? node16691 : node16688;
														assign node16688 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node16691 = (inp[4]) ? node16693 : 4'b0001;
															assign node16693 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node16696 = (inp[10]) ? node16702 : node16697;
														assign node16697 = (inp[2]) ? node16699 : 4'b0101;
															assign node16699 = (inp[4]) ? 4'b0101 : 4'b0000;
														assign node16702 = (inp[0]) ? 4'b0100 : node16703;
															assign node16703 = (inp[4]) ? 4'b0001 : 4'b0100;
											assign node16707 = (inp[0]) ? node16731 : node16708;
												assign node16708 = (inp[2]) ? node16718 : node16709;
													assign node16709 = (inp[1]) ? node16713 : node16710;
														assign node16710 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node16713 = (inp[10]) ? 4'b0000 : node16714;
															assign node16714 = (inp[4]) ? 4'b0001 : 4'b0001;
													assign node16718 = (inp[1]) ? node16724 : node16719;
														assign node16719 = (inp[10]) ? 4'b0101 : node16720;
															assign node16720 = (inp[4]) ? 4'b0000 : 4'b0101;
														assign node16724 = (inp[4]) ? node16728 : node16725;
															assign node16725 = (inp[10]) ? 4'b0101 : 4'b0000;
															assign node16728 = (inp[13]) ? 4'b0100 : 4'b0000;
												assign node16731 = (inp[13]) ? node16741 : node16732;
													assign node16732 = (inp[4]) ? node16736 : node16733;
														assign node16733 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node16736 = (inp[10]) ? node16738 : 4'b0100;
															assign node16738 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node16741 = (inp[2]) ? node16745 : node16742;
														assign node16742 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node16745 = (inp[4]) ? node16749 : node16746;
															assign node16746 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node16749 = (inp[1]) ? 4'b0101 : 4'b0100;
										assign node16752 = (inp[11]) ? node16784 : node16753;
											assign node16753 = (inp[10]) ? node16771 : node16754;
												assign node16754 = (inp[4]) ? node16764 : node16755;
													assign node16755 = (inp[13]) ? node16759 : node16756;
														assign node16756 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node16759 = (inp[1]) ? 4'b0100 : node16760;
															assign node16760 = (inp[0]) ? 4'b0100 : 4'b0000;
													assign node16764 = (inp[13]) ? 4'b0000 : node16765;
														assign node16765 = (inp[0]) ? 4'b0001 : node16766;
															assign node16766 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node16771 = (inp[1]) ? node16775 : node16772;
													assign node16772 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node16775 = (inp[13]) ? node16777 : 4'b0001;
														assign node16777 = (inp[4]) ? node16781 : node16778;
															assign node16778 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node16781 = (inp[2]) ? 4'b0001 : 4'b0101;
											assign node16784 = (inp[10]) ? node16800 : node16785;
												assign node16785 = (inp[0]) ? node16793 : node16786;
													assign node16786 = (inp[4]) ? node16790 : node16787;
														assign node16787 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node16790 = (inp[2]) ? 4'b0101 : 4'b0001;
													assign node16793 = (inp[4]) ? 4'b0101 : node16794;
														assign node16794 = (inp[13]) ? node16796 : 4'b0000;
															assign node16796 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node16800 = (inp[1]) ? node16804 : node16801;
													assign node16801 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node16804 = (inp[2]) ? 4'b0000 : 4'b0100;
							assign node16807 = (inp[4]) ? node17015 : node16808;
								assign node16808 = (inp[15]) ? node16914 : node16809;
									assign node16809 = (inp[10]) ? node16859 : node16810;
										assign node16810 = (inp[2]) ? node16840 : node16811;
											assign node16811 = (inp[13]) ? node16823 : node16812;
												assign node16812 = (inp[5]) ? 4'b0001 : node16813;
													assign node16813 = (inp[1]) ? node16819 : node16814;
														assign node16814 = (inp[11]) ? node16816 : 4'b0100;
															assign node16816 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node16819 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node16823 = (inp[11]) ? node16831 : node16824;
													assign node16824 = (inp[9]) ? 4'b0101 : node16825;
														assign node16825 = (inp[1]) ? node16827 : 4'b0101;
															assign node16827 = (inp[5]) ? 4'b0100 : 4'b0100;
													assign node16831 = (inp[1]) ? node16835 : node16832;
														assign node16832 = (inp[5]) ? 4'b0100 : 4'b0000;
														assign node16835 = (inp[0]) ? 4'b0100 : node16836;
															assign node16836 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node16840 = (inp[13]) ? node16850 : node16841;
												assign node16841 = (inp[0]) ? 4'b0101 : node16842;
													assign node16842 = (inp[1]) ? node16846 : node16843;
														assign node16843 = (inp[5]) ? 4'b0100 : 4'b0000;
														assign node16846 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node16850 = (inp[5]) ? 4'b0000 : node16851;
													assign node16851 = (inp[1]) ? 4'b0000 : node16852;
														assign node16852 = (inp[0]) ? node16854 : 4'b0100;
															assign node16854 = (inp[9]) ? 4'b0100 : 4'b0100;
										assign node16859 = (inp[1]) ? node16885 : node16860;
											assign node16860 = (inp[11]) ? node16868 : node16861;
												assign node16861 = (inp[9]) ? node16863 : 4'b0001;
													assign node16863 = (inp[5]) ? node16865 : 4'b0101;
														assign node16865 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node16868 = (inp[0]) ? node16872 : node16869;
													assign node16869 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node16872 = (inp[2]) ? node16880 : node16873;
														assign node16873 = (inp[9]) ? node16877 : node16874;
															assign node16874 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node16877 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node16880 = (inp[5]) ? node16882 : 4'b0101;
															assign node16882 = (inp[13]) ? 4'b0000 : 4'b0100;
											assign node16885 = (inp[0]) ? node16895 : node16886;
												assign node16886 = (inp[13]) ? node16892 : node16887;
													assign node16887 = (inp[2]) ? node16889 : 4'b0000;
														assign node16889 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node16892 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node16895 = (inp[9]) ? node16907 : node16896;
													assign node16896 = (inp[2]) ? node16904 : node16897;
														assign node16897 = (inp[13]) ? node16901 : node16898;
															assign node16898 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node16901 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node16904 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node16907 = (inp[5]) ? node16909 : 4'b0000;
														assign node16909 = (inp[11]) ? node16911 : 4'b0001;
															assign node16911 = (inp[13]) ? 4'b0101 : 4'b0001;
									assign node16914 = (inp[0]) ? node16968 : node16915;
										assign node16915 = (inp[5]) ? node16951 : node16916;
											assign node16916 = (inp[11]) ? node16940 : node16917;
												assign node16917 = (inp[1]) ? node16925 : node16918;
													assign node16918 = (inp[13]) ? node16922 : node16919;
														assign node16919 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node16922 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node16925 = (inp[9]) ? node16933 : node16926;
														assign node16926 = (inp[10]) ? node16930 : node16927;
															assign node16927 = (inp[2]) ? 4'b0010 : 4'b0111;
															assign node16930 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node16933 = (inp[2]) ? node16937 : node16934;
															assign node16934 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node16937 = (inp[13]) ? 4'b0011 : 4'b0110;
												assign node16940 = (inp[2]) ? node16946 : node16941;
													assign node16941 = (inp[9]) ? 4'b0110 : node16942;
														assign node16942 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node16946 = (inp[9]) ? 4'b0110 : node16947;
														assign node16947 = (inp[1]) ? 4'b0110 : 4'b0010;
											assign node16951 = (inp[10]) ? node16959 : node16952;
												assign node16952 = (inp[1]) ? node16956 : node16953;
													assign node16953 = (inp[13]) ? 4'b0111 : 4'b0010;
													assign node16956 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node16959 = (inp[2]) ? node16965 : node16960;
													assign node16960 = (inp[13]) ? 4'b0111 : node16961;
														assign node16961 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node16965 = (inp[13]) ? 4'b0011 : 4'b0111;
										assign node16968 = (inp[10]) ? node16994 : node16969;
											assign node16969 = (inp[9]) ? node16981 : node16970;
												assign node16970 = (inp[11]) ? node16972 : 4'b0110;
													assign node16972 = (inp[2]) ? node16978 : node16973;
														assign node16973 = (inp[13]) ? node16975 : 4'b0011;
															assign node16975 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node16978 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node16981 = (inp[13]) ? node16985 : node16982;
													assign node16982 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node16985 = (inp[2]) ? node16989 : node16986;
														assign node16986 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node16989 = (inp[1]) ? node16991 : 4'b0111;
															assign node16991 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node16994 = (inp[11]) ? node17000 : node16995;
												assign node16995 = (inp[9]) ? node16997 : 4'b0011;
													assign node16997 = (inp[5]) ? 4'b0111 : 4'b0011;
												assign node17000 = (inp[1]) ? node17008 : node17001;
													assign node17001 = (inp[9]) ? node17005 : node17002;
														assign node17002 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node17005 = (inp[5]) ? 4'b0011 : 4'b0111;
													assign node17008 = (inp[9]) ? 4'b0011 : node17009;
														assign node17009 = (inp[5]) ? 4'b0110 : node17010;
															assign node17010 = (inp[13]) ? 4'b0111 : 4'b0110;
								assign node17015 = (inp[1]) ? node17131 : node17016;
									assign node17016 = (inp[5]) ? node17080 : node17017;
										assign node17017 = (inp[10]) ? node17041 : node17018;
											assign node17018 = (inp[2]) ? node17032 : node17019;
												assign node17019 = (inp[13]) ? node17027 : node17020;
													assign node17020 = (inp[15]) ? 4'b0110 : node17021;
														assign node17021 = (inp[11]) ? node17023 : 4'b0010;
															assign node17023 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node17027 = (inp[15]) ? 4'b0010 : node17028;
														assign node17028 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node17032 = (inp[9]) ? 4'b0110 : node17033;
													assign node17033 = (inp[13]) ? node17035 : 4'b0111;
														assign node17035 = (inp[0]) ? 4'b0010 : node17036;
															assign node17036 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node17041 = (inp[9]) ? node17065 : node17042;
												assign node17042 = (inp[0]) ? node17054 : node17043;
													assign node17043 = (inp[2]) ? node17051 : node17044;
														assign node17044 = (inp[13]) ? node17048 : node17045;
															assign node17045 = (inp[15]) ? 4'b0111 : 4'b0011;
															assign node17048 = (inp[15]) ? 4'b0011 : 4'b0111;
														assign node17051 = (inp[15]) ? 4'b0011 : 4'b0110;
													assign node17054 = (inp[15]) ? node17060 : node17055;
														assign node17055 = (inp[11]) ? node17057 : 4'b0110;
															assign node17057 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node17060 = (inp[11]) ? node17062 : 4'b0011;
															assign node17062 = (inp[2]) ? 4'b0010 : 4'b0010;
												assign node17065 = (inp[2]) ? node17077 : node17066;
													assign node17066 = (inp[11]) ? node17072 : node17067;
														assign node17067 = (inp[15]) ? 4'b0010 : node17068;
															assign node17068 = (inp[13]) ? 4'b0110 : 4'b0010;
														assign node17072 = (inp[0]) ? node17074 : 4'b0010;
															assign node17074 = (inp[15]) ? 4'b0111 : 4'b0011;
													assign node17077 = (inp[11]) ? 4'b0011 : 4'b0111;
										assign node17080 = (inp[2]) ? node17106 : node17081;
											assign node17081 = (inp[15]) ? node17097 : node17082;
												assign node17082 = (inp[13]) ? 4'b0010 : node17083;
													assign node17083 = (inp[10]) ? node17091 : node17084;
														assign node17084 = (inp[0]) ? node17088 : node17085;
															assign node17085 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node17088 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node17091 = (inp[0]) ? node17093 : 4'b0110;
															assign node17093 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node17097 = (inp[13]) ? 4'b0111 : node17098;
													assign node17098 = (inp[10]) ? 4'b0010 : node17099;
														assign node17099 = (inp[9]) ? node17101 : 4'b0011;
															assign node17101 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node17106 = (inp[0]) ? node17124 : node17107;
												assign node17107 = (inp[9]) ? node17117 : node17108;
													assign node17108 = (inp[13]) ? node17114 : node17109;
														assign node17109 = (inp[15]) ? 4'b0111 : node17110;
															assign node17110 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node17114 = (inp[15]) ? 4'b0011 : 4'b0111;
													assign node17117 = (inp[13]) ? 4'b0110 : node17118;
														assign node17118 = (inp[11]) ? 4'b0110 : node17119;
															assign node17119 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node17124 = (inp[11]) ? node17126 : 4'b0010;
													assign node17126 = (inp[15]) ? node17128 : 4'b0011;
														assign node17128 = (inp[10]) ? 4'b0111 : 4'b0011;
									assign node17131 = (inp[11]) ? node17199 : node17132;
										assign node17132 = (inp[0]) ? node17168 : node17133;
											assign node17133 = (inp[15]) ? node17155 : node17134;
												assign node17134 = (inp[10]) ? node17144 : node17135;
													assign node17135 = (inp[9]) ? 4'b0011 : node17136;
														assign node17136 = (inp[5]) ? node17140 : node17137;
															assign node17137 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node17140 = (inp[2]) ? 4'b0111 : 4'b0011;
													assign node17144 = (inp[2]) ? node17150 : node17145;
														assign node17145 = (inp[13]) ? 4'b0011 : node17146;
															assign node17146 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node17150 = (inp[13]) ? 4'b0111 : node17151;
															assign node17151 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node17155 = (inp[5]) ? 4'b0010 : node17156;
													assign node17156 = (inp[9]) ? node17162 : node17157;
														assign node17157 = (inp[10]) ? 4'b0011 : node17158;
															assign node17158 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node17162 = (inp[10]) ? node17164 : 4'b0011;
															assign node17164 = (inp[13]) ? 4'b0110 : 4'b0010;
											assign node17168 = (inp[5]) ? node17186 : node17169;
												assign node17169 = (inp[15]) ? node17175 : node17170;
													assign node17170 = (inp[2]) ? node17172 : 4'b0010;
														assign node17172 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node17175 = (inp[10]) ? node17179 : node17176;
														assign node17176 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node17179 = (inp[9]) ? node17183 : node17180;
															assign node17180 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node17183 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node17186 = (inp[2]) ? node17192 : node17187;
													assign node17187 = (inp[9]) ? 4'b0010 : node17188;
														assign node17188 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node17192 = (inp[10]) ? 4'b0111 : node17193;
														assign node17193 = (inp[9]) ? node17195 : 4'b0010;
															assign node17195 = (inp[13]) ? 4'b0011 : 4'b0011;
										assign node17199 = (inp[9]) ? node17227 : node17200;
											assign node17200 = (inp[15]) ? node17212 : node17201;
												assign node17201 = (inp[5]) ? 4'b0110 : node17202;
													assign node17202 = (inp[10]) ? node17208 : node17203;
														assign node17203 = (inp[13]) ? 4'b0111 : node17204;
															assign node17204 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node17208 = (inp[2]) ? 4'b0110 : 4'b0011;
												assign node17212 = (inp[0]) ? node17218 : node17213;
													assign node17213 = (inp[10]) ? node17215 : 4'b0010;
														assign node17215 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node17218 = (inp[5]) ? node17222 : node17219;
														assign node17219 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node17222 = (inp[13]) ? node17224 : 4'b0011;
															assign node17224 = (inp[2]) ? 4'b0010 : 4'b0110;
											assign node17227 = (inp[13]) ? node17241 : node17228;
												assign node17228 = (inp[2]) ? node17236 : node17229;
													assign node17229 = (inp[15]) ? node17231 : 4'b0110;
														assign node17231 = (inp[5]) ? 4'b0010 : node17232;
															assign node17232 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node17236 = (inp[15]) ? 4'b0110 : node17237;
														assign node17237 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node17241 = (inp[0]) ? node17245 : node17242;
													assign node17242 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node17245 = (inp[10]) ? node17249 : node17246;
														assign node17246 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node17249 = (inp[15]) ? node17251 : 4'b0111;
															assign node17251 = (inp[2]) ? 4'b0011 : 4'b0111;
						assign node17254 = (inp[15]) ? node17620 : node17255;
							assign node17255 = (inp[13]) ? node17473 : node17256;
								assign node17256 = (inp[4]) ? node17362 : node17257;
									assign node17257 = (inp[0]) ? node17305 : node17258;
										assign node17258 = (inp[5]) ? node17282 : node17259;
											assign node17259 = (inp[12]) ? node17271 : node17260;
												assign node17260 = (inp[1]) ? node17264 : node17261;
													assign node17261 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node17264 = (inp[2]) ? node17268 : node17265;
														assign node17265 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node17268 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node17271 = (inp[1]) ? node17277 : node17272;
													assign node17272 = (inp[10]) ? node17274 : 4'b0110;
														assign node17274 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node17277 = (inp[9]) ? node17279 : 4'b0011;
														assign node17279 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node17282 = (inp[2]) ? node17294 : node17283;
												assign node17283 = (inp[9]) ? node17291 : node17284;
													assign node17284 = (inp[10]) ? node17286 : 4'b0010;
														assign node17286 = (inp[11]) ? node17288 : 4'b0010;
															assign node17288 = (inp[1]) ? 4'b0010 : 4'b0010;
													assign node17291 = (inp[11]) ? 4'b0011 : 4'b0111;
												assign node17294 = (inp[9]) ? node17300 : node17295;
													assign node17295 = (inp[1]) ? 4'b0011 : node17296;
														assign node17296 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node17300 = (inp[12]) ? 4'b0010 : node17301;
														assign node17301 = (inp[10]) ? 4'b0010 : 4'b0110;
										assign node17305 = (inp[12]) ? node17335 : node17306;
											assign node17306 = (inp[1]) ? node17320 : node17307;
												assign node17307 = (inp[2]) ? node17313 : node17308;
													assign node17308 = (inp[11]) ? node17310 : 4'b0010;
														assign node17310 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node17313 = (inp[5]) ? node17317 : node17314;
														assign node17314 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node17317 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node17320 = (inp[10]) ? node17328 : node17321;
													assign node17321 = (inp[9]) ? 4'b0110 : node17322;
														assign node17322 = (inp[5]) ? 4'b0111 : node17323;
															assign node17323 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node17328 = (inp[2]) ? node17330 : 4'b0110;
														assign node17330 = (inp[5]) ? node17332 : 4'b0110;
															assign node17332 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node17335 = (inp[1]) ? node17355 : node17336;
												assign node17336 = (inp[5]) ? node17344 : node17337;
													assign node17337 = (inp[10]) ? node17341 : node17338;
														assign node17338 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node17341 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node17344 = (inp[10]) ? node17350 : node17345;
														assign node17345 = (inp[9]) ? node17347 : 4'b0110;
															assign node17347 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node17350 = (inp[2]) ? node17352 : 4'b0110;
															assign node17352 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node17355 = (inp[2]) ? node17359 : node17356;
													assign node17356 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node17359 = (inp[9]) ? 4'b0011 : 4'b0010;
									assign node17362 = (inp[10]) ? node17408 : node17363;
										assign node17363 = (inp[1]) ? node17383 : node17364;
											assign node17364 = (inp[5]) ? node17374 : node17365;
												assign node17365 = (inp[9]) ? node17371 : node17366;
													assign node17366 = (inp[0]) ? node17368 : 4'b0010;
														assign node17368 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node17371 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node17374 = (inp[12]) ? 4'b0011 : node17375;
													assign node17375 = (inp[9]) ? node17379 : node17376;
														assign node17376 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node17379 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node17383 = (inp[11]) ? node17399 : node17384;
												assign node17384 = (inp[12]) ? node17392 : node17385;
													assign node17385 = (inp[9]) ? node17389 : node17386;
														assign node17386 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node17389 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node17392 = (inp[9]) ? node17394 : 4'b0011;
														assign node17394 = (inp[5]) ? 4'b0011 : node17395;
															assign node17395 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node17399 = (inp[12]) ? node17403 : node17400;
													assign node17400 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node17403 = (inp[9]) ? node17405 : 4'b0010;
														assign node17405 = (inp[0]) ? 4'b0011 : 4'b0010;
										assign node17408 = (inp[0]) ? node17434 : node17409;
											assign node17409 = (inp[1]) ? node17421 : node17410;
												assign node17410 = (inp[11]) ? 4'b0010 : node17411;
													assign node17411 = (inp[2]) ? node17415 : node17412;
														assign node17412 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node17415 = (inp[5]) ? node17417 : 4'b0010;
															assign node17417 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node17421 = (inp[11]) ? node17429 : node17422;
													assign node17422 = (inp[9]) ? node17426 : node17423;
														assign node17423 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node17426 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node17429 = (inp[5]) ? 4'b0011 : node17430;
														assign node17430 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node17434 = (inp[12]) ? node17454 : node17435;
												assign node17435 = (inp[11]) ? node17445 : node17436;
													assign node17436 = (inp[9]) ? 4'b0011 : node17437;
														assign node17437 = (inp[2]) ? node17441 : node17438;
															assign node17438 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node17441 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node17445 = (inp[5]) ? node17447 : 4'b0010;
														assign node17447 = (inp[1]) ? node17451 : node17448;
															assign node17448 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node17451 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node17454 = (inp[2]) ? node17466 : node17455;
													assign node17455 = (inp[1]) ? node17461 : node17456;
														assign node17456 = (inp[11]) ? 4'b0011 : node17457;
															assign node17457 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node17461 = (inp[5]) ? node17463 : 4'b0010;
															assign node17463 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node17466 = (inp[9]) ? node17468 : 4'b0011;
														assign node17468 = (inp[5]) ? 4'b0011 : node17469;
															assign node17469 = (inp[1]) ? 4'b0010 : 4'b0011;
								assign node17473 = (inp[4]) ? node17557 : node17474;
									assign node17474 = (inp[1]) ? node17518 : node17475;
										assign node17475 = (inp[12]) ? node17499 : node17476;
											assign node17476 = (inp[11]) ? node17484 : node17477;
												assign node17477 = (inp[10]) ? 4'b0111 : node17478;
													assign node17478 = (inp[0]) ? 4'b0111 : node17479;
														assign node17479 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node17484 = (inp[10]) ? node17494 : node17485;
													assign node17485 = (inp[0]) ? node17491 : node17486;
														assign node17486 = (inp[2]) ? 4'b0111 : node17487;
															assign node17487 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node17491 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node17494 = (inp[5]) ? 4'b0110 : node17495;
														assign node17495 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node17499 = (inp[9]) ? node17509 : node17500;
												assign node17500 = (inp[5]) ? 4'b0011 : node17501;
													assign node17501 = (inp[11]) ? node17503 : 4'b0011;
														assign node17503 = (inp[0]) ? node17505 : 4'b0010;
															assign node17505 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node17509 = (inp[2]) ? node17513 : node17510;
													assign node17510 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node17513 = (inp[5]) ? 4'b0011 : node17514;
														assign node17514 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node17518 = (inp[12]) ? node17542 : node17519;
											assign node17519 = (inp[11]) ? node17537 : node17520;
												assign node17520 = (inp[9]) ? node17526 : node17521;
													assign node17521 = (inp[5]) ? node17523 : 4'b0011;
														assign node17523 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node17526 = (inp[2]) ? node17532 : node17527;
														assign node17527 = (inp[0]) ? node17529 : 4'b0010;
															assign node17529 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node17532 = (inp[0]) ? node17534 : 4'b0011;
															assign node17534 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node17537 = (inp[5]) ? node17539 : 4'b0010;
													assign node17539 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node17542 = (inp[2]) ? node17552 : node17543;
												assign node17543 = (inp[9]) ? node17547 : node17544;
													assign node17544 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node17547 = (inp[0]) ? node17549 : 4'b0111;
														assign node17549 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node17552 = (inp[0]) ? 4'b0110 : node17553;
													assign node17553 = (inp[9]) ? 4'b0110 : 4'b0111;
									assign node17557 = (inp[10]) ? node17581 : node17558;
										assign node17558 = (inp[5]) ? node17572 : node17559;
											assign node17559 = (inp[9]) ? node17565 : node17560;
												assign node17560 = (inp[12]) ? 4'b0110 : node17561;
													assign node17561 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node17565 = (inp[0]) ? 4'b0111 : node17566;
													assign node17566 = (inp[12]) ? node17568 : 4'b0110;
														assign node17568 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node17572 = (inp[9]) ? node17574 : 4'b0111;
												assign node17574 = (inp[0]) ? 4'b0110 : node17575;
													assign node17575 = (inp[1]) ? node17577 : 4'b0111;
														assign node17577 = (inp[11]) ? 4'b0111 : 4'b0110;
										assign node17581 = (inp[5]) ? node17601 : node17582;
											assign node17582 = (inp[9]) ? node17592 : node17583;
												assign node17583 = (inp[0]) ? 4'b0110 : node17584;
													assign node17584 = (inp[12]) ? node17588 : node17585;
														assign node17585 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node17588 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node17592 = (inp[0]) ? 4'b0111 : node17593;
													assign node17593 = (inp[2]) ? node17595 : 4'b0111;
														assign node17595 = (inp[12]) ? node17597 : 4'b0110;
															assign node17597 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node17601 = (inp[9]) ? node17611 : node17602;
												assign node17602 = (inp[1]) ? node17608 : node17603;
													assign node17603 = (inp[0]) ? 4'b0111 : node17604;
														assign node17604 = (inp[12]) ? 4'b0110 : 4'b0111;
													assign node17608 = (inp[12]) ? 4'b0111 : 4'b0110;
												assign node17611 = (inp[0]) ? 4'b0110 : node17612;
													assign node17612 = (inp[11]) ? 4'b0110 : node17613;
														assign node17613 = (inp[1]) ? 4'b0111 : node17614;
															assign node17614 = (inp[12]) ? 4'b0111 : 4'b0110;
							assign node17620 = (inp[13]) ? node17792 : node17621;
								assign node17621 = (inp[12]) ? node17723 : node17622;
									assign node17622 = (inp[4]) ? node17672 : node17623;
										assign node17623 = (inp[11]) ? node17647 : node17624;
											assign node17624 = (inp[9]) ? node17638 : node17625;
												assign node17625 = (inp[5]) ? node17631 : node17626;
													assign node17626 = (inp[10]) ? 4'b0010 : node17627;
														assign node17627 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node17631 = (inp[0]) ? 4'b0011 : node17632;
														assign node17632 = (inp[10]) ? node17634 : 4'b0011;
															assign node17634 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node17638 = (inp[5]) ? node17642 : node17639;
													assign node17639 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node17642 = (inp[10]) ? node17644 : 4'b0010;
														assign node17644 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node17647 = (inp[9]) ? node17659 : node17648;
												assign node17648 = (inp[0]) ? 4'b0010 : node17649;
													assign node17649 = (inp[5]) ? node17651 : 4'b0011;
														assign node17651 = (inp[1]) ? node17655 : node17652;
															assign node17652 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node17655 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node17659 = (inp[2]) ? node17667 : node17660;
													assign node17660 = (inp[5]) ? 4'b0011 : node17661;
														assign node17661 = (inp[1]) ? node17663 : 4'b0010;
															assign node17663 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node17667 = (inp[1]) ? 4'b0011 : node17668;
														assign node17668 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node17672 = (inp[10]) ? node17700 : node17673;
											assign node17673 = (inp[1]) ? node17679 : node17674;
												assign node17674 = (inp[0]) ? node17676 : 4'b0110;
													assign node17676 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node17679 = (inp[2]) ? node17689 : node17680;
													assign node17680 = (inp[9]) ? node17682 : 4'b0111;
														assign node17682 = (inp[0]) ? node17686 : node17683;
															assign node17683 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node17686 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node17689 = (inp[5]) ? node17695 : node17690;
														assign node17690 = (inp[9]) ? 4'b0111 : node17691;
															assign node17691 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node17695 = (inp[0]) ? node17697 : 4'b0110;
															assign node17697 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node17700 = (inp[2]) ? node17710 : node17701;
												assign node17701 = (inp[1]) ? 4'b0110 : node17702;
													assign node17702 = (inp[9]) ? 4'b0111 : node17703;
														assign node17703 = (inp[11]) ? node17705 : 4'b0110;
															assign node17705 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node17710 = (inp[1]) ? node17712 : 4'b0111;
													assign node17712 = (inp[9]) ? node17718 : node17713;
														assign node17713 = (inp[0]) ? 4'b0111 : node17714;
															assign node17714 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node17718 = (inp[5]) ? node17720 : 4'b0110;
															assign node17720 = (inp[0]) ? 4'b0110 : 4'b0111;
									assign node17723 = (inp[1]) ? node17753 : node17724;
										assign node17724 = (inp[2]) ? node17740 : node17725;
											assign node17725 = (inp[9]) ? node17733 : node17726;
												assign node17726 = (inp[4]) ? node17730 : node17727;
													assign node17727 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node17730 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node17733 = (inp[10]) ? node17735 : 4'b0111;
													assign node17735 = (inp[4]) ? 4'b0111 : node17736;
														assign node17736 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node17740 = (inp[9]) ? node17748 : node17741;
												assign node17741 = (inp[5]) ? 4'b0111 : node17742;
													assign node17742 = (inp[11]) ? node17744 : 4'b0110;
														assign node17744 = (inp[4]) ? 4'b0110 : 4'b0111;
												assign node17748 = (inp[5]) ? 4'b0110 : node17749;
													assign node17749 = (inp[0]) ? 4'b0111 : 4'b0110;
										assign node17753 = (inp[11]) ? node17773 : node17754;
											assign node17754 = (inp[9]) ? node17766 : node17755;
												assign node17755 = (inp[5]) ? node17761 : node17756;
													assign node17756 = (inp[4]) ? 4'b0110 : node17757;
														assign node17757 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node17761 = (inp[4]) ? 4'b0111 : node17762;
														assign node17762 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node17766 = (inp[5]) ? node17768 : 4'b0111;
													assign node17768 = (inp[2]) ? 4'b0110 : node17769;
														assign node17769 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node17773 = (inp[2]) ? node17781 : node17774;
												assign node17774 = (inp[10]) ? node17776 : 4'b0110;
													assign node17776 = (inp[4]) ? node17778 : 4'b0110;
														assign node17778 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node17781 = (inp[5]) ? node17789 : node17782;
													assign node17782 = (inp[9]) ? 4'b0111 : node17783;
														assign node17783 = (inp[10]) ? node17785 : 4'b0110;
															assign node17785 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node17789 = (inp[9]) ? 4'b0110 : 4'b0111;
								assign node17792 = (inp[12]) ? node17896 : node17793;
									assign node17793 = (inp[4]) ? node17857 : node17794;
										assign node17794 = (inp[11]) ? node17838 : node17795;
											assign node17795 = (inp[9]) ? node17817 : node17796;
												assign node17796 = (inp[5]) ? node17806 : node17797;
													assign node17797 = (inp[0]) ? node17799 : 4'b0111;
														assign node17799 = (inp[10]) ? node17803 : node17800;
															assign node17800 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node17803 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node17806 = (inp[10]) ? node17812 : node17807;
														assign node17807 = (inp[2]) ? 4'b0110 : node17808;
															assign node17808 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node17812 = (inp[2]) ? node17814 : 4'b0111;
															assign node17814 = (inp[0]) ? 4'b0110 : 4'b0110;
												assign node17817 = (inp[5]) ? node17829 : node17818;
													assign node17818 = (inp[0]) ? node17824 : node17819;
														assign node17819 = (inp[10]) ? node17821 : 4'b0111;
															assign node17821 = (inp[2]) ? 4'b0110 : 4'b0110;
														assign node17824 = (inp[1]) ? node17826 : 4'b0110;
															assign node17826 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node17829 = (inp[10]) ? 4'b0111 : node17830;
														assign node17830 = (inp[2]) ? node17834 : node17831;
															assign node17831 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node17834 = (inp[1]) ? 4'b0110 : 4'b0110;
											assign node17838 = (inp[0]) ? node17844 : node17839;
												assign node17839 = (inp[10]) ? node17841 : 4'b0110;
													assign node17841 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node17844 = (inp[10]) ? 4'b0110 : node17845;
													assign node17845 = (inp[1]) ? node17851 : node17846;
														assign node17846 = (inp[2]) ? 4'b0110 : node17847;
															assign node17847 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node17851 = (inp[5]) ? 4'b0111 : node17852;
															assign node17852 = (inp[2]) ? 4'b0111 : 4'b0110;
										assign node17857 = (inp[10]) ? node17869 : node17858;
											assign node17858 = (inp[9]) ? 4'b0011 : node17859;
												assign node17859 = (inp[11]) ? node17861 : 4'b0011;
													assign node17861 = (inp[1]) ? node17863 : 4'b0010;
														assign node17863 = (inp[0]) ? node17865 : 4'b0010;
															assign node17865 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node17869 = (inp[0]) ? node17887 : node17870;
												assign node17870 = (inp[9]) ? node17876 : node17871;
													assign node17871 = (inp[1]) ? 4'b0011 : node17872;
														assign node17872 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node17876 = (inp[2]) ? node17882 : node17877;
														assign node17877 = (inp[1]) ? 4'b0011 : node17878;
															assign node17878 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node17882 = (inp[5]) ? 4'b0010 : node17883;
															assign node17883 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node17887 = (inp[5]) ? node17889 : 4'b0010;
													assign node17889 = (inp[2]) ? 4'b0011 : node17890;
														assign node17890 = (inp[9]) ? node17892 : 4'b0010;
															assign node17892 = (inp[1]) ? 4'b0010 : 4'b0011;
									assign node17896 = (inp[9]) ? node17912 : node17897;
										assign node17897 = (inp[5]) ? node17907 : node17898;
											assign node17898 = (inp[4]) ? 4'b0010 : node17899;
												assign node17899 = (inp[0]) ? node17903 : node17900;
													assign node17900 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node17903 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node17907 = (inp[2]) ? 4'b0011 : node17908;
												assign node17908 = (inp[0]) ? 4'b0011 : 4'b0010;
										assign node17912 = (inp[5]) ? node17926 : node17913;
											assign node17913 = (inp[4]) ? 4'b0011 : node17914;
												assign node17914 = (inp[11]) ? 4'b0010 : node17915;
													assign node17915 = (inp[1]) ? 4'b0011 : node17916;
														assign node17916 = (inp[10]) ? node17920 : node17917;
															assign node17917 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node17920 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node17926 = (inp[4]) ? 4'b0010 : node17927;
												assign node17927 = (inp[2]) ? 4'b0010 : 4'b0011;
					assign node17931 = (inp[6]) ? node18927 : node17932;
						assign node17932 = (inp[12]) ? node18452 : node17933;
							assign node17933 = (inp[15]) ? node18171 : node17934;
								assign node17934 = (inp[4]) ? node18054 : node17935;
									assign node17935 = (inp[2]) ? node18003 : node17936;
										assign node17936 = (inp[13]) ? node17976 : node17937;
											assign node17937 = (inp[1]) ? node17955 : node17938;
												assign node17938 = (inp[5]) ? node17948 : node17939;
													assign node17939 = (inp[0]) ? node17941 : 4'b0100;
														assign node17941 = (inp[11]) ? node17945 : node17942;
															assign node17942 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node17945 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node17948 = (inp[9]) ? node17952 : node17949;
														assign node17949 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node17952 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node17955 = (inp[9]) ? node17967 : node17956;
													assign node17956 = (inp[0]) ? node17962 : node17957;
														assign node17957 = (inp[10]) ? 4'b0000 : node17958;
															assign node17958 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node17962 = (inp[10]) ? 4'b0001 : node17963;
															assign node17963 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node17967 = (inp[11]) ? node17971 : node17968;
														assign node17968 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node17971 = (inp[10]) ? 4'b0001 : node17972;
															assign node17972 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node17976 = (inp[1]) ? node17988 : node17977;
												assign node17977 = (inp[5]) ? node17985 : node17978;
													assign node17978 = (inp[10]) ? node17980 : 4'b0001;
														assign node17980 = (inp[9]) ? node17982 : 4'b0000;
															assign node17982 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node17985 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node17988 = (inp[10]) ? node17996 : node17989;
													assign node17989 = (inp[5]) ? node17991 : 4'b0100;
														assign node17991 = (inp[0]) ? 4'b0100 : node17992;
															assign node17992 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node17996 = (inp[0]) ? 4'b0101 : node17997;
														assign node17997 = (inp[11]) ? 4'b0100 : node17998;
															assign node17998 = (inp[9]) ? 4'b0100 : 4'b0100;
										assign node18003 = (inp[13]) ? node18035 : node18004;
											assign node18004 = (inp[1]) ? node18022 : node18005;
												assign node18005 = (inp[5]) ? node18013 : node18006;
													assign node18006 = (inp[10]) ? 4'b0000 : node18007;
														assign node18007 = (inp[11]) ? 4'b0001 : node18008;
															assign node18008 = (inp[0]) ? 4'b0000 : 4'b0000;
													assign node18013 = (inp[11]) ? node18017 : node18014;
														assign node18014 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node18017 = (inp[0]) ? 4'b0100 : node18018;
															assign node18018 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node18022 = (inp[9]) ? node18030 : node18023;
													assign node18023 = (inp[0]) ? node18025 : 4'b0101;
														assign node18025 = (inp[5]) ? 4'b0101 : node18026;
															assign node18026 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node18030 = (inp[5]) ? node18032 : 4'b0100;
														assign node18032 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node18035 = (inp[11]) ? node18043 : node18036;
												assign node18036 = (inp[5]) ? node18040 : node18037;
													assign node18037 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node18040 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node18043 = (inp[1]) ? node18047 : node18044;
													assign node18044 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node18047 = (inp[9]) ? 4'b0000 : node18048;
														assign node18048 = (inp[10]) ? 4'b0000 : node18049;
															assign node18049 = (inp[5]) ? 4'b0000 : 4'b0001;
									assign node18054 = (inp[2]) ? node18122 : node18055;
										assign node18055 = (inp[13]) ? node18087 : node18056;
											assign node18056 = (inp[5]) ? node18072 : node18057;
												assign node18057 = (inp[1]) ? 4'b0011 : node18058;
													assign node18058 = (inp[9]) ? node18064 : node18059;
														assign node18059 = (inp[10]) ? 4'b0111 : node18060;
															assign node18060 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node18064 = (inp[10]) ? node18068 : node18065;
															assign node18065 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node18068 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node18072 = (inp[1]) ? node18080 : node18073;
													assign node18073 = (inp[11]) ? 4'b0011 : node18074;
														assign node18074 = (inp[0]) ? node18076 : 4'b0011;
															assign node18076 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node18080 = (inp[0]) ? node18082 : 4'b0010;
														assign node18082 = (inp[10]) ? 4'b0011 : node18083;
															assign node18083 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node18087 = (inp[5]) ? node18107 : node18088;
												assign node18088 = (inp[1]) ? node18098 : node18089;
													assign node18089 = (inp[9]) ? node18091 : 4'b0011;
														assign node18091 = (inp[11]) ? node18095 : node18092;
															assign node18092 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node18095 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node18098 = (inp[9]) ? node18102 : node18099;
														assign node18099 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node18102 = (inp[0]) ? node18104 : 4'b0110;
															assign node18104 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node18107 = (inp[11]) ? node18117 : node18108;
													assign node18108 = (inp[0]) ? node18112 : node18109;
														assign node18109 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node18112 = (inp[10]) ? 4'b0111 : node18113;
															assign node18113 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node18117 = (inp[0]) ? 4'b0110 : node18118;
														assign node18118 = (inp[9]) ? 4'b0111 : 4'b0110;
										assign node18122 = (inp[13]) ? node18152 : node18123;
											assign node18123 = (inp[5]) ? node18139 : node18124;
												assign node18124 = (inp[1]) ? node18136 : node18125;
													assign node18125 = (inp[9]) ? node18131 : node18126;
														assign node18126 = (inp[10]) ? node18128 : 4'b0011;
															assign node18128 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node18131 = (inp[11]) ? 4'b0011 : node18132;
															assign node18132 = (inp[10]) ? 4'b0010 : 4'b0010;
													assign node18136 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node18139 = (inp[1]) ? node18145 : node18140;
													assign node18140 = (inp[0]) ? 4'b0110 : node18141;
														assign node18141 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node18145 = (inp[11]) ? 4'b0111 : node18146;
														assign node18146 = (inp[10]) ? node18148 : 4'b0111;
															assign node18148 = (inp[0]) ? 4'b0110 : 4'b0110;
											assign node18152 = (inp[10]) ? node18158 : node18153;
												assign node18153 = (inp[9]) ? node18155 : 4'b0010;
													assign node18155 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node18158 = (inp[9]) ? node18164 : node18159;
													assign node18159 = (inp[1]) ? 4'b0011 : node18160;
														assign node18160 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node18164 = (inp[5]) ? node18168 : node18165;
														assign node18165 = (inp[1]) ? 4'b0011 : 4'b0110;
														assign node18168 = (inp[11]) ? 4'b0011 : 4'b0010;
								assign node18171 = (inp[1]) ? node18315 : node18172;
									assign node18172 = (inp[4]) ? node18242 : node18173;
										assign node18173 = (inp[11]) ? node18207 : node18174;
											assign node18174 = (inp[0]) ? node18192 : node18175;
												assign node18175 = (inp[13]) ? node18179 : node18176;
													assign node18176 = (inp[5]) ? 4'b0010 : 4'b0110;
													assign node18179 = (inp[9]) ? node18185 : node18180;
														assign node18180 = (inp[10]) ? 4'b0010 : node18181;
															assign node18181 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node18185 = (inp[2]) ? node18189 : node18186;
															assign node18186 = (inp[5]) ? 4'b0010 : 4'b0110;
															assign node18189 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node18192 = (inp[9]) ? node18202 : node18193;
													assign node18193 = (inp[13]) ? node18197 : node18194;
														assign node18194 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node18197 = (inp[10]) ? node18199 : 4'b0111;
															assign node18199 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node18202 = (inp[10]) ? node18204 : 4'b0011;
														assign node18204 = (inp[13]) ? 4'b0010 : 4'b0111;
											assign node18207 = (inp[9]) ? node18223 : node18208;
												assign node18208 = (inp[2]) ? node18212 : node18209;
													assign node18209 = (inp[13]) ? 4'b0010 : 4'b0111;
													assign node18212 = (inp[0]) ? node18218 : node18213;
														assign node18213 = (inp[10]) ? 4'b0110 : node18214;
															assign node18214 = (inp[5]) ? 4'b0010 : 4'b0010;
														assign node18218 = (inp[10]) ? 4'b0010 : node18219;
															assign node18219 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node18223 = (inp[10]) ? node18231 : node18224;
													assign node18224 = (inp[2]) ? node18228 : node18225;
														assign node18225 = (inp[0]) ? 4'b0110 : 4'b0010;
														assign node18228 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node18231 = (inp[5]) ? node18239 : node18232;
														assign node18232 = (inp[2]) ? node18236 : node18233;
															assign node18233 = (inp[13]) ? 4'b0111 : 4'b0010;
															assign node18236 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node18239 = (inp[2]) ? 4'b0111 : 4'b0110;
										assign node18242 = (inp[10]) ? node18284 : node18243;
											assign node18243 = (inp[11]) ? node18261 : node18244;
												assign node18244 = (inp[5]) ? node18250 : node18245;
													assign node18245 = (inp[2]) ? node18247 : 4'b0011;
														assign node18247 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node18250 = (inp[0]) ? node18258 : node18251;
														assign node18251 = (inp[2]) ? node18255 : node18252;
															assign node18252 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node18255 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node18258 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node18261 = (inp[9]) ? node18273 : node18262;
													assign node18262 = (inp[5]) ? node18268 : node18263;
														assign node18263 = (inp[0]) ? 4'b0111 : node18264;
															assign node18264 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node18268 = (inp[2]) ? 4'b0011 : node18269;
															assign node18269 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node18273 = (inp[13]) ? node18277 : node18274;
														assign node18274 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node18277 = (inp[5]) ? node18281 : node18278;
															assign node18278 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node18281 = (inp[2]) ? 4'b0010 : 4'b0110;
											assign node18284 = (inp[13]) ? node18298 : node18285;
												assign node18285 = (inp[9]) ? node18293 : node18286;
													assign node18286 = (inp[0]) ? node18288 : 4'b0011;
														assign node18288 = (inp[11]) ? node18290 : 4'b0110;
															assign node18290 = (inp[2]) ? 4'b0010 : 4'b0010;
													assign node18293 = (inp[2]) ? 4'b0010 : node18294;
														assign node18294 = (inp[0]) ? 4'b0010 : 4'b0110;
												assign node18298 = (inp[9]) ? node18304 : node18299;
													assign node18299 = (inp[5]) ? node18301 : 4'b0010;
														assign node18301 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node18304 = (inp[11]) ? node18310 : node18305;
														assign node18305 = (inp[0]) ? node18307 : 4'b0010;
															assign node18307 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node18310 = (inp[2]) ? 4'b0111 : node18311;
															assign node18311 = (inp[5]) ? 4'b0111 : 4'b0011;
									assign node18315 = (inp[0]) ? node18395 : node18316;
										assign node18316 = (inp[5]) ? node18350 : node18317;
											assign node18317 = (inp[11]) ? node18329 : node18318;
												assign node18318 = (inp[9]) ? node18324 : node18319;
													assign node18319 = (inp[10]) ? node18321 : 4'b0011;
														assign node18321 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node18324 = (inp[2]) ? 4'b0110 : node18325;
														assign node18325 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node18329 = (inp[4]) ? node18339 : node18330;
													assign node18330 = (inp[9]) ? node18334 : node18331;
														assign node18331 = (inp[2]) ? 4'b0011 : 4'b0110;
														assign node18334 = (inp[13]) ? node18336 : 4'b0011;
															assign node18336 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node18339 = (inp[9]) ? node18343 : node18340;
														assign node18340 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node18343 = (inp[10]) ? node18347 : node18344;
															assign node18344 = (inp[2]) ? 4'b0111 : 4'b0010;
															assign node18347 = (inp[2]) ? 4'b0010 : 4'b0110;
											assign node18350 = (inp[13]) ? node18372 : node18351;
												assign node18351 = (inp[10]) ? node18367 : node18352;
													assign node18352 = (inp[11]) ? node18360 : node18353;
														assign node18353 = (inp[2]) ? node18357 : node18354;
															assign node18354 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node18357 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node18360 = (inp[2]) ? node18364 : node18361;
															assign node18361 = (inp[4]) ? 4'b0011 : 4'b0110;
															assign node18364 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node18367 = (inp[9]) ? 4'b0011 : node18368;
														assign node18368 = (inp[2]) ? 4'b0010 : 4'b0111;
												assign node18372 = (inp[10]) ? node18386 : node18373;
													assign node18373 = (inp[9]) ? node18379 : node18374;
														assign node18374 = (inp[4]) ? node18376 : 4'b0010;
															assign node18376 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node18379 = (inp[11]) ? node18383 : node18380;
															assign node18380 = (inp[4]) ? 4'b0010 : 4'b0011;
															assign node18383 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node18386 = (inp[11]) ? 4'b0010 : node18387;
														assign node18387 = (inp[4]) ? node18391 : node18388;
															assign node18388 = (inp[2]) ? 4'b0111 : 4'b0010;
															assign node18391 = (inp[2]) ? 4'b0010 : 4'b0110;
										assign node18395 = (inp[13]) ? node18431 : node18396;
											assign node18396 = (inp[10]) ? node18414 : node18397;
												assign node18397 = (inp[9]) ? node18411 : node18398;
													assign node18398 = (inp[2]) ? node18406 : node18399;
														assign node18399 = (inp[4]) ? node18403 : node18400;
															assign node18400 = (inp[11]) ? 4'b0110 : 4'b0110;
															assign node18403 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node18406 = (inp[4]) ? 4'b0110 : node18407;
															assign node18407 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node18411 = (inp[11]) ? 4'b0011 : 4'b0111;
												assign node18414 = (inp[11]) ? node18424 : node18415;
													assign node18415 = (inp[5]) ? node18417 : 4'b0111;
														assign node18417 = (inp[2]) ? node18421 : node18418;
															assign node18418 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node18421 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node18424 = (inp[9]) ? 4'b0110 : node18425;
														assign node18425 = (inp[4]) ? 4'b0111 : node18426;
															assign node18426 = (inp[5]) ? 4'b0110 : 4'b0010;
											assign node18431 = (inp[10]) ? node18439 : node18432;
												assign node18432 = (inp[9]) ? 4'b0111 : node18433;
													assign node18433 = (inp[11]) ? 4'b0010 : node18434;
														assign node18434 = (inp[4]) ? 4'b0110 : 4'b0111;
												assign node18439 = (inp[9]) ? node18447 : node18440;
													assign node18440 = (inp[4]) ? node18444 : node18441;
														assign node18441 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node18444 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node18447 = (inp[4]) ? 4'b0010 : node18448;
														assign node18448 = (inp[5]) ? 4'b0011 : 4'b0010;
							assign node18452 = (inp[4]) ? node18670 : node18453;
								assign node18453 = (inp[15]) ? node18569 : node18454;
									assign node18454 = (inp[2]) ? node18504 : node18455;
										assign node18455 = (inp[13]) ? node18477 : node18456;
											assign node18456 = (inp[5]) ? node18468 : node18457;
												assign node18457 = (inp[10]) ? node18463 : node18458;
													assign node18458 = (inp[9]) ? node18460 : 4'b0111;
														assign node18460 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node18463 = (inp[1]) ? node18465 : 4'b0110;
														assign node18465 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node18468 = (inp[1]) ? node18472 : node18469;
													assign node18469 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node18472 = (inp[11]) ? node18474 : 4'b0011;
														assign node18474 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node18477 = (inp[5]) ? node18489 : node18478;
												assign node18478 = (inp[0]) ? node18482 : node18479;
													assign node18479 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node18482 = (inp[10]) ? node18484 : 4'b0010;
														assign node18484 = (inp[11]) ? node18486 : 4'b0011;
															assign node18486 = (inp[9]) ? 4'b0010 : 4'b0011;
												assign node18489 = (inp[1]) ? node18493 : node18490;
													assign node18490 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node18493 = (inp[0]) ? node18499 : node18494;
														assign node18494 = (inp[11]) ? node18496 : 4'b0111;
															assign node18496 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node18499 = (inp[9]) ? node18501 : 4'b0110;
															assign node18501 = (inp[10]) ? 4'b0111 : 4'b0110;
										assign node18504 = (inp[13]) ? node18542 : node18505;
											assign node18505 = (inp[1]) ? node18527 : node18506;
												assign node18506 = (inp[5]) ? node18514 : node18507;
													assign node18507 = (inp[0]) ? 4'b0010 : node18508;
														assign node18508 = (inp[11]) ? 4'b0011 : node18509;
															assign node18509 = (inp[10]) ? 4'b0010 : 4'b0010;
													assign node18514 = (inp[0]) ? node18520 : node18515;
														assign node18515 = (inp[9]) ? 4'b0011 : node18516;
															assign node18516 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node18520 = (inp[9]) ? node18524 : node18521;
															assign node18521 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node18524 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node18527 = (inp[5]) ? 4'b0110 : node18528;
													assign node18528 = (inp[11]) ? node18534 : node18529;
														assign node18529 = (inp[0]) ? node18531 : 4'b0010;
															assign node18531 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node18534 = (inp[9]) ? node18538 : node18535;
															assign node18535 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node18538 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node18542 = (inp[5]) ? node18548 : node18543;
												assign node18543 = (inp[10]) ? node18545 : 4'b0110;
													assign node18545 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node18548 = (inp[1]) ? node18556 : node18549;
													assign node18549 = (inp[11]) ? 4'b0110 : node18550;
														assign node18550 = (inp[9]) ? node18552 : 4'b0111;
															assign node18552 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node18556 = (inp[11]) ? node18564 : node18557;
														assign node18557 = (inp[9]) ? node18561 : node18558;
															assign node18558 = (inp[0]) ? 4'b0010 : 4'b0010;
															assign node18561 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node18564 = (inp[0]) ? node18566 : 4'b0010;
															assign node18566 = (inp[10]) ? 4'b0011 : 4'b0010;
									assign node18569 = (inp[13]) ? node18607 : node18570;
										assign node18570 = (inp[2]) ? node18582 : node18571;
											assign node18571 = (inp[5]) ? node18575 : node18572;
												assign node18572 = (inp[1]) ? 4'b0000 : 4'b0100;
												assign node18575 = (inp[9]) ? node18579 : node18576;
													assign node18576 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node18579 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node18582 = (inp[1]) ? node18596 : node18583;
												assign node18583 = (inp[5]) ? 4'b0101 : node18584;
													assign node18584 = (inp[0]) ? node18590 : node18585;
														assign node18585 = (inp[11]) ? node18587 : 4'b0001;
															assign node18587 = (inp[9]) ? 4'b0000 : 4'b0000;
														assign node18590 = (inp[10]) ? 4'b0000 : node18591;
															assign node18591 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node18596 = (inp[10]) ? node18602 : node18597;
													assign node18597 = (inp[5]) ? 4'b0100 : node18598;
														assign node18598 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node18602 = (inp[11]) ? 4'b0101 : node18603;
														assign node18603 = (inp[9]) ? 4'b0101 : 4'b0100;
										assign node18607 = (inp[2]) ? node18633 : node18608;
											assign node18608 = (inp[5]) ? node18622 : node18609;
												assign node18609 = (inp[1]) ? node18617 : node18610;
													assign node18610 = (inp[11]) ? node18612 : 4'b0001;
														assign node18612 = (inp[10]) ? 4'b0000 : node18613;
															assign node18613 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node18617 = (inp[9]) ? node18619 : 4'b0101;
														assign node18619 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node18622 = (inp[10]) ? node18628 : node18623;
													assign node18623 = (inp[9]) ? node18625 : 4'b0101;
														assign node18625 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node18628 = (inp[9]) ? node18630 : 4'b0100;
														assign node18630 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node18633 = (inp[5]) ? node18649 : node18634;
												assign node18634 = (inp[1]) ? node18642 : node18635;
													assign node18635 = (inp[11]) ? 4'b0100 : node18636;
														assign node18636 = (inp[10]) ? node18638 : 4'b0101;
															assign node18638 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node18642 = (inp[10]) ? 4'b0000 : node18643;
														assign node18643 = (inp[0]) ? node18645 : 4'b0000;
															assign node18645 = (inp[11]) ? 4'b0000 : 4'b0000;
												assign node18649 = (inp[0]) ? node18659 : node18650;
													assign node18650 = (inp[11]) ? node18654 : node18651;
														assign node18651 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node18654 = (inp[10]) ? 4'b0000 : node18655;
															assign node18655 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node18659 = (inp[1]) ? node18665 : node18660;
														assign node18660 = (inp[10]) ? node18662 : 4'b0001;
															assign node18662 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node18665 = (inp[11]) ? 4'b0001 : node18666;
															assign node18666 = (inp[9]) ? 4'b0001 : 4'b0000;
								assign node18670 = (inp[0]) ? node18816 : node18671;
									assign node18671 = (inp[10]) ? node18751 : node18672;
										assign node18672 = (inp[11]) ? node18712 : node18673;
											assign node18673 = (inp[9]) ? node18695 : node18674;
												assign node18674 = (inp[15]) ? node18686 : node18675;
													assign node18675 = (inp[13]) ? node18679 : node18676;
														assign node18676 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node18679 = (inp[2]) ? node18683 : node18680;
															assign node18680 = (inp[1]) ? 4'b0101 : 4'b0000;
															assign node18683 = (inp[1]) ? 4'b0001 : 4'b0101;
													assign node18686 = (inp[13]) ? node18692 : node18687;
														assign node18687 = (inp[5]) ? 4'b0001 : node18688;
															assign node18688 = (inp[2]) ? 4'b0001 : 4'b0001;
														assign node18692 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node18695 = (inp[2]) ? node18705 : node18696;
													assign node18696 = (inp[1]) ? 4'b0100 : node18697;
														assign node18697 = (inp[15]) ? node18701 : node18698;
															assign node18698 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node18701 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node18705 = (inp[5]) ? node18709 : node18706;
														assign node18706 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node18709 = (inp[15]) ? 4'b0100 : 4'b0101;
											assign node18712 = (inp[9]) ? node18732 : node18713;
												assign node18713 = (inp[2]) ? node18723 : node18714;
													assign node18714 = (inp[13]) ? node18720 : node18715;
														assign node18715 = (inp[15]) ? node18717 : 4'b0000;
															assign node18717 = (inp[5]) ? 4'b0001 : 4'b0001;
														assign node18720 = (inp[15]) ? 4'b0100 : 4'b0101;
													assign node18723 = (inp[13]) ? node18729 : node18724;
														assign node18724 = (inp[15]) ? 4'b0100 : node18725;
															assign node18725 = (inp[5]) ? 4'b0100 : 4'b0000;
														assign node18729 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node18732 = (inp[15]) ? node18742 : node18733;
													assign node18733 = (inp[2]) ? node18737 : node18734;
														assign node18734 = (inp[5]) ? 4'b0001 : 4'b0101;
														assign node18737 = (inp[5]) ? node18739 : 4'b0001;
															assign node18739 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node18742 = (inp[5]) ? 4'b0101 : node18743;
														assign node18743 = (inp[13]) ? node18747 : node18744;
															assign node18744 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node18747 = (inp[2]) ? 4'b0101 : 4'b0000;
										assign node18751 = (inp[9]) ? node18781 : node18752;
											assign node18752 = (inp[11]) ? node18766 : node18753;
												assign node18753 = (inp[15]) ? node18759 : node18754;
													assign node18754 = (inp[2]) ? 4'b0101 : node18755;
														assign node18755 = (inp[13]) ? 4'b0100 : 4'b0000;
													assign node18759 = (inp[5]) ? node18761 : 4'b0000;
														assign node18761 = (inp[2]) ? node18763 : 4'b0100;
															assign node18763 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node18766 = (inp[1]) ? node18776 : node18767;
													assign node18767 = (inp[5]) ? node18773 : node18768;
														assign node18768 = (inp[13]) ? 4'b0000 : node18769;
															assign node18769 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node18773 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node18776 = (inp[5]) ? 4'b0001 : node18777;
														assign node18777 = (inp[13]) ? 4'b0101 : 4'b0000;
											assign node18781 = (inp[15]) ? node18801 : node18782;
												assign node18782 = (inp[1]) ? node18798 : node18783;
													assign node18783 = (inp[2]) ? node18791 : node18784;
														assign node18784 = (inp[5]) ? node18788 : node18785;
															assign node18785 = (inp[13]) ? 4'b0000 : 4'b0101;
															assign node18788 = (inp[13]) ? 4'b0101 : 4'b0000;
														assign node18791 = (inp[5]) ? node18795 : node18792;
															assign node18792 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node18795 = (inp[13]) ? 4'b0001 : 4'b0100;
													assign node18798 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node18801 = (inp[13]) ? node18809 : node18802;
													assign node18802 = (inp[5]) ? 4'b0001 : node18803;
														assign node18803 = (inp[11]) ? 4'b0101 : node18804;
															assign node18804 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node18809 = (inp[11]) ? node18813 : node18810;
														assign node18810 = (inp[5]) ? 4'b0101 : 4'b0001;
														assign node18813 = (inp[1]) ? 4'b0100 : 4'b0000;
									assign node18816 = (inp[9]) ? node18872 : node18817;
										assign node18817 = (inp[10]) ? node18847 : node18818;
											assign node18818 = (inp[11]) ? node18832 : node18819;
												assign node18819 = (inp[2]) ? node18825 : node18820;
													assign node18820 = (inp[13]) ? node18822 : 4'b0001;
														assign node18822 = (inp[1]) ? 4'b0100 : 4'b0001;
													assign node18825 = (inp[1]) ? 4'b0000 : node18826;
														assign node18826 = (inp[5]) ? node18828 : 4'b0000;
															assign node18828 = (inp[15]) ? 4'b0000 : 4'b0001;
												assign node18832 = (inp[1]) ? node18840 : node18833;
													assign node18833 = (inp[15]) ? 4'b0100 : node18834;
														assign node18834 = (inp[5]) ? 4'b0000 : node18835;
															assign node18835 = (inp[2]) ? 4'b0100 : 4'b0000;
													assign node18840 = (inp[15]) ? node18842 : 4'b0001;
														assign node18842 = (inp[2]) ? 4'b0000 : node18843;
															assign node18843 = (inp[13]) ? 4'b0100 : 4'b0000;
											assign node18847 = (inp[15]) ? node18863 : node18848;
												assign node18848 = (inp[2]) ? node18858 : node18849;
													assign node18849 = (inp[5]) ? node18853 : node18850;
														assign node18850 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node18853 = (inp[1]) ? 4'b0000 : node18854;
															assign node18854 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node18858 = (inp[13]) ? 4'b0001 : node18859;
														assign node18859 = (inp[1]) ? 4'b0100 : 4'b0001;
												assign node18863 = (inp[1]) ? 4'b0001 : node18864;
													assign node18864 = (inp[2]) ? node18866 : 4'b0100;
														assign node18866 = (inp[5]) ? node18868 : 4'b0101;
															assign node18868 = (inp[13]) ? 4'b0001 : 4'b0101;
										assign node18872 = (inp[10]) ? node18894 : node18873;
											assign node18873 = (inp[11]) ? node18885 : node18874;
												assign node18874 = (inp[5]) ? node18878 : node18875;
													assign node18875 = (inp[2]) ? 4'b0100 : 4'b0000;
													assign node18878 = (inp[13]) ? node18882 : node18879;
														assign node18879 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node18882 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node18885 = (inp[2]) ? node18887 : 4'b0101;
													assign node18887 = (inp[1]) ? 4'b0101 : node18888;
														assign node18888 = (inp[5]) ? 4'b0001 : node18889;
															assign node18889 = (inp[15]) ? 4'b0101 : 4'b0001;
											assign node18894 = (inp[15]) ? node18912 : node18895;
												assign node18895 = (inp[1]) ? node18909 : node18896;
													assign node18896 = (inp[13]) ? node18902 : node18897;
														assign node18897 = (inp[2]) ? node18899 : 4'b0100;
															assign node18899 = (inp[5]) ? 4'b0100 : 4'b0000;
														assign node18902 = (inp[11]) ? node18906 : node18903;
															assign node18903 = (inp[5]) ? 4'b0001 : 4'b0101;
															assign node18906 = (inp[2]) ? 4'b0000 : 4'b0000;
													assign node18909 = (inp[2]) ? 4'b0101 : 4'b0000;
												assign node18912 = (inp[5]) ? node18918 : node18913;
													assign node18913 = (inp[1]) ? 4'b0000 : node18914;
														assign node18914 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node18918 = (inp[11]) ? node18922 : node18919;
														assign node18919 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node18922 = (inp[13]) ? 4'b0100 : node18923;
															assign node18923 = (inp[2]) ? 4'b0100 : 4'b0000;
						assign node18927 = (inp[13]) ? node19161 : node18928;
							assign node18928 = (inp[4]) ? node19098 : node18929;
								assign node18929 = (inp[12]) ? node19013 : node18930;
									assign node18930 = (inp[1]) ? node18972 : node18931;
										assign node18931 = (inp[15]) ? node18953 : node18932;
											assign node18932 = (inp[0]) ? node18948 : node18933;
												assign node18933 = (inp[9]) ? node18935 : 4'b0100;
													assign node18935 = (inp[10]) ? node18941 : node18936;
														assign node18936 = (inp[11]) ? node18938 : 4'b0100;
															assign node18938 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node18941 = (inp[5]) ? node18945 : node18942;
															assign node18942 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node18945 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node18948 = (inp[9]) ? node18950 : 4'b0101;
													assign node18950 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node18953 = (inp[2]) ? node18959 : node18954;
												assign node18954 = (inp[10]) ? node18956 : 4'b0000;
													assign node18956 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node18959 = (inp[11]) ? node18967 : node18960;
													assign node18960 = (inp[5]) ? node18962 : 4'b0000;
														assign node18962 = (inp[10]) ? node18964 : 4'b0001;
															assign node18964 = (inp[9]) ? 4'b0000 : 4'b0000;
													assign node18967 = (inp[9]) ? node18969 : 4'b0001;
														assign node18969 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node18972 = (inp[2]) ? node18986 : node18973;
											assign node18973 = (inp[15]) ? node18981 : node18974;
												assign node18974 = (inp[9]) ? node18976 : 4'b0000;
													assign node18976 = (inp[5]) ? node18978 : 4'b0001;
														assign node18978 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node18981 = (inp[5]) ? 4'b0001 : node18982;
													assign node18982 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node18986 = (inp[10]) ? node19002 : node18987;
												assign node18987 = (inp[11]) ? node18995 : node18988;
													assign node18988 = (inp[0]) ? node18992 : node18989;
														assign node18989 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node18992 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node18995 = (inp[0]) ? node18997 : 4'b0000;
														assign node18997 = (inp[5]) ? 4'b0000 : node18998;
															assign node18998 = (inp[15]) ? 4'b0001 : 4'b0000;
												assign node19002 = (inp[15]) ? 4'b0000 : node19003;
													assign node19003 = (inp[0]) ? node19005 : 4'b0001;
														assign node19005 = (inp[11]) ? node19009 : node19006;
															assign node19006 = (inp[5]) ? 4'b0000 : 4'b0000;
															assign node19009 = (inp[9]) ? 4'b0000 : 4'b0000;
									assign node19013 = (inp[1]) ? node19055 : node19014;
										assign node19014 = (inp[15]) ? node19040 : node19015;
											assign node19015 = (inp[11]) ? node19033 : node19016;
												assign node19016 = (inp[9]) ? node19022 : node19017;
													assign node19017 = (inp[0]) ? node19019 : 4'b0001;
														assign node19019 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node19022 = (inp[2]) ? node19028 : node19023;
														assign node19023 = (inp[5]) ? 4'b0001 : node19024;
															assign node19024 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node19028 = (inp[5]) ? 4'b0000 : node19029;
															assign node19029 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node19033 = (inp[5]) ? 4'b0000 : node19034;
													assign node19034 = (inp[10]) ? 4'b0001 : node19035;
														assign node19035 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node19040 = (inp[0]) ? node19050 : node19041;
												assign node19041 = (inp[5]) ? 4'b0100 : node19042;
													assign node19042 = (inp[11]) ? 4'b0100 : node19043;
														assign node19043 = (inp[2]) ? node19045 : 4'b0101;
															assign node19045 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node19050 = (inp[9]) ? 4'b0101 : node19051;
													assign node19051 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node19055 = (inp[2]) ? node19069 : node19056;
											assign node19056 = (inp[5]) ? node19062 : node19057;
												assign node19057 = (inp[9]) ? 4'b0100 : node19058;
													assign node19058 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node19062 = (inp[9]) ? node19066 : node19063;
													assign node19063 = (inp[15]) ? 4'b0100 : 4'b0101;
													assign node19066 = (inp[15]) ? 4'b0101 : 4'b0100;
											assign node19069 = (inp[5]) ? node19083 : node19070;
												assign node19070 = (inp[15]) ? node19078 : node19071;
													assign node19071 = (inp[9]) ? node19075 : node19072;
														assign node19072 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node19075 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node19078 = (inp[9]) ? node19080 : 4'b0101;
														assign node19080 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node19083 = (inp[11]) ? node19093 : node19084;
													assign node19084 = (inp[10]) ? 4'b0100 : node19085;
														assign node19085 = (inp[15]) ? node19089 : node19086;
															assign node19086 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node19089 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node19093 = (inp[0]) ? node19095 : 4'b0101;
														assign node19095 = (inp[9]) ? 4'b0101 : 4'b0100;
								assign node19098 = (inp[15]) ? node19150 : node19099;
									assign node19099 = (inp[9]) ? node19123 : node19100;
										assign node19100 = (inp[1]) ? 4'b0100 : node19101;
											assign node19101 = (inp[5]) ? node19115 : node19102;
												assign node19102 = (inp[11]) ? node19108 : node19103;
													assign node19103 = (inp[0]) ? 4'b0101 : node19104;
														assign node19104 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node19108 = (inp[0]) ? node19112 : node19109;
														assign node19109 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node19112 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node19115 = (inp[11]) ? 4'b0100 : node19116;
													assign node19116 = (inp[10]) ? node19118 : 4'b0100;
														assign node19118 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node19123 = (inp[1]) ? 4'b0101 : node19124;
											assign node19124 = (inp[5]) ? node19134 : node19125;
												assign node19125 = (inp[10]) ? 4'b0100 : node19126;
													assign node19126 = (inp[0]) ? node19130 : node19127;
														assign node19127 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node19130 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node19134 = (inp[2]) ? node19136 : 4'b0101;
													assign node19136 = (inp[10]) ? node19142 : node19137;
														assign node19137 = (inp[0]) ? 4'b0100 : node19138;
															assign node19138 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node19142 = (inp[11]) ? node19146 : node19143;
															assign node19143 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node19146 = (inp[0]) ? 4'b0100 : 4'b0101;
									assign node19150 = (inp[9]) ? node19156 : node19151;
										assign node19151 = (inp[12]) ? 4'b0101 : node19152;
											assign node19152 = (inp[1]) ? 4'b0101 : 4'b0100;
										assign node19156 = (inp[12]) ? 4'b0100 : node19157;
											assign node19157 = (inp[1]) ? 4'b0100 : 4'b0101;
							assign node19161 = (inp[4]) ? node19375 : node19162;
								assign node19162 = (inp[12]) ? node19280 : node19163;
									assign node19163 = (inp[15]) ? node19215 : node19164;
										assign node19164 = (inp[1]) ? node19190 : node19165;
											assign node19165 = (inp[9]) ? node19179 : node19166;
												assign node19166 = (inp[10]) ? node19172 : node19167;
													assign node19167 = (inp[2]) ? 4'b0001 : node19168;
														assign node19168 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node19172 = (inp[5]) ? 4'b0001 : node19173;
														assign node19173 = (inp[2]) ? node19175 : 4'b0001;
															assign node19175 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node19179 = (inp[2]) ? node19185 : node19180;
													assign node19180 = (inp[0]) ? 4'b0001 : node19181;
														assign node19181 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node19185 = (inp[0]) ? 4'b0000 : node19186;
														assign node19186 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node19190 = (inp[5]) ? node19202 : node19191;
												assign node19191 = (inp[2]) ? 4'b0100 : node19192;
													assign node19192 = (inp[10]) ? node19198 : node19193;
														assign node19193 = (inp[11]) ? node19195 : 4'b0101;
															assign node19195 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node19198 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node19202 = (inp[11]) ? 4'b0100 : node19203;
													assign node19203 = (inp[10]) ? node19209 : node19204;
														assign node19204 = (inp[0]) ? 4'b0101 : node19205;
															assign node19205 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node19209 = (inp[0]) ? 4'b0100 : node19210;
															assign node19210 = (inp[9]) ? 4'b0100 : 4'b0100;
										assign node19215 = (inp[0]) ? node19245 : node19216;
											assign node19216 = (inp[2]) ? node19224 : node19217;
												assign node19217 = (inp[11]) ? node19219 : 4'b0101;
													assign node19219 = (inp[10]) ? node19221 : 4'b0101;
														assign node19221 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node19224 = (inp[10]) ? node19240 : node19225;
													assign node19225 = (inp[1]) ? node19233 : node19226;
														assign node19226 = (inp[11]) ? node19230 : node19227;
															assign node19227 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node19230 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node19233 = (inp[9]) ? node19237 : node19234;
															assign node19234 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node19237 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node19240 = (inp[11]) ? node19242 : 4'b0101;
														assign node19242 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node19245 = (inp[11]) ? node19265 : node19246;
												assign node19246 = (inp[2]) ? node19256 : node19247;
													assign node19247 = (inp[5]) ? 4'b0100 : node19248;
														assign node19248 = (inp[10]) ? node19252 : node19249;
															assign node19249 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node19252 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node19256 = (inp[5]) ? 4'b0101 : node19257;
														assign node19257 = (inp[10]) ? node19261 : node19258;
															assign node19258 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node19261 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node19265 = (inp[1]) ? node19271 : node19266;
													assign node19266 = (inp[5]) ? 4'b0100 : node19267;
														assign node19267 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node19271 = (inp[5]) ? node19273 : 4'b0100;
														assign node19273 = (inp[10]) ? node19277 : node19274;
															assign node19274 = (inp[2]) ? 4'b0100 : 4'b0100;
															assign node19277 = (inp[9]) ? 4'b0100 : 4'b0101;
									assign node19280 = (inp[15]) ? node19322 : node19281;
										assign node19281 = (inp[1]) ? node19299 : node19282;
											assign node19282 = (inp[2]) ? node19292 : node19283;
												assign node19283 = (inp[9]) ? node19289 : node19284;
													assign node19284 = (inp[5]) ? node19286 : 4'b0101;
														assign node19286 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node19289 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node19292 = (inp[9]) ? node19294 : 4'b0100;
													assign node19294 = (inp[5]) ? node19296 : 4'b0101;
														assign node19296 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node19299 = (inp[11]) ? node19315 : node19300;
												assign node19300 = (inp[10]) ? node19302 : 4'b0001;
													assign node19302 = (inp[0]) ? node19308 : node19303;
														assign node19303 = (inp[5]) ? node19305 : 4'b0000;
															assign node19305 = (inp[9]) ? 4'b0000 : 4'b0000;
														assign node19308 = (inp[2]) ? node19312 : node19309;
															assign node19309 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node19312 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node19315 = (inp[5]) ? 4'b0000 : node19316;
													assign node19316 = (inp[2]) ? 4'b0000 : node19317;
														assign node19317 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node19322 = (inp[11]) ? node19352 : node19323;
											assign node19323 = (inp[5]) ? node19345 : node19324;
												assign node19324 = (inp[1]) ? node19338 : node19325;
													assign node19325 = (inp[2]) ? node19333 : node19326;
														assign node19326 = (inp[0]) ? node19330 : node19327;
															assign node19327 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node19330 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node19333 = (inp[0]) ? node19335 : 4'b0001;
															assign node19335 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node19338 = (inp[2]) ? 4'b0000 : node19339;
														assign node19339 = (inp[10]) ? node19341 : 4'b0001;
															assign node19341 = (inp[9]) ? 4'b0000 : 4'b0000;
												assign node19345 = (inp[1]) ? node19349 : node19346;
													assign node19346 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node19349 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node19352 = (inp[1]) ? node19366 : node19353;
												assign node19353 = (inp[0]) ? node19357 : node19354;
													assign node19354 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node19357 = (inp[5]) ? node19361 : node19358;
														assign node19358 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node19361 = (inp[2]) ? 4'b0000 : node19362;
															assign node19362 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node19366 = (inp[9]) ? 4'b0000 : node19367;
													assign node19367 = (inp[10]) ? node19369 : 4'b0000;
														assign node19369 = (inp[0]) ? 4'b0001 : node19370;
															assign node19370 = (inp[2]) ? 4'b0000 : 4'b0001;
								assign node19375 = (inp[9]) ? node19389 : node19376;
									assign node19376 = (inp[1]) ? 4'b0001 : node19377;
										assign node19377 = (inp[12]) ? node19383 : node19378;
											assign node19378 = (inp[15]) ? 4'b0000 : node19379;
												assign node19379 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node19383 = (inp[0]) ? 4'b0001 : node19384;
												assign node19384 = (inp[15]) ? 4'b0001 : 4'b0000;
									assign node19389 = (inp[1]) ? 4'b0000 : node19390;
										assign node19390 = (inp[12]) ? node19396 : node19391;
											assign node19391 = (inp[15]) ? 4'b0001 : node19392;
												assign node19392 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node19396 = (inp[0]) ? 4'b0000 : node19397;
												assign node19397 = (inp[15]) ? 4'b0000 : 4'b0001;
			assign node19402 = (inp[6]) ? node22006 : node19403;
				assign node19403 = (inp[12]) ? node20825 : node19404;
					assign node19404 = (inp[15]) ? node20150 : node19405;
						assign node19405 = (inp[14]) ? node19839 : node19406;
							assign node19406 = (inp[1]) ? node19648 : node19407;
								assign node19407 = (inp[4]) ? node19519 : node19408;
									assign node19408 = (inp[5]) ? node19466 : node19409;
										assign node19409 = (inp[0]) ? node19435 : node19410;
											assign node19410 = (inp[13]) ? node19420 : node19411;
												assign node19411 = (inp[9]) ? 4'b0000 : node19412;
													assign node19412 = (inp[11]) ? node19414 : 4'b0101;
														assign node19414 = (inp[10]) ? 4'b0001 : node19415;
															assign node19415 = (inp[7]) ? 4'b0001 : 4'b0100;
												assign node19420 = (inp[10]) ? node19426 : node19421;
													assign node19421 = (inp[9]) ? 4'b0101 : node19422;
														assign node19422 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node19426 = (inp[2]) ? node19430 : node19427;
														assign node19427 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node19430 = (inp[7]) ? node19432 : 4'b0100;
															assign node19432 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node19435 = (inp[9]) ? node19449 : node19436;
												assign node19436 = (inp[7]) ? node19442 : node19437;
													assign node19437 = (inp[2]) ? 4'b0100 : node19438;
														assign node19438 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node19442 = (inp[2]) ? 4'b0000 : node19443;
														assign node19443 = (inp[13]) ? 4'b0100 : node19444;
															assign node19444 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node19449 = (inp[7]) ? node19459 : node19450;
													assign node19450 = (inp[2]) ? node19452 : 4'b0000;
														assign node19452 = (inp[13]) ? node19456 : node19453;
															assign node19453 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node19456 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node19459 = (inp[2]) ? node19463 : node19460;
														assign node19460 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node19463 = (inp[10]) ? 4'b0001 : 4'b0000;
										assign node19466 = (inp[13]) ? node19482 : node19467;
											assign node19467 = (inp[2]) ? node19475 : node19468;
												assign node19468 = (inp[7]) ? node19472 : node19469;
													assign node19469 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node19472 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node19475 = (inp[7]) ? node19477 : 4'b0100;
													assign node19477 = (inp[11]) ? 4'b0000 : node19478;
														assign node19478 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node19482 = (inp[0]) ? node19498 : node19483;
												assign node19483 = (inp[9]) ? node19493 : node19484;
													assign node19484 = (inp[7]) ? node19490 : node19485;
														assign node19485 = (inp[10]) ? 4'b0100 : node19486;
															assign node19486 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node19490 = (inp[2]) ? 4'b0001 : 4'b0100;
													assign node19493 = (inp[10]) ? 4'b0101 : node19494;
														assign node19494 = (inp[2]) ? 4'b0101 : 4'b0001;
												assign node19498 = (inp[11]) ? node19508 : node19499;
													assign node19499 = (inp[2]) ? node19505 : node19500;
														assign node19500 = (inp[7]) ? 4'b0100 : node19501;
															assign node19501 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node19505 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node19508 = (inp[9]) ? node19514 : node19509;
														assign node19509 = (inp[2]) ? node19511 : 4'b0100;
															assign node19511 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node19514 = (inp[2]) ? node19516 : 4'b0101;
															assign node19516 = (inp[10]) ? 4'b0100 : 4'b0101;
									assign node19519 = (inp[11]) ? node19589 : node19520;
										assign node19520 = (inp[0]) ? node19554 : node19521;
											assign node19521 = (inp[9]) ? node19537 : node19522;
												assign node19522 = (inp[7]) ? node19524 : 4'b0101;
													assign node19524 = (inp[13]) ? node19530 : node19525;
														assign node19525 = (inp[5]) ? 4'b0100 : node19526;
															assign node19526 = (inp[2]) ? 4'b0001 : 4'b0100;
														assign node19530 = (inp[5]) ? node19534 : node19531;
															assign node19531 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node19534 = (inp[2]) ? 4'b0100 : 4'b0000;
												assign node19537 = (inp[7]) ? node19545 : node19538;
													assign node19538 = (inp[13]) ? 4'b0100 : node19539;
														assign node19539 = (inp[10]) ? 4'b0001 : node19540;
															assign node19540 = (inp[5]) ? 4'b0100 : 4'b0000;
													assign node19545 = (inp[10]) ? 4'b0100 : node19546;
														assign node19546 = (inp[13]) ? node19550 : node19547;
															assign node19547 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node19550 = (inp[2]) ? 4'b0000 : 4'b0101;
											assign node19554 = (inp[5]) ? node19566 : node19555;
												assign node19555 = (inp[10]) ? 4'b0101 : node19556;
													assign node19556 = (inp[2]) ? node19562 : node19557;
														assign node19557 = (inp[13]) ? 4'b0101 : node19558;
															assign node19558 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node19562 = (inp[13]) ? 4'b0000 : 4'b0101;
												assign node19566 = (inp[9]) ? node19578 : node19567;
													assign node19567 = (inp[13]) ? node19573 : node19568;
														assign node19568 = (inp[10]) ? node19570 : 4'b0000;
															assign node19570 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node19573 = (inp[2]) ? node19575 : 4'b0101;
															assign node19575 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node19578 = (inp[7]) ? node19584 : node19579;
														assign node19579 = (inp[2]) ? node19581 : 4'b0101;
															assign node19581 = (inp[13]) ? 4'b0000 : 4'b0000;
														assign node19584 = (inp[2]) ? 4'b0100 : node19585;
															assign node19585 = (inp[13]) ? 4'b0000 : 4'b0000;
										assign node19589 = (inp[7]) ? node19615 : node19590;
											assign node19590 = (inp[2]) ? node19602 : node19591;
												assign node19591 = (inp[5]) ? node19597 : node19592;
													assign node19592 = (inp[13]) ? 4'b0000 : node19593;
														assign node19593 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node19597 = (inp[9]) ? 4'b0101 : node19598;
														assign node19598 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node19602 = (inp[5]) ? node19610 : node19603;
													assign node19603 = (inp[13]) ? node19607 : node19604;
														assign node19604 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node19607 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node19610 = (inp[10]) ? 4'b0001 : node19611;
														assign node19611 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node19615 = (inp[9]) ? node19637 : node19616;
												assign node19616 = (inp[10]) ? node19626 : node19617;
													assign node19617 = (inp[5]) ? node19623 : node19618;
														assign node19618 = (inp[13]) ? 4'b0001 : node19619;
															assign node19619 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node19623 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node19626 = (inp[13]) ? node19632 : node19627;
														assign node19627 = (inp[5]) ? node19629 : 4'b0001;
															assign node19629 = (inp[0]) ? 4'b0001 : 4'b0100;
														assign node19632 = (inp[5]) ? 4'b0000 : node19633;
															assign node19633 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node19637 = (inp[10]) ? node19641 : node19638;
													assign node19638 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node19641 = (inp[13]) ? 4'b0000 : node19642;
														assign node19642 = (inp[0]) ? node19644 : 4'b0101;
															assign node19644 = (inp[5]) ? 4'b0000 : 4'b0001;
								assign node19648 = (inp[10]) ? node19744 : node19649;
									assign node19649 = (inp[11]) ? node19691 : node19650;
										assign node19650 = (inp[13]) ? node19672 : node19651;
											assign node19651 = (inp[0]) ? node19665 : node19652;
												assign node19652 = (inp[2]) ? node19658 : node19653;
													assign node19653 = (inp[5]) ? node19655 : 4'b0000;
														assign node19655 = (inp[9]) ? 4'b0101 : 4'b0000;
													assign node19658 = (inp[5]) ? node19660 : 4'b0101;
														assign node19660 = (inp[7]) ? 4'b0101 : node19661;
															assign node19661 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node19665 = (inp[4]) ? node19669 : node19666;
													assign node19666 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node19669 = (inp[2]) ? 4'b0000 : 4'b0100;
											assign node19672 = (inp[7]) ? node19678 : node19673;
												assign node19673 = (inp[2]) ? node19675 : 4'b0001;
													assign node19675 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node19678 = (inp[2]) ? node19684 : node19679;
													assign node19679 = (inp[5]) ? node19681 : 4'b0101;
														assign node19681 = (inp[4]) ? 4'b0001 : 4'b0100;
													assign node19684 = (inp[4]) ? node19688 : node19685;
														assign node19685 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node19688 = (inp[5]) ? 4'b0100 : 4'b0001;
										assign node19691 = (inp[13]) ? node19717 : node19692;
											assign node19692 = (inp[2]) ? node19704 : node19693;
												assign node19693 = (inp[7]) ? node19699 : node19694;
													assign node19694 = (inp[4]) ? node19696 : 4'b0001;
														assign node19696 = (inp[5]) ? 4'b0101 : 4'b0001;
													assign node19699 = (inp[5]) ? node19701 : 4'b0101;
														assign node19701 = (inp[4]) ? 4'b0001 : 4'b0100;
												assign node19704 = (inp[7]) ? node19710 : node19705;
													assign node19705 = (inp[5]) ? 4'b0001 : node19706;
														assign node19706 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node19710 = (inp[4]) ? node19714 : node19711;
														assign node19711 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node19714 = (inp[5]) ? 4'b0100 : 4'b0000;
											assign node19717 = (inp[7]) ? node19727 : node19718;
												assign node19718 = (inp[2]) ? node19724 : node19719;
													assign node19719 = (inp[9]) ? 4'b0000 : node19720;
														assign node19720 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node19724 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node19727 = (inp[0]) ? node19735 : node19728;
													assign node19728 = (inp[2]) ? 4'b0101 : node19729;
														assign node19729 = (inp[4]) ? node19731 : 4'b0101;
															assign node19731 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node19735 = (inp[2]) ? node19737 : 4'b0000;
														assign node19737 = (inp[4]) ? node19741 : node19738;
															assign node19738 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node19741 = (inp[5]) ? 4'b0101 : 4'b0001;
									assign node19744 = (inp[2]) ? node19796 : node19745;
										assign node19745 = (inp[7]) ? node19763 : node19746;
											assign node19746 = (inp[4]) ? node19754 : node19747;
												assign node19747 = (inp[11]) ? node19751 : node19748;
													assign node19748 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node19751 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node19754 = (inp[5]) ? node19760 : node19755;
													assign node19755 = (inp[11]) ? node19757 : 4'b0001;
														assign node19757 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node19760 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node19763 = (inp[4]) ? node19787 : node19764;
												assign node19764 = (inp[0]) ? node19778 : node19765;
													assign node19765 = (inp[5]) ? node19771 : node19766;
														assign node19766 = (inp[11]) ? 4'b0101 : node19767;
															assign node19767 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node19771 = (inp[11]) ? node19775 : node19772;
															assign node19772 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node19775 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node19778 = (inp[9]) ? node19780 : 4'b0100;
														assign node19780 = (inp[5]) ? node19784 : node19781;
															assign node19781 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node19784 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node19787 = (inp[5]) ? node19793 : node19788;
													assign node19788 = (inp[9]) ? 4'b0101 : node19789;
														assign node19789 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node19793 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node19796 = (inp[7]) ? node19816 : node19797;
											assign node19797 = (inp[5]) ? node19807 : node19798;
												assign node19798 = (inp[13]) ? 4'b0101 : node19799;
													assign node19799 = (inp[0]) ? 4'b0101 : node19800;
														assign node19800 = (inp[9]) ? node19802 : 4'b0100;
															assign node19802 = (inp[4]) ? 4'b0100 : 4'b0100;
												assign node19807 = (inp[4]) ? node19811 : node19808;
													assign node19808 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node19811 = (inp[9]) ? node19813 : 4'b0001;
														assign node19813 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node19816 = (inp[5]) ? node19828 : node19817;
												assign node19817 = (inp[0]) ? 4'b0001 : node19818;
													assign node19818 = (inp[9]) ? node19820 : 4'b0001;
														assign node19820 = (inp[4]) ? node19824 : node19821;
															assign node19821 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node19824 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node19828 = (inp[4]) ? node19832 : node19829;
													assign node19829 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node19832 = (inp[9]) ? 4'b0100 : node19833;
														assign node19833 = (inp[11]) ? 4'b0101 : node19834;
															assign node19834 = (inp[13]) ? 4'b0101 : 4'b0100;
							assign node19839 = (inp[10]) ? node20013 : node19840;
								assign node19840 = (inp[13]) ? node19928 : node19841;
									assign node19841 = (inp[11]) ? node19875 : node19842;
										assign node19842 = (inp[7]) ? node19860 : node19843;
											assign node19843 = (inp[5]) ? node19853 : node19844;
												assign node19844 = (inp[2]) ? node19846 : 4'b0010;
													assign node19846 = (inp[0]) ? 4'b0111 : node19847;
														assign node19847 = (inp[4]) ? 4'b0110 : node19848;
															assign node19848 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node19853 = (inp[4]) ? node19857 : node19854;
													assign node19854 = (inp[2]) ? 4'b0011 : 4'b0110;
													assign node19857 = (inp[2]) ? 4'b0110 : 4'b0011;
											assign node19860 = (inp[2]) ? node19868 : node19861;
												assign node19861 = (inp[4]) ? 4'b0110 : node19862;
													assign node19862 = (inp[5]) ? node19864 : 4'b0110;
														assign node19864 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node19868 = (inp[5]) ? node19872 : node19869;
													assign node19869 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node19872 = (inp[4]) ? 4'b0010 : 4'b0110;
										assign node19875 = (inp[0]) ? node19903 : node19876;
											assign node19876 = (inp[4]) ? node19892 : node19877;
												assign node19877 = (inp[1]) ? node19881 : node19878;
													assign node19878 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node19881 = (inp[2]) ? node19887 : node19882;
														assign node19882 = (inp[9]) ? 4'b0110 : node19883;
															assign node19883 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node19887 = (inp[5]) ? node19889 : 4'b0011;
															assign node19889 = (inp[7]) ? 4'b0110 : 4'b0011;
												assign node19892 = (inp[7]) ? node19900 : node19893;
													assign node19893 = (inp[2]) ? node19897 : node19894;
														assign node19894 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node19897 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node19900 = (inp[2]) ? 4'b0010 : 4'b0110;
											assign node19903 = (inp[1]) ? node19909 : node19904;
												assign node19904 = (inp[2]) ? node19906 : 4'b0111;
													assign node19906 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node19909 = (inp[4]) ? node19923 : node19910;
													assign node19910 = (inp[2]) ? node19916 : node19911;
														assign node19911 = (inp[5]) ? 4'b0110 : node19912;
															assign node19912 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node19916 = (inp[9]) ? node19920 : node19917;
															assign node19917 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node19920 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node19923 = (inp[5]) ? node19925 : 4'b0111;
														assign node19925 = (inp[2]) ? 4'b0010 : 4'b0011;
									assign node19928 = (inp[2]) ? node19972 : node19929;
										assign node19929 = (inp[7]) ? node19953 : node19930;
											assign node19930 = (inp[4]) ? node19942 : node19931;
												assign node19931 = (inp[5]) ? node19937 : node19932;
													assign node19932 = (inp[1]) ? 4'b0011 : node19933;
														assign node19933 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node19937 = (inp[11]) ? node19939 : 4'b0111;
														assign node19939 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node19942 = (inp[5]) ? node19948 : node19943;
													assign node19943 = (inp[1]) ? 4'b0011 : node19944;
														assign node19944 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node19948 = (inp[1]) ? 4'b0010 : node19949;
														assign node19949 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node19953 = (inp[5]) ? node19959 : node19954;
												assign node19954 = (inp[1]) ? 4'b0111 : node19955;
													assign node19955 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node19959 = (inp[4]) ? node19967 : node19960;
													assign node19960 = (inp[0]) ? 4'b0010 : node19961;
														assign node19961 = (inp[1]) ? node19963 : 4'b0010;
															assign node19963 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node19967 = (inp[1]) ? 4'b0111 : node19968;
														assign node19968 = (inp[11]) ? 4'b0110 : 4'b0111;
										assign node19972 = (inp[7]) ? node19994 : node19973;
											assign node19973 = (inp[11]) ? node19985 : node19974;
												assign node19974 = (inp[5]) ? node19982 : node19975;
													assign node19975 = (inp[4]) ? node19979 : node19976;
														assign node19976 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node19979 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node19982 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node19985 = (inp[4]) ? node19991 : node19986;
													assign node19986 = (inp[5]) ? node19988 : 4'b0111;
														assign node19988 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node19991 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node19994 = (inp[5]) ? node20004 : node19995;
												assign node19995 = (inp[4]) ? node20001 : node19996;
													assign node19996 = (inp[1]) ? 4'b0010 : node19997;
														assign node19997 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node20001 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node20004 = (inp[4]) ? node20010 : node20005;
													assign node20005 = (inp[1]) ? 4'b0111 : node20006;
														assign node20006 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node20010 = (inp[1]) ? 4'b0011 : 4'b0010;
								assign node20013 = (inp[13]) ? node20077 : node20014;
									assign node20014 = (inp[7]) ? node20052 : node20015;
										assign node20015 = (inp[2]) ? node20031 : node20016;
											assign node20016 = (inp[5]) ? node20022 : node20017;
												assign node20017 = (inp[11]) ? node20019 : 4'b0011;
													assign node20019 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node20022 = (inp[4]) ? node20028 : node20023;
													assign node20023 = (inp[1]) ? 4'b0111 : node20024;
														assign node20024 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node20028 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node20031 = (inp[11]) ? node20045 : node20032;
												assign node20032 = (inp[4]) ? node20038 : node20033;
													assign node20033 = (inp[5]) ? 4'b0010 : node20034;
														assign node20034 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node20038 = (inp[9]) ? 4'b0111 : node20039;
														assign node20039 = (inp[0]) ? node20041 : 4'b0110;
															assign node20041 = (inp[1]) ? 4'b0110 : 4'b0110;
												assign node20045 = (inp[4]) ? node20049 : node20046;
													assign node20046 = (inp[5]) ? 4'b0011 : 4'b0111;
													assign node20049 = (inp[5]) ? 4'b0111 : 4'b0110;
										assign node20052 = (inp[2]) ? node20064 : node20053;
											assign node20053 = (inp[5]) ? node20059 : node20054;
												assign node20054 = (inp[4]) ? node20056 : 4'b0111;
													assign node20056 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node20059 = (inp[4]) ? 4'b0111 : node20060;
													assign node20060 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node20064 = (inp[4]) ? node20072 : node20065;
												assign node20065 = (inp[5]) ? node20069 : node20066;
													assign node20066 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node20069 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node20072 = (inp[11]) ? node20074 : 4'b0011;
													assign node20074 = (inp[0]) ? 4'b0011 : 4'b0010;
									assign node20077 = (inp[4]) ? node20111 : node20078;
										assign node20078 = (inp[5]) ? node20092 : node20079;
											assign node20079 = (inp[2]) ? node20083 : node20080;
												assign node20080 = (inp[7]) ? 4'b0110 : 4'b0010;
												assign node20083 = (inp[7]) ? node20087 : node20084;
													assign node20084 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node20087 = (inp[11]) ? node20089 : 4'b0011;
														assign node20089 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node20092 = (inp[11]) ? node20106 : node20093;
												assign node20093 = (inp[0]) ? node20101 : node20094;
													assign node20094 = (inp[7]) ? node20096 : 4'b0011;
														assign node20096 = (inp[2]) ? 4'b0110 : node20097;
															assign node20097 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node20101 = (inp[7]) ? node20103 : 4'b0110;
														assign node20103 = (inp[2]) ? 4'b0110 : 4'b0011;
												assign node20106 = (inp[1]) ? node20108 : 4'b0111;
													assign node20108 = (inp[7]) ? 4'b0110 : 4'b0011;
										assign node20111 = (inp[11]) ? node20125 : node20112;
											assign node20112 = (inp[7]) ? node20122 : node20113;
												assign node20113 = (inp[2]) ? node20117 : node20114;
													assign node20114 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node20117 = (inp[5]) ? 4'b0111 : node20118;
														assign node20118 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node20122 = (inp[2]) ? 4'b0010 : 4'b0110;
											assign node20125 = (inp[1]) ? node20135 : node20126;
												assign node20126 = (inp[7]) ? node20132 : node20127;
													assign node20127 = (inp[5]) ? node20129 : 4'b0011;
														assign node20129 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node20132 = (inp[2]) ? 4'b0011 : 4'b0111;
												assign node20135 = (inp[9]) ? node20143 : node20136;
													assign node20136 = (inp[2]) ? node20140 : node20137;
														assign node20137 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node20140 = (inp[7]) ? 4'b0010 : 4'b0110;
													assign node20143 = (inp[0]) ? 4'b0011 : node20144;
														assign node20144 = (inp[5]) ? node20146 : 4'b0110;
															assign node20146 = (inp[2]) ? 4'b0110 : 4'b0011;
						assign node20150 = (inp[13]) ? node20470 : node20151;
							assign node20151 = (inp[10]) ? node20319 : node20152;
								assign node20152 = (inp[1]) ? node20240 : node20153;
									assign node20153 = (inp[14]) ? node20189 : node20154;
										assign node20154 = (inp[0]) ? node20172 : node20155;
											assign node20155 = (inp[2]) ? node20159 : node20156;
												assign node20156 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node20159 = (inp[4]) ? node20169 : node20160;
													assign node20160 = (inp[9]) ? 4'b0110 : node20161;
														assign node20161 = (inp[5]) ? node20165 : node20162;
															assign node20162 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node20165 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node20169 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node20172 = (inp[11]) ? node20182 : node20173;
												assign node20173 = (inp[7]) ? 4'b0011 : node20174;
													assign node20174 = (inp[4]) ? node20176 : 4'b0110;
														assign node20176 = (inp[2]) ? node20178 : 4'b0110;
															assign node20178 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node20182 = (inp[5]) ? 4'b0010 : node20183;
													assign node20183 = (inp[2]) ? 4'b0010 : node20184;
														assign node20184 = (inp[4]) ? 4'b0110 : 4'b0010;
										assign node20189 = (inp[7]) ? node20231 : node20190;
											assign node20190 = (inp[0]) ? node20214 : node20191;
												assign node20191 = (inp[9]) ? node20203 : node20192;
													assign node20192 = (inp[5]) ? node20200 : node20193;
														assign node20193 = (inp[11]) ? node20197 : node20194;
															assign node20194 = (inp[2]) ? 4'b0010 : 4'b0010;
															assign node20197 = (inp[2]) ? 4'b0110 : 4'b0011;
														assign node20200 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node20203 = (inp[2]) ? node20209 : node20204;
														assign node20204 = (inp[4]) ? node20206 : 4'b0011;
															assign node20206 = (inp[11]) ? 4'b0110 : 4'b0110;
														assign node20209 = (inp[4]) ? node20211 : 4'b0110;
															assign node20211 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node20214 = (inp[9]) ? node20222 : node20215;
													assign node20215 = (inp[11]) ? node20219 : node20216;
														assign node20216 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node20219 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node20222 = (inp[11]) ? 4'b0111 : node20223;
														assign node20223 = (inp[5]) ? node20227 : node20224;
															assign node20224 = (inp[2]) ? 4'b0010 : 4'b0010;
															assign node20227 = (inp[4]) ? 4'b0111 : 4'b0010;
											assign node20231 = (inp[2]) ? node20235 : node20232;
												assign node20232 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node20235 = (inp[4]) ? 4'b0010 : node20236;
													assign node20236 = (inp[5]) ? 4'b0110 : 4'b0111;
									assign node20240 = (inp[14]) ? node20280 : node20241;
										assign node20241 = (inp[7]) ? node20261 : node20242;
											assign node20242 = (inp[9]) ? node20256 : node20243;
												assign node20243 = (inp[2]) ? node20251 : node20244;
													assign node20244 = (inp[4]) ? node20246 : 4'b0011;
														assign node20246 = (inp[11]) ? node20248 : 4'b0111;
															assign node20248 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node20251 = (inp[4]) ? node20253 : 4'b0111;
														assign node20253 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node20256 = (inp[2]) ? node20258 : 4'b0011;
													assign node20258 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node20261 = (inp[4]) ? node20269 : node20262;
												assign node20262 = (inp[2]) ? node20264 : 4'b0010;
													assign node20264 = (inp[9]) ? 4'b0111 : node20265;
														assign node20265 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node20269 = (inp[2]) ? node20275 : node20270;
													assign node20270 = (inp[11]) ? node20272 : 4'b0111;
														assign node20272 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node20275 = (inp[11]) ? 4'b0011 : node20276;
														assign node20276 = (inp[9]) ? 4'b0010 : 4'b0011;
										assign node20280 = (inp[7]) ? node20306 : node20281;
											assign node20281 = (inp[9]) ? node20295 : node20282;
												assign node20282 = (inp[11]) ? node20290 : node20283;
													assign node20283 = (inp[4]) ? node20287 : node20284;
														assign node20284 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node20287 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node20290 = (inp[2]) ? 4'b0010 : node20291;
														assign node20291 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node20295 = (inp[11]) ? node20301 : node20296;
													assign node20296 = (inp[5]) ? node20298 : 4'b0111;
														assign node20298 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node20301 = (inp[2]) ? 4'b0111 : node20302;
														assign node20302 = (inp[4]) ? 4'b0111 : 4'b0010;
											assign node20306 = (inp[4]) ? node20316 : node20307;
												assign node20307 = (inp[2]) ? node20311 : node20308;
													assign node20308 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node20311 = (inp[5]) ? 4'b0111 : node20312;
														assign node20312 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node20316 = (inp[2]) ? 4'b0011 : 4'b0111;
								assign node20319 = (inp[1]) ? node20391 : node20320;
									assign node20320 = (inp[7]) ? node20348 : node20321;
										assign node20321 = (inp[2]) ? node20341 : node20322;
											assign node20322 = (inp[4]) ? node20330 : node20323;
												assign node20323 = (inp[0]) ? 4'b0011 : node20324;
													assign node20324 = (inp[14]) ? node20326 : 4'b0011;
														assign node20326 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node20330 = (inp[9]) ? node20332 : 4'b0111;
													assign node20332 = (inp[5]) ? node20334 : 4'b0111;
														assign node20334 = (inp[14]) ? node20338 : node20335;
															assign node20335 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node20338 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node20341 = (inp[4]) ? node20343 : 4'b0111;
												assign node20343 = (inp[5]) ? 4'b0011 : node20344;
													assign node20344 = (inp[0]) ? 4'b0011 : 4'b0010;
										assign node20348 = (inp[4]) ? node20376 : node20349;
											assign node20349 = (inp[2]) ? node20361 : node20350;
												assign node20350 = (inp[5]) ? node20352 : 4'b0011;
													assign node20352 = (inp[0]) ? node20356 : node20353;
														assign node20353 = (inp[14]) ? 4'b0010 : 4'b0011;
														assign node20356 = (inp[11]) ? 4'b0010 : node20357;
															assign node20357 = (inp[14]) ? 4'b0011 : 4'b0010;
												assign node20361 = (inp[5]) ? node20371 : node20362;
													assign node20362 = (inp[0]) ? 4'b0110 : node20363;
														assign node20363 = (inp[11]) ? node20367 : node20364;
															assign node20364 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node20367 = (inp[14]) ? 4'b0111 : 4'b0110;
													assign node20371 = (inp[11]) ? 4'b0111 : node20372;
														assign node20372 = (inp[14]) ? 4'b0111 : 4'b0110;
											assign node20376 = (inp[2]) ? node20386 : node20377;
												assign node20377 = (inp[0]) ? node20379 : 4'b0111;
													assign node20379 = (inp[5]) ? 4'b0111 : node20380;
														assign node20380 = (inp[14]) ? 4'b0111 : node20381;
															assign node20381 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node20386 = (inp[14]) ? 4'b0011 : node20387;
													assign node20387 = (inp[5]) ? 4'b0010 : 4'b0011;
									assign node20391 = (inp[11]) ? node20433 : node20392;
										assign node20392 = (inp[2]) ? node20406 : node20393;
											assign node20393 = (inp[4]) ? node20399 : node20394;
												assign node20394 = (inp[5]) ? node20396 : 4'b0010;
													assign node20396 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node20399 = (inp[5]) ? node20401 : 4'b0110;
													assign node20401 = (inp[14]) ? node20403 : 4'b0110;
														assign node20403 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node20406 = (inp[4]) ? node20426 : node20407;
												assign node20407 = (inp[14]) ? node20415 : node20408;
													assign node20408 = (inp[0]) ? 4'b0110 : node20409;
														assign node20409 = (inp[5]) ? node20411 : 4'b0110;
															assign node20411 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node20415 = (inp[0]) ? node20421 : node20416;
														assign node20416 = (inp[5]) ? 4'b0110 : node20417;
															assign node20417 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node20421 = (inp[7]) ? node20423 : 4'b0111;
															assign node20423 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node20426 = (inp[14]) ? node20428 : 4'b0011;
													assign node20428 = (inp[7]) ? 4'b0010 : node20429;
														assign node20429 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node20433 = (inp[2]) ? node20453 : node20434;
											assign node20434 = (inp[4]) ? node20444 : node20435;
												assign node20435 = (inp[5]) ? 4'b0010 : node20436;
													assign node20436 = (inp[0]) ? 4'b0011 : node20437;
														assign node20437 = (inp[14]) ? node20439 : 4'b0010;
															assign node20439 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node20444 = (inp[9]) ? node20446 : 4'b0111;
													assign node20446 = (inp[0]) ? node20448 : 4'b0110;
														assign node20448 = (inp[5]) ? node20450 : 4'b0111;
															assign node20450 = (inp[7]) ? 4'b0110 : 4'b0110;
											assign node20453 = (inp[4]) ? node20461 : node20454;
												assign node20454 = (inp[14]) ? 4'b0110 : node20455;
													assign node20455 = (inp[0]) ? 4'b0110 : node20456;
														assign node20456 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node20461 = (inp[14]) ? node20463 : 4'b0010;
													assign node20463 = (inp[9]) ? node20465 : 4'b0011;
														assign node20465 = (inp[7]) ? 4'b0010 : node20466;
															assign node20466 = (inp[5]) ? 4'b0010 : 4'b0011;
							assign node20470 = (inp[1]) ? node20626 : node20471;
								assign node20471 = (inp[10]) ? node20549 : node20472;
									assign node20472 = (inp[5]) ? node20502 : node20473;
										assign node20473 = (inp[4]) ? node20491 : node20474;
											assign node20474 = (inp[2]) ? node20482 : node20475;
												assign node20475 = (inp[0]) ? node20477 : 4'b0010;
													assign node20477 = (inp[11]) ? node20479 : 4'b0010;
														assign node20479 = (inp[14]) ? 4'b0011 : 4'b0010;
												assign node20482 = (inp[7]) ? node20484 : 4'b0110;
													assign node20484 = (inp[9]) ? 4'b0110 : node20485;
														assign node20485 = (inp[14]) ? node20487 : 4'b0111;
															assign node20487 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node20491 = (inp[2]) ? node20495 : node20492;
												assign node20492 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node20495 = (inp[7]) ? 4'b0010 : node20496;
													assign node20496 = (inp[14]) ? node20498 : 4'b0011;
														assign node20498 = (inp[11]) ? 4'b0011 : 4'b0010;
										assign node20502 = (inp[11]) ? node20524 : node20503;
											assign node20503 = (inp[2]) ? node20513 : node20504;
												assign node20504 = (inp[4]) ? node20508 : node20505;
													assign node20505 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node20508 = (inp[14]) ? node20510 : 4'b0110;
														assign node20510 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node20513 = (inp[4]) ? node20515 : 4'b0111;
													assign node20515 = (inp[9]) ? node20517 : 4'b0011;
														assign node20517 = (inp[7]) ? node20521 : node20518;
															assign node20518 = (inp[14]) ? 4'b0011 : 4'b0010;
															assign node20521 = (inp[14]) ? 4'b0010 : 4'b0011;
											assign node20524 = (inp[0]) ? node20540 : node20525;
												assign node20525 = (inp[7]) ? node20531 : node20526;
													assign node20526 = (inp[2]) ? node20528 : 4'b0010;
														assign node20528 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node20531 = (inp[14]) ? 4'b0110 : node20532;
														assign node20532 = (inp[2]) ? node20536 : node20533;
															assign node20533 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node20536 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node20540 = (inp[7]) ? node20546 : node20541;
													assign node20541 = (inp[14]) ? 4'b0110 : node20542;
														assign node20542 = (inp[4]) ? 4'b0111 : 4'b0010;
													assign node20546 = (inp[2]) ? 4'b0010 : 4'b0011;
									assign node20549 = (inp[2]) ? node20587 : node20550;
										assign node20550 = (inp[4]) ? node20564 : node20551;
											assign node20551 = (inp[11]) ? node20553 : 4'b0011;
												assign node20553 = (inp[14]) ? node20555 : 4'b0011;
													assign node20555 = (inp[9]) ? node20557 : 4'b0010;
														assign node20557 = (inp[5]) ? node20561 : node20558;
															assign node20558 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node20561 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node20564 = (inp[0]) ? node20582 : node20565;
												assign node20565 = (inp[7]) ? node20577 : node20566;
													assign node20566 = (inp[14]) ? node20572 : node20567;
														assign node20567 = (inp[5]) ? node20569 : 4'b0111;
															assign node20569 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node20572 = (inp[11]) ? 4'b0110 : node20573;
															assign node20573 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node20577 = (inp[5]) ? 4'b0111 : node20578;
														assign node20578 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node20582 = (inp[11]) ? node20584 : 4'b0111;
													assign node20584 = (inp[9]) ? 4'b0110 : 4'b0111;
										assign node20587 = (inp[4]) ? node20603 : node20588;
											assign node20588 = (inp[0]) ? 4'b0111 : node20589;
												assign node20589 = (inp[9]) ? node20597 : node20590;
													assign node20590 = (inp[11]) ? 4'b0111 : node20591;
														assign node20591 = (inp[7]) ? node20593 : 4'b0111;
															assign node20593 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node20597 = (inp[5]) ? 4'b0110 : node20598;
														assign node20598 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node20603 = (inp[7]) ? node20619 : node20604;
												assign node20604 = (inp[14]) ? node20610 : node20605;
													assign node20605 = (inp[11]) ? 4'b0011 : node20606;
														assign node20606 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node20610 = (inp[9]) ? 4'b0011 : node20611;
														assign node20611 = (inp[5]) ? node20615 : node20612;
															assign node20612 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node20615 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node20619 = (inp[11]) ? 4'b0011 : node20620;
													assign node20620 = (inp[5]) ? node20622 : 4'b0011;
														assign node20622 = (inp[14]) ? 4'b0011 : 4'b0010;
								assign node20626 = (inp[10]) ? node20710 : node20627;
									assign node20627 = (inp[5]) ? node20663 : node20628;
										assign node20628 = (inp[14]) ? node20640 : node20629;
											assign node20629 = (inp[2]) ? node20633 : node20630;
												assign node20630 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node20633 = (inp[4]) ? node20635 : 4'b0111;
													assign node20635 = (inp[11]) ? 4'b0011 : node20636;
														assign node20636 = (inp[7]) ? 4'b0011 : 4'b0010;
											assign node20640 = (inp[11]) ? node20650 : node20641;
												assign node20641 = (inp[4]) ? node20647 : node20642;
													assign node20642 = (inp[2]) ? node20644 : 4'b0011;
														assign node20644 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node20647 = (inp[2]) ? 4'b0011 : 4'b0111;
												assign node20650 = (inp[7]) ? node20658 : node20651;
													assign node20651 = (inp[2]) ? node20655 : node20652;
														assign node20652 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node20655 = (inp[4]) ? 4'b0010 : 4'b0111;
													assign node20658 = (inp[9]) ? node20660 : 4'b0111;
														assign node20660 = (inp[2]) ? 4'b0111 : 4'b0011;
										assign node20663 = (inp[11]) ? node20695 : node20664;
											assign node20664 = (inp[0]) ? node20680 : node20665;
												assign node20665 = (inp[4]) ? node20673 : node20666;
													assign node20666 = (inp[2]) ? 4'b0110 : node20667;
														assign node20667 = (inp[14]) ? 4'b0011 : node20668;
															assign node20668 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node20673 = (inp[2]) ? 4'b0011 : node20674;
														assign node20674 = (inp[7]) ? 4'b0111 : node20675;
															assign node20675 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node20680 = (inp[4]) ? node20686 : node20681;
													assign node20681 = (inp[2]) ? node20683 : 4'b0010;
														assign node20683 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node20686 = (inp[2]) ? node20690 : node20687;
														assign node20687 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node20690 = (inp[7]) ? node20692 : 4'b0010;
															assign node20692 = (inp[14]) ? 4'b0011 : 4'b0010;
											assign node20695 = (inp[2]) ? node20707 : node20696;
												assign node20696 = (inp[4]) ? node20702 : node20697;
													assign node20697 = (inp[7]) ? node20699 : 4'b0011;
														assign node20699 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node20702 = (inp[14]) ? 4'b0111 : node20703;
														assign node20703 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node20707 = (inp[4]) ? 4'b0011 : 4'b0111;
									assign node20710 = (inp[9]) ? node20762 : node20711;
										assign node20711 = (inp[11]) ? node20733 : node20712;
											assign node20712 = (inp[5]) ? node20724 : node20713;
												assign node20713 = (inp[2]) ? node20717 : node20714;
													assign node20714 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node20717 = (inp[4]) ? 4'b0010 : node20718;
														assign node20718 = (inp[14]) ? node20720 : 4'b0110;
															assign node20720 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node20724 = (inp[4]) ? node20728 : node20725;
													assign node20725 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node20728 = (inp[14]) ? node20730 : 4'b0010;
														assign node20730 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node20733 = (inp[2]) ? node20751 : node20734;
												assign node20734 = (inp[4]) ? node20744 : node20735;
													assign node20735 = (inp[7]) ? node20737 : 4'b0010;
														assign node20737 = (inp[14]) ? node20741 : node20738;
															assign node20738 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node20741 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node20744 = (inp[14]) ? 4'b0110 : node20745;
														assign node20745 = (inp[5]) ? node20747 : 4'b0110;
															assign node20747 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node20751 = (inp[4]) ? node20757 : node20752;
													assign node20752 = (inp[14]) ? 4'b0110 : node20753;
														assign node20753 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node20757 = (inp[7]) ? 4'b0010 : node20758;
														assign node20758 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node20762 = (inp[0]) ? node20792 : node20763;
											assign node20763 = (inp[11]) ? node20779 : node20764;
												assign node20764 = (inp[5]) ? node20772 : node20765;
													assign node20765 = (inp[4]) ? node20769 : node20766;
														assign node20766 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node20769 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node20772 = (inp[4]) ? node20774 : 4'b0111;
														assign node20774 = (inp[2]) ? node20776 : 4'b0110;
															assign node20776 = (inp[14]) ? 4'b0011 : 4'b0010;
												assign node20779 = (inp[4]) ? 4'b0111 : node20780;
													assign node20780 = (inp[2]) ? node20786 : node20781;
														assign node20781 = (inp[5]) ? 4'b0010 : node20782;
															assign node20782 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node20786 = (inp[14]) ? 4'b0110 : node20787;
															assign node20787 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node20792 = (inp[14]) ? node20808 : node20793;
												assign node20793 = (inp[7]) ? node20803 : node20794;
													assign node20794 = (inp[4]) ? node20798 : node20795;
														assign node20795 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node20798 = (inp[2]) ? node20800 : 4'b0111;
															assign node20800 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node20803 = (inp[2]) ? node20805 : 4'b0011;
														assign node20805 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node20808 = (inp[7]) ? node20818 : node20809;
													assign node20809 = (inp[4]) ? node20813 : node20810;
														assign node20810 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node20813 = (inp[2]) ? node20815 : 4'b0111;
															assign node20815 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node20818 = (inp[4]) ? node20822 : node20819;
														assign node20819 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node20822 = (inp[2]) ? 4'b0010 : 4'b0110;
					assign node20825 = (inp[14]) ? node21505 : node20826;
						assign node20826 = (inp[15]) ? node21198 : node20827;
							assign node20827 = (inp[4]) ? node20977 : node20828;
								assign node20828 = (inp[2]) ? node20902 : node20829;
									assign node20829 = (inp[7]) ? node20859 : node20830;
										assign node20830 = (inp[13]) ? node20842 : node20831;
											assign node20831 = (inp[10]) ? node20837 : node20832;
												assign node20832 = (inp[11]) ? 4'b0010 : node20833;
													assign node20833 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node20837 = (inp[1]) ? node20839 : 4'b0011;
													assign node20839 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node20842 = (inp[9]) ? node20848 : node20843;
												assign node20843 = (inp[1]) ? node20845 : 4'b0011;
													assign node20845 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node20848 = (inp[11]) ? node20856 : node20849;
													assign node20849 = (inp[10]) ? node20853 : node20850;
														assign node20850 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node20853 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node20856 = (inp[1]) ? 4'b0011 : 4'b0010;
										assign node20859 = (inp[13]) ? node20883 : node20860;
											assign node20860 = (inp[9]) ? node20868 : node20861;
												assign node20861 = (inp[10]) ? node20863 : 4'b0110;
													assign node20863 = (inp[5]) ? node20865 : 4'b0111;
														assign node20865 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node20868 = (inp[1]) ? node20876 : node20869;
													assign node20869 = (inp[0]) ? 4'b0111 : node20870;
														assign node20870 = (inp[11]) ? 4'b0111 : node20871;
															assign node20871 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node20876 = (inp[10]) ? node20880 : node20877;
														assign node20877 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node20880 = (inp[5]) ? 4'b0110 : 4'b0111;
											assign node20883 = (inp[5]) ? node20895 : node20884;
												assign node20884 = (inp[10]) ? node20890 : node20885;
													assign node20885 = (inp[1]) ? 4'b0111 : node20886;
														assign node20886 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node20890 = (inp[11]) ? node20892 : 4'b0110;
														assign node20892 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node20895 = (inp[0]) ? 4'b0111 : node20896;
													assign node20896 = (inp[11]) ? 4'b0110 : node20897;
														assign node20897 = (inp[10]) ? 4'b0111 : 4'b0110;
									assign node20902 = (inp[7]) ? node20928 : node20903;
										assign node20903 = (inp[11]) ? node20921 : node20904;
											assign node20904 = (inp[1]) ? node20912 : node20905;
												assign node20905 = (inp[0]) ? 4'b0110 : node20906;
													assign node20906 = (inp[13]) ? node20908 : 4'b0111;
														assign node20908 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node20912 = (inp[9]) ? 4'b0111 : node20913;
													assign node20913 = (inp[5]) ? node20915 : 4'b0111;
														assign node20915 = (inp[13]) ? node20917 : 4'b0110;
															assign node20917 = (inp[10]) ? 4'b0111 : 4'b0110;
											assign node20921 = (inp[13]) ? node20925 : node20922;
												assign node20922 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node20925 = (inp[10]) ? 4'b0110 : 4'b0111;
										assign node20928 = (inp[13]) ? node20954 : node20929;
											assign node20929 = (inp[10]) ? node20943 : node20930;
												assign node20930 = (inp[9]) ? 4'b0011 : node20931;
													assign node20931 = (inp[5]) ? node20937 : node20932;
														assign node20932 = (inp[1]) ? node20934 : 4'b0011;
															assign node20934 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node20937 = (inp[1]) ? node20939 : 4'b0010;
															assign node20939 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node20943 = (inp[5]) ? node20949 : node20944;
													assign node20944 = (inp[11]) ? 4'b0010 : node20945;
														assign node20945 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node20949 = (inp[11]) ? 4'b0011 : node20950;
														assign node20950 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node20954 = (inp[5]) ? node20966 : node20955;
												assign node20955 = (inp[10]) ? node20961 : node20956;
													assign node20956 = (inp[1]) ? node20958 : 4'b0010;
														assign node20958 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node20961 = (inp[1]) ? node20963 : 4'b0011;
														assign node20963 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node20966 = (inp[10]) ? node20970 : node20967;
													assign node20967 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node20970 = (inp[9]) ? node20972 : 4'b0010;
														assign node20972 = (inp[1]) ? node20974 : 4'b0010;
															assign node20974 = (inp[11]) ? 4'b0010 : 4'b0011;
								assign node20977 = (inp[11]) ? node21093 : node20978;
									assign node20978 = (inp[0]) ? node21038 : node20979;
										assign node20979 = (inp[7]) ? node21003 : node20980;
											assign node20980 = (inp[5]) ? node20988 : node20981;
												assign node20981 = (inp[2]) ? node20983 : 4'b0110;
													assign node20983 = (inp[13]) ? node20985 : 4'b0010;
														assign node20985 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node20988 = (inp[2]) ? node21000 : node20989;
													assign node20989 = (inp[10]) ? node20995 : node20990;
														assign node20990 = (inp[1]) ? 4'b0010 : node20991;
															assign node20991 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node20995 = (inp[9]) ? node20997 : 4'b0010;
															assign node20997 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node21000 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node21003 = (inp[5]) ? node21019 : node21004;
												assign node21004 = (inp[2]) ? node21006 : 4'b0011;
													assign node21006 = (inp[9]) ? node21014 : node21007;
														assign node21007 = (inp[10]) ? node21011 : node21008;
															assign node21008 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node21011 = (inp[13]) ? 4'b0110 : 4'b0110;
														assign node21014 = (inp[13]) ? node21016 : 4'b0111;
															assign node21016 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node21019 = (inp[2]) ? node21027 : node21020;
													assign node21020 = (inp[9]) ? 4'b0111 : node21021;
														assign node21021 = (inp[13]) ? node21023 : 4'b0110;
															assign node21023 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node21027 = (inp[1]) ? node21033 : node21028;
														assign node21028 = (inp[10]) ? node21030 : 4'b0010;
															assign node21030 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node21033 = (inp[9]) ? 4'b0011 : node21034;
															assign node21034 = (inp[10]) ? 4'b0010 : 4'b0010;
										assign node21038 = (inp[13]) ? node21064 : node21039;
											assign node21039 = (inp[2]) ? node21053 : node21040;
												assign node21040 = (inp[5]) ? node21048 : node21041;
													assign node21041 = (inp[7]) ? 4'b0011 : node21042;
														assign node21042 = (inp[10]) ? node21044 : 4'b0111;
															assign node21044 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node21048 = (inp[7]) ? node21050 : 4'b0010;
														assign node21050 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node21053 = (inp[7]) ? node21061 : node21054;
													assign node21054 = (inp[10]) ? node21058 : node21055;
														assign node21055 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node21058 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node21061 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node21064 = (inp[7]) ? node21078 : node21065;
												assign node21065 = (inp[1]) ? node21069 : node21066;
													assign node21066 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node21069 = (inp[2]) ? node21075 : node21070;
														assign node21070 = (inp[5]) ? 4'b0010 : node21071;
															assign node21071 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node21075 = (inp[5]) ? 4'b0110 : 4'b0010;
												assign node21078 = (inp[2]) ? node21086 : node21079;
													assign node21079 = (inp[5]) ? node21083 : node21080;
														assign node21080 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node21083 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node21086 = (inp[5]) ? 4'b0010 : node21087;
														assign node21087 = (inp[1]) ? node21089 : 4'b0111;
															assign node21089 = (inp[10]) ? 4'b0111 : 4'b0110;
									assign node21093 = (inp[5]) ? node21145 : node21094;
										assign node21094 = (inp[9]) ? node21128 : node21095;
											assign node21095 = (inp[0]) ? node21113 : node21096;
												assign node21096 = (inp[2]) ? node21102 : node21097;
													assign node21097 = (inp[7]) ? 4'b0011 : node21098;
														assign node21098 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node21102 = (inp[7]) ? node21110 : node21103;
														assign node21103 = (inp[13]) ? node21107 : node21104;
															assign node21104 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node21107 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node21110 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node21113 = (inp[1]) ? node21121 : node21114;
													assign node21114 = (inp[2]) ? node21118 : node21115;
														assign node21115 = (inp[7]) ? 4'b0010 : 4'b0110;
														assign node21118 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node21121 = (inp[7]) ? node21123 : 4'b0010;
														assign node21123 = (inp[10]) ? 4'b0011 : node21124;
															assign node21124 = (inp[13]) ? 4'b0010 : 4'b0011;
											assign node21128 = (inp[10]) ? node21138 : node21129;
												assign node21129 = (inp[13]) ? 4'b0010 : node21130;
													assign node21130 = (inp[1]) ? node21132 : 4'b0010;
														assign node21132 = (inp[7]) ? node21134 : 4'b0110;
															assign node21134 = (inp[0]) ? 4'b0110 : 4'b0011;
												assign node21138 = (inp[13]) ? node21140 : 4'b0010;
													assign node21140 = (inp[2]) ? node21142 : 4'b0110;
														assign node21142 = (inp[1]) ? 4'b0110 : 4'b0010;
										assign node21145 = (inp[1]) ? node21165 : node21146;
											assign node21146 = (inp[7]) ? node21156 : node21147;
												assign node21147 = (inp[2]) ? node21153 : node21148;
													assign node21148 = (inp[10]) ? node21150 : 4'b0011;
														assign node21150 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node21153 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node21156 = (inp[2]) ? 4'b0010 : node21157;
													assign node21157 = (inp[0]) ? 4'b0111 : node21158;
														assign node21158 = (inp[9]) ? 4'b0111 : node21159;
															assign node21159 = (inp[13]) ? 4'b0110 : 4'b0110;
											assign node21165 = (inp[10]) ? node21185 : node21166;
												assign node21166 = (inp[9]) ? node21176 : node21167;
													assign node21167 = (inp[0]) ? node21173 : node21168;
														assign node21168 = (inp[2]) ? 4'b0011 : node21169;
															assign node21169 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node21173 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node21176 = (inp[13]) ? node21180 : node21177;
														assign node21177 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node21180 = (inp[7]) ? node21182 : 4'b0111;
															assign node21182 = (inp[2]) ? 4'b0011 : 4'b0111;
												assign node21185 = (inp[7]) ? node21193 : node21186;
													assign node21186 = (inp[2]) ? node21190 : node21187;
														assign node21187 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node21190 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node21193 = (inp[2]) ? 4'b0010 : node21194;
														assign node21194 = (inp[13]) ? 4'b0110 : 4'b0111;
							assign node21198 = (inp[2]) ? node21358 : node21199;
								assign node21199 = (inp[5]) ? node21273 : node21200;
									assign node21200 = (inp[4]) ? node21232 : node21201;
										assign node21201 = (inp[13]) ? node21217 : node21202;
											assign node21202 = (inp[9]) ? node21210 : node21203;
												assign node21203 = (inp[7]) ? node21207 : node21204;
													assign node21204 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node21207 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node21210 = (inp[1]) ? node21212 : 4'b0001;
													assign node21212 = (inp[7]) ? 4'b0000 : node21213;
														assign node21213 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node21217 = (inp[9]) ? node21225 : node21218;
												assign node21218 = (inp[0]) ? 4'b0000 : node21219;
													assign node21219 = (inp[10]) ? node21221 : 4'b0000;
														assign node21221 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node21225 = (inp[7]) ? node21229 : node21226;
													assign node21226 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node21229 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node21232 = (inp[9]) ? node21250 : node21233;
											assign node21233 = (inp[10]) ? node21243 : node21234;
												assign node21234 = (inp[1]) ? node21240 : node21235;
													assign node21235 = (inp[7]) ? node21237 : 4'b0000;
														assign node21237 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node21240 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node21243 = (inp[13]) ? node21245 : 4'b0001;
													assign node21245 = (inp[11]) ? node21247 : 4'b0001;
														assign node21247 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node21250 = (inp[7]) ? node21268 : node21251;
												assign node21251 = (inp[13]) ? node21261 : node21252;
													assign node21252 = (inp[1]) ? node21254 : 4'b0000;
														assign node21254 = (inp[0]) ? node21258 : node21255;
															assign node21255 = (inp[11]) ? 4'b0000 : 4'b0000;
															assign node21258 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node21261 = (inp[1]) ? node21263 : 4'b0001;
														assign node21263 = (inp[11]) ? node21265 : 4'b0001;
															assign node21265 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node21268 = (inp[11]) ? node21270 : 4'b0000;
													assign node21270 = (inp[13]) ? 4'b0001 : 4'b0000;
									assign node21273 = (inp[13]) ? node21319 : node21274;
										assign node21274 = (inp[1]) ? node21302 : node21275;
											assign node21275 = (inp[9]) ? node21287 : node21276;
												assign node21276 = (inp[0]) ? node21278 : 4'b0101;
													assign node21278 = (inp[7]) ? node21282 : node21279;
														assign node21279 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node21282 = (inp[10]) ? node21284 : 4'b0100;
															assign node21284 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node21287 = (inp[7]) ? node21295 : node21288;
													assign node21288 = (inp[0]) ? 4'b0100 : node21289;
														assign node21289 = (inp[4]) ? 4'b0101 : node21290;
															assign node21290 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node21295 = (inp[11]) ? node21297 : 4'b0101;
														assign node21297 = (inp[0]) ? node21299 : 4'b0100;
															assign node21299 = (inp[10]) ? 4'b0100 : 4'b0100;
											assign node21302 = (inp[9]) ? node21308 : node21303;
												assign node21303 = (inp[4]) ? 4'b0100 : node21304;
													assign node21304 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node21308 = (inp[0]) ? node21310 : 4'b0100;
													assign node21310 = (inp[11]) ? node21316 : node21311;
														assign node21311 = (inp[7]) ? 4'b0101 : node21312;
															assign node21312 = (inp[10]) ? 4'b0100 : 4'b0100;
														assign node21316 = (inp[10]) ? 4'b0101 : 4'b0100;
										assign node21319 = (inp[11]) ? node21337 : node21320;
											assign node21320 = (inp[7]) ? node21328 : node21321;
												assign node21321 = (inp[10]) ? node21325 : node21322;
													assign node21322 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node21325 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node21328 = (inp[0]) ? node21330 : 4'b0101;
													assign node21330 = (inp[10]) ? node21334 : node21331;
														assign node21331 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node21334 = (inp[4]) ? 4'b0100 : 4'b0101;
											assign node21337 = (inp[7]) ? node21345 : node21338;
												assign node21338 = (inp[10]) ? node21342 : node21339;
													assign node21339 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node21342 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node21345 = (inp[0]) ? node21353 : node21346;
													assign node21346 = (inp[10]) ? node21350 : node21347;
														assign node21347 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node21350 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node21353 = (inp[4]) ? 4'b0100 : node21354;
														assign node21354 = (inp[10]) ? 4'b0101 : 4'b0100;
								assign node21358 = (inp[5]) ? node21448 : node21359;
									assign node21359 = (inp[9]) ? node21395 : node21360;
										assign node21360 = (inp[11]) ? node21382 : node21361;
											assign node21361 = (inp[4]) ? node21369 : node21362;
												assign node21362 = (inp[10]) ? node21366 : node21363;
													assign node21363 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node21366 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node21369 = (inp[1]) ? node21375 : node21370;
													assign node21370 = (inp[13]) ? node21372 : 4'b0101;
														assign node21372 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node21375 = (inp[13]) ? 4'b0101 : node21376;
														assign node21376 = (inp[10]) ? node21378 : 4'b0100;
															assign node21378 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node21382 = (inp[0]) ? node21388 : node21383;
												assign node21383 = (inp[10]) ? node21385 : 4'b0101;
													assign node21385 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node21388 = (inp[10]) ? node21392 : node21389;
													assign node21389 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node21392 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node21395 = (inp[0]) ? node21423 : node21396;
											assign node21396 = (inp[13]) ? node21414 : node21397;
												assign node21397 = (inp[11]) ? node21407 : node21398;
													assign node21398 = (inp[7]) ? 4'b0100 : node21399;
														assign node21399 = (inp[4]) ? node21403 : node21400;
															assign node21400 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node21403 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node21407 = (inp[7]) ? node21411 : node21408;
														assign node21408 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node21411 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node21414 = (inp[7]) ? 4'b0101 : node21415;
													assign node21415 = (inp[1]) ? node21417 : 4'b0100;
														assign node21417 = (inp[11]) ? 4'b0101 : node21418;
															assign node21418 = (inp[4]) ? 4'b0100 : 4'b0100;
											assign node21423 = (inp[13]) ? node21437 : node21424;
												assign node21424 = (inp[1]) ? node21432 : node21425;
													assign node21425 = (inp[11]) ? node21427 : 4'b0101;
														assign node21427 = (inp[7]) ? 4'b0101 : node21428;
															assign node21428 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node21432 = (inp[10]) ? node21434 : 4'b0101;
														assign node21434 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node21437 = (inp[10]) ? node21441 : node21438;
													assign node21438 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node21441 = (inp[1]) ? 4'b0100 : node21442;
														assign node21442 = (inp[7]) ? node21444 : 4'b0101;
															assign node21444 = (inp[4]) ? 4'b0100 : 4'b0100;
									assign node21448 = (inp[1]) ? node21456 : node21449;
										assign node21449 = (inp[10]) ? node21453 : node21450;
											assign node21450 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node21453 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node21456 = (inp[0]) ? node21476 : node21457;
											assign node21457 = (inp[7]) ? node21463 : node21458;
												assign node21458 = (inp[10]) ? node21460 : 4'b0001;
													assign node21460 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node21463 = (inp[4]) ? node21471 : node21464;
													assign node21464 = (inp[13]) ? 4'b0000 : node21465;
														assign node21465 = (inp[11]) ? 4'b0001 : node21466;
															assign node21466 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node21471 = (inp[10]) ? 4'b0001 : node21472;
														assign node21472 = (inp[13]) ? 4'b0001 : 4'b0000;
											assign node21476 = (inp[13]) ? node21490 : node21477;
												assign node21477 = (inp[4]) ? node21485 : node21478;
													assign node21478 = (inp[10]) ? node21482 : node21479;
														assign node21479 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node21482 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node21485 = (inp[9]) ? node21487 : 4'b0000;
														assign node21487 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node21490 = (inp[9]) ? node21496 : node21491;
													assign node21491 = (inp[11]) ? node21493 : 4'b0001;
														assign node21493 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node21496 = (inp[4]) ? node21500 : node21497;
														assign node21497 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node21500 = (inp[7]) ? 4'b0001 : node21501;
															assign node21501 = (inp[11]) ? 4'b0000 : 4'b0001;
						assign node21505 = (inp[2]) ? node21801 : node21506;
							assign node21506 = (inp[15]) ? node21664 : node21507;
								assign node21507 = (inp[7]) ? node21581 : node21508;
									assign node21508 = (inp[4]) ? node21536 : node21509;
										assign node21509 = (inp[5]) ? node21527 : node21510;
											assign node21510 = (inp[10]) ? node21522 : node21511;
												assign node21511 = (inp[0]) ? 4'b0100 : node21512;
													assign node21512 = (inp[9]) ? 4'b0101 : node21513;
														assign node21513 = (inp[13]) ? node21517 : node21514;
															assign node21514 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node21517 = (inp[1]) ? 4'b0100 : 4'b0100;
												assign node21522 = (inp[1]) ? node21524 : 4'b0101;
													assign node21524 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node21527 = (inp[10]) ? node21531 : node21528;
												assign node21528 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node21531 = (inp[1]) ? 4'b0000 : node21532;
													assign node21532 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node21536 = (inp[10]) ? node21564 : node21537;
											assign node21537 = (inp[9]) ? node21549 : node21538;
												assign node21538 = (inp[11]) ? 4'b0001 : node21539;
													assign node21539 = (inp[1]) ? 4'b0000 : node21540;
														assign node21540 = (inp[0]) ? node21544 : node21541;
															assign node21541 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node21544 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node21549 = (inp[0]) ? node21557 : node21550;
													assign node21550 = (inp[5]) ? node21552 : 4'b0000;
														assign node21552 = (inp[1]) ? 4'b0000 : node21553;
															assign node21553 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node21557 = (inp[5]) ? 4'b0000 : node21558;
														assign node21558 = (inp[13]) ? 4'b0001 : node21559;
															assign node21559 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node21564 = (inp[13]) ? node21570 : node21565;
												assign node21565 = (inp[5]) ? node21567 : 4'b0001;
													assign node21567 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node21570 = (inp[5]) ? node21576 : node21571;
													assign node21571 = (inp[1]) ? node21573 : 4'b0000;
														assign node21573 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node21576 = (inp[1]) ? node21578 : 4'b0001;
														assign node21578 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node21581 = (inp[4]) ? node21627 : node21582;
										assign node21582 = (inp[5]) ? node21614 : node21583;
											assign node21583 = (inp[0]) ? node21599 : node21584;
												assign node21584 = (inp[10]) ? node21592 : node21585;
													assign node21585 = (inp[13]) ? 4'b0001 : node21586;
														assign node21586 = (inp[1]) ? 4'b0000 : node21587;
															assign node21587 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node21592 = (inp[13]) ? 4'b0000 : node21593;
														assign node21593 = (inp[1]) ? 4'b0001 : node21594;
															assign node21594 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node21599 = (inp[11]) ? node21607 : node21600;
													assign node21600 = (inp[13]) ? 4'b0001 : node21601;
														assign node21601 = (inp[1]) ? 4'b0001 : node21602;
															assign node21602 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node21607 = (inp[10]) ? node21611 : node21608;
														assign node21608 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node21611 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node21614 = (inp[13]) ? node21620 : node21615;
												assign node21615 = (inp[10]) ? node21617 : 4'b0101;
													assign node21617 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node21620 = (inp[0]) ? 4'b0101 : node21621;
													assign node21621 = (inp[1]) ? 4'b0101 : node21622;
														assign node21622 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node21627 = (inp[11]) ? node21643 : node21628;
											assign node21628 = (inp[1]) ? node21638 : node21629;
												assign node21629 = (inp[9]) ? node21631 : 4'b0100;
													assign node21631 = (inp[13]) ? node21635 : node21632;
														assign node21632 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node21635 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node21638 = (inp[10]) ? node21640 : 4'b0101;
													assign node21640 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node21643 = (inp[9]) ? node21657 : node21644;
												assign node21644 = (inp[1]) ? node21650 : node21645;
													assign node21645 = (inp[13]) ? node21647 : 4'b0101;
														assign node21647 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node21650 = (inp[13]) ? node21654 : node21651;
														assign node21651 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node21654 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node21657 = (inp[10]) ? node21661 : node21658;
													assign node21658 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node21661 = (inp[13]) ? 4'b0100 : 4'b0101;
								assign node21664 = (inp[9]) ? node21742 : node21665;
									assign node21665 = (inp[13]) ? node21709 : node21666;
										assign node21666 = (inp[0]) ? node21684 : node21667;
											assign node21667 = (inp[11]) ? node21673 : node21668;
												assign node21668 = (inp[10]) ? 4'b0100 : node21669;
													assign node21669 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node21673 = (inp[7]) ? node21681 : node21674;
													assign node21674 = (inp[4]) ? node21676 : 4'b0100;
														assign node21676 = (inp[5]) ? node21678 : 4'b0100;
															assign node21678 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node21681 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node21684 = (inp[1]) ? node21696 : node21685;
												assign node21685 = (inp[11]) ? 4'b0101 : node21686;
													assign node21686 = (inp[7]) ? node21692 : node21687;
														assign node21687 = (inp[5]) ? 4'b0101 : node21688;
															assign node21688 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node21692 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node21696 = (inp[5]) ? node21704 : node21697;
													assign node21697 = (inp[4]) ? 4'b0101 : node21698;
														assign node21698 = (inp[11]) ? node21700 : 4'b0100;
															assign node21700 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node21704 = (inp[10]) ? 4'b0100 : node21705;
														assign node21705 = (inp[4]) ? 4'b0101 : 4'b0100;
										assign node21709 = (inp[10]) ? node21727 : node21710;
											assign node21710 = (inp[4]) ? node21722 : node21711;
												assign node21711 = (inp[5]) ? 4'b0100 : node21712;
													assign node21712 = (inp[0]) ? node21716 : node21713;
														assign node21713 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node21716 = (inp[1]) ? 4'b0101 : node21717;
															assign node21717 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node21722 = (inp[7]) ? 4'b0101 : node21723;
													assign node21723 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node21727 = (inp[4]) ? node21737 : node21728;
												assign node21728 = (inp[5]) ? 4'b0101 : node21729;
													assign node21729 = (inp[7]) ? node21733 : node21730;
														assign node21730 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node21733 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node21737 = (inp[7]) ? 4'b0100 : node21738;
													assign node21738 = (inp[5]) ? 4'b0100 : 4'b0101;
									assign node21742 = (inp[11]) ? node21766 : node21743;
										assign node21743 = (inp[13]) ? node21759 : node21744;
											assign node21744 = (inp[10]) ? node21756 : node21745;
												assign node21745 = (inp[4]) ? node21751 : node21746;
													assign node21746 = (inp[7]) ? node21748 : 4'b0100;
														assign node21748 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node21751 = (inp[7]) ? 4'b0101 : node21752;
														assign node21752 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node21756 = (inp[4]) ? 4'b0100 : 4'b0101;
											assign node21759 = (inp[10]) ? node21761 : 4'b0100;
												assign node21761 = (inp[5]) ? node21763 : 4'b0101;
													assign node21763 = (inp[4]) ? 4'b0100 : 4'b0101;
										assign node21766 = (inp[0]) ? node21776 : node21767;
											assign node21767 = (inp[10]) ? node21771 : node21768;
												assign node21768 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node21771 = (inp[4]) ? node21773 : 4'b0101;
													assign node21773 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node21776 = (inp[4]) ? node21786 : node21777;
												assign node21777 = (inp[10]) ? node21781 : node21778;
													assign node21778 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node21781 = (inp[5]) ? 4'b0101 : node21782;
														assign node21782 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node21786 = (inp[1]) ? node21796 : node21787;
													assign node21787 = (inp[10]) ? node21793 : node21788;
														assign node21788 = (inp[7]) ? 4'b0101 : node21789;
															assign node21789 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node21793 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node21796 = (inp[5]) ? 4'b0100 : node21797;
														assign node21797 = (inp[10]) ? 4'b0101 : 4'b0100;
							assign node21801 = (inp[15]) ? node21979 : node21802;
								assign node21802 = (inp[7]) ? node21896 : node21803;
									assign node21803 = (inp[5]) ? node21851 : node21804;
										assign node21804 = (inp[4]) ? node21830 : node21805;
											assign node21805 = (inp[1]) ? node21823 : node21806;
												assign node21806 = (inp[9]) ? node21814 : node21807;
													assign node21807 = (inp[10]) ? 4'b0000 : node21808;
														assign node21808 = (inp[11]) ? node21810 : 4'b0000;
															assign node21810 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node21814 = (inp[10]) ? node21816 : 4'b0000;
														assign node21816 = (inp[13]) ? node21820 : node21817;
															assign node21817 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node21820 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node21823 = (inp[13]) ? node21827 : node21824;
													assign node21824 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node21827 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node21830 = (inp[10]) ? node21836 : node21831;
												assign node21831 = (inp[13]) ? 4'b0100 : node21832;
													assign node21832 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node21836 = (inp[0]) ? node21844 : node21837;
													assign node21837 = (inp[11]) ? node21841 : node21838;
														assign node21838 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node21841 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node21844 = (inp[11]) ? 4'b0101 : node21845;
														assign node21845 = (inp[1]) ? 4'b0101 : node21846;
															assign node21846 = (inp[13]) ? 4'b0100 : 4'b0101;
										assign node21851 = (inp[0]) ? node21873 : node21852;
											assign node21852 = (inp[13]) ? node21866 : node21853;
												assign node21853 = (inp[10]) ? node21861 : node21854;
													assign node21854 = (inp[9]) ? node21856 : 4'b0100;
														assign node21856 = (inp[1]) ? 4'b0100 : node21857;
															assign node21857 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node21861 = (inp[11]) ? 4'b0101 : node21862;
														assign node21862 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node21866 = (inp[10]) ? 4'b0100 : node21867;
													assign node21867 = (inp[1]) ? 4'b0101 : node21868;
														assign node21868 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node21873 = (inp[1]) ? node21883 : node21874;
												assign node21874 = (inp[10]) ? node21876 : 4'b0101;
													assign node21876 = (inp[9]) ? node21878 : 4'b0100;
														assign node21878 = (inp[11]) ? 4'b0101 : node21879;
															assign node21879 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node21883 = (inp[4]) ? node21891 : node21884;
													assign node21884 = (inp[10]) ? node21888 : node21885;
														assign node21885 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node21888 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node21891 = (inp[13]) ? 4'b0100 : node21892;
														assign node21892 = (inp[9]) ? 4'b0100 : 4'b0101;
									assign node21896 = (inp[4]) ? node21936 : node21897;
										assign node21897 = (inp[5]) ? node21923 : node21898;
											assign node21898 = (inp[9]) ? node21914 : node21899;
												assign node21899 = (inp[1]) ? node21905 : node21900;
													assign node21900 = (inp[10]) ? node21902 : 4'b0100;
														assign node21902 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node21905 = (inp[13]) ? 4'b0100 : node21906;
														assign node21906 = (inp[10]) ? node21910 : node21907;
															assign node21907 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node21910 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node21914 = (inp[13]) ? node21916 : 4'b0101;
													assign node21916 = (inp[10]) ? 4'b0101 : node21917;
														assign node21917 = (inp[1]) ? node21919 : 4'b0100;
															assign node21919 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node21923 = (inp[11]) ? 4'b0000 : node21924;
												assign node21924 = (inp[0]) ? node21932 : node21925;
													assign node21925 = (inp[13]) ? 4'b0000 : node21926;
														assign node21926 = (inp[1]) ? 4'b0000 : node21927;
															assign node21927 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node21932 = (inp[13]) ? 4'b0001 : 4'b0000;
										assign node21936 = (inp[0]) ? node21962 : node21937;
											assign node21937 = (inp[9]) ? node21949 : node21938;
												assign node21938 = (inp[13]) ? node21946 : node21939;
													assign node21939 = (inp[10]) ? node21943 : node21940;
														assign node21940 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node21943 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node21946 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node21949 = (inp[1]) ? node21955 : node21950;
													assign node21950 = (inp[10]) ? node21952 : 4'b0000;
														assign node21952 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node21955 = (inp[13]) ? node21959 : node21956;
														assign node21956 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node21959 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node21962 = (inp[10]) ? node21968 : node21963;
												assign node21963 = (inp[13]) ? 4'b0001 : node21964;
													assign node21964 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node21968 = (inp[13]) ? node21974 : node21969;
													assign node21969 = (inp[11]) ? 4'b0001 : node21970;
														assign node21970 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node21974 = (inp[1]) ? 4'b0000 : node21975;
														assign node21975 = (inp[5]) ? 4'b0000 : 4'b0001;
								assign node21979 = (inp[10]) ? node21993 : node21980;
									assign node21980 = (inp[5]) ? 4'b0001 : node21981;
										assign node21981 = (inp[7]) ? node21987 : node21982;
											assign node21982 = (inp[4]) ? 4'b0000 : node21983;
												assign node21983 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node21987 = (inp[11]) ? 4'b0001 : node21988;
												assign node21988 = (inp[4]) ? 4'b0001 : 4'b0000;
									assign node21993 = (inp[5]) ? 4'b0000 : node21994;
										assign node21994 = (inp[7]) ? node22000 : node21995;
											assign node21995 = (inp[4]) ? 4'b0001 : node21996;
												assign node21996 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node22000 = (inp[11]) ? 4'b0000 : node22001;
												assign node22001 = (inp[4]) ? 4'b0000 : 4'b0001;
				assign node22006 = (inp[15]) ? node22886 : node22007;
					assign node22007 = (inp[14]) ? node22641 : node22008;
						assign node22008 = (inp[9]) ? node22374 : node22009;
							assign node22009 = (inp[10]) ? node22195 : node22010;
								assign node22010 = (inp[11]) ? node22100 : node22011;
									assign node22011 = (inp[13]) ? node22071 : node22012;
										assign node22012 = (inp[4]) ? node22040 : node22013;
											assign node22013 = (inp[1]) ? node22023 : node22014;
												assign node22014 = (inp[7]) ? node22018 : node22015;
													assign node22015 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node22018 = (inp[5]) ? 4'b0011 : node22019;
														assign node22019 = (inp[12]) ? 4'b0111 : 4'b0110;
												assign node22023 = (inp[7]) ? node22031 : node22024;
													assign node22024 = (inp[0]) ? 4'b0110 : node22025;
														assign node22025 = (inp[2]) ? node22027 : 4'b0111;
															assign node22027 = (inp[12]) ? 4'b0110 : 4'b0111;
													assign node22031 = (inp[5]) ? node22035 : node22032;
														assign node22032 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node22035 = (inp[2]) ? 4'b0010 : node22036;
															assign node22036 = (inp[12]) ? 4'b0011 : 4'b0010;
											assign node22040 = (inp[0]) ? node22056 : node22041;
												assign node22041 = (inp[1]) ? node22049 : node22042;
													assign node22042 = (inp[5]) ? node22044 : 4'b0010;
														assign node22044 = (inp[7]) ? 4'b0011 : node22045;
															assign node22045 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node22049 = (inp[7]) ? node22053 : node22050;
														assign node22050 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node22053 = (inp[5]) ? 4'b0010 : 4'b0110;
												assign node22056 = (inp[5]) ? node22064 : node22057;
													assign node22057 = (inp[7]) ? node22061 : node22058;
														assign node22058 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node22061 = (inp[12]) ? 4'b0111 : 4'b0110;
													assign node22064 = (inp[7]) ? 4'b0010 : node22065;
														assign node22065 = (inp[12]) ? 4'b0110 : node22066;
															assign node22066 = (inp[2]) ? 4'b0110 : 4'b0110;
										assign node22071 = (inp[2]) ? node22087 : node22072;
											assign node22072 = (inp[5]) ? node22076 : node22073;
												assign node22073 = (inp[7]) ? 4'b0111 : 4'b0011;
												assign node22076 = (inp[7]) ? node22082 : node22077;
													assign node22077 = (inp[12]) ? node22079 : 4'b0111;
														assign node22079 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node22082 = (inp[12]) ? 4'b0011 : node22083;
														assign node22083 = (inp[4]) ? 4'b0011 : 4'b0010;
											assign node22087 = (inp[5]) ? node22097 : node22088;
												assign node22088 = (inp[7]) ? node22092 : node22089;
													assign node22089 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node22092 = (inp[1]) ? node22094 : 4'b0111;
														assign node22094 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node22097 = (inp[7]) ? 4'b0011 : 4'b0111;
									assign node22100 = (inp[13]) ? node22158 : node22101;
										assign node22101 = (inp[12]) ? node22127 : node22102;
											assign node22102 = (inp[4]) ? node22118 : node22103;
												assign node22103 = (inp[0]) ? node22113 : node22104;
													assign node22104 = (inp[2]) ? node22108 : node22105;
														assign node22105 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node22108 = (inp[7]) ? node22110 : 4'b0110;
															assign node22110 = (inp[5]) ? 4'b0011 : 4'b0110;
													assign node22113 = (inp[2]) ? 4'b0011 : node22114;
														assign node22114 = (inp[7]) ? 4'b0011 : 4'b0111;
												assign node22118 = (inp[1]) ? node22122 : node22119;
													assign node22119 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node22122 = (inp[0]) ? node22124 : 4'b0011;
														assign node22124 = (inp[7]) ? 4'b0011 : 4'b0111;
											assign node22127 = (inp[2]) ? node22143 : node22128;
												assign node22128 = (inp[7]) ? node22136 : node22129;
													assign node22129 = (inp[5]) ? node22131 : 4'b0011;
														assign node22131 = (inp[1]) ? 4'b0110 : node22132;
															assign node22132 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node22136 = (inp[5]) ? node22138 : 4'b0110;
														assign node22138 = (inp[4]) ? 4'b0011 : node22139;
															assign node22139 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node22143 = (inp[0]) ? node22149 : node22144;
													assign node22144 = (inp[4]) ? node22146 : 4'b0011;
														assign node22146 = (inp[7]) ? 4'b0011 : 4'b0111;
													assign node22149 = (inp[1]) ? 4'b0111 : node22150;
														assign node22150 = (inp[7]) ? node22154 : node22151;
															assign node22151 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node22154 = (inp[5]) ? 4'b0011 : 4'b0110;
										assign node22158 = (inp[5]) ? node22174 : node22159;
											assign node22159 = (inp[7]) ? node22171 : node22160;
												assign node22160 = (inp[0]) ? 4'b0010 : node22161;
													assign node22161 = (inp[12]) ? node22165 : node22162;
														assign node22162 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node22165 = (inp[2]) ? 4'b0010 : node22166;
															assign node22166 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node22171 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node22174 = (inp[7]) ? node22186 : node22175;
												assign node22175 = (inp[4]) ? node22181 : node22176;
													assign node22176 = (inp[0]) ? 4'b0111 : node22177;
														assign node22177 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node22181 = (inp[1]) ? 4'b0110 : node22182;
														assign node22182 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node22186 = (inp[2]) ? 4'b0010 : node22187;
													assign node22187 = (inp[1]) ? 4'b0010 : node22188;
														assign node22188 = (inp[0]) ? 4'b0011 : node22189;
															assign node22189 = (inp[4]) ? 4'b0010 : 4'b0010;
								assign node22195 = (inp[5]) ? node22299 : node22196;
									assign node22196 = (inp[7]) ? node22254 : node22197;
										assign node22197 = (inp[0]) ? node22229 : node22198;
											assign node22198 = (inp[4]) ? node22218 : node22199;
												assign node22199 = (inp[1]) ? node22207 : node22200;
													assign node22200 = (inp[12]) ? 4'b0011 : node22201;
														assign node22201 = (inp[2]) ? node22203 : 4'b0011;
															assign node22203 = (inp[11]) ? 4'b0010 : 4'b0010;
													assign node22207 = (inp[2]) ? node22213 : node22208;
														assign node22208 = (inp[13]) ? 4'b0010 : node22209;
															assign node22209 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node22213 = (inp[12]) ? node22215 : 4'b0011;
															assign node22215 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node22218 = (inp[2]) ? 4'b0010 : node22219;
													assign node22219 = (inp[12]) ? 4'b0011 : node22220;
														assign node22220 = (inp[13]) ? node22224 : node22221;
															assign node22221 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node22224 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node22229 = (inp[4]) ? node22243 : node22230;
												assign node22230 = (inp[1]) ? 4'b0010 : node22231;
													assign node22231 = (inp[12]) ? node22237 : node22232;
														assign node22232 = (inp[11]) ? node22234 : 4'b0010;
															assign node22234 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node22237 = (inp[11]) ? 4'b0010 : node22238;
															assign node22238 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node22243 = (inp[1]) ? node22247 : node22244;
													assign node22244 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node22247 = (inp[11]) ? 4'b0011 : node22248;
														assign node22248 = (inp[2]) ? node22250 : 4'b0011;
															assign node22250 = (inp[13]) ? 4'b0010 : 4'b0011;
										assign node22254 = (inp[12]) ? node22274 : node22255;
											assign node22255 = (inp[2]) ? node22265 : node22256;
												assign node22256 = (inp[4]) ? 4'b0110 : node22257;
													assign node22257 = (inp[1]) ? node22261 : node22258;
														assign node22258 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node22261 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node22265 = (inp[11]) ? node22269 : node22266;
													assign node22266 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node22269 = (inp[4]) ? 4'b0111 : node22270;
														assign node22270 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node22274 = (inp[11]) ? node22288 : node22275;
												assign node22275 = (inp[13]) ? node22279 : node22276;
													assign node22276 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node22279 = (inp[1]) ? 4'b0111 : node22280;
														assign node22280 = (inp[0]) ? node22284 : node22281;
															assign node22281 = (inp[4]) ? 4'b0110 : 4'b0111;
															assign node22284 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node22288 = (inp[1]) ? node22296 : node22289;
													assign node22289 = (inp[4]) ? 4'b0110 : node22290;
														assign node22290 = (inp[0]) ? node22292 : 4'b0110;
															assign node22292 = (inp[2]) ? 4'b0110 : 4'b0110;
													assign node22296 = (inp[13]) ? 4'b0110 : 4'b0111;
									assign node22299 = (inp[7]) ? node22339 : node22300;
										assign node22300 = (inp[4]) ? node22320 : node22301;
											assign node22301 = (inp[1]) ? node22309 : node22302;
												assign node22302 = (inp[13]) ? node22306 : node22303;
													assign node22303 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node22306 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node22309 = (inp[0]) ? 4'b0110 : node22310;
													assign node22310 = (inp[2]) ? node22314 : node22311;
														assign node22311 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node22314 = (inp[11]) ? node22316 : 4'b0110;
															assign node22316 = (inp[12]) ? 4'b0110 : 4'b0110;
											assign node22320 = (inp[12]) ? node22334 : node22321;
												assign node22321 = (inp[1]) ? node22327 : node22322;
													assign node22322 = (inp[2]) ? 4'b0110 : node22323;
														assign node22323 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node22327 = (inp[2]) ? 4'b0111 : node22328;
														assign node22328 = (inp[13]) ? 4'b0110 : node22329;
															assign node22329 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node22334 = (inp[2]) ? node22336 : 4'b0110;
													assign node22336 = (inp[1]) ? 4'b0111 : 4'b0110;
										assign node22339 = (inp[13]) ? node22355 : node22340;
											assign node22340 = (inp[11]) ? node22350 : node22341;
												assign node22341 = (inp[1]) ? 4'b0010 : node22342;
													assign node22342 = (inp[12]) ? 4'b0010 : node22343;
														assign node22343 = (inp[4]) ? 4'b0011 : node22344;
															assign node22344 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node22350 = (inp[1]) ? 4'b0011 : node22351;
													assign node22351 = (inp[4]) ? 4'b0010 : 4'b0011;
											assign node22355 = (inp[11]) ? 4'b0010 : node22356;
												assign node22356 = (inp[1]) ? node22368 : node22357;
													assign node22357 = (inp[0]) ? node22363 : node22358;
														assign node22358 = (inp[2]) ? node22360 : 4'b0010;
															assign node22360 = (inp[12]) ? 4'b0011 : 4'b0010;
														assign node22363 = (inp[2]) ? 4'b0010 : node22364;
															assign node22364 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node22368 = (inp[12]) ? node22370 : 4'b0011;
														assign node22370 = (inp[2]) ? 4'b0011 : 4'b0010;
							assign node22374 = (inp[13]) ? node22500 : node22375;
								assign node22375 = (inp[11]) ? node22435 : node22376;
									assign node22376 = (inp[2]) ? node22398 : node22377;
										assign node22377 = (inp[12]) ? node22385 : node22378;
											assign node22378 = (inp[7]) ? node22382 : node22379;
												assign node22379 = (inp[5]) ? 4'b0110 : 4'b0010;
												assign node22382 = (inp[5]) ? 4'b0010 : 4'b0110;
											assign node22385 = (inp[5]) ? node22395 : node22386;
												assign node22386 = (inp[7]) ? node22392 : node22387;
													assign node22387 = (inp[10]) ? 4'b0010 : node22388;
														assign node22388 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node22392 = (inp[4]) ? 4'b0111 : 4'b0110;
												assign node22395 = (inp[7]) ? 4'b0011 : 4'b0111;
										assign node22398 = (inp[5]) ? node22420 : node22399;
											assign node22399 = (inp[7]) ? node22405 : node22400;
												assign node22400 = (inp[4]) ? 4'b0011 : node22401;
													assign node22401 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node22405 = (inp[12]) ? 4'b0110 : node22406;
													assign node22406 = (inp[10]) ? node22412 : node22407;
														assign node22407 = (inp[4]) ? 4'b0111 : node22408;
															assign node22408 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node22412 = (inp[0]) ? node22416 : node22413;
															assign node22413 = (inp[4]) ? 4'b0110 : 4'b0110;
															assign node22416 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node22420 = (inp[7]) ? node22428 : node22421;
												assign node22421 = (inp[1]) ? node22423 : 4'b0110;
													assign node22423 = (inp[4]) ? 4'b0110 : node22424;
														assign node22424 = (inp[12]) ? 4'b0110 : 4'b0111;
												assign node22428 = (inp[0]) ? node22430 : 4'b0010;
													assign node22430 = (inp[4]) ? node22432 : 4'b0010;
														assign node22432 = (inp[12]) ? 4'b0010 : 4'b0011;
									assign node22435 = (inp[12]) ? node22475 : node22436;
										assign node22436 = (inp[2]) ? node22452 : node22437;
											assign node22437 = (inp[5]) ? node22441 : node22438;
												assign node22438 = (inp[7]) ? 4'b0111 : 4'b0011;
												assign node22441 = (inp[7]) ? node22449 : node22442;
													assign node22442 = (inp[0]) ? 4'b0111 : node22443;
														assign node22443 = (inp[10]) ? 4'b0111 : node22444;
															assign node22444 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node22449 = (inp[4]) ? 4'b0011 : 4'b0010;
											assign node22452 = (inp[4]) ? node22466 : node22453;
												assign node22453 = (inp[1]) ? node22459 : node22454;
													assign node22454 = (inp[7]) ? 4'b0111 : node22455;
														assign node22455 = (inp[0]) ? 4'b0011 : 4'b0111;
													assign node22459 = (inp[5]) ? node22463 : node22460;
														assign node22460 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node22463 = (inp[7]) ? 4'b0011 : 4'b0110;
												assign node22466 = (inp[0]) ? 4'b0111 : node22467;
													assign node22467 = (inp[1]) ? node22469 : 4'b0010;
														assign node22469 = (inp[10]) ? 4'b0111 : node22470;
															assign node22470 = (inp[7]) ? 4'b0111 : 4'b0011;
										assign node22475 = (inp[2]) ? node22493 : node22476;
											assign node22476 = (inp[1]) ? node22486 : node22477;
												assign node22477 = (inp[7]) ? node22481 : node22478;
													assign node22478 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node22481 = (inp[5]) ? node22483 : 4'b0110;
														assign node22483 = (inp[4]) ? 4'b0010 : 4'b0011;
												assign node22486 = (inp[4]) ? 4'b0111 : node22487;
													assign node22487 = (inp[5]) ? node22489 : 4'b0010;
														assign node22489 = (inp[7]) ? 4'b0010 : 4'b0110;
											assign node22493 = (inp[5]) ? node22497 : node22494;
												assign node22494 = (inp[7]) ? 4'b0111 : 4'b0011;
												assign node22497 = (inp[7]) ? 4'b0011 : 4'b0111;
								assign node22500 = (inp[11]) ? node22560 : node22501;
									assign node22501 = (inp[5]) ? node22527 : node22502;
										assign node22502 = (inp[7]) ? node22514 : node22503;
											assign node22503 = (inp[10]) ? 4'b0011 : node22504;
												assign node22504 = (inp[1]) ? node22510 : node22505;
													assign node22505 = (inp[0]) ? node22507 : 4'b0011;
														assign node22507 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node22510 = (inp[12]) ? 4'b0010 : 4'b0011;
											assign node22514 = (inp[2]) ? node22516 : 4'b0111;
												assign node22516 = (inp[4]) ? node22522 : node22517;
													assign node22517 = (inp[1]) ? 4'b0110 : node22518;
														assign node22518 = (inp[12]) ? 4'b0110 : 4'b0111;
													assign node22522 = (inp[12]) ? 4'b0111 : node22523;
														assign node22523 = (inp[1]) ? 4'b0111 : 4'b0110;
										assign node22527 = (inp[7]) ? node22537 : node22528;
											assign node22528 = (inp[10]) ? node22530 : 4'b0111;
												assign node22530 = (inp[2]) ? 4'b0111 : node22531;
													assign node22531 = (inp[1]) ? node22533 : 4'b0111;
														assign node22533 = (inp[12]) ? 4'b0111 : 4'b0110;
											assign node22537 = (inp[1]) ? node22553 : node22538;
												assign node22538 = (inp[12]) ? node22548 : node22539;
													assign node22539 = (inp[10]) ? 4'b0010 : node22540;
														assign node22540 = (inp[4]) ? node22544 : node22541;
															assign node22541 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node22544 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node22548 = (inp[2]) ? 4'b0011 : node22549;
														assign node22549 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node22553 = (inp[2]) ? 4'b0011 : node22554;
													assign node22554 = (inp[4]) ? 4'b0011 : node22555;
														assign node22555 = (inp[0]) ? 4'b0010 : 4'b0011;
									assign node22560 = (inp[2]) ? node22598 : node22561;
										assign node22561 = (inp[12]) ? node22575 : node22562;
											assign node22562 = (inp[5]) ? node22566 : node22563;
												assign node22563 = (inp[7]) ? 4'b0110 : 4'b0010;
												assign node22566 = (inp[7]) ? node22570 : node22567;
													assign node22567 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node22570 = (inp[1]) ? 4'b0010 : node22571;
														assign node22571 = (inp[4]) ? 4'b0010 : 4'b0011;
											assign node22575 = (inp[5]) ? node22589 : node22576;
												assign node22576 = (inp[7]) ? node22584 : node22577;
													assign node22577 = (inp[0]) ? node22579 : 4'b0011;
														assign node22579 = (inp[4]) ? 4'b0010 : node22580;
															assign node22580 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node22584 = (inp[10]) ? node22586 : 4'b0110;
														assign node22586 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node22589 = (inp[7]) ? node22593 : node22590;
													assign node22590 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node22593 = (inp[1]) ? 4'b0011 : node22594;
														assign node22594 = (inp[4]) ? 4'b0011 : 4'b0010;
										assign node22598 = (inp[4]) ? node22618 : node22599;
											assign node22599 = (inp[12]) ? node22605 : node22600;
												assign node22600 = (inp[1]) ? 4'b0111 : node22601;
													assign node22601 = (inp[7]) ? 4'b0110 : 4'b0010;
												assign node22605 = (inp[1]) ? node22613 : node22606;
													assign node22606 = (inp[7]) ? node22610 : node22607;
														assign node22607 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node22610 = (inp[0]) ? 4'b0111 : 4'b0010;
													assign node22613 = (inp[5]) ? node22615 : 4'b0110;
														assign node22615 = (inp[7]) ? 4'b0010 : 4'b0110;
											assign node22618 = (inp[1]) ? node22632 : node22619;
												assign node22619 = (inp[12]) ? node22627 : node22620;
													assign node22620 = (inp[5]) ? node22624 : node22621;
														assign node22621 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node22624 = (inp[7]) ? 4'b0011 : 4'b0110;
													assign node22627 = (inp[0]) ? 4'b0110 : node22628;
														assign node22628 = (inp[5]) ? 4'b0010 : 4'b0110;
												assign node22632 = (inp[0]) ? node22634 : 4'b0010;
													assign node22634 = (inp[7]) ? 4'b0110 : node22635;
														assign node22635 = (inp[12]) ? 4'b0011 : node22636;
															assign node22636 = (inp[5]) ? 4'b0110 : 4'b0010;
						assign node22641 = (inp[7]) ? node22827 : node22642;
							assign node22642 = (inp[12]) ? node22674 : node22643;
								assign node22643 = (inp[4]) ? node22667 : node22644;
									assign node22644 = (inp[2]) ? node22656 : node22645;
										assign node22645 = (inp[13]) ? node22651 : node22646;
											assign node22646 = (inp[5]) ? node22648 : 4'b0000;
												assign node22648 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node22651 = (inp[1]) ? node22653 : 4'b0001;
												assign node22653 = (inp[5]) ? 4'b0000 : 4'b0001;
										assign node22656 = (inp[13]) ? node22662 : node22657;
											assign node22657 = (inp[1]) ? node22659 : 4'b0001;
												assign node22659 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node22662 = (inp[1]) ? node22664 : 4'b0000;
												assign node22664 = (inp[5]) ? 4'b0001 : 4'b0000;
									assign node22667 = (inp[13]) ? node22671 : node22668;
										assign node22668 = (inp[5]) ? 4'b0101 : 4'b0100;
										assign node22671 = (inp[5]) ? 4'b0100 : 4'b0101;
								assign node22674 = (inp[9]) ? node22756 : node22675;
									assign node22675 = (inp[1]) ? node22733 : node22676;
										assign node22676 = (inp[11]) ? node22700 : node22677;
											assign node22677 = (inp[10]) ? node22689 : node22678;
												assign node22678 = (inp[4]) ? node22682 : node22679;
													assign node22679 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node22682 = (inp[0]) ? node22684 : 4'b0101;
														assign node22684 = (inp[2]) ? 4'b0101 : node22685;
															assign node22685 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node22689 = (inp[5]) ? node22695 : node22690;
													assign node22690 = (inp[13]) ? 4'b0101 : node22691;
														assign node22691 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node22695 = (inp[2]) ? node22697 : 4'b0100;
														assign node22697 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node22700 = (inp[0]) ? node22716 : node22701;
												assign node22701 = (inp[5]) ? node22707 : node22702;
													assign node22702 = (inp[13]) ? node22704 : 4'b0100;
														assign node22704 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node22707 = (inp[2]) ? node22713 : node22708;
														assign node22708 = (inp[10]) ? node22710 : 4'b0100;
															assign node22710 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node22713 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node22716 = (inp[10]) ? node22728 : node22717;
													assign node22717 = (inp[2]) ? node22723 : node22718;
														assign node22718 = (inp[4]) ? node22720 : 4'b0100;
															assign node22720 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node22723 = (inp[13]) ? 4'b0100 : node22724;
															assign node22724 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node22728 = (inp[2]) ? 4'b0101 : node22729;
														assign node22729 = (inp[4]) ? 4'b0100 : 4'b0101;
										assign node22733 = (inp[13]) ? node22745 : node22734;
											assign node22734 = (inp[5]) ? node22740 : node22735;
												assign node22735 = (inp[2]) ? 4'b0100 : node22736;
													assign node22736 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node22740 = (inp[2]) ? 4'b0101 : node22741;
													assign node22741 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node22745 = (inp[5]) ? node22751 : node22746;
												assign node22746 = (inp[2]) ? 4'b0101 : node22747;
													assign node22747 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node22751 = (inp[2]) ? 4'b0100 : node22752;
													assign node22752 = (inp[4]) ? 4'b0100 : 4'b0101;
									assign node22756 = (inp[1]) ? node22796 : node22757;
										assign node22757 = (inp[11]) ? node22775 : node22758;
											assign node22758 = (inp[2]) ? node22766 : node22759;
												assign node22759 = (inp[13]) ? node22761 : 4'b0100;
													assign node22761 = (inp[0]) ? 4'b0101 : node22762;
														assign node22762 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node22766 = (inp[13]) ? node22772 : node22767;
													assign node22767 = (inp[10]) ? 4'b0101 : node22768;
														assign node22768 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node22772 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node22775 = (inp[4]) ? node22783 : node22776;
												assign node22776 = (inp[13]) ? node22780 : node22777;
													assign node22777 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node22780 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node22783 = (inp[2]) ? node22789 : node22784;
													assign node22784 = (inp[0]) ? node22786 : 4'b0101;
														assign node22786 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node22789 = (inp[10]) ? 4'b0100 : node22790;
														assign node22790 = (inp[0]) ? 4'b0100 : node22791;
															assign node22791 = (inp[13]) ? 4'b0100 : 4'b0101;
										assign node22796 = (inp[10]) ? node22810 : node22797;
											assign node22797 = (inp[5]) ? node22803 : node22798;
												assign node22798 = (inp[13]) ? node22800 : 4'b0100;
													assign node22800 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node22803 = (inp[13]) ? 4'b0100 : node22804;
													assign node22804 = (inp[4]) ? 4'b0101 : node22805;
														assign node22805 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node22810 = (inp[13]) ? node22822 : node22811;
												assign node22811 = (inp[5]) ? node22817 : node22812;
													assign node22812 = (inp[2]) ? 4'b0100 : node22813;
														assign node22813 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node22817 = (inp[2]) ? 4'b0101 : node22818;
														assign node22818 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node22822 = (inp[5]) ? 4'b0100 : node22823;
													assign node22823 = (inp[2]) ? 4'b0101 : 4'b0100;
							assign node22827 = (inp[12]) ? node22859 : node22828;
								assign node22828 = (inp[4]) ? node22852 : node22829;
									assign node22829 = (inp[13]) ? node22841 : node22830;
										assign node22830 = (inp[2]) ? node22836 : node22831;
											assign node22831 = (inp[5]) ? node22833 : 4'b0100;
												assign node22833 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node22836 = (inp[5]) ? node22838 : 4'b0101;
												assign node22838 = (inp[1]) ? 4'b0101 : 4'b0100;
										assign node22841 = (inp[2]) ? node22847 : node22842;
											assign node22842 = (inp[5]) ? node22844 : 4'b0101;
												assign node22844 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node22847 = (inp[5]) ? node22849 : 4'b0100;
												assign node22849 = (inp[1]) ? 4'b0100 : 4'b0101;
									assign node22852 = (inp[13]) ? node22856 : node22853;
										assign node22853 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node22856 = (inp[1]) ? 4'b0000 : 4'b0001;
								assign node22859 = (inp[13]) ? node22873 : node22860;
									assign node22860 = (inp[4]) ? 4'b0001 : node22861;
										assign node22861 = (inp[2]) ? node22867 : node22862;
											assign node22862 = (inp[5]) ? 4'b0000 : node22863;
												assign node22863 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node22867 = (inp[5]) ? 4'b0001 : node22868;
												assign node22868 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node22873 = (inp[4]) ? 4'b0000 : node22874;
										assign node22874 = (inp[2]) ? node22880 : node22875;
											assign node22875 = (inp[5]) ? 4'b0001 : node22876;
												assign node22876 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node22880 = (inp[1]) ? 4'b0000 : node22881;
												assign node22881 = (inp[5]) ? 4'b0000 : 4'b0001;
					assign node22886 = (inp[5]) ? node23264 : node22887;
						assign node22887 = (inp[14]) ? node23177 : node22888;
							assign node22888 = (inp[12]) ? node23070 : node22889;
								assign node22889 = (inp[4]) ? node22999 : node22890;
									assign node22890 = (inp[9]) ? node22956 : node22891;
										assign node22891 = (inp[7]) ? node22927 : node22892;
											assign node22892 = (inp[0]) ? node22906 : node22893;
												assign node22893 = (inp[10]) ? node22901 : node22894;
													assign node22894 = (inp[11]) ? node22898 : node22895;
														assign node22895 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node22898 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node22901 = (inp[1]) ? node22903 : 4'b0001;
														assign node22903 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node22906 = (inp[10]) ? node22914 : node22907;
													assign node22907 = (inp[2]) ? node22909 : 4'b0001;
														assign node22909 = (inp[11]) ? node22911 : 4'b0000;
															assign node22911 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node22914 = (inp[2]) ? node22920 : node22915;
														assign node22915 = (inp[13]) ? node22917 : 4'b0000;
															assign node22917 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node22920 = (inp[1]) ? node22924 : node22921;
															assign node22921 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node22924 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node22927 = (inp[13]) ? node22943 : node22928;
												assign node22928 = (inp[10]) ? node22934 : node22929;
													assign node22929 = (inp[1]) ? 4'b0001 : node22930;
														assign node22930 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node22934 = (inp[1]) ? node22936 : 4'b0001;
														assign node22936 = (inp[2]) ? node22940 : node22937;
															assign node22937 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node22940 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node22943 = (inp[10]) ? node22951 : node22944;
													assign node22944 = (inp[11]) ? 4'b0000 : node22945;
														assign node22945 = (inp[0]) ? 4'b0001 : node22946;
															assign node22946 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node22951 = (inp[2]) ? node22953 : 4'b0001;
														assign node22953 = (inp[1]) ? 4'b0001 : 4'b0000;
										assign node22956 = (inp[0]) ? node22978 : node22957;
											assign node22957 = (inp[2]) ? 4'b0000 : node22958;
												assign node22958 = (inp[10]) ? node22968 : node22959;
													assign node22959 = (inp[13]) ? 4'b0001 : node22960;
														assign node22960 = (inp[1]) ? node22964 : node22961;
															assign node22961 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node22964 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node22968 = (inp[7]) ? 4'b0000 : node22969;
														assign node22969 = (inp[1]) ? node22973 : node22970;
															assign node22970 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node22973 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node22978 = (inp[11]) ? node22990 : node22979;
												assign node22979 = (inp[1]) ? node22985 : node22980;
													assign node22980 = (inp[7]) ? node22982 : 4'b0000;
														assign node22982 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node22985 = (inp[7]) ? node22987 : 4'b0001;
														assign node22987 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node22990 = (inp[1]) ? node22992 : 4'b0001;
													assign node22992 = (inp[13]) ? node22994 : 4'b0001;
														assign node22994 = (inp[2]) ? node22996 : 4'b0000;
															assign node22996 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node22999 = (inp[10]) ? node23035 : node23000;
										assign node23000 = (inp[0]) ? node23018 : node23001;
											assign node23001 = (inp[1]) ? node23007 : node23002;
												assign node23002 = (inp[11]) ? 4'b0101 : node23003;
													assign node23003 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node23007 = (inp[11]) ? node23013 : node23008;
													assign node23008 = (inp[2]) ? node23010 : 4'b0101;
														assign node23010 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node23013 = (inp[2]) ? node23015 : 4'b0100;
														assign node23015 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node23018 = (inp[7]) ? node23022 : node23019;
												assign node23019 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node23022 = (inp[13]) ? node23028 : node23023;
													assign node23023 = (inp[1]) ? 4'b0101 : node23024;
														assign node23024 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node23028 = (inp[2]) ? 4'b0101 : node23029;
														assign node23029 = (inp[9]) ? node23031 : 4'b0100;
															assign node23031 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node23035 = (inp[7]) ? node23063 : node23036;
											assign node23036 = (inp[9]) ? node23046 : node23037;
												assign node23037 = (inp[13]) ? node23041 : node23038;
													assign node23038 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node23041 = (inp[11]) ? node23043 : 4'b0101;
														assign node23043 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node23046 = (inp[13]) ? node23058 : node23047;
													assign node23047 = (inp[1]) ? node23053 : node23048;
														assign node23048 = (inp[0]) ? node23050 : 4'b0100;
															assign node23050 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node23053 = (inp[11]) ? node23055 : 4'b0101;
															assign node23055 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node23058 = (inp[2]) ? node23060 : 4'b0100;
														assign node23060 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node23063 = (inp[11]) ? node23067 : node23064;
												assign node23064 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node23067 = (inp[1]) ? 4'b0100 : 4'b0101;
								assign node23070 = (inp[13]) ? node23146 : node23071;
									assign node23071 = (inp[9]) ? node23107 : node23072;
										assign node23072 = (inp[0]) ? node23094 : node23073;
											assign node23073 = (inp[4]) ? node23081 : node23074;
												assign node23074 = (inp[11]) ? node23078 : node23075;
													assign node23075 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node23078 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node23081 = (inp[10]) ? node23089 : node23082;
													assign node23082 = (inp[11]) ? node23086 : node23083;
														assign node23083 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node23086 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node23089 = (inp[7]) ? 4'b0100 : node23090;
														assign node23090 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node23094 = (inp[1]) ? node23102 : node23095;
												assign node23095 = (inp[7]) ? node23099 : node23096;
													assign node23096 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node23099 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node23102 = (inp[7]) ? node23104 : 4'b0101;
													assign node23104 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node23107 = (inp[10]) ? node23125 : node23108;
											assign node23108 = (inp[2]) ? node23114 : node23109;
												assign node23109 = (inp[7]) ? 4'b0100 : node23110;
													assign node23110 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node23114 = (inp[1]) ? node23120 : node23115;
													assign node23115 = (inp[4]) ? node23117 : 4'b0100;
														assign node23117 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node23120 = (inp[0]) ? 4'b0101 : node23121;
														assign node23121 = (inp[4]) ? 4'b0101 : 4'b0100;
											assign node23125 = (inp[1]) ? node23139 : node23126;
												assign node23126 = (inp[2]) ? node23132 : node23127;
													assign node23127 = (inp[11]) ? node23129 : 4'b0100;
														assign node23129 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node23132 = (inp[11]) ? node23136 : node23133;
														assign node23133 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node23136 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node23139 = (inp[7]) ? node23143 : node23140;
													assign node23140 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node23143 = (inp[11]) ? 4'b0100 : 4'b0101;
									assign node23146 = (inp[0]) ? node23170 : node23147;
										assign node23147 = (inp[2]) ? node23155 : node23148;
											assign node23148 = (inp[7]) ? node23152 : node23149;
												assign node23149 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node23152 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node23155 = (inp[9]) ? 4'b0101 : node23156;
												assign node23156 = (inp[10]) ? node23164 : node23157;
													assign node23157 = (inp[11]) ? node23161 : node23158;
														assign node23158 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node23161 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node23164 = (inp[7]) ? node23166 : 4'b0101;
														assign node23166 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node23170 = (inp[11]) ? node23174 : node23171;
											assign node23171 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node23174 = (inp[7]) ? 4'b0100 : 4'b0101;
							assign node23177 = (inp[4]) ? node23253 : node23178;
								assign node23178 = (inp[12]) ? node23216 : node23179;
									assign node23179 = (inp[9]) ? node23209 : node23180;
										assign node23180 = (inp[7]) ? node23194 : node23181;
											assign node23181 = (inp[11]) ? node23189 : node23182;
												assign node23182 = (inp[2]) ? node23186 : node23183;
													assign node23183 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node23186 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node23189 = (inp[2]) ? node23191 : 4'b0100;
													assign node23191 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node23194 = (inp[10]) ? node23202 : node23195;
												assign node23195 = (inp[2]) ? node23199 : node23196;
													assign node23196 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node23199 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node23202 = (inp[2]) ? node23206 : node23203;
													assign node23203 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node23206 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node23209 = (inp[2]) ? node23213 : node23210;
											assign node23210 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node23213 = (inp[1]) ? 4'b0100 : 4'b0101;
									assign node23216 = (inp[13]) ? node23246 : node23217;
										assign node23217 = (inp[0]) ? node23239 : node23218;
											assign node23218 = (inp[11]) ? node23232 : node23219;
												assign node23219 = (inp[1]) ? node23227 : node23220;
													assign node23220 = (inp[7]) ? node23224 : node23221;
														assign node23221 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node23224 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node23227 = (inp[7]) ? node23229 : 4'b0001;
														assign node23229 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node23232 = (inp[9]) ? node23234 : 4'b0001;
													assign node23234 = (inp[10]) ? node23236 : 4'b0001;
														assign node23236 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node23239 = (inp[7]) ? node23243 : node23240;
												assign node23240 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node23243 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node23246 = (inp[2]) ? node23250 : node23247;
											assign node23247 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node23250 = (inp[7]) ? 4'b0000 : 4'b0001;
								assign node23253 = (inp[7]) ? node23259 : node23254;
									assign node23254 = (inp[12]) ? 4'b0001 : node23255;
										assign node23255 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node23259 = (inp[1]) ? 4'b0000 : node23260;
										assign node23260 = (inp[12]) ? 4'b0000 : 4'b0001;
						assign node23264 = (inp[4]) ? node23326 : node23265;
							assign node23265 = (inp[12]) ? node23315 : node23266;
								assign node23266 = (inp[11]) ? node23300 : node23267;
									assign node23267 = (inp[1]) ? node23291 : node23268;
										assign node23268 = (inp[13]) ? node23282 : node23269;
											assign node23269 = (inp[7]) ? node23275 : node23270;
												assign node23270 = (inp[14]) ? node23272 : 4'b0100;
													assign node23272 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node23275 = (inp[14]) ? node23279 : node23276;
													assign node23276 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node23279 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node23282 = (inp[2]) ? node23288 : node23283;
												assign node23283 = (inp[7]) ? node23285 : 4'b0100;
													assign node23285 = (inp[14]) ? 4'b0100 : 4'b0101;
												assign node23288 = (inp[14]) ? 4'b0101 : 4'b0100;
										assign node23291 = (inp[14]) ? node23297 : node23292;
											assign node23292 = (inp[2]) ? 4'b0101 : node23293;
												assign node23293 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node23297 = (inp[2]) ? 4'b0100 : 4'b0101;
									assign node23300 = (inp[1]) ? node23308 : node23301;
										assign node23301 = (inp[2]) ? 4'b0101 : node23302;
											assign node23302 = (inp[14]) ? 4'b0100 : node23303;
												assign node23303 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node23308 = (inp[2]) ? 4'b0100 : node23309;
											assign node23309 = (inp[7]) ? 4'b0101 : node23310;
												assign node23310 = (inp[14]) ? 4'b0101 : 4'b0100;
								assign node23315 = (inp[2]) ? node23321 : node23316;
									assign node23316 = (inp[14]) ? 4'b0001 : node23317;
										assign node23317 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node23321 = (inp[14]) ? 4'b0000 : node23322;
										assign node23322 = (inp[11]) ? 4'b0000 : 4'b0001;
							assign node23326 = (inp[1]) ? node23346 : node23327;
								assign node23327 = (inp[12]) ? node23341 : node23328;
									assign node23328 = (inp[14]) ? 4'b0001 : node23329;
										assign node23329 = (inp[11]) ? node23335 : node23330;
											assign node23330 = (inp[2]) ? 4'b0000 : node23331;
												assign node23331 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node23335 = (inp[7]) ? 4'b0001 : node23336;
												assign node23336 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node23341 = (inp[11]) ? 4'b0000 : node23342;
										assign node23342 = (inp[14]) ? 4'b0000 : 4'b0001;
								assign node23346 = (inp[14]) ? 4'b0000 : node23347;
									assign node23347 = (inp[11]) ? node23355 : node23348;
										assign node23348 = (inp[12]) ? 4'b0001 : node23349;
											assign node23349 = (inp[7]) ? 4'b0001 : node23350;
												assign node23350 = (inp[2]) ? 4'b0001 : 4'b0000;
										assign node23355 = (inp[12]) ? 4'b0000 : node23356;
											assign node23356 = (inp[7]) ? 4'b0000 : node23357;
												assign node23357 = (inp[2]) ? 4'b0000 : 4'b0001;

endmodule