module dtc_split05_bm15 (
	input  wire [15-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node6;
	wire [1-1:0] node8;
	wire [1-1:0] node10;
	wire [1-1:0] node12;
	wire [1-1:0] node15;
	wire [1-1:0] node16;
	wire [1-1:0] node18;
	wire [1-1:0] node20;
	wire [1-1:0] node21;
	wire [1-1:0] node23;
	wire [1-1:0] node27;
	wire [1-1:0] node28;
	wire [1-1:0] node30;
	wire [1-1:0] node32;
	wire [1-1:0] node34;
	wire [1-1:0] node35;
	wire [1-1:0] node39;
	wire [1-1:0] node40;
	wire [1-1:0] node41;
	wire [1-1:0] node43;
	wire [1-1:0] node46;
	wire [1-1:0] node47;
	wire [1-1:0] node51;
	wire [1-1:0] node52;
	wire [1-1:0] node56;
	wire [1-1:0] node57;
	wire [1-1:0] node58;
	wire [1-1:0] node60;
	wire [1-1:0] node62;
	wire [1-1:0] node64;
	wire [1-1:0] node67;
	wire [1-1:0] node68;
	wire [1-1:0] node70;
	wire [1-1:0] node71;
	wire [1-1:0] node73;
	wire [1-1:0] node76;
	wire [1-1:0] node79;
	wire [1-1:0] node80;
	wire [1-1:0] node81;
	wire [1-1:0] node83;
	wire [1-1:0] node85;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node93;
	wire [1-1:0] node94;
	wire [1-1:0] node96;
	wire [1-1:0] node100;
	wire [1-1:0] node101;
	wire [1-1:0] node102;
	wire [1-1:0] node104;
	wire [1-1:0] node105;
	wire [1-1:0] node107;
	wire [1-1:0] node110;
	wire [1-1:0] node113;
	wire [1-1:0] node114;
	wire [1-1:0] node116;
	wire [1-1:0] node117;
	wire [1-1:0] node119;
	wire [1-1:0] node121;
	wire [1-1:0] node122;
	wire [1-1:0] node127;
	wire [1-1:0] node128;
	wire [1-1:0] node129;
	wire [1-1:0] node131;
	wire [1-1:0] node136;
	wire [1-1:0] node137;
	wire [1-1:0] node138;
	wire [1-1:0] node140;
	wire [1-1:0] node143;
	wire [1-1:0] node144;
	wire [1-1:0] node148;
	wire [1-1:0] node149;
	wire [1-1:0] node150;
	wire [1-1:0] node151;
	wire [1-1:0] node153;
	wire [1-1:0] node159;
	wire [1-1:0] node160;
	wire [1-1:0] node161;
	wire [1-1:0] node162;
	wire [1-1:0] node164;
	wire [1-1:0] node166;
	wire [1-1:0] node168;
	wire [1-1:0] node171;
	wire [1-1:0] node172;
	wire [1-1:0] node174;
	wire [1-1:0] node175;
	wire [1-1:0] node176;
	wire [1-1:0] node178;
	wire [1-1:0] node182;
	wire [1-1:0] node183;
	wire [1-1:0] node184;
	wire [1-1:0] node189;
	wire [1-1:0] node190;
	wire [1-1:0] node192;
	wire [1-1:0] node193;
	wire [1-1:0] node195;
	wire [1-1:0] node199;
	wire [1-1:0] node200;
	wire [1-1:0] node201;
	wire [1-1:0] node206;
	wire [1-1:0] node207;
	wire [1-1:0] node208;
	wire [1-1:0] node210;
	wire [1-1:0] node212;
	wire [1-1:0] node213;
	wire [1-1:0] node217;
	wire [1-1:0] node218;
	wire [1-1:0] node220;
	wire [1-1:0] node223;
	wire [1-1:0] node224;
	wire [1-1:0] node226;
	wire [1-1:0] node230;
	wire [1-1:0] node231;
	wire [1-1:0] node232;
	wire [1-1:0] node234;
	wire [1-1:0] node235;
	wire [1-1:0] node237;
	wire [1-1:0] node240;
	wire [1-1:0] node241;
	wire [1-1:0] node245;
	wire [1-1:0] node246;
	wire [1-1:0] node248;
	wire [1-1:0] node249;
	wire [1-1:0] node254;
	wire [1-1:0] node255;
	wire [1-1:0] node256;
	wire [1-1:0] node261;
	wire [1-1:0] node262;
	wire [1-1:0] node263;
	wire [1-1:0] node264;
	wire [1-1:0] node266;
	wire [1-1:0] node268;
	wire [1-1:0] node270;
	wire [1-1:0] node272;
	wire [1-1:0] node275;
	wire [1-1:0] node276;
	wire [1-1:0] node278;
	wire [1-1:0] node280;
	wire [1-1:0] node283;
	wire [1-1:0] node284;
	wire [1-1:0] node286;
	wire [1-1:0] node287;
	wire [1-1:0] node292;
	wire [1-1:0] node293;
	wire [1-1:0] node294;
	wire [1-1:0] node296;
	wire [1-1:0] node298;
	wire [1-1:0] node299;
	wire [1-1:0] node303;
	wire [1-1:0] node304;
	wire [1-1:0] node306;
	wire [1-1:0] node307;
	wire [1-1:0] node311;
	wire [1-1:0] node312;
	wire [1-1:0] node316;
	wire [1-1:0] node317;
	wire [1-1:0] node318;
	wire [1-1:0] node319;
	wire [1-1:0] node321;
	wire [1-1:0] node327;
	wire [1-1:0] node328;
	wire [1-1:0] node329;
	wire [1-1:0] node330;
	wire [1-1:0] node332;
	wire [1-1:0] node335;
	wire [1-1:0] node336;
	wire [1-1:0] node338;
	wire [1-1:0] node342;
	wire [1-1:0] node343;
	wire [1-1:0] node347;
	wire [1-1:0] node348;
	wire [1-1:0] node349;
	wire [1-1:0] node351;
	wire [1-1:0] node352;
	wire [1-1:0] node358;
	wire [1-1:0] node359;
	wire [1-1:0] node360;
	wire [1-1:0] node361;
	wire [1-1:0] node362;
	wire [1-1:0] node364;
	wire [1-1:0] node366;
	wire [1-1:0] node368;
	wire [1-1:0] node370;
	wire [1-1:0] node373;
	wire [1-1:0] node374;
	wire [1-1:0] node376;
	wire [1-1:0] node378;
	wire [1-1:0] node379;
	wire [1-1:0] node383;
	wire [1-1:0] node384;
	wire [1-1:0] node386;
	wire [1-1:0] node389;
	wire [1-1:0] node390;
	wire [1-1:0] node394;
	wire [1-1:0] node395;
	wire [1-1:0] node396;
	wire [1-1:0] node398;
	wire [1-1:0] node399;
	wire [1-1:0] node401;
	wire [1-1:0] node404;
	wire [1-1:0] node405;
	wire [1-1:0] node407;
	wire [1-1:0] node410;
	wire [1-1:0] node411;
	wire [1-1:0] node415;
	wire [1-1:0] node416;
	wire [1-1:0] node417;
	wire [1-1:0] node419;
	wire [1-1:0] node422;
	wire [1-1:0] node423;
	wire [1-1:0] node425;
	wire [1-1:0] node429;
	wire [1-1:0] node430;
	wire [1-1:0] node431;
	wire [1-1:0] node433;
	wire [1-1:0] node438;
	wire [1-1:0] node439;
	wire [1-1:0] node441;
	wire [1-1:0] node442;
	wire [1-1:0] node444;
	wire [1-1:0] node448;
	wire [1-1:0] node449;
	wire [1-1:0] node450;
	wire [1-1:0] node452;
	wire [1-1:0] node453;
	wire [1-1:0] node457;
	wire [1-1:0] node458;
	wire [1-1:0] node459;
	wire [1-1:0] node465;
	wire [1-1:0] node466;
	wire [1-1:0] node467;
	wire [1-1:0] node468;
	wire [1-1:0] node470;
	wire [1-1:0] node471;
	wire [1-1:0] node473;
	wire [1-1:0] node476;
	wire [1-1:0] node479;
	wire [1-1:0] node480;
	wire [1-1:0] node481;
	wire [1-1:0] node482;
	wire [1-1:0] node486;
	wire [1-1:0] node487;
	wire [1-1:0] node492;
	wire [1-1:0] node493;
	wire [1-1:0] node494;
	wire [1-1:0] node496;
	wire [1-1:0] node499;
	wire [1-1:0] node500;
	wire [1-1:0] node501;
	wire [1-1:0] node503;
	wire [1-1:0] node508;
	wire [1-1:0] node510;
	wire [1-1:0] node511;
	wire [1-1:0] node513;
	wire [1-1:0] node515;
	wire [1-1:0] node519;
	wire [1-1:0] node520;
	wire [1-1:0] node521;
	wire [1-1:0] node522;
	wire [1-1:0] node524;
	wire [1-1:0] node526;
	wire [1-1:0] node529;
	wire [1-1:0] node530;
	wire [1-1:0] node532;
	wire [1-1:0] node535;
	wire [1-1:0] node536;
	wire [1-1:0] node540;
	wire [1-1:0] node541;
	wire [1-1:0] node542;
	wire [1-1:0] node544;
	wire [1-1:0] node548;
	wire [1-1:0] node550;
	wire [1-1:0] node551;
	wire [1-1:0] node555;
	wire [1-1:0] node556;
	wire [1-1:0] node557;
	wire [1-1:0] node559;
	wire [1-1:0] node560;
	wire [1-1:0] node566;
	wire [1-1:0] node567;
	wire [1-1:0] node568;
	wire [1-1:0] node569;
	wire [1-1:0] node570;
	wire [1-1:0] node572;
	wire [1-1:0] node574;
	wire [1-1:0] node576;
	wire [1-1:0] node577;
	wire [1-1:0] node581;
	wire [1-1:0] node582;
	wire [1-1:0] node584;
	wire [1-1:0] node587;
	wire [1-1:0] node589;
	wire [1-1:0] node590;
	wire [1-1:0] node594;
	wire [1-1:0] node595;
	wire [1-1:0] node596;
	wire [1-1:0] node597;
	wire [1-1:0] node599;
	wire [1-1:0] node602;
	wire [1-1:0] node603;
	wire [1-1:0] node607;
	wire [1-1:0] node608;
	wire [1-1:0] node609;
	wire [1-1:0] node611;
	wire [1-1:0] node614;
	wire [1-1:0] node615;
	wire [1-1:0] node620;
	wire [1-1:0] node621;
	wire [1-1:0] node622;
	wire [1-1:0] node627;
	wire [1-1:0] node628;
	wire [1-1:0] node629;
	wire [1-1:0] node630;
	wire [1-1:0] node632;
	wire [1-1:0] node635;
	wire [1-1:0] node636;
	wire [1-1:0] node637;
	wire [1-1:0] node639;
	wire [1-1:0] node644;
	wire [1-1:0] node645;
	wire [1-1:0] node646;
	wire [1-1:0] node652;
	wire [1-1:0] node653;
	wire [1-1:0] node654;
	wire [1-1:0] node655;
	wire [1-1:0] node656;
	wire [1-1:0] node658;
	wire [1-1:0] node661;
	wire [1-1:0] node662;
	wire [1-1:0] node666;
	wire [1-1:0] node667;
	wire [1-1:0] node668;
	wire [1-1:0] node673;
	wire [1-1:0] node674;
	wire [1-1:0] node675;
	wire [1-1:0] node676;
	wire [1-1:0] node682;
	wire [1-1:0] node683;
	wire [1-1:0] node684;
	wire [1-1:0] node685;
	wire [1-1:0] node686;
	wire [1-1:0] node688;
	wire [1-1:0] node689;
	wire [1-1:0] node691;
	wire [1-1:0] node696;
	wire [1-1:0] node697;
	wire [1-1:0] node698;

	assign outp = (inp[2]) ? node358 : node1;
		assign node1 = (inp[14]) ? node159 : node2;
			assign node2 = (inp[10]) ? node56 : node3;
				assign node3 = (inp[3]) ? node15 : node4;
					assign node4 = (inp[7]) ? node6 : 1'b1;
						assign node6 = (inp[8]) ? node8 : 1'b1;
							assign node8 = (inp[6]) ? node10 : 1'b1;
								assign node10 = (inp[4]) ? node12 : 1'b1;
									assign node12 = (inp[11]) ? 1'b0 : 1'b1;
					assign node15 = (inp[9]) ? node27 : node16;
						assign node16 = (inp[12]) ? node18 : 1'b1;
							assign node18 = (inp[8]) ? node20 : 1'b1;
								assign node20 = (inp[1]) ? 1'b0 : node21;
									assign node21 = (inp[13]) ? node23 : 1'b1;
										assign node23 = (inp[4]) ? 1'b0 : 1'b1;
						assign node27 = (inp[0]) ? node39 : node28;
							assign node28 = (inp[6]) ? node30 : 1'b1;
								assign node30 = (inp[7]) ? node32 : 1'b1;
									assign node32 = (inp[12]) ? node34 : 1'b1;
										assign node34 = (inp[1]) ? 1'b0 : node35;
											assign node35 = (inp[11]) ? 1'b0 : 1'b1;
							assign node39 = (inp[7]) ? node51 : node40;
								assign node40 = (inp[8]) ? node46 : node41;
									assign node41 = (inp[6]) ? node43 : 1'b1;
										assign node43 = (inp[12]) ? 1'b0 : 1'b1;
									assign node46 = (inp[11]) ? 1'b0 : node47;
										assign node47 = (inp[12]) ? 1'b0 : 1'b1;
								assign node51 = (inp[4]) ? 1'b0 : node52;
									assign node52 = (inp[5]) ? 1'b0 : 1'b1;
				assign node56 = (inp[0]) ? node100 : node57;
					assign node57 = (inp[4]) ? node67 : node58;
						assign node58 = (inp[6]) ? node60 : 1'b1;
							assign node60 = (inp[9]) ? node62 : 1'b1;
								assign node62 = (inp[7]) ? node64 : 1'b1;
									assign node64 = (inp[13]) ? 1'b0 : 1'b1;
						assign node67 = (inp[8]) ? node79 : node68;
							assign node68 = (inp[1]) ? node70 : 1'b1;
								assign node70 = (inp[3]) ? node76 : node71;
									assign node71 = (inp[7]) ? node73 : 1'b1;
										assign node73 = (inp[6]) ? 1'b0 : 1'b1;
									assign node76 = (inp[13]) ? 1'b0 : 1'b1;
							assign node79 = (inp[1]) ? node93 : node80;
								assign node80 = (inp[13]) ? node88 : node81;
									assign node81 = (inp[3]) ? node83 : 1'b1;
										assign node83 = (inp[12]) ? node85 : 1'b1;
											assign node85 = (inp[9]) ? 1'b0 : 1'b1;
									assign node88 = (inp[11]) ? 1'b0 : node89;
										assign node89 = (inp[9]) ? 1'b0 : 1'b1;
								assign node93 = (inp[11]) ? 1'b0 : node94;
									assign node94 = (inp[13]) ? node96 : 1'b1;
										assign node96 = (inp[9]) ? 1'b1 : 1'b0;
					assign node100 = (inp[3]) ? node136 : node101;
						assign node101 = (inp[5]) ? node113 : node102;
							assign node102 = (inp[12]) ? node104 : 1'b1;
								assign node104 = (inp[6]) ? node110 : node105;
									assign node105 = (inp[7]) ? node107 : 1'b1;
										assign node107 = (inp[1]) ? 1'b0 : 1'b1;
									assign node110 = (inp[13]) ? 1'b0 : 1'b1;
							assign node113 = (inp[4]) ? node127 : node114;
								assign node114 = (inp[1]) ? node116 : 1'b1;
									assign node116 = (inp[7]) ? 1'b0 : node117;
										assign node117 = (inp[11]) ? node119 : 1'b1;
											assign node119 = (inp[12]) ? node121 : 1'b1;
												assign node121 = (inp[6]) ? 1'b0 : node122;
													assign node122 = (inp[9]) ? 1'b0 : 1'b1;
								assign node127 = (inp[13]) ? 1'b0 : node128;
									assign node128 = (inp[1]) ? 1'b0 : node129;
										assign node129 = (inp[8]) ? node131 : 1'b1;
											assign node131 = (inp[12]) ? 1'b0 : 1'b1;
						assign node136 = (inp[11]) ? node148 : node137;
							assign node137 = (inp[12]) ? node143 : node138;
								assign node138 = (inp[1]) ? node140 : 1'b1;
									assign node140 = (inp[7]) ? 1'b0 : 1'b1;
								assign node143 = (inp[5]) ? 1'b0 : node144;
									assign node144 = (inp[13]) ? 1'b0 : 1'b1;
							assign node148 = (inp[4]) ? 1'b0 : node149;
								assign node149 = (inp[6]) ? 1'b0 : node150;
									assign node150 = (inp[13]) ? 1'b0 : node151;
										assign node151 = (inp[8]) ? node153 : 1'b1;
											assign node153 = (inp[12]) ? 1'b0 : 1'b1;
			assign node159 = (inp[5]) ? node261 : node160;
				assign node160 = (inp[12]) ? node206 : node161;
					assign node161 = (inp[8]) ? node171 : node162;
						assign node162 = (inp[10]) ? node164 : 1'b1;
							assign node164 = (inp[6]) ? node166 : 1'b1;
								assign node166 = (inp[7]) ? node168 : 1'b1;
									assign node168 = (inp[3]) ? 1'b0 : 1'b1;
						assign node171 = (inp[11]) ? node189 : node172;
							assign node172 = (inp[13]) ? node174 : 1'b1;
								assign node174 = (inp[7]) ? node182 : node175;
									assign node175 = (inp[3]) ? 1'b1 : node176;
										assign node176 = (inp[9]) ? node178 : 1'b1;
											assign node178 = (inp[0]) ? 1'b0 : 1'b1;
									assign node182 = (inp[3]) ? 1'b0 : node183;
										assign node183 = (inp[9]) ? 1'b0 : node184;
											assign node184 = (inp[0]) ? 1'b0 : 1'b1;
							assign node189 = (inp[1]) ? node199 : node190;
								assign node190 = (inp[9]) ? node192 : 1'b1;
									assign node192 = (inp[10]) ? 1'b1 : node193;
										assign node193 = (inp[3]) ? node195 : 1'b0;
											assign node195 = (inp[6]) ? 1'b0 : 1'b1;
								assign node199 = (inp[6]) ? 1'b0 : node200;
									assign node200 = (inp[4]) ? 1'b0 : node201;
										assign node201 = (inp[7]) ? 1'b0 : 1'b1;
					assign node206 = (inp[4]) ? node230 : node207;
						assign node207 = (inp[13]) ? node217 : node208;
							assign node208 = (inp[9]) ? node210 : 1'b1;
								assign node210 = (inp[6]) ? node212 : 1'b1;
									assign node212 = (inp[0]) ? 1'b0 : node213;
										assign node213 = (inp[8]) ? 1'b0 : 1'b1;
							assign node217 = (inp[11]) ? node223 : node218;
								assign node218 = (inp[9]) ? node220 : 1'b1;
									assign node220 = (inp[1]) ? 1'b0 : 1'b1;
								assign node223 = (inp[7]) ? 1'b0 : node224;
									assign node224 = (inp[0]) ? node226 : 1'b1;
										assign node226 = (inp[8]) ? 1'b0 : 1'b1;
						assign node230 = (inp[1]) ? node254 : node231;
							assign node231 = (inp[11]) ? node245 : node232;
								assign node232 = (inp[10]) ? node234 : 1'b1;
									assign node234 = (inp[7]) ? node240 : node235;
										assign node235 = (inp[6]) ? node237 : 1'b1;
											assign node237 = (inp[3]) ? 1'b0 : 1'b1;
										assign node240 = (inp[0]) ? 1'b0 : node241;
											assign node241 = (inp[6]) ? 1'b0 : 1'b1;
								assign node245 = (inp[3]) ? 1'b0 : node246;
									assign node246 = (inp[8]) ? node248 : 1'b1;
										assign node248 = (inp[10]) ? 1'b0 : node249;
											assign node249 = (inp[7]) ? 1'b0 : 1'b1;
							assign node254 = (inp[3]) ? 1'b0 : node255;
								assign node255 = (inp[10]) ? 1'b0 : node256;
									assign node256 = (inp[6]) ? 1'b0 : 1'b1;
				assign node261 = (inp[3]) ? node327 : node262;
					assign node262 = (inp[11]) ? node292 : node263;
						assign node263 = (inp[4]) ? node275 : node264;
							assign node264 = (inp[10]) ? node266 : 1'b1;
								assign node266 = (inp[12]) ? node268 : 1'b1;
									assign node268 = (inp[6]) ? node270 : 1'b1;
										assign node270 = (inp[13]) ? node272 : 1'b0;
											assign node272 = (inp[8]) ? 1'b0 : 1'b1;
							assign node275 = (inp[7]) ? node283 : node276;
								assign node276 = (inp[1]) ? node278 : 1'b1;
									assign node278 = (inp[13]) ? node280 : 1'b1;
										assign node280 = (inp[9]) ? 1'b0 : 1'b1;
								assign node283 = (inp[13]) ? 1'b0 : node284;
									assign node284 = (inp[9]) ? node286 : 1'b1;
										assign node286 = (inp[0]) ? 1'b0 : node287;
											assign node287 = (inp[8]) ? 1'b0 : 1'b1;
						assign node292 = (inp[6]) ? node316 : node293;
							assign node293 = (inp[10]) ? node303 : node294;
								assign node294 = (inp[13]) ? node296 : 1'b1;
									assign node296 = (inp[4]) ? node298 : 1'b1;
										assign node298 = (inp[8]) ? 1'b0 : node299;
											assign node299 = (inp[7]) ? 1'b0 : 1'b1;
								assign node303 = (inp[12]) ? node311 : node304;
									assign node304 = (inp[0]) ? node306 : 1'b1;
										assign node306 = (inp[1]) ? 1'b0 : node307;
											assign node307 = (inp[4]) ? 1'b0 : 1'b1;
									assign node311 = (inp[8]) ? 1'b0 : node312;
										assign node312 = (inp[13]) ? 1'b0 : 1'b1;
							assign node316 = (inp[9]) ? 1'b0 : node317;
								assign node317 = (inp[10]) ? 1'b0 : node318;
									assign node318 = (inp[7]) ? 1'b0 : node319;
										assign node319 = (inp[8]) ? node321 : 1'b1;
											assign node321 = (inp[0]) ? 1'b0 : 1'b1;
					assign node327 = (inp[13]) ? node347 : node328;
						assign node328 = (inp[4]) ? node342 : node329;
							assign node329 = (inp[11]) ? node335 : node330;
								assign node330 = (inp[1]) ? node332 : 1'b1;
									assign node332 = (inp[0]) ? 1'b0 : 1'b1;
								assign node335 = (inp[9]) ? 1'b0 : node336;
									assign node336 = (inp[0]) ? node338 : 1'b1;
										assign node338 = (inp[8]) ? 1'b0 : 1'b1;
							assign node342 = (inp[8]) ? 1'b0 : node343;
								assign node343 = (inp[7]) ? 1'b0 : 1'b1;
						assign node347 = (inp[9]) ? 1'b0 : node348;
							assign node348 = (inp[0]) ? 1'b0 : node349;
								assign node349 = (inp[11]) ? node351 : 1'b1;
									assign node351 = (inp[1]) ? 1'b0 : node352;
										assign node352 = (inp[6]) ? 1'b0 : 1'b1;
		assign node358 = (inp[7]) ? node566 : node359;
			assign node359 = (inp[4]) ? node465 : node360;
				assign node360 = (inp[10]) ? node394 : node361;
					assign node361 = (inp[11]) ? node373 : node362;
						assign node362 = (inp[0]) ? node364 : 1'b1;
							assign node364 = (inp[13]) ? node366 : 1'b1;
								assign node366 = (inp[8]) ? node368 : 1'b1;
									assign node368 = (inp[9]) ? node370 : 1'b1;
										assign node370 = (inp[12]) ? 1'b0 : 1'b1;
						assign node373 = (inp[8]) ? node383 : node374;
							assign node374 = (inp[12]) ? node376 : 1'b1;
								assign node376 = (inp[13]) ? node378 : 1'b1;
									assign node378 = (inp[0]) ? 1'b0 : node379;
										assign node379 = (inp[5]) ? 1'b0 : 1'b1;
							assign node383 = (inp[9]) ? node389 : node384;
								assign node384 = (inp[1]) ? node386 : 1'b1;
									assign node386 = (inp[6]) ? 1'b0 : 1'b1;
								assign node389 = (inp[3]) ? 1'b0 : node390;
									assign node390 = (inp[0]) ? 1'b1 : 1'b0;
					assign node394 = (inp[0]) ? node438 : node395;
						assign node395 = (inp[9]) ? node415 : node396;
							assign node396 = (inp[1]) ? node398 : 1'b1;
								assign node398 = (inp[13]) ? node404 : node399;
									assign node399 = (inp[3]) ? node401 : 1'b1;
										assign node401 = (inp[14]) ? 1'b0 : 1'b1;
									assign node404 = (inp[6]) ? node410 : node405;
										assign node405 = (inp[5]) ? node407 : 1'b1;
											assign node407 = (inp[12]) ? 1'b0 : 1'b1;
										assign node410 = (inp[12]) ? 1'b0 : node411;
											assign node411 = (inp[14]) ? 1'b0 : 1'b1;
							assign node415 = (inp[8]) ? node429 : node416;
								assign node416 = (inp[6]) ? node422 : node417;
									assign node417 = (inp[12]) ? node419 : 1'b1;
										assign node419 = (inp[3]) ? 1'b0 : 1'b1;
									assign node422 = (inp[1]) ? 1'b0 : node423;
										assign node423 = (inp[3]) ? node425 : 1'b1;
											assign node425 = (inp[13]) ? 1'b0 : 1'b1;
								assign node429 = (inp[11]) ? 1'b0 : node430;
									assign node430 = (inp[5]) ? 1'b0 : node431;
										assign node431 = (inp[3]) ? node433 : 1'b1;
											assign node433 = (inp[6]) ? 1'b0 : 1'b1;
						assign node438 = (inp[9]) ? node448 : node439;
							assign node439 = (inp[14]) ? node441 : 1'b1;
								assign node441 = (inp[11]) ? 1'b0 : node442;
									assign node442 = (inp[8]) ? node444 : 1'b1;
										assign node444 = (inp[5]) ? 1'b0 : 1'b1;
							assign node448 = (inp[12]) ? 1'b0 : node449;
								assign node449 = (inp[3]) ? node457 : node450;
									assign node450 = (inp[1]) ? node452 : 1'b1;
										assign node452 = (inp[8]) ? 1'b0 : node453;
											assign node453 = (inp[11]) ? 1'b0 : 1'b1;
									assign node457 = (inp[1]) ? 1'b0 : node458;
										assign node458 = (inp[8]) ? 1'b0 : node459;
											assign node459 = (inp[5]) ? 1'b0 : 1'b1;
				assign node465 = (inp[12]) ? node519 : node466;
					assign node466 = (inp[13]) ? node492 : node467;
						assign node467 = (inp[1]) ? node479 : node468;
							assign node468 = (inp[3]) ? node470 : 1'b1;
								assign node470 = (inp[14]) ? node476 : node471;
									assign node471 = (inp[8]) ? node473 : 1'b1;
										assign node473 = (inp[5]) ? 1'b0 : 1'b1;
									assign node476 = (inp[11]) ? 1'b0 : 1'b1;
							assign node479 = (inp[9]) ? 1'b0 : node480;
								assign node480 = (inp[6]) ? node486 : node481;
									assign node481 = (inp[10]) ? 1'b1 : node482;
										assign node482 = (inp[11]) ? 1'b0 : 1'b1;
									assign node486 = (inp[11]) ? 1'b0 : node487;
										assign node487 = (inp[3]) ? 1'b0 : 1'b1;
						assign node492 = (inp[3]) ? node508 : node493;
							assign node493 = (inp[14]) ? node499 : node494;
								assign node494 = (inp[8]) ? node496 : 1'b1;
									assign node496 = (inp[5]) ? 1'b0 : 1'b1;
								assign node499 = (inp[11]) ? 1'b0 : node500;
									assign node500 = (inp[1]) ? 1'b0 : node501;
										assign node501 = (inp[0]) ? node503 : 1'b1;
											assign node503 = (inp[9]) ? 1'b0 : 1'b1;
							assign node508 = (inp[14]) ? node510 : 1'b0;
								assign node510 = (inp[8]) ? 1'b0 : node511;
									assign node511 = (inp[10]) ? node513 : 1'b1;
										assign node513 = (inp[9]) ? node515 : 1'b0;
											assign node515 = (inp[6]) ? 1'b0 : 1'b1;
					assign node519 = (inp[9]) ? node555 : node520;
						assign node520 = (inp[10]) ? node540 : node521;
							assign node521 = (inp[5]) ? node529 : node522;
								assign node522 = (inp[3]) ? node524 : 1'b1;
									assign node524 = (inp[8]) ? node526 : 1'b1;
										assign node526 = (inp[0]) ? 1'b0 : 1'b1;
								assign node529 = (inp[0]) ? node535 : node530;
									assign node530 = (inp[8]) ? node532 : 1'b1;
										assign node532 = (inp[14]) ? 1'b0 : 1'b1;
									assign node535 = (inp[1]) ? 1'b0 : node536;
										assign node536 = (inp[6]) ? 1'b1 : 1'b0;
							assign node540 = (inp[8]) ? node548 : node541;
								assign node541 = (inp[0]) ? 1'b0 : node542;
									assign node542 = (inp[13]) ? node544 : 1'b1;
										assign node544 = (inp[6]) ? 1'b0 : 1'b1;
								assign node548 = (inp[6]) ? node550 : 1'b0;
									assign node550 = (inp[13]) ? 1'b0 : node551;
										assign node551 = (inp[14]) ? 1'b1 : 1'b0;
						assign node555 = (inp[0]) ? 1'b0 : node556;
							assign node556 = (inp[11]) ? 1'b0 : node557;
								assign node557 = (inp[8]) ? node559 : 1'b1;
									assign node559 = (inp[1]) ? 1'b0 : node560;
										assign node560 = (inp[6]) ? 1'b0 : 1'b1;
			assign node566 = (inp[10]) ? node652 : node567;
				assign node567 = (inp[14]) ? node627 : node568;
					assign node568 = (inp[5]) ? node594 : node569;
						assign node569 = (inp[13]) ? node581 : node570;
							assign node570 = (inp[4]) ? node572 : 1'b1;
								assign node572 = (inp[8]) ? node574 : 1'b1;
									assign node574 = (inp[6]) ? node576 : 1'b1;
										assign node576 = (inp[1]) ? 1'b0 : node577;
											assign node577 = (inp[12]) ? 1'b1 : 1'b0;
							assign node581 = (inp[1]) ? node587 : node582;
								assign node582 = (inp[3]) ? node584 : 1'b1;
									assign node584 = (inp[9]) ? 1'b1 : 1'b0;
								assign node587 = (inp[4]) ? node589 : 1'b0;
									assign node589 = (inp[11]) ? 1'b0 : node590;
										assign node590 = (inp[8]) ? 1'b0 : 1'b1;
						assign node594 = (inp[0]) ? node620 : node595;
							assign node595 = (inp[4]) ? node607 : node596;
								assign node596 = (inp[9]) ? node602 : node597;
									assign node597 = (inp[11]) ? node599 : 1'b1;
										assign node599 = (inp[1]) ? 1'b0 : 1'b1;
									assign node602 = (inp[1]) ? 1'b0 : node603;
										assign node603 = (inp[6]) ? 1'b1 : 1'b0;
								assign node607 = (inp[3]) ? 1'b0 : node608;
									assign node608 = (inp[6]) ? node614 : node609;
										assign node609 = (inp[13]) ? node611 : 1'b1;
											assign node611 = (inp[9]) ? 1'b0 : 1'b1;
										assign node614 = (inp[12]) ? 1'b0 : node615;
											assign node615 = (inp[13]) ? 1'b0 : 1'b1;
							assign node620 = (inp[8]) ? 1'b0 : node621;
								assign node621 = (inp[11]) ? 1'b0 : node622;
									assign node622 = (inp[13]) ? 1'b0 : 1'b1;
					assign node627 = (inp[11]) ? 1'b0 : node628;
						assign node628 = (inp[6]) ? node644 : node629;
							assign node629 = (inp[8]) ? node635 : node630;
								assign node630 = (inp[3]) ? node632 : 1'b1;
									assign node632 = (inp[5]) ? 1'b0 : 1'b1;
								assign node635 = (inp[4]) ? 1'b0 : node636;
									assign node636 = (inp[9]) ? 1'b0 : node637;
										assign node637 = (inp[1]) ? node639 : 1'b1;
											assign node639 = (inp[3]) ? 1'b0 : 1'b1;
							assign node644 = (inp[4]) ? 1'b0 : node645;
								assign node645 = (inp[12]) ? 1'b0 : node646;
									assign node646 = (inp[8]) ? 1'b0 : 1'b1;
				assign node652 = (inp[1]) ? node682 : node653;
					assign node653 = (inp[0]) ? node673 : node654;
						assign node654 = (inp[13]) ? node666 : node655;
							assign node655 = (inp[3]) ? node661 : node656;
								assign node656 = (inp[8]) ? node658 : 1'b1;
									assign node658 = (inp[5]) ? 1'b0 : 1'b1;
								assign node661 = (inp[11]) ? 1'b0 : node662;
									assign node662 = (inp[14]) ? 1'b0 : 1'b1;
							assign node666 = (inp[12]) ? 1'b0 : node667;
								assign node667 = (inp[9]) ? 1'b0 : node668;
									assign node668 = (inp[11]) ? 1'b0 : 1'b1;
						assign node673 = (inp[9]) ? 1'b0 : node674;
							assign node674 = (inp[14]) ? 1'b0 : node675;
								assign node675 = (inp[5]) ? 1'b0 : node676;
									assign node676 = (inp[11]) ? 1'b0 : 1'b1;
					assign node682 = (inp[5]) ? 1'b0 : node683;
						assign node683 = (inp[14]) ? 1'b0 : node684;
							assign node684 = (inp[8]) ? node696 : node685;
								assign node685 = (inp[12]) ? 1'b0 : node686;
									assign node686 = (inp[3]) ? node688 : 1'b1;
										assign node688 = (inp[9]) ? 1'b0 : node689;
											assign node689 = (inp[6]) ? node691 : 1'b1;
												assign node691 = (inp[11]) ? 1'b0 : 1'b1;
								assign node696 = (inp[0]) ? 1'b0 : node697;
									assign node697 = (inp[13]) ? 1'b0 : node698;
										assign node698 = (inp[4]) ? 1'b0 : 1'b1;

endmodule